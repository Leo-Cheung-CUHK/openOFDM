

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AI/QYvIliftnts5RXJGSrvg1TqYlL1M8wkSkOysRy8qWhfFWX9W1xaSkDevDviK+T20QHIVswpRp
G3PxYrONyw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lcNSrBM5nZvebPMGfAhvveep3H2yp0xsJcnB/qgeE5Sw94DPwEi/hlIGiNmn91r7c/rFTFG2m6j/
OnLuDWVKIVwwho73ocsN9+50LHkM0cKu1GiustXe1f3YExMUto/ukPDu4kmiixZ/QIkacPiGVc1e
cm6Xt/p4HNnFVTBHiBw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ppV7NrZvES3FTndBUxfHhqP76gqXY1k19OOlSILrN8WL7Dx7d7FVhtBkYwhDt9mL37+q6bd+sAs7
esyMCtC23zwaExSjDLhWE401J6Y7XgHuQ1+X35empoRwYsCJon/ReuUrZUu/NhcuvQy89LPduLaI
9a4mTRM3mgkNSsUzQ7xtxG6hPZ1VJt4sv8rZJVuto75quXVzToLO7Hi4XzWKm465Imrw9AmPleEd
DWhWlLgkaJIQKaDrGi8z1E2Kux6+EkyqJLQNUXrJ6BzZC7AnfKr3prjBYSPHgPpnjkVVX0iWTrpx
jOGuzcA3SuTXzNbBWZTqeVa3NczuYHD123KGsg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ad2A31XTXhVTCJ9eadjDPSFLiQOU7kQCFrrvlT76B7jHPnj7AmPJHDzot+XvDqU/R/D+zBwgaX/q
knabzUxzgdF+6WhDjw606R1RzVqNaoaE27+iW47dc+hozwLtoULSCm0nEBgV72PqMZeefPOoNKM6
Unk3Qy1cGQyPIVpg773LFBurdQx0B/y1jkw2JtTsnMeAWYriqS6AxKRV7cAwsaaQtyzkajpCMoCj
J9vDknZvJMNo5Ld5gTku4sogBuV9BHIxmFsF8SaD9sEFBtTD3Ssfk0lwf7aPSv7kRCiNpQ7wR/rn
Akbnw6ozUL8xeQLG/sI8gBUMPp6C1Y+Ms/MsHw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T66zwGU+r7Zb8iQViuiAdMbNazUQK7tTMIsW16GHXERHg6l56Xu4ZWzOOT3fgFN4wsOsU44v3qvn
cMNuAzEraaUaZMKLuLl1yUP1XwaQ80akKCF4TkJ3jMhaYvNkGbShACRPSjaePfpPFIoiOLkNl7gV
UyqcQIuqSlHRWVtBcL4gaMUkm3GNKbbL5Ur5eKjb3/JPRBxTqFVIgY6/UZajmQscjCsafAhrS7Pn
OJM8pQhBZgNHkZeXyUpV+xm3ddAHsIAPB3al2zBrc4PTu5Z/o4b9h1d59C6EbXorRhLIrw7jtzHQ
M2Y//XIorBVTqWUr+pmv/GYgSYKDht071w55Bw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YWR4lyiIWUAWOF8rOP2f4Afhpj8nObUtQU9ayadIKSNXVdxIA2h5E64tEjyOD/ZyBikekCB2HMGQ
ZlARJZXwcc29nem76cQK3EE03HoDH6hc+3Muq0k2X9DhQzvOjSdvwX7zHwCBrflXaiLXtnVvf7Mk
VpNIZ8yKERWGhRLn2Bo=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QYwS4pvvDfxzvD1lMHTUJ037/1WsdgxRV/iyeTfMTemYhD/apC2iSahtdAVmD/EzhGmBF9JMKUgI
DsLYyXDLhZuT8lvZzK+rQxSBvz4GjKBxvBMtX4bS5jEDHCBXyorqh9PngqBIyrY2tgpSzsxwW0ee
Ztshh0LEg8k+mMBH+6xRcyOqAdM2Ko4fPZdTQ38AzxpVCC9BXSrv4w1H7+BOS1CC8I4JkFTyT3v/
X2DGaPv35nIT4C+/6cWZu756vzyRHwjagJdN9pjfBMI7cOKyOqg+/+hXd6z/zrILdPcMY6I52fxI
NnxVZzIdq956MKI5tG647NXndb6W/RJMWxqpFQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 99632)
`protect data_block
+XG4O21zpz+JxW4xBX290Y8DHTwL5hZ/JC1StlepY0X+6v0niJMJGEvWXE4wgBQduOv6eu5u9+t9
n/dFXJbqafAjbxnZxtfyQrPQk7O6CDEthRkMlLiXriO0Zjir6Y8LkiA+ieHC1cNcwTts5u5vu0Rj
sib2lMrHqo5txmt4iWaaujwiAzMHWJpgFiajmhdhVXeuiGaUYzSAAP+P2NI9X1ZpxK30dvHwyMqd
YcQcV3Oi9UsY4tqjdBqfHozyaBAE69xTnfdSbLz4TWxGDsII9JWISkrti/BaEi+w++6xm+5Za5ND
4tyHXvp0JHEhWjhebm/siEPovijiBsDBr48sodCoK1ucXBdvpawdxGZsfLRuyKaoALGZxdzHGZdC
rnLJYSXP3zzITKoUeRdWJjeiqsZt+MJyKDhUEfDZ5Cua6QN/8Q27sSVMaTgaBOFBJdjy8WD9QrpK
E/I5JFW5BtIIbhQmTtC+hCQTutmprF+W/vwp0EoVaGc7WOLGExVKabdoN5EtP1jOA2oh+Ela06lE
viXqLy04EBTwuggCzLs2Ocl/mTYsvQI8Vk8kgEXZ9eHi2/kbxAwd15Xgvog1jj0VznDFNmgZQBum
VrIksTT38rLxgy4zVIN0Gx/4T3FUT7TLheO7CKRUu4WVD9o8exzF/0zq9Mz3anFXOorduot6Y6EL
2uVLIftVAI8wEaPRVhoE94g10pYGS9PAw5t2hzqn833+JKFxMPxzZ+C/4Rln0V8yE7dmkY3q2y5p
pET8gUifvmYhkjYibdz9ynoCHcb5LbsQatk89NM1kl6+bQVdqbko/o3KA9gT7Q0lkLUfqhMvuWX5
b8hJq93WWzTXtJ5WzS5KkLubiwIt+xLYFfskgGG2U42wCIkWGnpTUgze4xf3m3A6M7ZW80GlRtDw
kgiXYfqRS1/eeG3DFiBxLhht2FBgXGO56tsJeb9meLmTD8BvTX+M0yN/K0piWP9Yi0pTW/sng8rO
aX0UwWJ19YTgk/DvZmpHzQF8bbhyoAEn71klzx1HSqcqoIRyF14Uzabd4f0Xvui4dUdkYkGhH17U
itoQ7AiiKVQ3OA0yAyXFm2nwOk5NFPQq6e9ARJdJcq5J3vyPFRK6pplf2lGO74bXyC4s7vCYU/6O
kLKrwjcsV1diP8mEQJG/1qIiw7ePzZJN0AbTtZVxZj0NpoIiGGnR0dULqGgP7g7e0yCF3yTBvaqS
MUmxSBvEFtM07qe8G7yhaW9GsOFvW0NwrDTWUJuZUitSnEW8zUo4RkCHNScUappJ/ZmvUuRi+6FH
VJvYOgi3hUori0HanXxNAv3LoFXAnPPPq832WkkMm7NHiQl0+FjiwZQS86tJLFtbn8JzO+0g5c8H
fb+Utxzh1KcfyPtCRT1h4n16NlNOnlgjv4DZ3nsx71GqbCJrbPUH+QrhpnjM/srnIu0niNQC1cWR
2yGDi0czsK+LYjm1qHKhE3XLQhWKNxjh2wNRrRYWW2/DozGJ9jKup/dw2gJyJ1uBAkC7Tk87TMea
ECt78qhdNUpDjkyMCIvDogsYXgrOP1Fe9swqk43PuoGbvmz4YnnC3QZc3IqG4QCQeA7TDWIovpI5
zH+Tkp+/o9jP7ENzaYE6un/DhL/uN5kY2PNgEKFR5HiN89IFDukFMii/ZQYgpFLHWHOlrDMXwF4h
kFPs1HZ3OGZRWHGHgiyYfGwc4Bi0/Rsa2W+5GByKPQlcCk7AdC7wjVPCsAktcnQd06O2ahAa78JD
iCbmfH8TVmYwr9nDhzAeiJJgdxOOy6x7wd8Lszd2P1sbilfbycCwlY4dGbwaqcEGJoWjhNAcmqW3
TS9cmbqbj1Jt2nd1QVclqQ6u+4jz+dSUHcIqLgGF4A+dRGbJ2NpqhlKHpdf6jtv1Hpwdj/Lb6o9K
wwAKBI0EzFztOf0A0bBt/PX0QxbdONvQ0hXbZlFEUlEwsgPApZC1rqMjruDBRR35hg4wFquuNE85
7+H2Nwc0vXWGaKfvLQjQLqagoEgjd1AnulIHB+YYRrxDQZ7iIU0iyzPy3uRYPdsnCxBLvVFHypqx
laMYwnUN4ME92Iy/h5zX8raEtt/AtZNjE9cRpGDCiUkJvyH5EUZFF5irGuzeGyeSY2gyxrbrBvA8
iAoW8vAgkRC2ttIAOlwFHUzIxOrt+vL5PMx6ie/h0UmHh1i463S0/w/9JzZfHiOLN4Rl+K7dG30g
3YsegGxuoa5lfBVA23NlLWG6SewtoksOHw09qEYNmw7O8SwR4ykJ3l68K04dnT1SRRIdkjg6yeEU
JUxol4RkacWW9RZ40zqbOS4Oj+aHRMYUClkAcBAh+pzFqpbPbtB1H13YgEE1Go07yEQJ/UhL05Tb
awCGc6lfHf3fXCsiw9pn2D0vC0nYkSOP3hRz8l0ztCHBn5/PswZ4p6srjgLBM8CSRTkJnHVAuSpp
epBTzadLVYet7RJNxrQ/Gz7WBS66CFcHquoKuM0TZFYsPjEE4z94KBK/axprYFEprtTRfFAosk2l
B8PnjN8B8GOUWV9+oD7EWCe+cqEPpfvXG0fFSK0kfgafbGjPRvmdw7/mztjXd+vZ+aI9j1lHtnkV
a52SmVTBr/MYGml+0qZUV1G0Ivw9Y14VKNEEF0vjb19huVsqw+p8+DRDe/8KwAuTUbaY/BBrEghi
jg4EThhxVuW/rWami7bR3iLJgEtvSmKXH9fRU+YlMggcUsHYGojg0R2F8HWAgd21j16YdWOhLWnd
oijIJw50rgtIO7tyFzSdOqmBLHzZ+9wJ2mVK97lnoQNq656gpVt0oW2JPVfgv6kzhDuKnN/fbbkY
Sx19DBzvIqix5Wazn8Kfl5U6JQSQwV5dTYMcotTBWG2m0X/gxJrPjnKFRa1/4lQZy+xDDWvFoSvz
99qMObAqPWU3OI1UmHsne9NpcXsBnJyDeBuUloqg+09ejcdqV/2mHCy+Wjt+IfW0/LxRm9FtjXsF
2OAvFZ4+QDpjmK3nkC5akI1Am/GyOSjQ9cJjnnfFdTpNVCr3L1qaZAsRULDCR36t68GUImHVIJsK
2SH8YodOzDsx3AVJeLD+Mt5MJSiYr+MhZhDIzg8fBHvBY718GHOKdY1GczfBMNIPqaYd8MooFJws
+xmhwCnUdFlubp9M0UC8sHylXbX7Hgi6C5JmI4BFpfoTD94i0bFK2HQttopHgB/SfG7RVliDHyTT
DXFk93vA3M0b4pJw6hsy/48imoHJZvct7uOm0EIIhoc3YeX5KUPqJQLNcNhqFtVuXLMLJK+tCwTM
oK40ua12kWOe+tRguOz/zyb6Emz0R5ZqD6KOh67GdCRBoLU6lqsG8QdwRSfX8NqHfLggLuujDEQ0
QosZpMGercordCyvlZYWn1XAtVK3b11QUjfXUWX0y2xzLYl2EhQHQm02YxvYrQf/dyjAZjhQXSmZ
+oFYwlIkpX6UjGpoe9ZEt1E/uV/WD/hwfC5fqEddPPleqXydsd8lGhdpyhVa0IQvE1bjyH2PupJy
+DQDWcAv9xmTAt8ms8NuOR1TY0dFUeneVqWNoKeouL6kd2kaJWDyYq6Y/cfldF5e3DwNEOYWSfuM
z3RA71GHxQFV6Bw4CQs5M+u2wkXd+hF74NZQ8Sz8BnV5kchTjh7jBVZnapXX1dpGSh4xaS4u56GW
xSsa5zU0ZMO3jF0b1sWmH7MLJMvVwOJpqyoIpCw2ToMmYX0Nlaad0XXOab0rGDSleRyYk2loHrkD
+zoHmynq60AerikcVnyK3nsdmyKENUHCVnAX2bXa/cGtPZhfUMWoM91OcuQq+xzpl945dP5guwAM
2S1EPGoJrd/o1YgaBr3uubeMlnQTbqjnJ5OL+b2lpWi/C0GGk9qCdnFk86xHblYHPN3pPhcbJzs5
/JojSIS5hBze7knrxHxpOJzyzI67oPlrdOMhndXLPxy5N5XMjo9pTDTaBRGhtlFDMBzH4Y2JhErh
SU6wIgKX2kTBwOi/M1MVOaMVh/7FlJUlkEVcnvOGR0LNCvfk/5jI5m9xGjE8slj+IDBLps0QQdl8
pTLQxMvYSyA0su8AJBE5S1LWQXp9VJ8iyKyjfuKchPCNBcKB3yZb/pBDGKLuMgg4VbSGv8h4djZd
Twri0dXxyx7aeLY9O5aqUAO/DornvHCcGhr9b3MWBmLAKFGkvwn+P6HSkWlFTRbbfA7OZUj1GUeA
+64zi3eTtvb1K+vEOYHJQ/F8Skdrm4pyspOobYa1ge7VKyzPHg4/MGS5t7L6AvEXiTghUQb72y1N
GpkqaTwXZCdmCWfOf2C6YJTPasx0/wp2mQkedgH+aaecOhDzlMR+Umj3UYmueFX1qpjwKrUddcOR
zXeNQriXJN8rVm2iEn5uI4X/TuQPav7TYbehrQx/u2e3Gg8kWqbgyWDd+HKQMUCC4qmRY87cEnim
ettqhLyFOeN1CB+e1MLvYx66d/nq1Rcumd7eERp7sLTTdLnJQcBKTcWzks4IlV0pXrtpglrwMSj8
ZaaKZqkoVXYyUA9B2DfuiL1ZwEmYGnNNTuZcxUtzRBknxQXyMA+FSoVxPx6O1785c0WXbncFxDCa
lMSExceut4QqTT6vNGENuX4Mhny2rfbrb1FJzV8MUV3t+e5mys3TpfRqeSy4nwQrjASP+/PCWQER
UFYrHtuBaGpPt/B8jEjVKepnycgHQhcI0GeQKnPOEoZRRLx0C9vdJ3atIm5YrChNql+TfYYKRs1B
f7oGBSp4Qj0Eb1X1oGjR7gRc5nDOrVt/s+nfUZ7H0B8KRsKANd1ZjvlYdFGXto0YtF3KkH709VOu
0iDJXEQalomOGxyaBQIdOl6pdzf1h5a8FbFLBo3qsmKrqxTAKMb68Wis3TbKg2mSLKd9yf80Jw6d
hrCjC+pY+Jk9+OJZa5u4Nld8U1YYpZBcJEwLhWseiCz6Ffok5PNa586HULi9z6Nt8UiX7t78skYK
Lfg2UOWtxr6MBpxt5RX/J7zBo2x5fAaUfNu7LhE1yafmE90wrGwmEbEuILpooLVCkvkJCNa88KPJ
EStjIohkLpZFQkdb4Py34z/gdadqVU2J69mZS78QoteoRlrJnduWCsWTQ8EitkpsDm30Q/+fpl4h
Lwt+90aK65OnlgTb4gve4R/f0Z4doAaav9zA9EHV0+1/0wsjP42cPHEH1yO6u6U1XfgTBPb12PSD
wDlQfMqUnQE5Z/gD90vdN7gYa7tlnmotAbLGcRwDU8HX0c2QCJR3UgS4ljtR01ivAy8FNYIJKdRt
0bIrApgiQXOD1dudPX28Nnixapj80S38aiiZDdlwTjLlqIaqtoskJ6eEIugTON4oCZm1E7AFIxkt
pHpQgl+CAcNl7kFdiUGKTtBbVO20t6OynccA0NVtym7OOv7PVinjhwtADAANo48DlLTAQobTPN6d
MZKSrSgDifC2a5Q4bN/98978VT46ypLTEf5p8Pt3lWjZYesRDBnkHjZDkdViShBRVMagjvHdBf1i
W+L15I8x+5aRBQzUaDzZfWrK7irM0GwlN5sZUwrsmDVfymCU0Ht763Lpm/nvdOFkPT2xgAVGfPBH
g9H5/MnJtgFw8lrCubMS37zHv0XXX7wq8MUO6e1iLGVJh6Af1tGdIAL7jwB0JlieiDo0fREjbViY
uQUvAe+igz/8VjrN0qQzniHzlAvGgGvWyvu7VvcsypT9zG1LHN4DJLJ/bRF3WYu2CTYHXtsWH9PK
D+RrQ47o8+VGX5arx6bVIQAU3U3iTWWhPVKBnYqvM9gVipYvUx3crjgxzsfS40fauy1XHqQOG0/H
oJDRBS/0O1Ayjc/tYMLjL9Sa2A3H6L6l8WSG3b/r80SnIypMcJmWwpbwtS/O/vpMWkXEnxzpRDf2
N8VQ65cyKQwhGiepX31YltdYP7He6joGKMNNF8mQuT0SrhuMqxhNzLRTdixou9MwdwfGauZGjW4A
RdMAyHGa1Zj5HuLnqpnCXwzbxOVB8GMxz+VFlsou5qZnY3e5eOOLoqm4/lX/PkWDnu2QzZSblcjI
SRUxqpFL3sa/S7OPYiYecq5o66IYzl0d5h6DA/ZAvy60WzediwPHMm1+mbfABblQSLUWV5ITCIXI
Q63yb1VyZjZMhBySkfAv6+lWHJBv2NxHQCp2Kpx6YvhfQe4yGuF9lCkKsuVQYUFYSHnmYFT5Y4lx
htx9ocIJ8vAD8y6r8Q7lXgt7y6zGSiUAJxRtjfL67QTQlt8+5Ba/8SU4e+UNdd46XkW19WERl46r
X1fOag86asTSmSrDlai/nonk5JCv/2jleGH5Rf6lAVNVhCQJPKCNnXyEOvJmGQtdF+OyQcJUZ4Iz
BagGq5E9rchL3Jf4LZxDY/8AfSp688BFPraz8NEArNnH3GLa5uASMnstuOkHOW6xjytjEeVCaRH9
mOjhe3sTcR1znEdOLLypILZ8fX1sQsfvV8agEPBPLB/LemdeZUEvUmkATKoR2x/urc/L4F2eWpQp
Q6z25HDgY/7fvGRQuX4w7VYox58lp+NIJb+goJfi+NgHms+WfORVOPEZ8JuAZGJ1MUYFg0W4qFmq
mxs+yWqzTV64S0sFKjGixa9aYxM36YPDkpCxqOCBU/aEhVCIBhhg1Jyhj9bfD664dugW04t/gjc/
OuQYv5g6Dcn4HvEJ3MvwjAjJ7fkk3aYVhe7P2k1qrUDELwlXpcASH+4aNrMR2ngCvtShZv3Jc2Py
hsIB2bIa6Dnan5U0gyNw6YlXM87kTHMFF1XuUdHK4E32y5NmOfmpIE8e9LFem/QSXbheczYNbTBs
XgOGYmVOmiQpqSDrJJMlEYr2WRzgI5+qE4GE0Z5HAo3daQh0ndDphQ/d080Yi2LHqRLbrqzWSwCn
52UjP/rvn3xMxqfC6iR+D5kjF7OgFEV9nClzL75jNovWs1lZiEg33gU3+L0r533w6leC0/xl9Qtf
S8gvI2LgbBDQkO46oEQ7DVy+oty/IZ8HEouuP774ygGEf+L0A/57co4bqwcLNlbNcoRrdoJGq3W/
dsvy1wW0GLVOd/CEySRCWwCvVZf2Vx8TtwWguw7MiOhtxzpRU1JCaNsSA+Xr+xDdvQ02y3Rh89gj
gZ0ziGwirobyTleO272XIxvJO0WPrbUBOF8VMh1//VGi7SB7IlGm5XBh9Pgm+bkju7YS0U6ZmGrg
wQ/4Nvff0/O6HMpP7KibeGFUgxaX1kBj6HPfwp6KfCTAlG1/uKPsjFkBFDhb07gYqY4eKB8vTuA1
ekJq63rvUYikOy9eo0DPMGOMbAprO6px52wVo5uuysMbYX/Lpnrt4OwHmCVnsb0Tft7dWdlSKLLy
OJsMxZYYe1khLgUGlyibcSXDNAjXHPXil5lwA6kwlO/DbRi8paSIWpaIjamQYSgw+geQuEJFPgxz
b3YdJgKZSYR+J0upw4DVxHrpZB9CL5YspvdLl0GmGm5RLIz4Rl8Tp2Iq02FABRSCycKbzA27c5UD
PY7acBwy0QrY3KdGmvE1iF4yiVHzR3U8ba1r4zhom5HLzrdEgnSJLuOUU8y95UugYdsXthw5uzFf
TLFAhueBijWgQR/lQDYatdFy+rPacq4/nDnsbX+IgeTRAVCtLrz9DQkSiiZEhnj0qojPWU/LsDq3
c6b/vD3rdhaL11SbVZG4hefr3Cvj0yuOIAEYhluOs+RSX7BgIas6VnkBiw2nS3teNAQ32u679ctc
8C/3/sZ10N6JTUTHCZPzWyRfcoNVQgmqIXJou3XLQa/xOFQvRgNCSCSFXNoUzKFYD13PRr5CBMr0
MEAPr7F+5tnnIWbq3teDgb0PX5uGUW8qO2SxbPwELt4zh2x29sQ7yTmRwuV0YFeQzAHHSColavdy
9JhE61X6SOq+So1UQlF3sA159w6wAL97cEEw5U0PNbsmAs7QInf1gZFTpewme2dpK+2BHCgAaGbE
+AahoxTKpJrV20bt8REdfkYkTP1JPzI9arhOlxedUKoinHuz9eXUIrY0JiLtHgF4reZuYUH+O/mP
0Yy8Z5Oz4lXV+5SV9XSv16/H/lx0hX+/+zEqrfdQ7Xc4FOa9neN5HlXuKAzzbX8JRZgH5Ty/xC2t
GIyxpIvFuLSS9LlXRZnl/0xutH8yYSCS7fSrNbBSFj7LZWSATSdUdQxzlh3+kQJgTjFmzgc4NMbY
QD9prictkXqQ3YOTS+FHo9EoF3y8RD6Gf+4lD2atL/+0MqwY5l/oxlQS8uWJJtSSNBmGQMJq6INh
ck0/RQfQ03yzyCkEiUvPx1Bcrk/6nVt8RqZiz3y/PhWsNWRHRm5XrdVg3dDoD54YB0O42wgJPS63
+AG/KtNtIwJu/ShHvUAIcb8zB9ArMdBLUipvFPkChpLrgkAtGRFKYFOHszoKHxUbyf3HQWngm4Xx
evyeSkSVBRJZCENU1TjG7kuXsqieamqK95vQwFpJ3Wa+TFdySrNlTHLavMXXfRnp2WHm5Xv+J551
wIuCyec1A036Pb8ZGd8NgJktuNv6EuEJGGVhhiWlaWWFyCO8Fa9bDdRKlSK4dYjiPO4S8Zq37wkh
gvcbH+Ns/xobeauMmhzfEDsoKMwkm2cmR/TkJx7rmmfjfkqJRGX5osCFerMw2g+vBDs1/UMz/83i
O+8Y51kFwKKuo+AZqL9g9/SR+ZKSJ390ajTKf4rbHC1X38Uo+GhmL3xH/61BaFFm6D/t5PhHT3U2
vvHoIZI1135hAcuXXq2iHR5eO1AOone78Zs93ysXN8ixt2vkb+8uZ9PrUxrPHwPcgX6f7u+DNdvj
M8kCANvVv45bbWV8yNGnur5z0VoEHnkFZ5Fl2CjF8kMROYWspJFGLUkH3ss83bD1PO930KiXTIgt
LB3onA9UYyGKqOJDqQGkT5WRexnSCos9zToNW4LlobzzdlaWu4+LA7aZylsxsyiUj2j5yw57iQ1Q
SGvTlLn2cM+HdKQox91YT73sqZa1DfGo2DMG6vtOL75X7Yv+hrhl551ihiIjxs7sBjULTtl1eSCS
BuIy9aeCcxYEa2x7kQhM8/aZGh0C0OIt3Sfr+yxWENqCJuIADe641gNjjq8825mqgchdYLFCwIOi
PfxM0GzG/e1IaotUZbPLWEd6rX171nFjMOqFINu9jhFrrjYCRG2VcRG6irdyvAbz+H0nds1hagp/
DaAirvxvPxXYioAU50HaYC/JLcvmxsMjawoy41HJY/GhTo8/33NMtCGa2daKQsVN1sI9RUch/+7M
sWIefl5tPR6kUJWz1VKdOzkhFdiuz9nax2dUo0hXzcdaE/9Ql4aRDjdDAz3QJmhZj0PHGsIpkynt
SHSAWEG85uboH7Z74rOqKAa9RrPz9x8r9y8edYtx71br8ZrLDvE8NouI6UBliLAsl8lkxulGI9NO
EYcr644kp+1Fm2Cx8YNTgHJRzVMbV9SVsxkwZyuhOm1AzqChb2rDDqy3nKPJ5wFMUhDos7ha3dWt
GeaCboGPdK/P4qqO05orUio9ttfxWl+j0BDyQkio5EQAly8NLp76IWdWWFS157FNr8ZT9ips2A8n
1Jy1cqrP9UTXmnXRsRnQIWR+V5P1qJEV3oj1Xy4HmKrEThgN8zRj3aBs9gNgPE2fi+Ndn580iWkw
pN8+0GCVJYuDTa5/7RyJqHX9qxRRPfuyQZ4+I161ueqztA8UrlLTMEB45CHz0ZVzjZEj+PPFqeCO
aGkQ+KQS6rvTcdLTZ8skS5LFdMnlBoJL/pNTERTnn+RWHUnntVpM6au+pmASsrXs1HSLutoq5rjC
N/XMZXJhk7Npe65gbkssil6v28yPFl7t4cc85WaMTKsKTEsiZEJT3xYM9mQgUN7dY+asTYL6roLs
7TusOZgryXBWX9peqf+weBS635whJoo9k/xPUCWXt4w4YvtzgQG2XdFD7Y3quZsJHSLaYDGJrWHw
+He5cHuw+CPjFSRKoD9lF6AJcbO/2dlgeIzTB7FWQuI5Sz68EzNV8LO1fzSFCeBcrdKQvGQcB6lE
3Jw5z/u065NPUUDK10Rfe2ZkJpcxVplQfV9Ze0qO+7iQtTG+VS8PJM3w8Y+uKOIEARmNe1VE8RY2
Wnn6ITS8oeT35ZqkgO2AEvx8S0WJX4EbUDcmtUa8jtGwWkTJj/8KBCC1UoU9FjwJb3xCdB/+R+LA
iVuo13O6LCMEi8iXItcpHuZdVPVFPLQGFQ4M8E6QGnvucxHP7LMkOC+Zi0iDsKe5QNDVT12a1TR2
xDLnJxoUI8CCi+9W85aLpYdQICeU5Qb1evVNzb0KhWl+Jdw5FoGKd9dazIWF8/eqsd2c00xRKz6c
MmMzvic6uh/Lh248d+qU2Z+Xm5kxrPkAoBut+TBZsrTeHTSDmp3D2DAUKpIvUzC6sB/oTbiwlPgo
ziduVWOvt6jBJhwYIbNSvc03PDnlDGJ5ZbvREtCUIf9baTy+cFcPMJjDO1xcUK2+6N6ZRIwKs/cB
v/UoUWSFx9oxBDpeaA6FirMdjBOTj8Y967iVb70Rv/ligqiPnl84QNznHPEkkUzZISQYeF3Rb6ed
lWD114oaQ9CtiQYN5rcbONDwuljdNUx0WjgWMmEG0tfyP2f5uAZ/72KONkF3TjmmkqHUCX5ueUNd
5UB+ri9wGP+03VsW7iHGk6S/wpmZc0NX16NG/YFz/DRWA8vBLcyO1swCLJivTvUJYhfGuaMO3uMa
Den8EnE3ilyiMVFNYkKlK+DNScE/h8i01kW2sn+ve17N0S3cw9Xss+XNetdV/MekLE3w/K0S62ga
W4ndRNkeONUnfDktqTF3SAdIXJFMmQNd1vsW00lXmSH4Mlb5xpBpCIpym3bIppSTqq1yiPO8FB3W
aff4hHXcJ5RR3M8gaeS1Mgkxirk/HfkzjSeCEML0lTe/OyMoAH670Pl+8oSDr04u6OTNdeNlki11
GrILR04OPhNXExvX9UPMi9qTK+TTqUw7Dgf6SKbuHLYNb89a3OneCjLlGBK+NrgkUlmaCaNAB3JI
Xli02RNMBsGQI4IzbAZdsvK0AcJ/3sVPiI8oY/84D8ZhP3GHAVTtIqsDRUdquZB6g40URPeOQhaC
rFNWa7OYfja/YHXZbQmoooLqOahIdEBl7lCjtxYDFkuP6ut0duETWridhc7Fntsrh3wDiXNbDvGH
+iGW4xgyrx4XHWIpZf3AiSgHP6ETASoS0OfyF7IejR664sn+yGtn+LBFIaRUj3AhGPxpkjQ91AzC
37oucGCBb9ObJuqZQkSJVLJVk6cgX0yzjcryjg+6q0oK2Ec6hq+efrASDaTv6NcEEAcK4PxTYLHp
CKy5AeEngnPRMGpH1VaLr8FI1ES/VD01WWWF6/IvJfWwSMTkYJP2gYE8H48Wp95BlNOpN6zIYAeZ
4pOAbUyApob0pqrbspt1BoJWK7DfLdZPWeK6cc0CS5scRi2jtvakInTK6BBx/ZwyPiKVeEFyUZDy
YsRmLbpek97/Nl1kufQuevKEvN4UL0RKO+kmYaGUefjEut49qyxFbq2hknAJqLyS2n/GIC65XYUT
OtBImsmftLhZZrNLOlYq/hzb/LiMgtvKm38R2hzlbM4sGOO44ymp73MOgJ9uknhxKNGxMz+DGkb7
qIsX6eW3oC0OTNjb5X/L9DFnbUK9VWvX0vfoMHjUiRaM/HfFz4vMDQjXftzLKkcnJhJ/LfnVAux5
nSkNVpbfUyC4Juf4rWbBioZOESfWQlOlbGbYjUwH6VSkyx//Cnia4c8snOqjwznt31NIq9nzhrwc
w8h604iU8s58gPU4rmLq9cITLgjqaHV8JuJCUEfdFVLShz9OCxPhwyOnyqVI1vOWpbCir4ZkVmcw
0p+UMjg0pVJJLho0F0ez5SGe0+MTyDEDgRqUHwqLeDVb0wo8fR6zjuDX5/+zLSDGFiOfbrNbmI+t
iRqLYG6O5PFdn1Cp3UVwmHMVdeS8MJW0S14Pf/9AEu7ElRkfrtQi0v1tCud2qRjUm5rkMHBul3+4
DyooE97CAG8ZVnnWJ+elR6a1xRxBZe9TzCQ0/bK4jFtR3FfjA3IblblEVhR1qHdz4/A/1KBzS+wF
4dSFsH6MVJcf2bQdHsbD9JTmGzTN9U4gVxTKVGYtlHapfIF+QeQ4gZz4xHnxHJ0PFsqPhebztj5j
sYYNIKf5J6JXiibkCulDHNULLO3o+W+Cz1hiPCxltV9TX0M7M/9GZyAP4nbGe6CmDDR1L8le3dvl
MuCVVVbFMPT4C14/F8yBVN6zcoPjqGjnJNayd9/mr5yioDpxOUAxc2vwN0X7MQ/zdh7Yk3wYetzk
ZEx5VqJeYmtOOPrMj3NG4c9frTobNqTzzC4ZlBUdLyJq3q23UvZBiVJz2zX5HJ5Zl70xrWZGrb5I
pJCY93dNT/vB6fGJTaTuHnK31LizEfPyUhPPOJFZkIMwxjSnKMDq9nn/R8i/MpEFLOuG1xRIUWVr
mLFRCaLZ5/w/cVVKMW4Y8tgSEXUYS/HFLYWni6ue5+L8uaPIijbqdlYkNvtYiMqR+4B87ocObyCE
r16ajBhOa5wi0YUQUiKJopZUSi6tmRj+d6raZF4fj2ANupo9fMcEv3RAra6SDwEUbYVQtu+wHzPT
i87GpXGqX7uzMQS5HJPSauocwDjvITBUm1AOEIMyik5t4dD3lKGlf+YKEpukxRPVy//lKJzpRN0K
daD/0FRSU7X06e3E1Em5c+MYjZX+h17GualkNdNobGFybziZoFsn/cp3EzG3Zy/AIiHSOSSuRMEC
/6SORJNYjPCMihEqZqL5rCJu5nRu8MZSEQO7jriohbJcq4L3OOaQhIw25+4kpZaTZtO9H096mNDH
5vzXdOZU+vuJYYSYR0sWiD8U9J36UU25EI+UbPdLKC/hZ2PmUSJQ53nFSrvrcgMMxB9ei2MINAF8
M7OX7xCB8kcR8kHx1U+C8GWN0jgwRJqW+HrfWEuyOQmQpe25iMJRgTxGs9JUIYaSyyFbTMSRB7nb
hhugzaPMNldvZGNu0e8XCqazzp+gO0utasZqXZzB8++acFrX0dGUDuyvbC+04qTcPiUKhUXSVZOS
qVS3Qgh7R2YAhnPV9iDoe6u0yxlDZqDXnGqFQxwgJ2uaovkhofnmqawbgNj6sjcYu0fRM99EnvCi
QxJj7FCywjopM6n8BAw8qYe0/UGDLanZ8OonK4zcLm77HhuWqjuKxibh1Y/S8vjSAhWOF3idgiGg
HqvfMDw9TezzMxt3d7l92HdofYYMFLy8sY/hiylEZArRZqp7MP37HUpJ8e053gpY/6gJ061TuU23
HhzCf7ruYu8btGgpVGqzahMo1uTTv6DwKEEIq7bbZbvV1FDzPgMQQOEGOu18p+D0Z+xtSlaKg9i6
l4d3BxoehgpUjw9jZq3E9X52WbFHr5qlGLXrlNtob8aBC/kYcRXyScmSHsFntKIkBBMHFu6HN+7Q
YWJ3RfgXcUv3dvTU28ZN9htjyqy+7WFOTPGe2T21zshetXX9aFvN8mMgIWkye9dKkO3N+jdMu3b6
J+KwS1NQIfjm/b9VpKjqmCohXacugq52f6RGl1IQtxDGzgUgGqLRY/ik+XwPCtEmZW8suTmR3S+/
Aoqod2+ADldl1LwfPun5ObKVSlRlVBg70TV/umNIQPdSzw+0WOrpGnd7OSGXrwbFJOsOXFhd5c4Y
zVp6U/LRvCct4fN/cbZ5P+qd6c8Xppcx0bn8XIu66piVw9gridhHwPSbYQccI/mStOSEz0Yc/baY
Sa4brDNZgwHB55ev72Ggk1pad41rY3v/k+IJb6mHRL8aripJtutfHOHqdkt9ZyyZ7/q00keuLk87
WGiJiyMK6fTDGW658kOqvWo29GL8J/zYZ/f9SFhn0KvTzhER/54DvdhS4aRkqZabe8A/DpMlmvUK
CDPq6ozxUlnrTWelTzLpwX+sbhegeqYSP0kj1aDeegCRJ03mT5wUutiIow0G2UpMFtgPHnhVCuKx
PQjPJBul4bcTt+LeCLkjX9Elt9XR5ecJhiNljXwjqAqLrciWJqOwLPE02DQ9D9PFV/q1Q+H9JZtb
N2YApbC8yc3eRWLhBYTUEe7GHWaqbtNkkzQuWZJMEHtze91aT6MF/7OykKGxx7TTvc4SVvA9CY6S
11tDp6vB9YHjUpeJKA+FsiGWDJm8wNbYSvhjgpg8tC6Lb0C4k5HoC5WIV8fMurldCHoQN3wpbCdZ
v8CMyuwrTvC+s4ZKSxC3cJj7hxcFsZz0Is2PQqWDkfBWHZzD3KfDFCaqa7lADaEdWhzEybKm5N+W
sCbUIYQlviSDo6PE/7AB3RqoWf+cJCcOoAW5gndHIYoATEoLDontgsotkjdFV/SEYIAlY0P7Bf00
UB4ZpqwiVxQJiZUigWtvCTSZ5Wm6t5go1vZppLX3HOBzvk0e6Q5xDuZTSyqBKuWHSbOUI97DdTRv
zd2h3wIh2ClDezyksf5cY8nlp/apcmtbygGUAds8gT4XhLsh50dZL0m6MXY/tim9Wy2o4Fpgn8gA
pF4XxNUYcb8cGEkJ5bFN7rbJj5UGcEEU8BED02MS9YK2TRqOT3o3ZLFr2oI+TinJosnWzoSf8gv4
dOvgbe0jSCU4CTb4QBWxVLq4Bag/ZgB8VOtUhVmK6B6+3z8rIVxXcpvlKMfOstb8sTbXLqXV6j8t
HjOJm8z3FNXRAsnAHkuun5ObtKuTi2wZC3/dHNQV5z3lrbdTyzleQ+9oVS5A82aHt8VOOUz16w2y
mIwkgReOhgXkkYvNtRlFxzkb9Ri92oDhSml3+u9aLUjPxJjFUmmprUAjrISHeUdzEsCKvre4k3Z0
FqnmEnimqhEQWBxfy/Z0vGUcFtacTcaW0WKtxodabskWvgctFp4Qz1bz64KqVdsPcEJNoweXFyO+
UhJCC5WLESaU3lloyZQf9Bo8iLHUhfstT0H4cKubIMX/x1Q8E/Xmpg0pgatyYvqI/HNz/fDwqlID
QewSTC8UX7JIeqINXJVTSwUebKGwgv0IIkht+F3FleNEfGA3Phv2g35xhKdZ6aqb8BDw8GIps9yx
8dFWh35b5sM9PFpwvMhrozMjaGJWLKV99cTVJJcl4gRfEEsh70hXOkJUReOSO2xzlVONOjHyAdih
fPOVG+2EjdU9aeiSFW/sfnJ0TqaAKtEOHVqVZMlMtSJFgxe9qoJuGHCFsor/xlBZgSX4zBMX8t/7
Wp9Q9aeFSmF6Y31Vq4rn9zCzlR6koAE4s1cgRnsPPfauOZV+89bJHcbQ5ug2V/eYOCbjNmqqsMM7
pKSjSWtsQz4W/s02w0Vt5c054ihPTN0kBi9+9KumJngdH5vQ8EI5B3MGhRTKV4pjJWycy+nc2aSU
Uf8m/xJWYYZtTGwUiq2pe1ba6vK+t+EoW3tIiaTdChQVSxgdIKHxJDKjvWGS+sfXVgYNej3ErsOL
MxhdyhcUFt58QYlKvPlFJPsUwnBYtcsxG7DXTEiIzS+19nXAMh6ieUtmZNowTpWz8vCRPbhHFbE0
atp90xMn2X77Nye8Ar1fF61uQWF7HX4SqbzAFmeEcLjwBs8VuHK8sckJBEAjkH5CDMs52ctSSgRf
9EIT5RoXMtBERLlamCf07tuSzaYu4GZHpV6FldawPm7DcIZJEc01tpgsP5WV1j8Y787LCQXtKrxW
I5FbMx/zROvw8lvTduCvzn/lQvzv9VqjpSYTBhmEdfZFUxVwOoRPBAzYUlSclgD9O8+BMF79vvEw
WuE6XDjf0wGLYDOEG5l7r8bRUSEDlHPr/ZVrRAOXgzXMqlW9RVmlJPVBoe2TzN2LWnB8GRKEm9a3
pIjPexjAkCYdRNxSqh4XI02PJO2mTB3hPwLSMYvde91SmTMRmbbb/dVm1eAMpHvCh/ECzkb6Hpuf
5jkYBFc5DHGRRFL/bru2qhd+5rxymR6/fS2375z+nFtiom6HQk4ty+Lhy9ZWLoN+Lv42pA5C5S/V
jvKdqfAd/x7S1niJ1T921pXXz6e0BT5kS4VnMC4OClr+yrZuWI3cmjuxr18RttZe5jdnRa7WoWrn
C0L4pPCJQcd5WD8ND+eqFySXrcJBjXwTUWIKB0j6ZBiv7iRMs+nb+hvhiF8dl4tiupFAPqCQKnFK
exNG4a0xxhZjhkulY7yiBNITMRBKOQ5OuSM78P9mMZkHqkrTtpiNgiQc28iJNZoPHq2XmkRQbZbN
6SR3Jc/xRFcWrpfF+UHtUXJduBO/Z0mkKGfMxsq/x6IPI/ZYW8R1aIzxJUiodTEa5Q5IBhTR9z+8
Yp9c1mgM7ZIE8KI/J9WfBG+Z0j4czFiVuMjPB3N4GL4y2bv/TvPCYXxH5Q1oflW10aLxzx0zlhHn
apLgULxYS8vnIlaL51LuwpXqCI4xvGUa3LcdOyelwZ9Iyg2OW0BNMHAenYLej/msMjprCOm/ZGw6
N6WA7fxjtoB8J3Y0XnnPEmde3yR0vZ1+xZPIj2coc1p6GdcWArBLEegIm4ZKfsLaVQXs0sDohkcn
xeXbqll6KSBdpnoWrZawA/rKfnnwfqRglPBQLUiTic75kj3niU6bw5Tor0cmC+aCALFSqSEbp2KW
YdAxPVwbSOyoIk6LB6YAJfK53Ef79jmE6elRsMHhi1F3GZz0XtW7cHMoZ9aKLV2iO7VD3N0KFkhZ
V1HMF0l2BiJRR7w3RMaLwr9782Pef97Z3OY+0mQnn9frUzWbxoIIgYZB7ZefUfjb0mBBxzR5VCkG
v4NL+ufyeH7ReVm1CsXGa1W6r2Sc6fbbYt4WGqpdGGKKk7MVxCD9xlMvzU7GKpTOvpy/8XgTY6v4
Nw3lnBfSIEEjOgNxQhdQjUhYKRzgmMw1HmRRJzRpspVPYDmBm2jukCeTDE0ygaUg3aPP0NzYYRzC
rmwLvhj/ZSNLJT8cgZtcIRzhMzGK50FzHJNAVOvKLekQBc3oyUD7IEU84GIeyu50bhL3MuMSD3Wu
X0ExsDzqRGPX0lBSQYMj9O3yWZAWMzkQj4sj/qEUx7Sdb9jCHdfen+HyPgZw/HYW0Uh8gbSKwCDX
MNHUj//0wvA1vSeJHtmNjwZMwuuWKsCWrysRabhczKhTGt4zDq0fKooSAOWew5d4XYOLiwbTMCRT
AkIpD3Y4zENShwQHX5XPZ6S801rqx1DWrJNCM2BG5bD3vliEUKDdCdTUS3BzL1C28I1vkv6qGXTs
L7aZZqTdGtH/Ao1o/ySlyT7ZQ6/7mEfE+S6NJycv5fGpZe6r/5ofr5jpaPtSJ/u+0BDKA1je4ffw
35qaw+twaUhX9SFsoBntwpfbqTpsSQcI4u8ahBU45vFnpIvtKOR3f9B6jFBG2oe4TWk1qCwvXgAP
2Cr3VSV5jlO2G0HiISuwI6DxUQpVihWZj216+Wu1c6chhnxcOUy0c1iFnRtcXY2gGEsuvFVzAsbj
joVY6mJ9xKi+0/psEy40LZvMMyL7sKuJ3dshycbC5kubs6IuHHiOtPoLnoUjFGlCcxZQn0V0cw3u
6xSuShxnrmZspcMmmPJ01mfj5XjmNrqIZ4H9+vvaJtT3RLeWKApLysH1mb/lDmwGty+UWuf6x6FY
9OyTuzZkVwxCWUk8D7ArGq0NMjbjOHciLZnxcKew7TU7G29HD/1g8BnYLLtYaw/lmJ+OHUGm9Qhd
0HpA8HRaroAMDLXybCVb/KjQCrC8QVoZSEAs3RRs2YwrF6URcCM7iRkaD311+U9GYjuS7VV9whKF
3WubjCgPyd89HVFjoAnqVPgGhNludlfm+IwYeD9owrjs7xT7yD/iXXoQOxpFLT0un61Yz82GiNNc
VU3+mvr85F3w2qNEME0Qgq3y6EvwOEKhruEPeFJjUNTCVJpWVUk7Y+z9Z/MMczSJvTG91An5FeJ1
VVS+Navyu4Rd9c+4dcJ1+LaF1jKLGcQTpRMKvK2g0u4XjDSlUbVaUDkn4HYTU+zFUjL5nv59ryKR
znD6oTcaPAOlHrGlDReJdJEHjqVAzCAmo4SzKS10pjS+Kbr5HH+XUj6GB1sl9OsHpAXT9B2WYhHW
9hqKUDmHDKw9MBtWIpTrXzMIWIgonh9L6l7LpE2XwbfrFTT2o804jrVyH5UkgrFytlUCtOhqEawq
hh8ksFVlj6UJBqr2/RTMQ6E+osy4+h9uePiV+6/yrzfMPrRA9TmN2QF1FszP+mMZHwsgZZ05/PMv
LXuHmUMJjf15/Bec/lOpdiZDwI9CNFtGFAUaYp8WEyJNKy4yombiEbl1ei0FDgjK/+Du0rD+50cf
xTV34vUG5kKgwYRtjEuK7I/Ca+PBxf+A/w6Y6EBe0R8oadq9cLFdB1n/qgBEvJaKezzzuhEBgZ1N
hezKTGxO4+wkV1U144itNYmtFy2DBy+rBH3PgQs3qzrwFpfEGehE4RjbRS4U99Hx0znk/q28jyB+
HNGsZsmUaZu3Q/89v3E9nPUxXmhJ3B4LET6rtq4IMTD3zviu6crvVunqXnRQBS3qGA5nPuRxXaQR
h130YWX6gzvnU0WS8TnKSYUHiAnn+pksZQYsrryzqadukoXxqLf9AexQvYWM9RrNp35O8uVJ3FET
21XeXmxh8sOpjPu6TjvxEkqyRMHrSjzyJGlJr/1ueREP+yy8lm4X8AiUFy7MVc9HHNTjSDUA+Eu0
jnouhjX14TABDfPFXE8Wh3wuP6ikCJCckieahgQKx0LxpzM3yejHMafcUdeH725uyMw0mZLzDmzR
pKHrpYTgFaeMsPiA6sMJ2byaO6SahrUPXUIkrdGGTj6A2U+SiljOf6r/X+OvhPgFfBc0fux8vCoq
Hj55JO+XQqRnOXfjZAX35aPGXil/KATjRMLVoVCk/MyursYRC2+5eW8r57MZSbIKbtLbtIZvLCGP
INPIsv199WH1zgkhBDtZ4SOD787d7U9lgEe5xdcDGs1lJZEXt2zdyAAhljExJkwUY4gIxQlUyb2v
ryx22qdzIUQMPkDnh9f8Sj9XCMcx1R3L5tv7rha2GMTXbSrHi3GTyTVvXEvX4H2dchBE2O9DIe69
vQVoXo2GTpcMNPDRJB6OeusznKeN+hFLiPVt5pSAM/cg+O/YHYrSoi3mN+o9IG7FHrsTZxROUokX
4IGULvq7MEuxdLLubKdD5Tjw3np7g1PmTC6ViFrNmhN3I65Wtq5+O4jozNEOU3GIGoMfECS3MD8T
Txede/Bk64J+wYD/CFrD+5/PTBHC5fhWI/MwK7vYaONloUE1b4b839Cm7drWb3CdvuEQ8AuxRr6N
xWvuFc2/FqloZ13trhyTilWsllkYI15sh0a0tIXpCZ3oVJhY08w2loa4WB8qaoHAO7y2s5dFgkzj
ms9hq6QdK+3unO9E2VyN4dhApWtUF4XNuQ97HVV/tC1nyHBVSZJL+7vIlz16nXwWmzdSRkAnjz0l
RRmxmVE2wGoSxN04OVccmYwRI2cyitw53Nac4KuHEopM/yxqUUlYu652zbAv4qRrfeLndcIe4448
JISUp46HpoX6inxKTf8QbuDicNrF99TVKOxr1K7O63xB8c4xv3ASoFjd8X51rqUUXvfJx6Wtzall
mQm+q2OZHuDdmnaqhRdH/R9FkrTnhycRvrggc8ldBCYKVflVOlrXgLZCXLyyJnK/fZWVuDlx/Gkj
3qTXZ2crsA77EJWGME8kJkmVe3MCwF+BqnjEDturaz0ceaOnMWeZR5CPyUrrkmIjl371BBlW76Rh
gPwCJX2Yl2gACHEEyECqucftSRyPmSeHkjbHpa8vZtdZA1esWlFGTuFe1k+7DPr/9+CTFE3GYZf+
DsKKK2OgTTO5o/QeOSIwT9BnNpKGn/asJeFp2l+Ms6ZRc3JBZfDDizWCeIMc/NOmBbwKCiLHvDW2
GcGIgLAuE0LfOd1JXKtMfrmlPGkMKg3DLcrcpDjqHCJo4WNRnGckcpEJi5BqBk/yvLFXgwuO2VV1
+ucpKDv/Su+g2ernCJXtreJ7vas3Kni8yRVAYFzU6x1HHoYgKl0wRFyMi1sT132bIeAbsqBZOjev
ApSKC56CCyEdKFqjhjZvyQood9nqgVHiacoP7egvaPxCzp+4+4hIKC3hONj5XjgHg+vUj8RQQnsB
BdPhxcePasHUldbIIFS2qhNA6uoOo1l7NSsnyC48NhNj81Pw66l0taxhl7PORqXNWIkfLp5tKBUE
Xh0RWC3IcJg34EqWFhw9c+CGyziSyp62HxKTX0Ibu0RNTbHsg2UDFwVjqq7Tje5jZN3L9Rh9ZzWh
A2HYuGCkcd5xogcOCMM1HgQQd+PMuQCBVm+OFupZACf8hj1eoQvjQT1K1rMQAmWp+z1h6VHJ+DNu
MO3IxGy/p3elrt5gxMod0c7W7npBcoUs6/jEhBciN/E5l3a5yaWFHVFzZdJqHX+OYyPJ7o4iCvZB
Uild4MWNmBW82O5EHBQrjsrel468AMtvveey84nPu/G7c1Q8oD9xW/0t7NeaXbw6F2RtL6xxwhM8
EH6bOpvzb2Utmy60iMua39GJt1KKPwgMdDTkBA+apyT3H0QTzU1QW2fE8Zx0XQzkkqgoFMzdqcIG
vV2BFOhx8CT0QkVNv2TU8h9kgUP9petF52y4onEEvODwUuTTL0LYTgPTWGTEYdVwx6aBQcNcGVfx
/J+HQjFAy9j4Hdnn1f+Tq+or8TND0lhVJW4pKgwmKeeJf/gZ8xW8GZUwqD4f8y2qgDZNLevZBSUM
lMkZYQvidMe/t9ZMn/ndueLnOXoMFNX2pFAP8kfw5BDw7PN7OkGDCYvSP/FfB0aFe9Nh7KV0fXv5
M5bGkrq4fCzgCoR5V5hAEDyffc3vt70dY7GowhdHkMNPh2DFa9ZEjX7bAJkMavpmeebwT5DfK1Yk
dXACj9Son3qsfbUdU1UAjijWYxcQlokwUoeTTFbMPB4OzAo0XXAobVw1KbKeeSOc7FjssirYVNEs
q1IzYdBszUrKOAG8aciI4K9pMsJBazWLMe1UwGjhKiPCxlYc218CYnK57a7Reo28KHMpSwJug1av
LxgX1w3Rb/flNEwCruZpij8GI4GrwGjs7Dgj6bTXin6mMWffqFbaHpPm1zt0vrrXRysXH6fuNdH7
jv+hpWo7wd+VbPPSsxzK7SqqvsKqk+ulsjtqEmqCSI8Ua8lWRSta1vQC5VSZh+kwP4Rtobhvz0P0
0OTsDoObA3XNjgjQ9AOtyyhKOeXqO+n0+Eu4szswORTTbLXckAvw7gaOi9ZZfe+86DBbfqL59HqA
VgtylbH9UHTy2JSLlfA5eJMcSDYFJNgGPWmC/kgq7bcduLQpBPi9fvsXxG+nS4mgsfGwu/wPn+kW
B4ghrMSNXZksqGLrVuBwxY6IZx8w0ZhNN3cIvajmts5PKFoQZ++L/VfXfRnFrPIsazjAmHEtsaxd
ghWXUQkn2uvN94IrQuYdHoHe9ywc/JvdAZu4kT2JYL52lS7gD8UHXkcVTCPsCVfRe8gkurP1fMih
dvhIZ62+3bBsKSqeLZO0fhc7NqFWl7IVUrcTKxx4TJI5C8YlRs7CGv+xU/gU6oQKgZt/tpX+O7/z
n+79R6Z+cegRsbo1orzm2lz0PDYaEtXJd88qES+9QRqIjTpCxYWwKrXeqyB8QgHnvkUtP8r8XG1Q
gjT0OT3P5w8xJ0icz1MV8aRjJXkNjp3qhqPlnUWoDrR/XYQctsQUfB6gadptMQOTLkoa/87qoCoE
5PPIpbFoGuSWxC/CWZky6k3zm41ITUIMDKqOyYe9A7CnJlU41+ozUxquLALzzItkRsNXYeEhvSfa
EqK8eAEsG6s8j9m07Ja7ujvrX5lKk5WMDjtO5fBcdx7w9k9mIt6jjx0Hd73LaXva8isWE6uhoBkO
TFXZXREAgYwUzirT40qRBdwfaRDejlBn0jVrliSrkryhvOqh26RjIz8XGt3zZJPIO0OZ+htIioAd
RZjaMHE+ERu3Bm6K06xgohNC/YZWoCmmvHHQff33Dv1uImXBiPyjhZrxPF6SqLtvEwOXu7lNCgwE
NM8xxUBB+h7rz8kyczhZuJfiZAK2CcXW/EoIrexrgdVh6FgXShoh/KT9dYqnic+2+ohLTl35LyS9
vO76JGma/nxhlN8NkTptrpqXojCR/KbIzETVTwQ3eM6p8wBytpB70LkbDICd2eIX1O+ksAotOYg5
cgKS0AvSCDEYF7yzJ4y1lDrEPR91uqh6brKdU+yGEAPKa6MtJPRPKT9VSTkB/6uPpZIyT+M5wZvJ
lfr+hEc9ow5MvvEPFB6sSDFDGXUnFdMoy926Nbhbzrq1BT1pQ9E/o725xHW8jP4QK1ykxJbViDNa
EU+ZJJHYswPODf+oswh/LTcLBK6zfqHNyJ+naMk7X5IZB/40+HyZYurT1ia7eyLVj9+OYUfXOrAx
Gzdm7Ec3dZpuwdWLwrQDbG7azJDbLcfN/m/SMkp/3417d8Wva/7plGiOIWEORVvdA8ENrdCIOAYU
82aN37u0YELHAqcCNxiwM7lvB/Q5oZewkkamuovH8Prsi/sqpitl7KjI8kdtwowxBltGSEaDn6O6
GAbdna+z4ZWvQdcFf4odDoganqsTNWjl6rrc8ugT7A0oMBRE+Z26sj0jRHzwpEM3/Wae3Vcid4q/
WjLK5xtA55vbEuCTXK1/32ZeE+pzu8g+z4YgUrl4KnM+XMYmo+6UAa2VwOtv72JkDWLsw6tar7q+
cKjAesDc0OczQxNf4UAlvaZ9bZtVPi9iDwjiJ6cDAuGj126aZpDOTzm9qXJFlR6aJuXmHwFujk5M
oN2P7YBHL0Zo8gxrvhjXNU837ORIL6IbRfFn3LTBLF9yaiZa1JmnDbkUQL9iSqbxrEzD0SB7NzAd
07GvUj4PFm3XmZd5VIvJglQDZQ8QeDG8iS0CsCNXaiEVJhr9N/4CGZ3hg/uHkuQrnCFsRMh7uGll
VLrAzLzsyNGoqbVNnJCn+zZu9N5z4s8rjQjDBG5HCgV6QeXcj4QLwAehigzc+5Yc3tuiEnHYexPs
83m7eLWJPGtvI4bHdA/q96dqUqFy3Ou3aXXzxp3sssIqPVDKe2hIZO5bn9cfLCymzQ+bE6ucMIo2
/EIT9ITiZlQR/wpxLDFOuKP0P+T5PWxCKNnaGlHgGmNGF1wNo85ieLYg1gDU/j/n53Yosaca5v4z
4sfke8Gen8UjPcFf5mjWQciOVc/oOHh4S3vc/K+KO3xLBIInX2ZvvQGvKpHdWaTS540uXdild4hI
VPxKY4jZ4IlCWJyRE7mMK566dT2FJj+LhsB/TNC+fudmWOGUEqGCqtR2e7HUK8u73UXHeIFxTWxL
PPSpd2C/u7HM6c6AcTkpvnVXT+HCLUmAJM4sqJdUulqLnQsxyrsoP1USGX7nDS3laZvaILKZgDw1
a2IlNlRupCJgnm+R8dTQbnRD6NPoC/iq5RMoOgusnBapONrJv24W30wqhkRfyA6H13mAO7eSL/Gq
e2kEfZUP0L6y3WAMAn5BsANhAjqdywPDt7eVyEUSjtfWMGx9j2v+bTstduZGeCdHWn+AhZgTztFU
EMG858Ze6zjso8BV4KIhIKf+LCJPdliGvOAEK+5BZitsjy5HPUwhBPPCXMLmg7zPcO3ktzYMZTLE
miihkOX1kgS4Q+wmpPQWCk8tR3ycAkgsDE2rWbviMqQ/CKxD+QkVhsaH2LNjowvXUVsfXjQYzYmF
iqSeIXCUNY7gjzMtqrOJOzu7Q8KJ00P5Vosx1Dwt9N9ajuZEyCE5COax8Xishz8sLH1vYfSrSnfc
4OPU8CntQqb2pWIWrUeBu/f4s7QKeNK3w+vmXvPz2ANmmbhkXoq/fPGofNgd8Bu6lxYKigcxjIek
qvWzXoVHzve7cbPd86/JvYd3T3bPZQxz1FPKNqMEOJkR8DUN/aIrnOHqSF2c7ziEWDAel+MvOA+Y
jfOvAwgFrYtRO6Sx123y0d452AVipCDiimqK+Mns7/LJfRa43I9gkNpKMc0duvw086BqWyJzJOpE
IR1W09JztLhUAI690DdigZ5f9MS+NUKNz4BbSPaqIhQdypQBtt5ZciC3kceB4zfsH1SkL/L+q9Dz
FsGehz3XgLWEOGguWH9FQPpya3KkV6onko1EjaM3xrdbYuVBb2KKG/JjC44HHNWdulvPu5fq7pwc
6f7HEJm0Uor2U838/hoN+AcRlUS72Z3QDEJhCXxm6lhrUlETKRRX7/pT82lWauo5jv4yWABzQ6nW
uZjJcoiECYccqVPqLXBV78dOQE5Hw9y9NKaTrcG3ht45JbsZdfPx8Qm5dkcaG8gNZ911XqlQZBTg
fhhXWvELvW4MTrvcCIHDlxK1xPiSLponJ7bxwnGupxt10MGAwtLWek7/6abZkXnB7Ot4xpNZMv4b
H0Sm7+5MHPyG/dbNw+KHugR0D25igbzWBr9N0Nqln/DksJX/ZyflqTlHqwST+gNBo39yTfDFRfQz
VmpqCqbtQG/qUXplg9u1BJiedkpp3cIeTMviQzONppEBgYt+OXN9rKvLZ1gGALaQlNVeT6GThcAa
07bCCrpM+VF5xO4XJw2FZkKb389Op72t/TxXYu0RToU9jkK+vVy4rcR33U9k6XOO39aEjdAk9ew+
IYEFMNj5FJ5Q4oBwb/Qr47OiEUDOVuX51rTzN5Xj5yz7D6oPSAfA6Q57YsrEFrUw3YtQUB4bfa3k
RZzTBiM7bfkUG0Z8kD1MOFKQVsOw2Uew0MI1x/OzG0XmnmCPfHQBQcOUMmnAA/WvGqbZb+hETPWy
o5HtlLUjro9OjKcWjI5HHS2MRK+bjIlqGO8T/THrioxXjBZAEAE+s9VSkjuUdHhz/V8/D4s5uL0Z
kurPoMvFcm3GTr8kgeXKSeQaJYCiFpPWJPe/oCrpnXp5FkOItt7GPambfpTn1/mQhQkVtelujVDu
HahW59cHr5vB2UAmLij5bvnw8OZopOQh594S16DZ7mVSPmv5Cevs347U+9Im9PSxrfYezTR5Muhp
eRqzS/pZmNTxItGdIAS0f/e62FktN2iBDt3vLWWkyBppfZqq00SVp7RwdKMs3cHVKSAQOlDD5L54
seDjShlTXzsJ6qVZwQ+XQE5eKN9VOYsErlow3g008iOMmg8B5MNlM9nDYfgGol5HCA9zizBMYetU
tJ0/0PsVXc5O8AqrygddyXlzGfeCpmIiq3GPB4deV40SVTqqWNL7qyhaw/hM+ILIrRQIaazrVgmh
I/VHbGFmSrVsV456u/O6k1v6qo9YHyjKLD22qfUNQF1aInxrLlmmX3hgXChm3cajK9rUjzwYuK27
k3J86eQJA4sJI7ONJrMX+UhUNidGrZGGw++qGid1Wmscc9gcz7RnUuXF1bUPHgK1CWlbTX0MIZNA
/L3/dIZ/Uq1n7NOePjEMLSAk2Yy/bIQfQ0caezM0sWov6VSHZGFdGoCyLg4J4GNYIlNRPXfWTGJ+
xpPnnc5xmOtKO4jYVvCPnqWDru/zeeVoJh+H0eDSCf4ZQHbanNAVyDdjzF5YDB6PJo0sdVNkB85o
fgDrGAmGGg1YFoqOShuB7Q0Goc/MLbFCcnUu+yyO3f9HEuC8r2IlnBFo6j2tzpzXYkJvxX6w1rwU
BqMsYRzE+SjzhnYoVUQLXS7otaSsc3hjOMwuVevstVF78/CnHATTCMd29+3VSzpw8+w/1NL+PyG1
aaDrWcIE2cI0qBAG6FcK9zzubmYoJ4PvhUxdVcUmL+ASi14x0U86m7903n7c+UG+lEbrxvdxT3lh
A5YBh6Zy3t1oYlnH1VmkYE8Tn9ImBzHVki3mowyzQ1E3meKeSvxf68Lgi8Sor7xedouTQONY38MW
udRt7CO3/Xt8wao0H1LcyiL/2arwgfD36wgsyiwm/PE9MS7RQM4IcGfjV+VarXM2ubEz9rWyitr6
tVACRZ0TRclT2Yi0Qfzua+38oRSl154jFE9hrKvo8bHC173mw7XE/+rrptFRIDZUGFx5upNCTeW4
6pTuLgg0ibOiE0z9S5RbnMf1oS9iOVakwKR7PNLQZnQ8qhBx52YymWgoZJkbr6DwpoFHAkRitgiU
WywNGUgRiM4r86Hy6cAEHW3TrmkICVWsYLDQzZ8S2+dcURhjNFCAJYT4cqcZxmxWg6X3qYdLKeyJ
7ZiH3j/pK/QSpPH9P7/Kxym+sXYqTL8bRvdGoxUrsmbYYcL9KiB544bAqysM0eQmP+6AuYBxH24v
mDCNx2pUFqrooQULmdwIenZ0L1OsR8NZolGpbxvzCZFRtDHIYrD3VJaF5CJeOdPzgFh58B6b1wxF
rUUPcYd0nMOngnP4dtMdY3bditaL3/fuYE+cx/S2Gtod9WaNHXDFkaoEdZ5BeKTwzRZz4btMu42c
s2s7bhsX0zAJBW46ARZZF5q7ehvHJqFwRvcUfrcNGcui2sRDDmHK7Gq/PvCGrHe4335O1Kw0LWQK
3KrM2ayo1mfaplKIJ5gAok24w/2k1gX94Kwa+/Y5gluBaISi+FH6FxTRC8VRgfddelIz1ypf3dVL
DpYQx52XKZCrJfWrZtcZ1FWehuNcFU+5cv4ULqJdV97/M5rLh/OKYXQDNwWdtJU1I7wgtdJAiGhh
ukUy/2AqJQ/vuOeFArtQPvtoit+PtVQQnZnrU4tMyVYF2i8gc9LY8Dvxsw1cTuWsuVd4IVhoo5/d
Z3QGCdf7PdIiMOKZCNDAc8BZp3vS1MzLsJNINzfncvj2AFHPLc0xG14FkEsZ6pDRvpP8nuwVVfOc
kQcThNLOMaZkH0zGh+THbSzyultZKZvVkQzGqJLfrhAxToFmOo5x895VwRj0JCZEGNyYNciz15KG
HyM5EMRrZJXKrUVIWCvhT4e1v0fMWLSZLwr3odv3poDJZoHW5P83Eh4jsgWYgU0pFfF4i6F0BASx
484OGp/HUaDYkhezagJ23xZYztRyWkRqu90QanM1x3fXLEQucdqnE6vKTChQ7PSQaTD9DxMor6Te
pRn5zOWJsDc3FZIZsbxexaXfMirJ1dmrVkBwuW50K5vQBRot8MUB+h4aCi5VqpHpUAqTh9jW1yev
3QQ1NzN1I8ggaT73F6MTm1vs2ukMpubj5Cx2cSfgm90bV2T657g4J1oWg/h277EICeW4fxk0rKp6
iH1e8h1I72yO+I8Hv+/D+dKuq5c7h4kvJBMK7GJ7sdINuSdtT/otc+zgzbxMEOWwmufK5n0Afyfn
b8FvFvIPyndtsAG/NtdrVjF1UMTKaMZp/BA1roXiCh2JnBYyGQWZPty213VgXdBSxIxdte9vjP3R
B38rBkGOyT/b182JlReoGS2HY/diyJk++h/4F2YEbdYfWrZJGWUus4CthVzC84wn/83LnbI6xMZu
S0/8hOzNSikutm/CZtDJzAHnxNDWhnUdGpvWFrxZv3CscLG1kvQy+zuZVvy97GRCjKzeoAG2yTvx
C0BkXY3VSiObzmlQEDfpBVuDPVzdq0SKmzy4vCJejZy5BMdf1Bu5nvtCDiucdh95C/aOgFxQ/iek
Jp116wCiZryMRH7elQ2UP8CCVGro9JaFxTlIxg6ww4jBm8NTkM8dxOm6K7wtxiOne139T2EQQBbV
xGM0gB98vo/Jk5dS4H3+6i3KcXN5518vaIb11m0vBoop2WYlsX4hYYEpAXkiUbI3FLnhh0NVU8RD
fFELRNQ7kYY7D6uy9T8OUkX9EnJQHCLNomHNJAJyjzqvYTFtxujB7DUOBESf4soTKE55R5uQQXAK
y9/YVHnpzI5uEa7Mg+yvj3YbUzbzYuZ64tnPbCzo09Gs6FD96wRYEwEz3/t3UguTaqpmg+o5+48Q
JlbrPacdsSyGftd6c4gxpg+4j5hyEUWiQ2jJd/ItWG3lxD9DR9gdnFO4UfENYn1U4aoINmBSM2xX
/TsVPuBFCGCAXyhafz75dcJDmTDbT4kdZBbAeRu2MY9dMMdC2iMTo+v+tEZyBdCu0iozCc7tvIJX
/gJvRKUxkOGGGNEh8Z8Fv+aJEvFfA4KLUkTXOdyTAIvjWEnBotkr9ccqLrJ7TG3DQ+Swza5ad4Ux
XS6Jc76EUoMO7gdFoSdJwPz4i1o2a/8kyIzJxkrbwOOO2zA0yjpR/RcRtbXvl73dPdT+SZxnzkq5
KxDY++QLbuBojo2CBSCVj3BVzhkFiFQn2ZwsbUbFJqPJVSS/9eU8MO6TgcQRNt5n0wF70/mKuCQz
cqSJS83TybQhK4AnrC48J4ldlif1CBLLDfWuAL6taFH5+5odk7gAPhZI/ab+yKdsi5A3Ho3ORNoA
oH3w9xkjJ1uhkvxePOYmAalQPecT7T/1oP0fkTJdBGpmvxnkK3/KXPzuwzmQAOynppcAvrBoHySu
wkbDeEf2hC6wDrXSyFaxl+l5QPXXedzxNEJBQW47GJygo1W2vIqwFBmXP7HsxVxolHqF+SjMx4Ep
F7Os4Wos8mLLQYPsJdH4LYXLwOTgHVZnZqIw/rWhuFVvvxe1bFzZZ1B8tmTvx/0WpA1SSBtk8q4a
xK4WI3PqZY9BeyF/h/sdxcfSExFn92vGQI+Tk4zks+C1IyR3sENcTJsdNGvwwVBxargEQb8d4rcO
iX4LIt3YA/ub/iXz7NQI5sy32MglHvhWwAvkEF1jhPJoMzdo6O9nEOosHeElPHfBMNBjDkqSO86n
6lKgLqPdt9wjA+5zjCgzo18J5blzL6bNir8vjo6zfcgFibCrchf8uZTl7aDkjiBs0MXymlLadgT/
UFfCgPSQ0r51pja9GeMkd5zL7D5xFCV4hqvIml8GkiKMI1gyWq+wD6QRsp7AyMBCdT7fzx3xXwAv
LiPDPmX/AoM3wbs5FZsPuQI0XeipK6rGE/migK4jdjxLOOZSi6qkGp00frlmMgrQxZkyD3X3BMhe
FWc6Wuy08Oywx/ltWVVcl6H5TXPE8lN61cn/FFVltYVzFfH12IZlzorcMSkGfK7MsMjrJiDscRC5
Q6QsHZDNISmr55ieCsnZ99hFEigIOewgM6DWBMCpDkDw+uCKDD7SCaH4D+RgDTdgf78En6uufyK7
eR7qqaZnd+5+IbEYN+Mdms0oOtwfa0pajgO/S/cjRtMr/GfMPPlPnZBYFUVnuHLiVOWj4XM2Etml
bFY/OwisrFJO82Qh0sFP01jff+KQYg/y8XpZHL4Lq57QsVRLSlztfkGPrtfujrw3Io24ve0avbdX
WgvNuvpkP8+/8JdaPL/8xtaQmbaNK3X60IgzjFQFlV+EsNPCMzm0PSLI8pnfVvJLmGOE5O1cqDo1
HEDbL3ctH4F8KVH+Y+f+0ho5rAmDIaptOYWc5m+HCa152xVioIYvXPg1+MMfmDOK322e9dvKK8u2
Rwq5JltMETrCfjuljE68nPrB/8TM5O1wHCYiwkEkDhsmdnZam80n3WtgyfUGpuGCvfRDXHQ5Z1HL
sPUx6Q5IBN3+nrsMIvNxpN8NLOByhMbTbB5k6aWPy5WYCi8McTFKLxCOiusbgmMycSeUcmi452gV
2eAzWmYz0skpaQAgNV38a314KuhntCZB7JM37PvTu9vdImu3E0tjxaLtrmwNyRJg1BLUN1tGvTPS
A3yPKeOlspAxGFLWxkxzQcFejMpLVtvRznaBr0vAZf1Zbc0MZ7JnBQmwYr5H4UhGlsAmyoO+g1RZ
888M2maTlejg4OaBIbrGhaXcO2J6QuQ5ceNCUyXXsfvl2xs8UXAwReY7zzrH5n7Dy/4vsfaKL9cU
qSbAbZYmk9pQwicmmUosyBmMNooud+5g7ixaDWFjl3odk+wobXdjwSwGA1K+A9I9JnIEgymsHxjc
yE+Jr+kVALa1pDuqMoLgenOD6te2OkvO7nk737MWDlu/TaKsGGBByM40try4dyhXZ1KYj9cHbl50
RqxrqKljvIbf+K3CeYGWwUCh0HfCAiwa/MzImg6zsgqUfZ6EuCyQ9fbm//iA5DnCX1GIRygHNZdQ
hIKxi6hfLgIPRMpX6jpTC4HLB+lNLJ5ZA2dHJSmY8m25KuesVFjKzMkunGAfQrFJYijKJeL9lIB6
Qg86njXlVT9XyGIIbSI8fwG8L5u/HEQfdM09Fecd3mTB+XYYIOwYAV0pQokmejz0j1J6oLw2QjbZ
/I3Q3OnxHlGKRe85qHfW2/SjhFbduObn04uJFAJ1iRmhK0+ZLGxT3E8tQ7BnQIrtQ9Z2WcMEyjt0
qQcrAe+uVFntLAn6RhexzzlH9FkOyS5n5WNczA6qgEY488HXkZ2t1RavIMIIhMwEHu7w0Rp5/BtD
r3eXE9HUGPls4G0PMU0KNW7xtrc7VAZgskImkqVn2zyAuPYjO1u17vtzV6DuHtDq8YsSn6Y6p9f2
WiQxXIpfNqwAwIQTvjyQCReCqy0BIxCmbzGtv9xgCZhK3cV1hWIuUO+GuChAmdah0JphgqTv2ylC
SFKFOyXExuD++V8ioKpNQl6/ZxHUtAfE7r0dCFPG893od0so9xEOta1Fn7WbZUA/He7EUTrvPUNi
HsXy0eA7xXOws9WCI6ajwIBhAhPY8ENeBd1fccovbMbMehbEkoq4p3A/mXcvZzkIwWPuH9le8SAu
PkT7im0J6zafIkiyL7vLQX1Cp3pdoLNYbk6c2nevscpe7D1VX/AN5rdtMOiu0pbJQeDXJsmqLcms
hW9A3IXImEybBmuefeECUe/66tF/3FedXQBDzi4qaCrf/Cs3JA5SCrMmzSllYsJKkjx7/z9YxRdQ
KUf/rE1tGB+LtvxMOPGsLZwOogvqjAGjN61LR2tRVAygNJg+M+0AUmRcWB8DAiBykurOGQcyJWCI
3Opm9wAzusZzxa8jC9NXoy4HdXL5vkFnJyWeCDSk97tDV5EtYHGV7xCYRYdyVPaw6jc5Q/J7+kzn
i87G+UNpt6Q9Dx+twITieMo/4jElEKel6pKlB+UzY9eyZOPMW/Y0uqs79DdPCpRvL1I/zELcXRUL
nEZRurL7PrC89SXVYWzSDXmOgCS71AJ4EVPNSqxS3xOv+8tixmT80I81izrdncF9w5JjoeLXPv1j
780+4UUMYFcT8P85CfkJb50SMCETX2BFnPLn8muz8qqsl5lIO2lAhGk1QLgNKyZkU0aove9+S7e6
9rJYZmoRLcfTrAAbo/D9skI6GiI6VHtezpFtu+P2xAdnGwT1lreMjWu4xB+H6y87xuxlVO4BqKZ6
lfckNt39pRh/6Xwt2MrpzyzZzkAiv2dT6MpIMFG30kuOxfOeICGPruImVvPgj/XAnSSzG40aAgNs
KyFxblNrkPIoJCUmW+JGbB2YmSwafy1K9JjFOu4fPhHUWBW1ZDkLf6Y+/xvMOPLpCXHOK+XV0Qba
07Xu8TYXTnrHlMxl9xJgJYrM1nq/btwoJebysSKh5xCBe2GlEumvs8hge3TE9uBvuf62qLBAg6KV
eBeYAtz15rGadFYHKwFV5zALyGv+NH0NZxhNoNsb8LJtcGjs0ZwqNojIRgvwaH4+OZDZzwRvqjzW
o1x8ULQx35BeJeD2/2qClYK0wj0UBJgEWCpowmhGT3vVBFej7nPfyHMZ2nx3TMrPcf2iO/+wVfdT
pqSFwHFwKNfZHAk/dgum7wzrfQJyAlndLbmkPb+GaKA8Lapw65L4YOjAJDAmjB3XNCpqqTSp0jyM
UU8BKL/iOS9NHvVnvCDsmUD5HAmeThupVzo+x6fStCXBql76AIuaOFt9raRwwPAPKNXNK5ZJarXn
ZJo5mrWOBaogLmI4g0ZM5hBHfZb9IL8yd/JdG4XeKxOL7zUAd+elTaEvbP9P0xe7sqZI6Kq8BiJb
iJLqroKexTSCV88jy+kCOjeLqMrBCxnn35eh40tgBg1Wny3PY9Uuvkwhrd6B8drrkAi1agq+mqBy
bwmoOk1yZmSW5eiETUfXf9UFtmGIax3IhK/kWFF954rFPNhSM9YfbYfdsMrQQxJ9QROxWp3GzdkE
m0iQhEhqlSq4Y6T0bO01PLSToAauQXWhf1V96QX0mcRTTh7+ClIRgo2Qoe0W+d89Ts7Xf0DH/uvs
UbCiG+ZMr+PIQc7kcd5ypS5IXejIaW/GE46TzGbq7cKToF+hREUh3HhK9SdFzhDMIGKD0vffzzCb
EHRA3sHXfBWlIBZyaA3Iayr8FEkGvKLSrqBXauLAiI/8V0mq6xrhy7kvNEiYju8q956rOboyVT9M
evGff/In0wxBSuKwMHpA2DKg/oQIAKsn0DkhsBNaXpNHm6I/Qn9mVogFXZhnjCJL+6bxQJYkVKZP
3sy0QL61mLlKJQzb5bTL3WlDhZk3PH56+AnxyBmaQsJPWERCbn8N/SkHlk5C87FgkPaSCnWpQEsi
r0kfBK0/FmOjPOkXa8kKpeRDEhO9XKnct2vFJS+lhWcHYEfVP8lWCtOQ5Bddub82tz8/rdylKF+0
5AZ9Ph6t1S2GT4ljwunbfoQLDaaCI2kwIHRFTCRXZdgV9UFhrO4hm15WjHheA/x/0jpxPL0NKZco
Zaq/VnzCsAEw1b/quXR+33F+jYgxQ9+AJjTd28OxH1VvIQgI8ipmNWMxhgRQcjkhBbBrYAUQYii9
FU/GWMlzufjIM2ZOzAcdOXALXq0c+ATN34+LYr9w2YI7A0B83xjDGpakrifWelabTT4DAtX4oLs5
nYWguLkHj02VUxsagWt0N8l41XPZ9ZYOkTFDwib9amGMItsFPg4q7VpjUKlvNFjcUbZkFZqzWoDV
HUId8S419lGG4ITpWPAXDSPxV1nlFRFKoCETQXXz+zqMDt8DCFfRkzEpituaBIHx6JVnj6RxVzbW
VcGVPnaGHxhQUUV0TNgpHnVDBo9k5v5XxfL0hEyBTZQa1i8yrgor1GDiR4lhStQ9O3l6uP+To7pc
IgxTpQbK+kPvI8I0CGYIFx36yuNBFXZGXEm9yZ+x4ouHK41Rm7eo9ACcO2J+YTcaCTMsFT8A9NYb
IqyqiateyPlhOc+gDmSVjz0tLk7i1e2OBIx3Y7vrSM9rtwmCtQvlOeI+NV7ZFMMfUdC3Hnn0TxIf
adAVtEbvoA+l0q7cBxkUvZmwHagF1A+EyyptZxTpprzXeh1UwtSMSozUy6gYewQyDQf9QaMan/k2
BW8r9ciNeaqiDViUbtqnqA+dv4MoPbgIVAA6VSxuSUaAx9Y+pEfoQazZYkDcUir/pf9VQrxoqzKG
o76adqZGCrFrDatISon5yWe5sj1abKKrDd6a19l0wV+fXPrO32Mpv8pwW74LDvKg4sORDPiFB46x
31z8+IURCvEvg8q4xya3LtS4mRs93++sWHmPFhcFjoZmeVy4R52wRuPG5Tk7iXWxI8f8D5TBBszM
rEZlQ8SifXNiK1F2vubI/jSGHQwNkPDoH9rm2Ajq3CRdSr5w7G6/rsKioNQkzAnOEr+XcsKPRxaQ
sJ5KbP15lz2n/B7GiN5sywran0zsd+TeYl35dOd1uPSn3K/r/ZJVUx6A3VzLxFWce8Kab/JFGu6E
C7DdzN737Nah7Se5Hr6DY3H/5BLeew3a1DckbPUNoxzbyuW7Xjm7q+8EeQ6VdOOvLBEjEtiJsG6i
qmvJBDV+k5sOjZmRgMyzPkM86tJ8278lRZqRVVIoNarQ5NXtj5JZ8Suou4sHffdv4wLSrHz0eFL7
Q2tJQ8tQh2ylIXTQrqwL4SbPtWTpEEQ6NvnI9DXDVpi8weM7zvNu1CgSv8tcqPr++VSO04n5fzcq
Vq/9r4DghPwZ4Gsw6Q58bia4CPJ/wsf+2qpfcM0IT2CS+eHMMdiDAWyLg+BWPOC+3rBCQ8NNP4fT
psDmhouCz1l99OKDpHaOn8d87ScW8KAy4xWnPkGrXnfFCVKcAMfeAvklIe7J0btG/k3Yn9/DPvsS
RpTp2XKik4eDhgl7PrJxQ40UgK+T2TZHT+OYQF+7d5/AeNYfycZ3OHwpOGpIRgvW3N7HkJTq8oa3
pfu1G94/nw4JUytHO7x2d9V61sxQsO5MByz1ZigEOBD7WFdxrF5K6Ng7XhQ7Icq7qhpk/3lciABf
qgU/0dui2u+cHPtlGjWudpC7VnJ56iHIkrupCQWTlYqKbIwyD6uoXf7qD25HOEoAfLsUfQ0KNHGt
Nv+YnxjgNWuk2+2z281zGHQOfW7Lf2F+TmAaf5vsBhW+O1Mtk7zjRG3/QeMwsgny5jvgEz/ShEm0
n1wOoJlZGE6sVjSusaLUfFGiDeEmM/nwKCwFs79NaqS4Z9gM8Js15EVq1yBW3lclJPCwZkz8wE4Q
AwCRAlkXB3Xxe/ozWuEce4faxt81cz1UNmHafKtbSs1VxaDn5ZbTCSFTS2g6jgecAL0bupZKkMnh
Nx0ZmWdFkLEQJuTG1UdAcv2Y0PpYo5FuCHPOu5p+XgWz7pPk5Bboff56UmGCJJajQ33NEZFDwxFo
EyPf5wxcFClqLiuRH44g9z6nKGiwz5hMsGamY6xefJ0BuMiDuQQENDORPaS0HiFdys4gJhkTi/FW
FkvUbwWbumX5DvvUVYN1MyaNmObshGMY1vNP4QtUPp2/NMjS7txdgpWLMUukGJTtqTpP9w2ApHbl
QMM14+ssgTGWAtiDhx4t1vYG55neeF4ClGTbE3lUP/Eq7KOEJxzrkDAUPEV+3ThUdiPGVoKGhGq7
vjcBcOwocYLp+bOrzbOm1MkSDk5dbb2rgt4sHV+mjNs7sixX9Wss2lb5T9kwNZUEHU+IUHSFwb9y
wjsl2PhOhE6l5N3kf5jYofJRMyyX5Aisybz1yAVwPWgrzWpKVpEq2iEyVNqzF1sYwJkGWdUCERe2
bXT1AVg/LuGIo6qPMO4ornVk8UN5kuBek0SZZjGcPinu/dxqz2UwOqb9yJ0LHnTsHoLXOV1hYRFi
mKVPfp/KG8OwV25HqheX/B+0tVSVxeV7BVtv+7Q2ObXfjE0myZoZ1A52rmvnDPFScKDmNxOb5RgN
7kJq9hM4rGhT+403ocNLqMfvoSmPVKtqe6aQ5E2xZ74hCB7MsWciLwYIs20YNR2A+/cvI7dUbmor
dpzCYgEpdH/RBKaZ3agvinMryTNsTKUUmMBFnKvavwc48k38bz35EGH37Xyx46vNlGZ1SwQsm2Tb
fjnfffcmvRfZ0fWf+LCj85plvQEyGZIWFfpcqdftS0nRi9q50Uk9g4bCh9OCyCu5CHvA7iVct6PI
UW6HCxL20QC27GN9EOVK3wClcjN2i4YTxaJE5L8M/7YxzS3TYx42FfMtrJ9k+gBK++VPpoqLXa+8
5thrLh2OFhm32upX4F8w5vJ9+jr/Or0TOg7X02hVK+RZ7rvVn+MzD/BgRVvr+WnptEXfx4CBiu0V
KVem4XzXOsaB/cBRQMLDR3oaLj1OgWHzRnaS4E+7TINqwGQA5FiFEAy/tBQFcBQc80FHZH1d8VMg
6gVcNsHyqAZHL7JkqbXc+JzMBAKrN92NTQLntWHKgya/jWkN9AIjuQ1CAD2LIzSMzxdike7cY2Cu
0+9tPL7L0ev+n0LRrvKbNE4bctaxInFDRlIV+3kqp2CjnQxy+fmPjMeShLopmO8w8s+8cxuwpCcV
hGGVv2YGlGEJbWyVjLMoYraX1LGCD+DYRD4HijZnQ0IagN7p8z3uP2OU12/7B4G7r+BL/XZlNex9
LoHmJKBDX3Mwtp7479/q3mJjjUiJ3W1SGVdtNKP5+lEsY7FaynhhksxNP6+rlkfslCNiYeXFNRgn
JgzjhGaPDQ4HN+2sbt8RmHi6NaBSMmjNVSuRWMagQE9l0NlGz6gpqk9p3WcPxd0NDOcypCioP3y4
kAPmV7yKrLeYdIyKL1cGbA9q5kkRn8rE5R7JRpA9GrweUyNiQCPMvSVUQVb1mdIOOBGBsAdD1ehD
SXMwWxBSvJyaE8XsPVHOom2fKXx+Qxa8Gymu7XUoOJWaR8yzlI9csMgJH0RUC8oEz8hbiwi7ZzjR
vTg83B++TCg6hFxPsw2kbcxNJSDTybRFP8TVc0Z29bN8kc+TFzXakx/HGBRFzh23C11B3tuuVvah
1eR60APU1yeZYBdaMahSq+ay7kkPT6IKj0PNbZ3pzeCLR7aTtYXmKGETbnDPmFnwzaIduSpusNLt
HBdOCAlXlG9LU12AIPWHCve5zdvgCiLsafUxkRVR9MSA6V5QqnJ0cB08qzahMFo3j8KBd54LCeUH
BMKKnDIBIW5ws46rqVrRMZb+Vu9+8QBSY2CVK08Vmg+YXmwVZBWX1Hnky/5cgiNQS/bulnL3JhyU
4tm9vGJGARfC3y2daV1y0lsVxs4eJUi7L1afuGnV3UTh4YkI1m8r64c9kCR4lCkoT6QMsvvpERYL
zIl4v2bUzv4zjKrY38/HJlQPg6auRUHzhzTpdIXbXQhJ85ee+S0i0nsyMCBdLuEAxr9HZjmW4rsi
hXRWrwlHPleuSSK8aPJC6zRsphNaU8rl3UenCMZlBN3abnCMHlZbMgQ451eUUfZ0Hlw6Oe6gXTjL
uEy48zbNShw695v1JyF7wGXdu938GBnpPjZK2pfNYcZgHvdgOvXSO+XmB5bg/5vdWAsCswFTC2Ca
RpqpVGda3HUV0hkByB9Jvhd/aGe1lSTiujiXERTmuBX+LEib/cUatuvE+26kvy0bBkF3dQcb1lik
gXIYFtG28q1TDa8yqUaGQ5kcN74ejMUoe2Zmmx1OW+nrkEMDo60dR3ZIrSEoXinVl4BH0xAEOB3K
x5ZweGvJ9Y2C0R7OgdGiuJq+ezhG7UUSXTdiasL3ZPOBOkbroUg0KTb592YNGUxWERI9PEv0c/qW
163ELBeBq/aGCGphSPMF3CwK4H4NaEqfkHY5Py2ZQr3UKBpNFzqZJqfIO1JR1SKY/VDPxSV1DS81
kNyaAAW2cBrPGM7VGIBQrvyzuyZEVER4BpyqPcKgAaTvYTM+pMYlpudiYPOeQCAq+T2wRLvyDkmI
8kqDsAqpflzuj/cPZCw4AHiOh7VdeP8wPpnQVkxDxGLGe4qXTDbkqjD1xPcjRQf8g4uqsjwFr2vL
Qnv3qL6ZNqM7sCa3UN/OFnaLH7QeHN+Ue2xA1KFIrnYwzv3JegHTyTmGdcoTiJ13u9fjG2g3vvMs
gP0r/neJZjsQY4yvJsAX4G7VW3oKdqrsoQAcS4oNEJSI4MAJkE1FwfDVJ2iflWBaASv36hDz3RVk
6Llh069cOWKrqpySEvtzN6VToli4nDf6YX4DNTsZfxpI2MWgx8ijkQAzYh+0Io9gmP0BT7J+q3hd
RCOnxu4z3F3tVRbf1bqCxnGBwfosGjFux6unvo+NwPtxCFR0LDdLn/OKJKYf1ooGeM+XDJkqUSNS
SYeKln2T5e6VW/nYneB32REsSSCPHim7O0YUzLdXumLR0bBPDpNj5UN8bFWdACS8Tu2gDfEUyQtz
yXIpUxf1mj/EqcBsHFOaHyjXAGT0sYcsO0Wr46aMjyoYV3ihk+ctAOUtY2GuGbdGoUu131qfcS9y
7asERHJSVO1TSTf2EyiDrqYQQuYtfzc9syW0gmAoutR1ETuSnpKsENzJN803Lfp1Rf0eVwpbVgaH
YRSvQFHJ3EbT4X78jKu15hy2+YptB0h2Hro7zdX/Osaz540caQH2TPmhy7zHqbgQPAjaXdAs6r9Q
k7kPGJtxXZ29luBoLS7a6aEWYDF2jp03oMkPAF1IkqeyJuRbzHTOj8eA3Du7Py3LJxNSjeRCX+Zk
inNVcGo8erSPw5l7wJF5Imxghshcp0dz/q8ad/25fuKwKdTrpDHtIodCvy2Wki02zqpe2MVHQqDu
zAW5d5CB1ey62gsukfu+qVkKyT0rPAevLWG1qnRHU5AJdYpLSn0pqVkVj1JabOZXKmAL4+PsBzF4
U//KhD/bU7iOEHXWzrKLdqfH2u2UXL+qeFul9gEArYfrQdHtvr7iMFjJNVz5QiSKCNel5vJHejfo
/RGw2w5fd98kc8RD9e6hi64HajM0UEI4mGBqXJEHWPR0q4xAbB2MF4MMZtgTYEW11ouv+3l41wDC
Zc27wwbh/vPgu9wGccgJIST+P8qrFhVHJqiRosy8gN5DHO9qFfin46F3bs6QViPeTpXfLdXo4L+k
Qq2R92z+v253LgM7yTsxb8s+Be/rPt2UUkdMk6FAgVpqcyOtLZ9KHcl0h/OgJ4B78hUKP69A/rtd
3SCCXsnw6NSa1xRMdZpIHsBpqmrepQLC9F0FfePPHM/aDkXN9dUneOTKayashvpFslMt+CO4SHQ/
OH3gPUZDq6ZZInF6yOGrpl4+C2XLzzmUah0UMTUI1MvcAG3AlOunCod2SFQgmCfJmXTHLUAaHS6+
WE0LDtzFPyXp1BDMVuM5DNYeaJ1zUQLsFaKu4oaPrKlgNtogc5WsXoCxb1MRCpI1JKn2lLJnN5W1
JYDliy5as+zHPsdPlttCQKpwS7Lz66YbGHAwNT88wt0slUt/EX3bnAeG0BgT+oiQtj/sQU4Vy1TJ
HoN22LJEdTUKppRIfjWCNOWneTqNMkjRcYM5AeRN0Um2+V/GPWrPjLI3Fgdb1C3XYcYRlRxeeRpT
w/6w0nvn1c3dzEzVvp2OaBaBwP5Eb2IqaGW/RxIQLldxGVJt8x5B4+XOcmGC7qCZk2ozfOMLz9wH
GpZMLa20thhXp0om4oTZFVZtfu0zGVWhRRh1362oqNeHKggwMftQWPiiJaKETXiYnQhoVkzZ06AZ
ApX2GBsqQVnCDkaix5vm8ErITJmDzDaTzlzgIz/PgmSvwO9FDQOB/IGtJzhDd65b4lYuaCeCALRB
1OhNbDuNQuOx6alTqB+VCDzDMt83567R0QOY4kwQrkadaaCjHpAsza9ssXmnmFdHivq525kNOaEh
huEq69kYayQuozAv5jQjM166COJtOte6tCdBwuvALKcOe1zcKsAEyFjI6C8DDsBXrRynATo66t4c
5pqgdjsxfPt6+WpBLBkR6v0gu1cFHEDZb3w3VLtNxCLvFFr2udpvBNFLhkplWvhpmi1YLsAok9CH
EHJyYJpQV46lyeD9vJggt1jdL76/Jpz+rPFhZw4HykSkqa4NnNLKr3q3yiRewoFL8MxK30PsGzqO
MqmmaBNdmh+R+iFH6xfcwV8zIi9YPCRow/LiSrKrIn4ADide8i4nHpb/23ZIEGP2uSZ2/y58TrUt
BaxRppfKBrG2rOHGk1Jxpda8cXcU/UEa3BIEB/3hrE49krjXN1wXx42KNawyyt1BPV8zPLJJ1vFl
jV84ma8V4mWxOH+BP0Sl+eAi42RgANsW68tARw8WKI9lwDVaDb4FVGLqoIDs3feLtUm9ROmmSu2L
0sgb5pKe6fHWh66cjIhQtWXLpNSQuYAY4F0Oixfmpr+fF76i3MUyqmHe30cienhikBd1V6RzxBH2
NTI5mvry+Add/32mCynZxgOsRJpJTiwFK0hEACHM62P36JDYyRx/O+HPsMDqG7w+MUUVT4Ll9FuP
Yv7Lv9NaEbPloyWmRTG6UcuKmpJKYELX2SH64eNxZJXLwXpY7KBWsJrIvh5+gmuxtb1+KaS2DldI
0qIyrDdVhW5LSMS4skc5D9e8VxWB694Kr8mWfCdIrIRLHso+HPcn7jTow1Xr2iyDtsJmgToobIO5
TK2ONBDPFweLKDWDOFxzH1/et/baJzdgYbCPm74Xan1PG6lUFOcPm0u73t6AEMKXREAL/9d94VLf
MLD/Ttwbn438kV3Lsd0kWC13zZCmiwxLlSziaLtBokx2AwNF6fVd/QqHpefpXqwbyiR9m23lb9U/
6TUr5pRAVxHiemZ8J/+X6knArsNcylrOgGZi+E6alVQS1ic2d2xCJ1VslQpATqJtxooCLFlBFwFg
CpTAuVywuOey+qD8upd6pTpEKshf02fhvoW7yX92qJRhRS1uPM/6sHCxDgAvR5cxhJDvueXmHK1w
IngffshESSMVo8yXecBW3UdH40mry89pfT7V70Fq+3g5YLYkgKal2I+C2vY+ntDk6zZ5WM5Suz9w
hI8ZKBUMGn10sh2wudymbtw/teg+Hy7mb72xP4qcM0SY8QodDRyX3s1bj2MUz/WiiAqoI7ANqkvN
chg5+fl69qFTx+DZbLV4sJsCqM5/wmU85q89eJYXr46SPTPM8dk89DC7Wd2+qpO2OOTFC30iZlwA
uKuIGA09RI0nmtbPrQ0i2po0N6en7StxN41Ad/fk6utXEG43xS6Tn+F9Ba+OLm+0MipThNbLwFar
xvpZSgXEFP5EpTf78/rtb9CIRxxiEfbJnPL0UmmDdA5b684e1dTKosGwtOEM8GgAuoUtEM+z7tJe
3gUHBsCx/2Bwahjz2syoAaS2SaG4kuykOqfO2D4TCAh7OQ4cTfWxK3xQOvy29kac6zSe162cqwzi
egGcFDe0/Q8lKpFkRPuYwdDsmhDPrgItTugj+TtQVtv26863A/aqRzj6J9eozZzLnHW+Ml21cnuC
94I0Ir8KD9SGeUUE9vCSLlJuNgt7ig2BHTZXB6bopmUcOJMQ0sKF15obBUKQHs2Cnzrw2X0NFiLE
9lXUZgpj1QgIXB+6RZGlqWHTpy3G+eYn+LKcMHMdkKXtInsgGi0j1f38RN5Ilpd743nKFzz/FhZ8
Lo9+DoJTVP3+pOBrL5niUNcHlcdcd4RlhF9NWO1zgWWgiQJBS+uJymBx9pW5L6EMac7ji7tsLj7x
6ZAMFJirKzSuNUzxfrNmvUq3CKtw9quHJfd5gCqY83uiKoNz4R23LsO5zaz17F2gctsSjmi6GjHb
nYu5bq2Qk3+QIGoh0+qX+xyJoIEkTcARDdGc8jngH9NzYMmoTKoWQH5/kTmUgFwLbDlsMetvrZFd
3gLbWa0/TE2CRbZyu5RfGHUBGarJV0dFr8p3+pMlJjbqqOwBlPQc+WiDUyW3DvMmKr4ETTSeqcOA
2Js+SCLkYKP4QJ+++jkfWxvEW0Yrd5YLeoloZn5Mz4xyfBQohrtBjZfryzU4zr7iJCK3JSIwDlS9
r6PqicgaC6dWuhSr6qms0+D/xqtVJxshJiZMtQazQSdLUJmVSgXrXTvIQ6Pz4JJHjVJeM+Xnec94
ASZApl86OoviVq4QSzq7UduyePk9v++CIP+nTDETO/xkVIqHO2Q395eaN/JcWZZQf8Arh/3Nce13
1gt85BPoCT29uPZLEzMLgWTRs7WnZWrmKy4/x7vosYxQij4FtZfPPf4Q2jk3+iplA1/ebVnXTRVY
3/96rpWIAaOUgIVHZjtNVVd0YhxHXatm6i7oFGLvRamnbeD70eTBwx8XMZxiageCgjQfX83kgYxz
VV50PQvpADde2aROtu1OT24LcdVZa7/FSCMPxNei5G8EAOaGQ4mfsDtsbwhmesXBtcxSED8DiAOM
vx2+ycQ+yZfUNuJa6Z5X5It9FUmb3V5TJ7oHDJ/VawuZMqfb/Rt54ovDcui1fLo6oLAy7HoU7Pjh
5NVlxDP9/SjPDi8PJDdXFNz1PkyN1afP+MEcNvEKYSHQzv4mRDDiEYklfy48GXyHB7NuzdEjMWcH
Mp8QYNkpaF4VDJNLP56BOWDLS0HTuEKrn5/DisbSom39qoIHHrS0gyFK97EvKYOutO5ZwgcEItrV
ep0okxmzeKHg/LR556bX+vUGyB4lvPpWPuzkrBloj2sJYRMdYLB8f/8DYDDcFw6jrMgufMiF7GaT
dzTW5fh9HLb1JzN4YQkLwbtvwfT1StEnJTFTaad64b3MNVl8MZkPR/5NMyUHHu7cqn4ONuQ7zfbL
1Fxjbkpo+SqfDC41ISzNhY0/8tbA8Q2wRkWoHlXbqs2wCtQxaf7KmOv5U5wgJUX2eajgaYd3QMxt
sjANen2oLoX+OicO1fQS1v4L2H8mxO8fSyUa8/GeNyA2egKQZoEj0em4k0M9jgmAvCLIvo14vYq4
3CM1bVQddsmO8mY3PI8vuWVZLYoG4d8qU43/QCnpWkEhCPlqWJcMNZHEfMwcvFM+Az8ZCqBJFV+O
BJHfh2/dWpqViBhs3DKjtaxylYJXtGeot1YI7zWQkjOB/4azlEsEaveFrrZppo71hniZHld3Irv3
fYl9LuuS/oM9thTCP+uKCPxEHuG5aBkX2OJ3tgNpVlzN1a7cdoaJDyR+Abl1J1RvggMJQE6hr8LB
8c4YsRfUhWCRwiQ8ne4JaFk6iwNINvuu1fUFjdsy2tJyDiuabJ5pXyvgl2UNKVCwFIx0GsbMBvAw
qEWRSE8E5Kr5d7Ps24cZJsreU0ofNvwOcfXDnbrdqhq1gZiFPw+ocfUlgxt27Tm1DNeojHXc9be1
mSptcdEiiyXn1j4Sbr9x50x5adG8Fy8b6ly0XkQlkF4Mt8TDtYK28owGBWqmbIWx8WyqUfrzSjnx
LwmNEM0mV/exwxZ9NjRTkc9C9T0Ag7W/uv8A1Rs67NkJTWLM8LfazQ4FRuNVNGy6ej2QPO2VznmV
FKq/k9uFetFyJtp5ELwXCZnQpQYlgXFL73GETqmJDKrjEBOtN5UMW5YknnV4DeqCrkybQSfYAlqi
MM2r60X0kJSxU02NXO0uJ0pndKKqZE51XG0g+O1kMW7t3ljarTIYPfS+4nZnPCT+4BanJG0S9sKq
pmYivZ/2JjGWFFLUdE1YO3GVAN+hGAP1mi3NIrWS7NjeP0bSvX4rZhj8ai3j9wh/xAqDbker2fG/
u8jgsMrvYnC8E1m+Go8T1eVbJ+YoV1X7slhSVDdh4pM1XUM/2G3QsBII+5LNiCgzXmEEbFqOSp6M
IgR7xvN4FhuGzuaarVDEfaxwcOK5sP5b5xwCYgEs7P8XGf4uRIevDM5MITsusXc3VzDtRCF2XsyY
7P/Tw/nUh8doJXNV0AnHYueAvWmwWqL6n9fVYct3tKlSQztBNbroQTEnYnZK8G3Wcm6DfZWDQ2y9
/3OBIx0nU2iIdtaAEOL6w0rLtCE5kr2QV/ZorS/E1fTGU3j90+khxS0aQLeOTqgTpQw4La0m2gto
K22vyqCeOAdYXw06dse81yaPwzB4FcXMHjEQw4yZ5Lqu8w2Pol9qtyxcTrxFCPQZahMdVjf10xfx
ZYd3pIGivSYXXbXIdYg830+qahSduVTuSwUL+7NqRsgiCgGHUVferFZiuSWAYugs7/oisLyHA6S3
lbkuPMRxyb6jE1arYIX/uMbVDnz+qtt0jewIj5Zdb/p1Y+2L2Up/P8n0ecRDi2obrBmZbala48cI
yzBI4M9RSqf7+QJTY2vI2CrX8sK2f/tWx8Z5r5TrhoXsN0rMpR7iN/winSqYNmwq+L4wTGD6A1cY
t47zbkf2OiIRFSXhoMjnNFIy/mIvXp9cmLsBCh5Yxkzq2ZnXhu27RwpRhu8Tz3vEpbeuwbWq/nXx
7Il3GuQ7zmUUnmbxY4zOHgjOx3SEKQQgL80Pg41y0K+USF1C+onsFUYhqrYmxm9PnoWyFPCwpDTb
TeZOBEDqlSax33ZmE/aOdYaT74wJ/DzDMgCqvkb505MK7ty5j9J3Ky8F1GU8A6eMrO/mH2wkRTp9
Yk7rSUbR7RGiKCXGAAjN0BTpwALP5alsMzfkh1HYhRki0nnh0KuYAx394/G0PRaGfzIHKCkq1Fsx
AgnxpeH4v8CdJq76s8QaTkYwOJqUw9KRSp6A5XeqlSjrfjA5RGqEU5jCNsFV8r8mK6BGTEZWrTyE
cQyCYXHASCcPbsPBcWCPEXfGbJukEobsjlyfMi6GeJFcY4GPo7RwRJTKJWgcQTqdeTfp0NQa45wo
pzMCjFllIKBIiJCUPuUqsFpL3MBMJOb/hYqz9bRW6fX3Kd72Y7jjlruEx9+UcsalvmY+gIi0HlX6
tYR1oILsq8cc1QrD8TuH1aVh12ahFDoB7VnYpWKU3uj6k9skAEkngBJxEauUy9FFYidnQPQcNotk
XgZ63NsDadVYurWPxAuQExpkoLO4oi/ZbJiUvUN3KBRSh1XZ8oFnhLEFSLQt60oGDcf7J1ZmRB17
fb19XKTGSONakz0LWLom4O/2LMWfNvsQ/Y37ohKhlnZSY6CZOjqq8c0rGjlAcagkBhpUE98Xxz2V
p3pdo69KRdcv+92YfCBkcwpoHGMZ+a4s652z8IoTQrp3Yq6Fd2pX24CThQn3a72yuuPm3x8nsKbX
+snz+RJxLtvVAFGumhMpdxbno0J895paszv05g+mkEfqgdI3961oIKNvR1M6QjwqDpnqFJusKM1q
W/mIU2XyYewlfc6R6gRAJLprxgXyiyb9HVbpZ8bLo/h5DjLbO5oyWnjvyQ44E1BfPSLXDOK4bb6e
VtOQJKO5z3Nxn76aCz1uDQAzK68cdJ6ogK9uSQ/FdyfWVnuxwJrhSQ7jnhpEafUVvzxUXhg+4QGt
kbySBbDEjz3rxf7MexbJt3Lo9BkffMwP8y3+X4YGDm2LylX9mv+Rrl3fONeHt0nxSs2M5Q6cJGpe
rWV52rH8z5oVuCKU8rDgz96qeOUJs3eiaZpxQ5Dq6FfBr70m/N4d3uZbtPRuRCFjYZsIDYEHzi3G
2K1+p4Di3ISbYZNCKdNwyMfgRmwiWaDaDqEJr1pJHg5of6H9peMutj89Mp8FpcOosM8wGX491l8E
HBY0HjabrV58Ev9mJHLwcxkJybr6N5+p8eRPvKfrdJuqMBHVAkVO0p2oNcftXZEVcnwP4Sg5SJs3
MspoC+s28DuD2VFhj9h8vDbpjA23KAOw8kx5c+zBwVT9OJmqSSn6GhcvGJy2qHBe+dyFScTdL0Iy
Q7RdkiLkxA81zm2wDlu/IfadvvITwIfW5oLOtuV5TtZ9tIOwvFrA/8clBW0hkhrze0PkXa3KA/E1
7f5bESKkfp4nZQjifPSK3PUgkHLwoNcmWhSZDSA6kWWZZ8ON8vcPii66o52BoWrx++U4LslFwS5S
rwm/KbmLG8hUCqKABtlUFR5T2I/w4aEVRF2YI7Co36XUAO7yL/1LAdOZkwjGmAVNLM+3DkXxN7xp
pnBkej2uSTBL+nN+a0l/v5/2VPjltZftxiPkEqZNn8jK7HcdP0/09aQEoZTS5VuC+9GB/HrRoAbE
JZa4EMgv+gmECkM/+lzECT/1vwXBcn/zo/ucPUade8gtIClGB8BCzDNNN6Bga6Xj/w5i8tVXO2CH
nKQobAJpHwGpVOk6TF3sql+tr73zFuZi4QEBLdKcwKgOTtZ+4zSb961R7B9qfWaWtnvf3SUp1BzC
zdwETs+ztIYafPnfBgs2xdrGSaWowjc08EZvK3G3Yf+LomkJKjwK6aUsZVRCbKaUH9O52kX2R0ZK
gCWMQ9TMmhmtnQgST8ybmw+p5p+KMCE87EOjS0qYmjtQ9F05LzwAOfZtW65UIfXwbI5I2q8eax3m
1JRBDPpxpht7ijzN3bRrehBSp1CZVgMsY1Bg3lazxMlMxAjEAz277ekXOA+7UZqjtLKCcHcpQ0ru
LTMtD3qfZmouOscp6i9F3uHqZEANCE0f0FC243UUOARMBcdbEX3zRaTJkhzOSqPkzptWAC6i9hJ/
Sxf9/y7OvnWOU51kugU2w03Gc3ojmSY5BKod91ga2qJBXleltHtBl8WL6Jv2a6wyTuFYdVkir+b+
lFKJK2lEWzkVsvs1X/Q17sCKGZO6vuiZuMDn0ZjL4wq4stj62aK8hfjt/ygOnnkCfcewHEGQAID/
FGHRs2gaYtFFNhD7tjtva/XdNki2fP4Z1Uk91zsaEX2pNYdYIFJR0G/JpyV2VF+SsicN4mu15PAd
dh8cXP2vPP4wE6mFy8DHrwDtVCUz4AkIaSiEFzAiqsMgL7EPdanz4Q9LFzmfXikKkI/daFuJYaO2
j0CjBpoI5qkqecVkbFwhycnra49WxrjuMiSDYbRSRhJg0Nh+tU2GQbjF01ppekLkDGZR9zHQQiYs
SkLkHFAZMt5GMEsGhp/fSvommNX+XTPmnHapqVg9yulX9OlQUI7SJqdb52tDoKONXjOx3DDsflWE
v0W1KNjvrMdNlLr2HmA/fS0AjyfMmjPAYHv6ssih9Hk7nGvNE7IkYOcdA2a3IU+z/FLIQ+TjgVKY
iIZZefBBYNc2QcZh5cm5L3PHvWpK3BRPKKcxkQ4IBfPLstW5Sy6noxb6aFCR0j2a1+6sroLVfOp8
hd6HUK1CRCxEcR5jHMcN9jL6f9uAB/WOxiCY6ENfr3YPQs/D+glXGqnSdW19T8QMfpPM2ng71OFv
PbdksZ8Uz5bDbmHbIiUB/gwanxoHpiYpVvXz03sfU+DMXtuB4KvJDmZCSXY463h9KQWJqLu7O48s
anvd8+xHRzwZw1E2FV6x2U5gvpzOZ/auFYveRUjWrVu8fAStcMfu6C4pmzSFij6SvntcZLYk1aph
QhGz0v5CTk6GT2z0pb3wQn4J8iBoAUyiICimxFSKOx1L88xZ6P4iDRIAD6ifivQ6Y1j1yB42M1Rv
LS4HF2iR1F0S6v5A6fw5pU+xz6GJ1UqS9zSxvF1tHMUSb1VK0VGhFjsNezQgjMwg2aXK7zUt55na
23bylHb/AK5MV6DjgyAPYuqSFLbvrBRpe+4/y8HhG2w1mooIe2ZiUpuZw81QfMk5L/vSwTP4rw1D
naRVf+FqDVq5gUt73gfWKebATmiJqaGsRcQS0FAMGYZdzWSwqoeoankWiX1d6BZ9b17ktB97zOvn
756a2a9BK/HMW5hqnAdaE6dGJbw6Vhx3XBpr5AjKqrn+ySnPXCaKFIH4Bzlv+fde23AxrFXV1n7R
Dpb8U1dcZYA6bc1r4aGekAZsCjS1lLLBDxCmfqIDTdbgLLm4a3WUJoCv4c/u0gmkTJaTrBxmXLX3
dOW2dJAxbrKwOLk+4LLUR8+AT1pEfqH/DP53LyMPVpYsuO4TdDGLkB6DwHiKg7w1Rkzs5wz0NXLP
NSDbrDZ3tuUXv81HYwnt+vOw5mGumQm3eQX54kRjwvo8kkIYELGCFI29n06UKz+aXEbYQfRvp79U
A1YtQDLLnNnrazgdHw4S0i+s4kjZPs9/bmMHNDdS/drcBhUPr3Ek+QtpUTdgZvO1k/EpwSa0+k73
E1Y89jOHAtp72LUIst/J7dXHBSzX13M2zXqYNR4JkNxgmVQxyOWZjBeRzNDNVC6XvdsrTA4wfdV5
LDLpclLJqz88qFMQUzRRxVE1moA16qZ8ISLDMPeW+26x+/ALL3StIkEnPwRss15J8nvmHaatgA/Y
2uOEfVtaBkZO8KBMPh+dBj3NHEMeND88Is5FDq6VwmHN7w1zRQ0JS4Pyizsh9UsoXCHNrSwqlW0v
2EJZdqBnMUZtwqwNfSwQsItSMwtW/n0nwqOXYPfravCn0xMecBco/QMrMu2basbvzJA/AYSQaIWJ
svkm0Nn00xmTodK+r/R5UObl6fr7BBZIdOkM2KYpeRCtyJCeF/yvGghLA6rQxaYzOKGXFwhH/O8q
o4wwsiCdJu9X9nCPZHjfSy9Oa622E+LsOHU0XtAKdEbSb/hKT5BYRn7NFD/bNAr8/ZTr9eGxxo8B
KxGWZJAoPw/4gjrPUjupKwkp2n6SmmG8ObMel8vtyVGQLlJKWupHPxkqCTeHfMasuFqNZvFVLP8i
ZjFwhdI20Ph9cD7AM0ypnykCCKhFvYYnkwLW4zvS4daiNKTp0XO03fGNzY2JBTAy6r9Exa/schhy
xbHwi+TCpzw+zdVHlPph45CvHUXzeS747ZdlnJEDfkkFRImGKFg/qXDZbLPtCoM4CkDoExfYGbtv
znqlsPjbqhgwE4NpXZA6QM/0Pjj4gGkhKq88+8b9NMK3gL5fZOW1zdqw1llHBHTJ8MzMDz4hW9xu
m1zzZNni1Wy9wEaJSL3DZqv3eRlWFreSPhyCEKw2e7xitF49/gCQkB1j8KhHjnWLcAad1nKX+yTF
KBNAhz+/DwfF66N7PvpgVp+GCEB+nBg4nfiMarpwauYIYKCkhFHClBtcvccCYElJmY6imrtAS+D2
JEk5Yp69jsiCvQGQ0saa2ElV9EJZLyeu0qxo1MVtdqL459IY7meciYzRmF132GyUvKYfYz4mO0GS
5flPCD5qL7AnwxWIUK1D/SIzKjfiHp7sfaOQl1BN1QvXvZk77GQwwT5ktEtKwHKTXqYuTAxRE4H6
o88r6yzEey/uNxoZ1OUvqtdj6VGohOO7k7y5eNNeIqc61Jf0dSh0Vr/wCAhENrpZEvjyflOAXnhF
CWd5SCKPXVxt+WxhSq4XHJ3QN0iU4I4S4J7oy3V1mua5OsBeX1reyvOII3qWvSVP8sldsn7DWeOw
+8Hq7VOzJXgczTyhTLbAst7m44spW+O63K2CYIOgAnhfUWWik0+CYtSgfByZrfML0ORvpLza0ASU
T74tVa242uEjf4bPUDhWhBp9TQXum/Ly/9Www8g1xq4gp3wZePgutbXnC7v9KlKXgSMSOXtPRqVd
+dpi58AdvRrPwv4GkUfoRbOc5eUsFCJcA9cqdUBBGq/D/0kftH2CYtzINhMlfWi0MdVolCfKEI1t
vGoHa2sV/byLjbpWaQUyl6nS0HieXpUEYorkGd7t+kfwDeLOiHfvvdFQtqF1eKIYRzOVGdBkBMlK
DXyw0zjFelc/H86/gyyrmx3RjwNI+aCohR4eWGSXkI/mDy5roFQQXpPXhPxu1WJctHMrsNxpoeZs
AKUh3cLXm2Hgr8kiND56/ivPP7ESrI0oSMkWO7M8vg3m/tcyOGhNvcbafw9JPBWkNGYatd9oFjc7
yfE9rLIu8sZCuKt+0Z3AfNVDJNoRy/lRZ3CAA8umt1d7nzJ8hdUTedDe3yw4Aev4D6F7WxK1C7I8
PtoVQ/AEMVDa4D6G6rvrEKk95iyukGoMxQaAppUpjBcgTTOvqEnWfQCmLHreeCuvGwdRO92fBFJ1
EGl4UQAF5PpYThVEy/69TFYOTbK+vLY7otw/y3dti6/BFpbhrBiUXLaXbscMoq0pIn41aGK+MvuY
sJzk9SSb5mF7zKmuuuTyNFi7y6+Sol9QmKGgSyQfA7k/9DLS4rW06TNA0Alio53L2P1ETtZkOl6C
gWINVJ0SzAp/xlu37cctBMKBJdjlF7UQa1oBVVrNMhBrfF43VBieacoYLuCYCgX7DBzCQj+RZEBZ
RRpAirAMnkxwyVGtMbC4yDg0PYF5vL8tQyKwL3ZjegBdgeTyXB0SbbAc4koJuLUzTLcGh2MDWgt1
atLo5XEh9H5+GYSo3zZ+MF38ufrfqEcQ+FLU7LhPEkFNN4DAqypR4DUS4PB0znzG46yUyIyloBxH
4s8ijgukfrdQl5meKRqIBaSYi7aAlGauNPMXV5Jrc3MJhimkJ0wF2dD8DJAqpEysQ6osvUNwlwkJ
daAdCDr3t8eoX380sebfv4Eb3uMoECqpWQiHe+zHjw6OuJxKUSlDCZZ6z69rxDY8t7t36X2IJmGZ
ppYEZHPyViK3JdFWrfD5abD73bd9FS24KX6S0veknUSTLDk1nRoP9i6JywZGl/Qv3FR6FF9Afe7k
LMzeCvflBcsV8qN9fEzD+k9r82FdgnmqBUHIkSO1q+6EMKxy1A0CQ7pDWEKDw9GoZiqM8n7BpFsB
iDnoQrU0TjsgGSd45TYYbak/CItcJ9WqZOUcDhvkYOgrQcWI7CnVv3WIMtb9CMytnr+siaEvCjRK
xyU660MN+ujc2AN0E+DpN3nHivb4inAsEYdR/m+DpN5BUVtzY0R1LYyOq9Qk6jPXPmkEzZtth+rX
cled68hRABCyYepM7LgrBPLZF8FN+12lu10V3iBKr4CZZB/6UhLbv7ldFs3bMsD1XlbD34ARpjP7
F3czqmRZlVQAfDitTAkoY3edaM0IigqOgCtsYa3mTwsO3Ow81Bwbb+qbKElRO0HGwrjYPGyZ4Gxt
yC+1pC8lAg9BjmjeH6ewd1pbbVDDEm/MMjj5aWwip414Cu5+/oZOwvT5W7A5EXKmW1BASu5aO9eR
C5xHDRqYYzMRltimrjYXNOQsmTEh8I4ONU/Fa4ZxYU4T2uHU3ZQ+cH2f7gTi7juOsgZM0r9ScCNJ
/4rNWRKMqiqtzGpemmMfr4cCj+4Q8DPfDE3C3NdAuPGdJXtoG01P43y/HmjwejFowMB/NkqIgcHS
F38uLFsw9V2Yiohm2m3rOabxwoIHk9Bgj0mFC7wSTGL905DwsnLwnNUuC1o8/5jNAwu8Y0aovIby
joZeQwDx6LEYAS/ORvz++us3GxWt33WoVXO6p3ULZYfC2LRZyko3V87+6iQjqVXjS+cn5lyTq6Hd
6HjCFRiEVk8kU1N9GU7MQTQ4eh0+/zAUbAxzR2fLQiBklGsmkSvv6sdm4LMgtqJ6IqW+yp71V9LN
6CAI7w7uO3rpqiZGE74bzk6PcolzgNjHdrzp/yBalQm7Q9KsTmKvuFGeEVE9XBu2JDa02Q9SdnRr
nOwKWQl1tp4xtFCCkaimflAybDRinY7hbTLUMPeASzoalmYf2V1kj5z5FxSBymyXk4e/uGzaQU8Y
CBE5F/fjvWWKgB2shBmVNWbb/4JY24GETmbGOFmFxoyL1j1UJ7p/8bNOBXmeM3rwxt+kWnCxnVIl
r7HL32JShfPdduGFflJldgayBlKmjkK0PNEo3rq8ELycWRyyXrOcbi+3ZmwrgPMBb7ifC58BOTND
ravM0nX99WEWkwVXPW6hbrf4k9nXWHwn5QCyturSP2Tr87U7w0G65JscxmdJNf7+Anl/Ha44KTvJ
PsC39BEo2lwMQiMoODzw9gC6aJRg58iY+PayF+Io2IUHiuWaGxE3XyD4bVlz/UxOy8cwfENStzKg
33DqrwvFkhlfsJY3lQe/9p0zlIHkzDyYzi17sQW4+o+Vot+CkzSnjMFP5s29FpZ3S7r7STIXHPQH
zCR7h7fzgpAxXuUgSDhtzty46+nK8CN4W/OWqIpeL4s8CiisVTlJKyiojGBxiVL/5wdQzYSYSBDE
UK2cbW9/UGcPU9PDc/3ICXSSMhDwNxEfXevT4ObkCgTBctGatPUGEwuoYNDqCqMdyx1RpHgovwYY
NbNDTmY3PzeSsvh7EnvUW6twBS+JefOYSXWpT+P2J/Y/y0tneCxInyJmE1YLopeYo+ZUWjbaApeU
BaoshtBgRr9fycfjo+L9u5jTZijBEKTbpRM+qcgQiD0PBhfOvtc/F0+mfSPlzwgA7pOfTpcYCBc8
eiWKCbzYF5Ny2++Fb9WJbyVhgU8ait2S1t+oP+PSXm04OHKndvKPDA51DdT2ZvXyk4RieX4f7dfC
DM9/FViDkA0v6uNILYIFSbpdAnT3YjynMn+VMPR/q4Zve5gUTXdmqAprlDNkXwIdbhDR1CSMkb6b
dqLfnRa+coQc1mzMqUiJMNWuTXnTGi4K93Pk5olb1s/dZlNfOb2MN/eoDkcYubE6FGUUR+hu8BNL
ToUSaT2xUTf3L6aza9qgbImBSUbRUE+2fXNl8N4Z+a6v5Av6p/hsjf3vVNUB45KorcFpp81WHq0i
kOSpkcy2PlsmWgvcjkQcXn2b1rrZu6BuXxdlaopiVt/9bebPv2qXIa54UJ+h3xwWkYnoQC/B1bLs
R13pyhOl3dXWDlBTbrw9W0SjC9JczuLArw8np5k6WK7YFonpbm2PB5TBl3KC6QNnHKOawH8WPH+i
yzcXkHPflYXgwIong7Fv/BPI/wTLB7I6lKegor0rBzTUWa771yWhQdft9BxHbqOE8D7Yo1BA6SIh
qecyo8668T7GO3HIgkCbi6Q36rQNFZVnyyy/0qOi6JwY6K75aGFnjRHCEI1EDej7Irm3ilXcAocH
p126ByKyHQ5XklscIyesresUrcFovadPCImcKt075IypV4Kfbdw1X50hszv4geChyEtFpGnJvrVn
aNVMJWwFw8jupkyHWM1Nasu5jaySIKnMzBtR86kijgKa+MkiLa1vBZjTHVhPqWTUdI9H3Jv/FCjR
UOf0vkV4/cuXljqr2Rbv0F3zQLf/K1WUIHqxt7KJPjo5ckv0ovl1rtaFSqJCBTFH6o6I1P8sz4Hi
VHZW66tSKfnLW+1Utmvk3bDbKxqRHpsKF/1MW1xjdyOoiveKXYnjcJmf4v1mZG0QVTc3UgxV537V
+SUgKC73MvsWsQBed/AN4GFBsxapwXnaB3OHeGp1G7hStEWJwyUtco7EJiz1ReaOE1zrC4r1ZoCw
CGF12QxfN80z4rQNCR/uY3aAr1xY1hWvytqEAptGW8ndjrpJWZkMWpacQ3FcyG8Zd5djEJGo2yk6
mM4Sw4M4R5tSpQ14XwUGrVJQ2mLoXRfrQxCvnS720qz0vGkLs/9txP8N7Fxq0jRrnQkonK/QCPDM
/iG2bX0F5mcurP/lLrWE2f9eioG8UNLjiOdMzLaYYzKtunLcCpUq0gfxhbU03sZ/wUX5Xj1QlbLE
idmHaBykecfn7xFwKtocuy4OmIBb1zzdItJ/bAKbpt0+NFyurBX5JN/qZzKtF2Z4I9981qkOKHv/
yc42CKmJGAcxjai8vsMo8qZ4AGSS3B9T7D2yQPjKHf+xHCWhCVRI48FNdYTnpFUxlgiSf4ylOkNC
SxuADmwdviChzawlVw8O9h+/WgAMkG2CJ6m/ItItw5GuqOLhlAPeGYHiHUKDjA7EWYgLiX2zmR1e
1dMeDPPp5fJkK1KYNiXJ1q2ax5KsMk+wKm6LQRsr27idhz2eWfPfYJ2/9b4YfcHy5cLNeYurXFIX
PqFxJuGahqq59bNoa0/hqCFVvDqHhjh6E4wWI4w41CFC3jv3tLyR14FGOFFfPREM6iASqdzNQ/qh
L7l7Kld+VAKHupXE/C+rqyGIMrHF5jyNOfnlGF99zIdzP/UVKOvB+OJFNYiWaeq6guVjE4WEUF2U
9DugGRVDZKuDtEUBUBHpjWaB0bKhVAtDL5eXyfvz8sVAyrAFV0/KY1ldVjh+LQeuuywI1724fLeA
j4F5265kAOE+09rCXrNEuq953t4d+fWn16NbYYu/7KaVQDfH/NiaZuY8vdEovmAs2FwKmdI4pITR
tp9CCV+e5/n7x9KzAWlDAPBuPZTMWJTb2mwAnpECFNHhACUpo0Cw9wuUQT0zbfn8VMzubzOox1Do
+vPY4QQMUEggcICF+tttYwyE3GtTk7YNBZrCVFUwScSq4SqWIZAdVO3oLaEIjCK/zWukZpcpjY/Z
3L+bX09apPMRTb/xFTDY+4WSr88jTnmUZOkqa2HpUXQ38qIVjwaf124JFYiEabwCXqNuSyaNslZo
pHU6fcxQAH2Od+AtWfm4ZKU7duuquCDZdOdFPxaI1aJ2Dze/opsknsQi2W1c8UCptYd2YRR5ZUzz
gQrhJyJgXoMBZnqOJQKX8FPSmthXarXhL90LQv2E1Qeizqms9NnpPQZtsBjRJCgJXpBKVEHtZPI3
9gYQ+i5T+tyZ3mDNnCH16IzwVHMAVJ6q2xvQ+7CfQfDwDvXkmVsSMCjnaa616tDoGcQ3Fua1Gwhm
D6YfcB0m+IOlHpnF0TcaVIejor8U6hVp982YcG7O74q7XAYc1u/R11401o0TtEoyWUzsjL+Lu04G
wA5yxK0PwNtxk8rFS2K606kA9HDw/10P4mf2WHYX8ZuFy3PcoVxPN85Mm0HBWiNLHRnht8lZb+pe
hEEPavxDaZWbHWlnK067P4ui9iYRmArUb/xDx5nzlWLfuBCdFe5mlbgGF1238E33XOO89aVPIdOj
ZgI+DZM+u0opLq8tmkLqzCl6CV0swyAKCmX7gpZ1Z54k0hhUyG9n0h9xXRSbLHXxW2OWBgZxPNP2
ZvxPzZfaNH77CgR0HJWzD0qA6sUMJaEAWL0jQtc4egiH0lAD1IoOFa3No6hGgA/DvroPoG/5cshQ
pSCDHLONDHB0/DFUoQKg6hynUaf452IuZGBwKtolx8pIfQCknvRDpTfLnQUOfK/kGiWDRic01Uwi
p5KrchB8E7andP2cHq4FuC7VVptSxqkW0my1lSabDxahZV0/2lF/coNCd9rWiGskfcSiup98t7ON
sf8GuNj1vScVw6WSvGol7H2LXT+hO2dzenri3dxwBOPlHui0uCOtdf9lVAwSRXzysVkyQI4xe7A+
JS5agF7/12bBP2XdxFyAcLybuXvoEXh3g5dtLjdLSFCM//TPmAEFOI6ucQhSxFAmJ8OREyUTfLIh
rUBc/4Iph9pK2S6N1AVgiXwMUHii3S2OBMo8uZSLFmuznNUhzAWLELi+McVpxzNPL8vsyyokpYGP
deXsJEHW79d+0+dEwwMROVctJdo+gsNFcZ/+piBFJ2eWoRi4YPNyHAasmhsNLJjnVf3+yAE1gxpB
4txGvEQ3CUt/J9b3h3Y8Amf7eABNaNB2mJNU2gIzC34TxzN8oIgcOhojAQOkT9/d8yDTvvQRZq2u
/YhhUJScTFD3ASFW1QPOQbUzSEC04/TBGZmFmMZBI9tWhTyTvpyfXqy/F0AAj1hljPhKpDFyU5PH
wpPuuIwq3+InQlarX3mjlOzsIBhxoEuC1Fkt93anyV6+6NiPsMrujd+bV6YDmJvhKClIs4vqaDZW
TJL+syjEviw2qxWdUZKogQa9dBcf1NU/+YuWuAWMo95EHzAsnQJmk/rVJrgnZx0gOU5pv+wcyCIO
mSPlXVzZCw9PVFyZztTMpcz1TaPt5Rpw9KMcKp2N3fZr2kjrdOrqr9DG65kUxlOOccJHSrct6Aik
MtpVac70rfVF2cCUNQx9DruTAiz5d4yTLQhM3UrESlsF38ru/quS9NXlja0V2DAt6uSqdnQPYvt/
HIxmcGSobJB2ZyXrG126M4F/q3xmQL2+XuNHIV9C285L63l15fCyOgHkUFznCFPOMEq34RsG+jBE
nvCivySYfj0VHAwVh1NjL1BlCh9YygKfVw2aRPT2AWRLxLND+td2fQMXkK2jkphHtUpNnUY8Jvjz
l+zeYMdVs7cxwQg8Ygpu2ViIYFSMZ3Z5LrquO8CrJiZ/WHCxLwJEa2xqthwTCbbFS9i1zA84yZvp
XCdn6OG9Mdvs4seipnShirhaO0nuNCBOq3wXYBy7g3HoTAzp9snvmMnlM+MdH/WsdmvNwy78Qey+
cKso6HczggtaBFplCfdQxCR+gjphkr+xVQFptIO0TFc6zlbfPNmByHDKXLrrMdE8G185LhDuS+lw
+2l3XSasyFb/UHMaTGB8ylbbAJ4SPAC4BEihVXxUdr3Ol2MfSlIvYdJ5Amku7b2jF+ixPpgSEruc
iNZu8d3PV4y41KXljOdDh4KD1lSIXbMXfR561a2P8KyekmHZVxAxL4cnk9FKGVDBdpbzB9kFHl0l
+p+YDjSY8WtT8xMZRV0Iv83U45BNHMyEETlMWBAG2/HfYeVw+pg1BS61aSOd5SrcYrZhKplUyeba
GigoLEDYIUUtuTQq+alK/C6pZNVt9gsjwUXAWN9VNoY/IvL+2agg5Zf94QP9SKLnJiNc328Bmxvp
M5Sd6wnGckcyvpSWUOzuRJ01EjF3Xz+eJ5yEYnxCiDZUofQu+IObd1Vp8OnruVIl494GShJp1zoE
j+e3wJNK59KregUWQDiSMncpXnfduvKpw4uwEYs0ZSeCdRwHc4/eJug/9fPpYX2SwEHCPYOvG78d
AoFXsXGuV0lKfYis7DpvGAuW5a3bxGFLDCS2TO+JBD1B4kV5qqDEbXibtnpEyTW9cD0TwGankPdV
+QJTXBHZeTJiRc3zJvUsyITTzDv06wX82cz9Vqv+2fS4zuBkqJYwa4343cORuSwwCmp3ygzYu0KV
UeIlI1lcZFuL0ivqZ6j5ZbTjI6KYfkzv3lIYASdaIQLobwIB/Blo5JIBq8VZKcnetEgE2jxY9z04
8FJddB1xb3l5wncka9lC7IFtjv6erYZU3Nyh8vJT820G2ad/vcDdI4+dxkqSwGulpo9uQqfHy1Yc
hHLX6Ym1dbbJs9tV9Vqg9SdsclNAwS2WgzH+zwRMGgksIPqnZJR026krCwMVszVIetxLz1J92wQ7
DNfM+YHVXBupyF3Yl7/8Y1P22W7zTBmhXsTnGx/detPIMv0QPlHNHGAtofy3dQAKvVOD4u7rnOzL
Kp64Z9U4MxnxRSnqcMag0QMZls7R4Bo90dXqvIpD6AdAx4SvmDB3/kuaR7x1mkUVLMS5MsllF9lc
r8OzDtuumqABn2B8rR6cPGc/JDnW8wG22/IOuub8oQ3C7RadCw5o9XvykVzWwcrq3JPlsdM6q5cM
S1ZcM5BovJ5s1prMP4vT333G2RgFGuRsrxPsjBq/qXE9qdUxoAB6VSbtJzmEqHxczWYic7T8LWJz
9tr3vpa7pb5kEdvWaUczBSTzdanFZy6EgPvuJRQjmhNFUBxhr/pJ6zGH4qRFE9LoEEQvDPzngawU
s/gvFKgICNd3PrXY6tQcladKeAMOxZY9hcc/LEFiq7ZpFX24t+/UvQ6lgwfAUDEsHBZfaMTF+TlX
e4GhGMAQ+l8wdHWsQjzf2+OY0H25i9g/yUksiyZ+B20uQgorO+JgixPssijazl+PjrIFH8kE+cQv
ezK60NK6Fbpo57O/s385rMJevNdZxgRfc0vW5BqbMheU+sMypPAhsS/HkoGBf/S+Rtgmq05yMexm
8XxZcq7YbKhlFdrK3xyHfdN/W6xZGEsV0Skouc/ZRv7rgDxTuIda5i3/UM3iFnLIWwV5oA/FE55a
qUEKX8Bj9x1vRSWxN6g3PIs3PfA7bH05It1Z9AFmHNSyupITBTAIouIBU+9hPdg9fYDrfQYobyN4
OYTKqxu9SCLBWnlgifbIphOTcsjW844kbBsn+HiBqePgvgHt8KOyw2gljhLOF+2AXV0eLdkaeDc7
+cFKu0b/rGUb91uUjkhbLJGi+VNHDF4nH9mqnSPEbANUl1tPUuB9CnOeV7ALxIAUnsh++p7RMe2y
0M9DOSq1hHcgbLkPq8d49OqIKmFnivZr6id6KGHQfvKWQhJBHFe0yIacw3cJZAGwQCm0Qv2FWjBC
D6dY2KSdd53hKaAu/OcZ+9xz9wbk28tUHlnQD/4SiSapIRDNcjEIr2Nwp6x9txbkswPfx/kwafTI
IOIlZ3dOBasvStoG/eVhEChd7S4o9Yhs5R93Crb56yTHmlnOpTN7kjBbzVnUl0cZKLQEMAzeoEC4
hpcI9p7YPyiEoKBnxFpYbcM9W/o4JMrYAbn166O0Xlida4Ropc+JTxi/K6gHNUTn9I/mY5epqYly
Mau6LyocgiDAfUiAFSVy3xSFBiPyP3k2ZX6R9hVAsdMntX/t42eeLzRGrhylK5e3Qrb/T0Nx6bj3
N8+5MmMa/gT6PoxSbVR3aOAJm+UP7KVR3uWRlRnM5U81HdxNhF2DwqeJEIOJ1HRdNsB/8lx131xk
gda/8vJw7aNEtnNue1GjVN9Yo8gODEbl6jnW3TxSdxofJECpkgV9/JVjlL2dhaQYcQ7jg6guf+aH
Z0O7lZLKQqN1Lu1poZ+2rtk/F0JUR61eGxhf/FYMY5z5ePcRs2Dc23CNU6bZ/pFadkothG8J4nO7
YHW27d9WpTGpzGQFDMNSw66dyXbrLoexKOHgy+5r3Tz0jGVBXY54UM2iY0qyTzEokNl40i5SEv5/
pvLNJDJsP/q4ZHdQ8Iw7PaNk4lW4EtRAHi82ZLbWI8cgBmCoSCe0q/VNG5wfnVDNTj/qyYfAwfuQ
rN1hvBAOwj4x4NHxw75mPRAP/xHs+FRp9RqZGrnGM6bGcedcpxs3os9NbYG/NypwZNMBBAHjOa1u
sFlZf7d+AR28NBEGSs7RmPoeLTJ2xbVNBsEq7QFt8OYf82W7rgygv3ElMFbTIDhT62WCmuvquL2z
dFQGN6yN2PvY3xxqBsdJrzvCvWxv2h+QXCPG/zjVsLUo7pr9KcQB/QyOO5qc0y++U55RGfBbcR6X
3ZuKGBCrhdkqtLH+71osQcQw0O48fT7SSqSLN6LiLBykKaSjU2S9cEg0dq3QrFtNGO5jfLxEebI5
MD8wVe9gJ1RBMfd0z6F5WuXUrVz4E4b+PJEckrYPVwCxi2tIQ7mCsIBHG3F0hkW6Fkp3usTvNV2+
PobNGnItNgtFyjhyZuTX5PTjzOyJITAujfJQW6rsiFDCrlL8+RyrZ9pqSThK/y8DXYnYJOpDH4Mp
fwRrxty+57smrzuByf+7hQpG78jDAZ3B5tJKapkoiXKgppWzF6SCHMoo4O//CBA0LDkEUwRPbnmp
SnBt7Nvbzb4/40RWTy19faudXttpYPLmvlPHSp/57X+3FTP8OW0c1r3B9BxtM/V5TRm34oFBnbA0
dDi+2POVFIWgbpssXQkVtowctEY/fdDLMLiPgNTguUgjA5vf+cCARz7Somgp/9gp8udna1QfHF3F
xUXDstui0QUCVqKsgLO47sv+CCndAiAmHT5O2hv05mGY7caAJ3Na7ZtqRKSgm72k3Lz4PTukWuAj
PCQyfsk4KMQkrCTucaHaQ75TahJ/47uhorXGXCkmFAnxOSm+D4vQryLxU21H66d3iqiET5EeTcf5
1z//Cvde6BDRcwGMs4MEAiqNk6Hn2+LrbRjGz3a0hVbAo052pSEHVxqLoqOOMRapvg1/tSViZfKP
cl0HQXPsbUkysalxuJbRc3jBNcxvV9F50Ni/gjdA79X1g0ShXp6vRgP5PXhBoA8Ng6cZ2slcw8ze
8ui2Ga+lcBJ+OUVgcp6+ASeQzLJmMwLREYCxb51rbl4PCARWoTKIocnPJKWuuRMdN80/gJN8/idP
g83v/T2vi99CnFPmUNgkB8jkMkFgMoMpvzXVZi0CcQQmFnlt51XlCMJXxztY3HE6+YgTQwrhyI2/
/Ar4ySu1M2+3aSeUQCllUUHoj4yP4qr1XKyeOGGKyANLb7ysXiG9Cw8hKyxt+2C/Q12FmBYM8b5A
FEV5CMaeU2dwy55RbqVUY+wmv2unU5I4CmPUviTiRN1Pw9g39MsUq8qU1Zl0scEM3Mom8gbEpzgf
XCcT/2GW5qwLOWph5bBte5RGwUyVsxvBmHATwhb7hS2nJcyDve2SXwIkGoNuK97aw/NRDxih1XAP
3Swj80EjZTo04uyYLfo8Ys9Dy4qrYoRYGusY8KqVDbBcZOZifMRBuuWqtv2rlz8AA9V9XIdG7pvY
m58U/68MLJPV7E2IgRhpJVE6Q6OJW4SQtcA/cd3xeWoCj2W/RTSELJufhQfNXbpwhgfQAgFCd6Y7
wxNMsackCZU4VJfkiHHCrD4zWmcDH19VXJjCaXZqtjOPn+YDSUstTLIxohbQp5p8uhX37fBQU/lb
dW357JpFj0ATeSB3JItP1WqcrSPpxd2Hk/g7v8LXI3jiDEDf64rUgQUhpUX9koaEX2CQ4aXVMFZC
JOfw3HW2iRnG79tpx1VcC9YG3yLNtsXdimPTDwB5H1PRpCyhWEUukxIA0tsxjIIgeBlMKAojhVb2
yLTyzBd6DnXuOjc4EYhupwJ1P6p+qQ+g/pS/aHvPu7z+HWudyHRbNi4ayROUoaIH8EqA3KaZn802
gGI4kYM5Vjg5smk1hnpq044WuPhVY/mOVNszega+nZTgKqKopzYqhaeUYHrJJWxR3O+G5BatfD7C
IxDDwEZlpMdIBRrdvq5kNGXSrQwc9cLNIXvvf7qHnQ+VlbiyFiCENCqfof467VQfR+xBZj2+mmtl
dGY/6ckKAV08RQ5+p8H/K+N8PIISwyQcCLTGxRlOdnqSOQCEyOivMwNAnl3ussFbe7PZ2oZfdcGW
ImlH+gKDLsRoVaX68UA86cFSYbIlo6phatjSC0tliWp0q0xZ7QljhplMXSvZ1JKydB3AloMB4ZYk
8it1tI/S0aWR/s7HN4oCs7aTOTewojGkOwnkmXJ9uwz3vqUmGQRZM7rFNqgkvkDlJUKcwkVMfvii
Cje292x6WbD+GfrhBZYSjCioKkd4kNEuvV0Dv+MswMqPJz1XgZ8V9rCtzla0MtGO0CfMnUC6LNT4
m3BUls3AMp5z+0Ks7WvFCvH6oeDGKLsTL2yVFKu8gO/2kUxi7Ph59v2eIr5qBdJtqIfeP2p4FBjr
/sQxHeykyZXafn9/nHiR+U6U7RJv5IhrcnVNpRghfksjM0Qz9FRcns+xDx0KVFoyVYAuINX7Vyjg
T0120UncCkqwJhv4k63vaRQ8HxNGbjv/PagVecte0X2PgaP4lEZUV3s35W9e/woeRXZZCqHRbUxr
FZgX5b/BbaGiivXh39+YMhP7wTrjlxLEO6NtifrwmVhqTSWLd/zM+qzVprdbJwCN81MsiOkRn8At
dMVWlwtQc1B+mirlfKxl4oFVGXyZIq2T+8Mn8XljXWoIAss8bP3umpYBp6cgEbKfrvzgo4VURe5W
LTmq8QF+Hnl+5uO2ZAv6rczdKoqtNn2jPB07CG+L8zUjRuXVeHRbLTT1UWoc/62RfZFlvvQi58yw
lxAHKesD2eYgE4JLRWvvcWMyk3G0fGjFvzejg1wEkDTSaDHEtQW7ZvqPaZDNBJR01/7tUrCtBmAe
c2WAGZGKOYaCqdKY2YA5FNIbY6qdxz0IqAGx2l+0YUlAmMnrOJwyXrQv2I85KBGMFWT4z9Lf8NPB
QpYvdOGmxIK2U5FFJNolS4Q2M3ydr8Gr5nN+KTZIdApeXTN3QoK8kAspdgUAtGr8GAdlhCy5ltlk
zOnwkvIcPmOst2qb/6yVE0FUEWAYXnT8u5orCF0URceoL7TedIpDQ7n264A76hR5OOOhEPRnmfgp
KEfNiUVEigITOWnfgk4oVZxac4ZCriqRaZNrRLEnm/ChjmlmhKXvHTG6gHLT4CJ4Sf5sazm/eDFu
D9bkjR3tJ09uXFXXRjHNW0Qz5qFluWli/7imAtLkIBZVVivVOQu9zOMCV8J+eQRmtENUtlGdm7A4
hxqWARALI9QrP2dfF9/8YPCM+q4qUzvidSv69Wuq/jCQ296pD7U4Y4yj6zazsI5k/HJsHWnXXESp
F/IY8xtGI9fIdPdP/Cusp54MgDLx3bQJ9/K9VWItEZIohQIxtiGu3hml+ulOW6mIAE643k7XeVPT
frxXJpZGfmP83w7V+zHISioXz4qbCJKihKSa5aditvWB+SNWOHgW1fMFH2fGE7iLALtvnui1RTWK
B8NayfPudl1PqYZ7gwp1O+F4t3ah1Era5No9bBFwFlZ5MyPuaKfihS7JdXNIbwjtqApEMfClmFx6
Za0GlVP5EZmz+dS8rGnemn3jkNY7YHZE7rRNROy9MN4FZt7qXrftOEBnUrvUKJteyB/7pcf3liZk
GLYwCYVQrCzMgXuk0ltJQxTjMyp6DhF6Uxr0KBWLhkX2UBzGS/gP122syqiek6pEriZfttzuANoF
rA43o+cjhEuSOZrJ6eLgdcF9EMaZjiiIJUSsQjgamKLRl+F/rcPFmsITmgC7PfzBBExgtZZsEuJ2
DxnzpBRRcd2Ig5BF+/43n7g5C8+JApEx4ZP8GgqS+yaDHKecKJMA1x6qYi1b4pqix4BKW5zJaGY/
WoRvthJOpam+UL+wJ35OG5O3oofG3rw3U4lVjPYBmq/B3ZTM+PaN25IcCSu4jf1RCCTz407bVzSu
grXvnNyNPGuXZ/NF2dOcRc7DQOIYA9GxqtyRh1K4x3H1m7gZUMfORDc50M0ZK/AQzoT4YAVg+jey
8E2vujwmVek1HQP0d54uEqmJhsNc2Wt6WYABwKF4rUjHSUkcy6YAvG1Lt+7MTshf4+V+uvbJDYto
79lWsTHV1k/rF1XEME3yzitOnLH4T0Tq6DnbVhzJrFlqgwh+VYcKXz4Ql6sArU/2IM7RaVk8cETP
D5F/beEN+uS4QCs+93Ns3QffoW+oHiEBdVsybILP2JmCUc+EQ7ULa3bNKMgp+TKcGbN8i+sPLIp1
RdHXt1ZWyUCCkW07I7URDWeXRgQfAOdVRhxASwHgKkS9Y2cqKo8QwrKSj9/JeylmAVlU+YO3DX8j
hm9WVpDf8uEqO8tXzXtSzFLGtc8c30P0W8IHglYPw/fOPND22ZxpTtlQjPoR47n/VmbyurhQ3HQh
9DJc42ssfkHJMEMFP6UDacWDwrO2nYBShcqHAdFH6aQ8CjA8DoxNQK13wvuPIxRPm7SftkCDsvCf
sC3neDgwwa7ikCIhlMjPdDZH6Z1EWJ03L6svKLMfk1hUhgZ4K668SprinsNru6Z66Ceyhg8pomzf
0+8jsPU7RghoIqZE8lrZyra2F/VMdOMd1FOgndPxcy6SNIEt3HWM06n/sz1CtxXMUZ69jq1yxx96
IaYhyI8nXkK5r9LK5292rKSP+uBL5Pd/IDF1on1lYeUYhSyAlOMhZbKYcQw68Xkt2ZH3XBQVpPlU
7xW5YeuXDPFKKxMKBKH5xJcVfIsdSYIFUkQOZBy2TMHaWDsTy0wLZk9KD0WzabFcb9h0pMRy4Rph
z9hZMlHxmLIXfPH1lBjfKcVv5l1ZIO7cl/LZl7HqpdX5LcCwfkcpEs1BaKqxIUnN4p4UcrqJS1l0
Sp6I4at28tWmMyXUql6FPay3TrKTkoD921BAfoLCbDidS7j7vUe7DWJ7nxxbv6rCS8L9W6Pc1So4
gEVBEMBrCBsS0dPcSkGZNdgwhhk+ce2+3LvN41f4wY99CdWJjMMMFnjYXYDRv57CAGPPfAhlouhh
lKwZDm83gDJS+D07skSe5YoeAx9juNl/2kfs7v+/P623XlLirq1WiOhdxAhk97UOFL1Vjg0LwEI/
0jVk8gy80Si5Oj1xjSdjXnZ2QSw+Xmr5+pI4+FQEfBBTgCuodCiNcK3R53LtQsafiJBFvcqt9xJV
exXF0ftAHOW5lCyos4T5n2pBmNlNKfb4LDcx/i9Cay+JDW0wsB7jmFP27HGsi8th5DfHBTlUNcpN
liW+yGDasB1qlBzTJMQN4HBThus+/+MP0Sl+Gpnz/YgQZwmzaNEh7qrU9I/9wsjs5YVOJboD9HPt
yby+1OnySgnlfmihm5RZmeAQYEiwqfVPdPqWs7m33GVD1BR1kfMzT+0cQFkS38IKByf93IDxph4/
zsyw5rdljJyWDwW1NudIsACgkj+sZdLFnp+W//bOBToQ0h/heyEFjRUsl7ion3kX5D9mQfmdeMBs
ZaD0G2VkohSdypBIAOomgMG6p5PVNjQMcJ/yQKgHF53fE3P0gMaPFT8CVSt4C5421uhz0CGvXnDo
ZeEEUY9mvLSiDk8RME//9trx6GFsIirWdofIL/a7VTeBeDbB71nOiBh9AoH9fAcbcQqFJnEtUTEV
GiplmBQLyKoakkgHFY0xX1nDOTVFeccHXV60Jka+YCaaikYL6++7FLcOnOiPh5h4iMWNIdX12hng
7Az1m5ceQ2rDAzZ2TGRVH1EsjTc2wWkjAtdcqXq67y+6DuHl2gfcT4A7bDpIIVSu9CjSKzlp/rpl
kPOXJv1tLPz5eZhBORxatNZoJwEG8JRs2dmyAFcKclpUUdIeLitBKk69amLmH141sxtIQDkfrtTQ
G4wG2+ylXjuNDrbv16lH534nngzsjcRh8qE10FGSD2fi7AyyzNYlEamKQVNT8HYiI1BP65DPz0Hn
bw/cKkVgnWNeKMVubY0aRB7Mh17rLbdx+Iw/4g34ozL6S77tkwZYE8Mfy0JT/x2dwPQ6zoHNJ4Fj
ITQ8gqUg2Dl5kO00+BEnAjx59vf0bvNYrUkJGlK+mXul6D+RrJIkmIcWL1M0RDGT7BBqbTe170i7
w2nYVTidFCP8hK/pZ1P7ZRAluodQrVUDecFecEGtjdhCpB3dYxjM5b/3Ko0aMygNBG68gaaHtKw+
EnZnmaycnF446jWqbyIbwCwuEU0h6YdItVw4r0bmm4TgRAZsDYtSUVyfNtoeXi20EW5Ohy+SDf0h
ekfB0vutA/tRkq5JncK4Wiw2CxmF4rK/j47LukEQpmhzHWC2gB2qtsWHGb7V5DhWCFHU5FYH7Lw2
lAzhFc8NXIhe9seL8bAbOaBxG8nFqAb1gR4fGy3N6R7RQXkcOMGae9IjaVawgx4KBjHufmvZs/mn
4FW9HPbW61rS3oSOTDGKIcgD+7sK8nxBukUpMKS4nxyR++OFNj0YU3YA+mVnImVtGKYSrkQuPK1C
xtsD7sodlIQJhfzrO6TlARbevFVF3iJNeczKhj92Tsyafm3PPhiEPVMx2zXTZzFbqp5aIjLVz3Ij
HHopOMEz4hwEYlEJ86SksR9pTC7rtX9XWv4yw/y65kBvdM7BIWbr/22RRaUJqUe1LyIrpIUhcejT
0LhpnTtTdOdIwSPqhAR/WOgHTDGr92g/NMUQuU4kDW9kk1t2XYmz3F0ER3QknYKXZpwKXJbxWjkU
+0P5h+uta1Ix38NKelGOYGdnK3Q4LxcC9DSEWdIWDPUVbCK4glGkvd8bRw2t6MYCmzaLy0K1p3co
ExxeoW5KKHm6PwgDy1BjUH9in0xnSxlQGZP07BZfuqKFArZH6lwXWbZcWg1icsvNKToa9/jY5zye
LAMMpFqARXjVcn3aMV6QwCST2pCawy2LBgV7Wxq044OCTliMBk5EN9rnafRgdJWodZUNNjffXkte
KO/iolWfaYaT3brigXYPx7clAxCJ3NNN8obS4YtgREk4xwOip1+OQNPsJ0MdKusWzt8eieNCas0K
ojDJcYz52vRpERZ9MMBhAgQvZpZ5mbmQXlSFp9rRam4cU1mnZ8BObmAzS842+zU4Hj64K8nYQM65
OJiR8q8xgpVcKNtIZ2zdt0I+C87lNCj3p99Mp5+9NN7LR3xL/si4W2Ub58nhfI1522L+xCWhz9+9
eCSh+wrIdd8lloQZQYDfYYF/iXmcVTXHuZwtPYgjzWvTDTzF+Hu4rD3Sv8BnM34zrw8AlFpktEtJ
BToWXqvruEKv3gJDb9uGYt/I/9dOFOq4Mz2CsHzjq/IhWU64gy7x441jGZg2NUsc6KondrI66DCv
j88/ZZay93bNEPdeRHt/JNLyDgZ+ZPtO49tgIuBbE08XR5yDE92+ixDZuoy8lrXKTZKPu/uTspK8
Pe9z7VNvrXZWiP+QFww5/F7c5/9M0IkmP5xlL9E5cSfwv6qqYE5UHIEkettc1/FVxVJDHBnmZvDu
Mb07pF9dwZq0zWpk0zTxV7CCKdRKI3Kg2jaqeSiUmWvqYlvqqINsm8iPFvUGruP5H56TTffsh8Qt
qAR6EZ4Vb2e1e18KNmpeQwZUVGm5dci32VUUcTnGHU53LgCZtw9fe3Hysv2MQqASCcFcln+0okkF
ZI+q4DhYdIYDgVcTn18YtX2sZBataOZWy3v1Uci9O50jrU4+dPYYUymH5XPdBTZU2W7O+t91Orwl
hJF/+KCCH2YlTWtPMnULK2PCYyOTLFhSvYZauorxBY5mHjRc7md3NVT/C035ZgUiBsIDx2w09Hu8
+yi+o3D4zUqvfCfNVvA8C6G5KjzO5OTtFtqGrEUO8yJ6erFmwZUJnQCRzbcejA02SuJaAs6r+bhQ
SI9RoXEIdG5VYICmttUv4AsCnyrsZa7YEFDmdtwT5ZpoSw2kEVKQ/ZYcGsDbe8jrrqiuckCuGqtJ
duNAwovC9WHyCU3nzPAApEWrF0hIlxvTqwoscdHoKJs4g5rYyHwRNYFSJBZuI+LLNktuGQ335BHC
0fe4+WeX1vNpaPSI8uMlhytzdT+/IcOGQkGJ2Mgmeo5o3XXCLAZ9UydsrDJeKRca75b0FPgVFUwY
fbM0aJ6uLvcXu1wzEx7MD3exe5iCwC73SX0B4c6QjcoYPWMe9GX1X/szaz6PIOtrjvBqlPDrP2b2
VNDH8FbBIyzZhve+LUdBkG9shfXo9HYYr2Rw8WgpW0g+5tpPO5qkYFpEEHRtVajgq9ypR2zPljl6
KCe1Y6dnmyEX5oONCmyXgm3qcL97mO4OibyC6UsRnnDBW7fuXLHB47UpNCTMNFcXtdQ/27HTZB72
7urWvZgt7uSQjRWGAan5wFuge9v5iCqO6rWdyGBDVGX20EnMG70G3SVOPQO9WL4zf3TKen2Huc9j
TNz0HP9f2hq4phJotW9B3pLvnPO0YnRP+K3jiUpsM3GujI7Tkf0Px4eYImxJJwwxHJgzfDrygm1c
Fdoh1nfcIXCttdI62I1le3lnnecJhOMsr1m24rFVUuPQzNqhTbT0gPMpgFmETPjpDcNCQMmfjbqS
afkxwSyZjkBuFOApubc/eLpo7d3lQy1bO7/NYdFr75BBNun4p/+afuYQATKPbre4E47GYji4669j
/Ifzrb+OofIwOewuJqULnEmuDOdvAhPPlgdlLL3EmstHvxoOS8Y3R95Ten0t3bPwXRkQe99bNrgZ
NFXTZ2LCCsOsdgWWfQQj4EXS72t4zWw421Ab/oWQXH3kc9VG1c7xoeduQeB+LX66Ej4ZPy3GBDEa
w6aYnRaBCed5ST6MWVBkSEd+7+yQCeXjnJc0sYZIrWEAh9raGoesQalQTclS9BeKf73ibtU2KBMB
F5//wpSXzVGU2si7Ebx78JLDzSiEsA2G+S3CTr/Ahap51DiicuxpqxAK64J05TyyXgG7pkDW4T/7
yolVJE50IXRj9u7bgZ1XMXc9Wy0WlIYI0ZQJ3JJN2DaA22A05fjGs9Pq5YPz25DzQtyx5Jo9xpJh
AloX3sEAgvZg5HjwgG5j6lXBi/16lghyp68JMV8BNwR6ZdUSy29+RRMcZnvO4K0Ftc1wSHT0doCb
9Q52d5WSIKgL54XNXBg5GfU2iGlWQ9c2K+9MzfRo0QUo9AXymVXTtLjz4NSIMIdveSIuv3MEYHfv
ra9QqknHq0REF+LNC9aPXGXkxcudqpTKr2H4MTCEHlgRr5c+9holZakQYrEduhbq1iVrOixxgcA7
OGDCYB0ag43stIiMkeEgqcYi3DxongzNF8d7WqP0awDYLxkTVn+3m6S3mwgLHYc6UxjeFWWuBU5k
SGHTW0vBcUqr8wJX9U9IcposHk/qVLbM43vq1/ughJL5Yt5kKHfZy8HG0ewsakp5CewYCncACmVi
R2wJsQqOZZOHbDEeZYPLwPlLPY31ayy6CJtWQae1cI99DQUniTmC9pyrOnprm6VhIdIeTpEiWZ9w
buhcZ/afTUr+hPS91J0UUzRRBHNnm0gt34awRJfjnaa8RY/2pOYD1RYOG+Zb0SSBGVuuzNCJrpix
qlXSrX+dVrQBjw2MTCyOsdsBnSWDEUlsQqPoAW7r06cC+HTLmEiVJOZwOB5UUMkYw9swL+rXqsy9
VHQBPxbGxJGe78QOrErDz5Ze2K6QBN8PSaXuC09o3pt7kslPgAxqYpZ/Lp+oire8mwKWaFw+J2w4
QJvoJSCW8SNrCDk9HSeDFZxpZ5LqGh9Ja4enfdwbCIVEuu6f8IBk757M6FvqScFOi8zvTMVr0XeR
hM0hxbuAg3lq+N5VdH9baC8mwcncixYawFDRZcQFq4U+/v4pORaufmZgYYF+t3eBdY3YOQ6B7XND
4kDhIqYwTAbnY2ugutTB5wn/QHOBFpLtHaZQwUjg9EM6mNZvmlKq+WnqcWXo2or1kZjpRk1z5Yz/
a4nsDzQ+Z1dqbwRw7UpDjQkB5Oo/Y4YDo5rx6gI3fTarD8JUaB7w1YYLLvydoYZDBJKfDJuD8vOr
oeccGWHXbeOg+q8HGWcWdx0BvJYe0LYzb61bQmR3cP4vj9HEV42eF+/QuIQgaWGDWZPpXb8lv6XY
Yz3Ju3juPDHCSFt6uW98go7vLk4dYniv9MZNXYYpjtqYcr2ru7he7TTb6CyMjfN8E53lj4/slrIu
Kv/fS5pAQjapWS7W//Pjf3kD6gRbm8DNv38O1/YoMRwmwKKjS2goQKR3FZi8V070913fDHXMAoF9
1SpjJILZVJGmF3R0RPl/RWGZeK6a7rfphUO0n/Kjtn8wpbWp3fQKnzKj3gOS5wPOs+yaOXBl6Lpd
ZVM+hPRz/78NKk3yoAYS6zFdaiojQITc7yimWbsPCTLaqskeh2URHL8Pu+KXswM/xJwcAWLFGCM+
/zdC4og/ytljwNifYQIoS1gcKgeesKTq79VoCKJyGDXyyXFSvA5gePOY8UbRt33zp8YlXoEBt6We
5950D+A8sQGu7v3jU/qSJeEic+eYuTrebSfPRyPtCXcZTYnab7HkP4lpTr2o6oLzG+hPucCPnU0M
5lAoS+fHByQ1cW3TJu4MoeS+XafwTmzvjkZB/GDtbwnYIZhHegaaICUrFkcSpuK2eiFN83lGFEHF
qVqS1o9wIo4NlmYM1BbwKaZwvOS5Z4ROKsukylAnphdl92syvMaX4UOpLdnCtnzdcVj/Z5OUtS5z
GINNUttKbi8JYQ9feZn6Ser78KJOWo2ZYs55tLxr2UYE8PMHMRISyWMmnINqhDIHwWpLBNjy5Ru3
x/VwiWXUdD/Ue3qvch/gGGD5I8GpNoSZGMvnU4gQIow029Qd8AhviG3GU3DLCawxO1G/r3ocFY0d
nT168ftkjn0FlYynKKu2EGcC10aM3XN6hgWBuFFgFM5Kx8lPaIHQhidKRuqZym3Pk/rq45b3XBh3
JoB0i07oJoN4Cgl2BTDx+SvjfX7xkNVSjhyEeE7lq2wX/7695Hx+KUcOGzG+XEhqJXrRA/CluvQD
bc+aJLPO4x12tjZsBUMvICco3u6LI+sC0TyKVY1ddPXm7CwHKG2hJAFsuMr3VtCfc9/Ad7qSMah0
aK7nz3ANB2Ryxy67xT1Gi58kv2CLlNZACnxKp85N+P79NXb6tpd/KOoVhr7HVqiEZX6CcSXltxFM
r9aiQXRS5laMtEkig0ZWRSxibMDllRbqJUEFejW9SrBjBrG9bw73bVPH/qgWgf8zZzbOMTBqjgk9
E5/ZQ0d16YZUNzDMvDo0Bhs+alsACCvLyNflNUvzgzwziayp/G6/4L++OCNTfpB9UWXkFI1+ABv1
JMj9IdgH7GdEGsCXp+Ff38WpnJ3onwHTrZzrhaZ+REoOpKHD8BHXMcc0vA6MlRhKvjjcTLfiCIeK
iivZPzhjlxv5YZDpXBj+gOBOZRmz2sH3H1h5ZSwGlxfNqUhQW97Qnz3MHUWVzB/DKm+ILtzv/Awy
WTQeWVI3AkVgK8z6mqI59XmiBWrG4KOtUB3rz1Eo1GDpyhKjJIsuVvYgugGs7r3uPvcaecxDE0Wi
yjNk8ItBwSQSVH/Bm1c1zwEjwMDiwUAS3eQl0nQwZ/GwM+xdpT3i2HslGOG9i92KZF/qkG510jdv
6Ed89zQOxGzysm1cxmdb9ULStBsXb0aWZ/tu4veJDRTVgQt4JFBllrcbYd1Uul/PBSpUA0A9asuM
Tc0wUGbTemBeWQuzEupPCqRPG/+eTP5w+xvP0BTPTipfcv8nF/5x9O+iJ1Jk+Yqq5aYe+DO6ld33
oKezJj0MG7oysK0Hu71jExdcAacTrQExP43+Q8jmw/9BjJyVe9azQ4N6dY23PSkxyNbZOFPq8D4m
WTIMsegLDAqw+ef1Xx1bD9ZDvYNV70WJHmhnrm1T8GMdWForR5ROaEEGkymFhZ4DUu8ZqijNXwO6
mqZY4gA3uamautq0l1uXxYZXP2jc6CNRXFwHB1vnagPLEjVY4z+ia8jeO8Iuebps8CQEc2vuxj6A
EkE9Lplk9aFUrGUEV6GJ31AwAVmHpRgbOPi9/HsoJUyqzUZz7Ms+m70TLJF63v8W9fJCmGOo5N4+
S5UdwzFbLx/ohszFVvg1UoBd1U6UidymOdQ/mQZ0LSDPrkdP4yDvN9+oayz2VdPgt7WiidUPiBRl
Ymfv6wcP9FcsBrGCLaAMdRJiF3K8kSFdom9QnoNm7OkYUSe0p3Cy6B1tRAHI7ixbW1cDMb6HCRYm
e9UrnuBkUc1aFQxwBPJLLMN27J1Hhcbh3y6LdzSnyDCU0a5nJNpGfjMMnIdq3JTMH7FmCUcgXoEE
/FB0glhmkACAwfUIL9Z4mHqLdAYuCsJeLm9xDLNgHYYJfIEUvjKceoSfRsBqMQNKjNHk3NZXBefZ
6+kWsCaYoH+Vybgx0hNJrseroZM7HWbuALNQhif40h6jndsYGx9qQTbzDFRe6F1jlTxbi7l8FYXB
e+DT4Y7AQaEgX0XH24W1zGOHee7K+wqRKU/lFtgW9GJIAIxStt4kt800V+3b/kGesvB4fWuG/2MV
fLcRXEzsy/R5B9hXQGow44NRVAE0m5O7PS6yItmymink8GPMa0dJM3r9Hlfqel9hx3J09GpqEjFM
JBLoFxx7NT6KglsC2cpxTBHCoFAG0sFV+YaH6F6bDifNbcrVYOtLStYX2wKMjZYCVwTSTyO9Ftw6
D3yHLQ+rz8RtQ//zt5AMjT2C6A5PSd88SYAvo40oECURWqa53vKNVJD2mpDYlC0PF64x2NSCKLXL
qVtpUooMttYjHEwP9W/cN/SC6kERnD58o7mG6saAs62jvK2VABWUWlEyQr6tDLHOFI041wguPw6I
BSvCBIKtQY4KOab9HhJYQWfxCQBxHTmpnLKCuCXozXYppP50AnHy2D/EDJfRRFu27qneKRacx5BP
uzvMtgnW+Kl/UI27Fzazw1W8oMFclXWzWXCJWuVN1+QP0I9dkT/p3qCz+gf+4o5rVX103OneUoCA
SzV7kAwj+8DezojEnMZ057/2IlP3TenGhumZSgtp2IWLrB/RdjnQpdUqyXqx+jHXCm/6o3bW5jOO
g7J06lxA/SRRK/5raJQuzFcoTJZTZj/CvlHVEnT9fY9U0wOlwUXidEKRyA2uargX5EWECZXDNEWP
cFKYybPPAm/CWZ9ek3gnjc5DEEcEyYtl6/hQi7BnLgAuhDx78q0+QYawSn9HXiz3L6ASuYcq20C0
Ji7z83T6SMkjphApAPcSDGKBdlXDJhf0Ua1bLp/RvWhcTbJ7V7HWDOVwDGjANhxTnfcqCknkKdlT
y9Fo1cdw6R2fXCjlN1Jk3k44ciz4LWLus5S0vOUgcUN9uo56L8cB3Q0xqP6SsKKQL+SpLttx4HwO
KiBvBRFT5KRze3ATLv2RtHQFCG7zONnfPuu9kB4aGNvYGU2p9WoX5vJVPxTu6tlDbj8VmeEZuxdN
19w40/Mkx5lvcim1PRE8emcsm2e2lpextJd9Q4P8UhSPBB5WFjCZN1pvuXiAkKvW4YGKXwvPrA0u
WRlHDhOzTTfbDCjwFZcp8AskseVaEL3ClzH8I6HWBCcKDfrqSrhybHAZH+Iq06dCgI0EpDYRaHOw
oAEoNykmC8y4yjJsrq9ZGZLjVP31WUE5I+MvYlVI9CL4Z6BGbWBz58kMoQBdXMBwS+2aiJNyZKMy
+JVwjvPHKBYOz08X4GdiXhEwod0orLNhMYwqKNDg1+kLOGANvUtsNNH7BlGHY/BT+Kpv/Typ5vKC
bal/9TNnsmJ5A0YFkNzQkYCxbCMVaDC+WTa/XRZpFSksWffjVZ4FiV8GgHCHExeZk5xK7QquH8sT
9WA8Lifv8m3UIMVP0cMkClW07/Y3MigqiqnQZDesso+bEJG1wjqxPhUmmrnK4YcRmPYUzrnTJRBx
v8/D7uArnUlhjdtW1ZD5N/J71jiosOpvKFVEJFUxCCiouHKxLhjsx41Zn7Hw+BXfin5sCtyWAe9c
/cxEr2b+EtS/mZLkWlXQtZsbbwmTmjRqOM5iRQy3Ddbphc5uMSOsjXs6bw/ko1kFUx9wJFzhz3Ba
IMKlhT2RORwEue7iA3M9jl00JUR5eX7enFQn6Au0DXN8wpGqsfrjBJVxwTbkwR8FNiDQKOSv/YYs
fgGy8Ig0bZOx+FS8XtB5PrsrDLpH1E9FlwS/gHAEyVMvNqrJBGTqATHHDyj0DPjhGy7tIpDxwo3B
/PP95alcDXzpi6dM1nKrkgSjqlcUw9esxXIBBR8ji+x7OlMBekovOJTWSewT/Pm9uBZp5f5NdaB7
4j2kGScipwcApcXKAc/wp3TzQVZnmF3kbrEXUR/vUClMFQ4Ilt1otIMdPdAQ05F9xE3Gkwx/hDd8
k5yFpVsEsIeTz1mnu1jzWnJdG0KJxL39YOnq0cQbmKdrCPlHAGEEq9ZAHcg8OWrpgtKEpe3aXpHe
HaQG+h5qTuBdUQ4h5ZVmCS6itXorUnKGxAtEtXLwCATzegJ2g79XEHgkb1d7yMk37MswV5xPJ6tv
Ct61B4khj/h2Tle8XgiamvZxIWULFntVggdwLKsovvMjcswaYSgzQrBK/vfKafAuFokdtn0qyXLK
Lh1YqJt4MctylfPmXfm0Nw3fsSx8Ogca5Ef9r9ZxNywlGDUqpClIwdYqt+rnIvQnv5DcKasCat1+
1OFpENasIUQBjFvgEFB29F1zcKhr89dTT8wwylg1qhl0Ot4aYGLXGIhwpLZw7Qv9V4cd3gma/MWc
SN8bhBFPnWvEyD5RXt0X3zJGr+rBgTzI/K1kf43NJIVNQAkve5AHhHikIxdRbGCdvP3WRD71usc/
R/+rQftTZmrnb4GCJDqwrY8Gf3nROhMYmOIP4Je84YL/vHtl6UO1qEwVF4+W35ANhz8jXJBZaXwM
9y6L7c+2u+XqwxrxMxSDvq3/eXGc8YQlyJqQSqOf9DrKrt5M8rsL6fhExh31FA5VxrCHaG503n03
p/+rTUnDmaJwwBSvA5uLso5Uf1Y0r/RxoYD9YM0zyFxztSttTIgwYm/ABAZeRHCk6EgI1BsxARe3
PqzWgi3UI37JwK5mmqrz9g/gjcqp2jj0ODFOav+953AskePR1xgWmr9KKXS2erMTW/Ogr+rAI1gZ
7kb4bw7/pou1ezK4+qxhFk2Y6g8LqYy+CLXaTCCfkqJPuBuLi4FCCtEhMx7uXYlmcQhJ4j85Zqz/
bz1jYVzxONPwanplCgLidXEkdAGtDwGVMH4L5MhKzmsvDRBicodwveZBDMbej/DmLwQXGHLz0+bq
wuWgAegiwtzpW+DrRCpMscJtiRHpIi0+sFayfNiHz64ynZVHifXyiQMzy6u+ETWN6/q2btT3OIG5
OJshKKWiFMI2NX2sNp523WE6+y7EOhviFDUTH/WNkdf/a0HyJ3F+4PWhFPM/IFIMGrOCUb7jarmJ
OVqLi0Rgv08O60buUrFLS+q4DJs8ft8jAqZFuh3JVTll3v6o1n4O0qX+drdKLLwAoL2c4OFN9l7E
7hPjMOO8ZRhRA57YmWzfRCVad9q7+NMHp7/0XsY0ZjETRYnECcviMaDBwNprtdPtCXHV9PNAReKu
CzhMhSZpSGgn15AdubhoseowmvouWZQThgKEn4OmQGlUc4JHHSzToRdQFOEjay4dGRwxWpR/LKZh
V9kwHLw6kotQelTE77ePTcob1r95wkCsuN2kPhA1iYRHp4Bmj62SGmm7CuF6i60vWz7L8eDa5JnH
fm3kIbOdYEkjOnwIy6NT1OkgDicHp4aLDyieAZVYeIpeSP/lNYp04fB0phFU2RErcN6pYkP6p/g/
7td7cshblSgn1ezi2KHTSeEU8lyrV8o9WdCtXvXgJKW15VatszV+JmQVGlnTT6AYAZ+sbTP+84lD
w33Laa9Oyj50RRc7H7UKloTOtO17Rrcs/hQ6Y94KJxeFwqsF98RdZ+uN6wKxi1si1eRUyesC13PO
OLwG2uCgf7U9tlIpmmL9BFerWU+5j9IKFtrLFiiolk4yPgZcj5F9HatfUMZ4NKCg4c42c04hCs8C
4zTWt12Z7YkaUNMcuEA6z5qgvx0rJTJRTAacf79Vyja10jHxx7mqXAFlDDeEPcfIUO50oii7YRm1
e3rnsDbVI1ISTzqy3vCMtf7RsX1kcOjEa+cczwRfaLmSDSj2YRSl/Vm+/Q+sQFUmFE49+cUzNMgk
L1SaJSXxFiAzsxIVK2sKmDLuElGxRoF8NNnDO5lnwoX47463Z+XVXB8U5clO0pY40S8Eo1FO/nHs
UUAE/vGT9LNkoRxtwX8mXYGhdgPWhFfCFyQMBjYUwI1XrryjZoWyDB5+tZOm0RwygceXjiOofea+
Qm6fCcmrRawy9WzPOOHrlW4wKjb9nzLHmBAzABiOz42lDl/N9JHpRTvla7/s1mJ3QUg3ZL0Yv3DI
ktyYjxqqq6r1teEaXNaQ5OkKfLjAtz4yoY3DeHzFTXQCMHJcIGmmMe1TYNw4NN7yu/tzAUQCr+xE
piGtv9U5TWCOkhKT8nArknvZ4Ly+YHsEDojsXxQwwwrz0ICurT5PHhaHBT6GOAgGQVLtV64+Q82u
186dn6a/1ZHx2aDAobKCOJBDKdw5wLcsx2Ba2AOnfEsowc2juBZcEOvqVwYVrR3jFTzJxcaomHKL
h/BzdJz4+dpc6hx7MqmBzpjqg9dEfoit+dvWW8Qydp3Axl08q66i1O6ZqWbXmZnY6+FQ7jgsQMrf
ZmDIhEgmVGY15cItslEh3V1WTx7Et8sVzzqZ6WpFOH7bjQEjBXLxNrMoivdhbyADnJGKSN1xDgHA
lAPeb1hO8hEKuMm3oo24eebv+TXJeWOzaJDQKk8yELJK4pHeTkLcHshEphyz8YG7XXxRfSfbvAmF
Aem5xLxV9rMzXnasxBeWghmVyCwV/lpQU8Con8x5vGDrkLdGbd4WMzSkIluv/2VWo5AlWu9pr85Q
sE445lkx2Odb4BQyJKTvyE8RLNADUTawGNS4CKgmf3lGUdqJk5rmAve1BeWZukAr97S2fqDOET1F
FvLhEpy3JByvxrr2GOScwk9l78at+q856ZorfTX5Z2Bzv5oYfFXN0/xbOGbuQX8B4JXi5D46tc/V
LS+zGitUVGbe61ojp9PeTM+/iseNgtb99tnvewlE4bYOKNWHJ4H53wohpYenrTVDXVaZb/R/ucs+
q18p7T8DGESD6vUV57fF9x81YzKeiCrQiJPohOnYi5Vo1MNegq0ga2BeSyKShM2zVIIx9PD6rSUz
RhE5/GEV9QeR0l5NaDqMA4gJ2N0Dbh69R+d8zC7v0ks4jWDHzJkjM2LYQEgPk9XfMguYd5Npxo3O
D1WfTDpJryLOH9wa3huRd2mCAXjHzZV1RMAhBJwWYBxJnDyDIJmz7JYdKs+Ns+eLw6rM6/3cDZjs
hnLB/yJA6DnUmGnFQwa0BugO4HStAjDwBOY7Nxu3o/uUzVIHBe5iRj4wDE7RS40pFoEo5lGV1aO2
It/pdnaDs6xD7fc0LNvkgq2PIsKV9LYahzhAUnLZTMaJC3/UkGVOeCTPlWvyx6FKdga3PAX0O/EC
uGqvyn8cAT3mFuoIS/fnrzBZnPhafbg4DlawRfRNyGLkjpq7EvpHlHSlNfbeeESjPf/cOgRgLFt0
5XIfhJPg3l8rae42UfQjKVhtCOszfd+edW8Rl84+aIR1M5tRQb4BPadV540Wr6WlWFiRaf24wlFa
Nw4/0UE6jiF1sWAxGBzIWltBNKPgGnyg9bNgT0mONi+rcP1OVHLD7LUadSDW33PXO6SadtMPr0Ev
q0zyrTzIcat4YWh3qmPVHEd4S+BpFiwsjAA7W9XGUuMDD9dUAsZL1B24WeMWMM+gNtLudhjr17Hx
/hEcAsKr8hFVO6olhSBg432wQIsKTMomcQTpAYL2RJozesh9U+lnzN8hKgI0wvOddN/05j1Aq32Q
+HFWeoNevPZZTZ4lHLfOi8BOsJLxevhafLbtP2jaStMI87Du/9xkaRPA9WqWopacaRnExw3UAN1l
FGFgX0kd/uYDauZ9yK4K06YblwiZ3n5b0aR3sXizF2/naxB+LHqOm61jNFalyNo/gmQEqQQCkKs7
Mxs5VA5pOcGdah5q4llROpBcfUH46hJ1Ua88g4FWdCVSE1BZAOdquaqzw4tUNOIRHnLet1L5QAcq
kle28cneRt2hbPbfZsigcH5Egnqw6hKWHyf5+LvpZrTxV+bty9RBHgY9ZzdqY+4hUOE4mZgDClA9
OQz+8iUYITVj+UscSmChy4Aj2fXXTesaNOTYCtgR7QS52NaoHfUzf/l35AtIp3QlXdDZIboDE1z+
r9ROBIjUba4S65caUtqkwWmwRyCfrGfwsR/N9JkYvvSEy0Iu9p5nuqvQzatouGFScg7+H+6OrDLl
DXvaxRRE/pMRk9oCA7lav0ulRZlFI3vkFWeM1Oy3cT9xfiWlgpYgzpm8XT6XmwMDJyub+EvjWiEc
EgHvStTJa6MH/+jeZruOi2bygDzEcdmDvZaAn5z3v9X0PoHscvudBWPa5Na5G/oSs/5C8PovkSeE
qHHv1y5zdnK44t0A9MMYpJguIQEpz6pXZyKjZ6/47Pr0qAp24QiP1LxmaRCLP30oitg7FHb72Bhq
hKR6GkWCklrAuaFGyf2UaKnXCrgO3VIxpC1Ir4dLHwd3cGZSdrSTO5rGRvpdVm+Go/PsFe6TVHrA
PbKWYKk6B9M3n4CxCNDaS9aRuFwr1CQxvvNrYTLpPoKtymwjpJ6m81BWQ4S7fvaGXdgyC5/8QzsD
iL9g7ZO3EE/THthrG470D4Ea3Eq7msPmGIAk666qRuYsW3ooEzJhKWTDhvWQcWKZQD5HTP1mPyD1
BoNtWlPuH8voa1HwxIHdu2+hQFgE53bUlZ0uswfZ18QPlj2igjoWxpT70U09KYXm7j5b16WqAlpY
l/I6MUcSSMLSdiDWJ88Hs6nRBkm86+bfqtEmcvRw3xmesrlmjiKItmSEbY3hyJglUCZr/m0wuDKP
1iB18QceunasRSWSnmM6QdV9omcQ+FUsX16RBzIT95RhZpcnUX5Qr891FHXfDzS42fy2hsERWvmB
fQRAxoNMRa2UCHLap2jn5n0vU5eYXsLBYy814WnjfGSKgzNDOxjPTZkUebGBoSj8YeBdoRF12dbP
/8qFEgj6JypRYkcJLFjbPkhUqoTKqkkBL8H4Ff8OXO4B6l6TixPtivIvVHMCjWOGjD1k3SWnmmQz
577k5EhQb/aU1lgLRMLMGglV2NiUUyUm2MKHrrb380H13uAUlJt+tkphvdu+f378F90Jq/lybvOb
3eO1sOio2jPj8ptcsqZqgFZYVeolzzPKJtsZcI9bAphTzJhwR0w6vsmUX5LDBqwDcwAafRWaTFk3
YvUubd9UPfnMSJ8/qeaMRhDGtD6eQWLiz8IbLLw59gEr0A6DIqXOqqBb6VeaNJqZXt80UtistHHR
1eEL5br6nQeXPl9QaP81FSIRSx6ehJf1uMJHSJr+EWoeMQS4jXShgaEMnfz1c/JDgHQxUnmbD6Ua
iJax281Kyvuw98shE3PwzitimhBmnfTCm/QvnBpb1ElPpqQ8DNynoLbx3IRdCiVppfVjKRNvQED7
N9v2TdZwkIdoAkm47fAzcqGrGgEY3V4vs7x2vCajaQqyOBPb5ZRH80gJy56MYTDGSjo4qRv0VIqP
8TNbxZxnavgQ7QYqJkNa4ASqlKvj4DwRsYS5t4lnPxyjfzvWV1Cnfra6kqFbS4w0Zd5tDdgb4BAu
+Mv6M863u/FuLjmZPYe9+gMBX3VopDb0RlCvRiOhoTYBoAkuQUJY2SdRcDwifrZK7HH0tCysAjtT
oUor1+H+tWtMHgGDPFv8blsHRTRL0fyb8OgT0zjSKTGnw3hhDZcW4YKO6nwc3W6Xy4hpzCn4Zev+
moTw2IVLe4epUZdslaqA1jTejK3nV/jgzEg7uiZ/zZ5CndH936drv3o18qg1b8kxCTk3w5hjlV2Y
WU7Z5HPyy5/L6BvImujjF9JF3ATlt9cublk+VaQh6ySKESc4JBq6MfxoMAi6Q0MUrzXWzILobcRB
4O9t2IqYt4G1SlHXDbLQNT67ItA4pYuCm5ftTvYou76+SeoqBIXvzrxU7i1+jXYtATm0AAHr60Gd
kiqF5tSd8i25h5htf/qVt5+ekdOYVaxLmgWud46qlzYiNGNIwyZxL0mL5UyLLgvCiVMTVpXpmaDX
4Ps08cB4G//PV1xcmqh/OknAz3ALnH/2mEWYew3XObJkY3aRqwcTO9XgY0IRgigUjJRV62r8hUUi
prDs15e22yR6OOWKFosP+P0fxcvKNZxG8gab/4AbbX/AwV7hbNPGxopTrPmjnO5g4m8pRKM9g0X9
4u0ML5WbWkmrmnuQMTWH9Jm7/NI76p6PMzUmhm7pj3D9y9LnBtt6n3NG0UeHe5jQ+tqgb3+8eBRv
WbCrkAlr61+PCRkCalk6aarwuPX5HldGrtxig8EtFRi2c758KxED27cP3xCWuJMFnzQqFvQ85sgi
IOzLEUEhdupUZzrUMbBwvwzpNaRK+IbtT7qF0FF5S2WSsxyqCG+AiZaCKEaMjvyTDsXa1K3iAZTw
zN6Sc+IBKbTSArCNSsXW/cpuC5XqIPmxGmnJbnd1pagW38omCgZMQos854s0dlnTRqjOPHGCYEes
qa4tXyCxmca6ElgX/AkN8oUbFazrMxM9c+NwXiCKkAsgX4AGKmzZNq5pFWghNtmF2c9FIfHnvW7N
FX+Py2aYzU9o2Qwyp96GqufQJOdIwU9imYCTXYYdGZjHDl2CQCGuTkMoEJwC/9lUpttKiMtCZ1as
sq0wCFZblrp5zPLp56tt5cPqzMOM/q65KD5QlLHrKuGZnJfUu9lscYmOfGnp7C20iqnl5ACaXMCN
Ivo0mQXbiEb30ZuXFF4ESY+AtxvSNLP08u/OdSE9hxJozaWjIUgqiCUgw09/xkIrTLaThlK3C+l4
ZPmPngu/xO3cf//33Wf+8+w8uH2zBcHHZYrWpj1Yr7L59m7P45sGhRW3Hy+rYyYsOq3PRa0EBXe4
c5tAmjICd0BcwlPMeuws8tH6eExWEoq+g9ALuMwDjYZbVgHFyAcKq+331ogouKVieJ5y2oYwoS13
/4bcAfp+4RB3H5oLjetF4VSFjqRD53B5sqklzhRk7UIDlhiejQIo8+qKC8d/0wBG4X68o+uHVUcZ
uoemrx7n7Yb5duc3BE2vQi8WveJCgWrwT5Qb4ZDFxqUcYqvSeAMAcgg75FfwUV/DJjmz+onH/2jk
FhqEau09WNtEw6PbZXoW+YleA/nKhW5eq0WqgoMAVMoyxdqSxd0QJ5lDiWQaj1arkvmEQ2DS5yf9
fyoPs/mJL0eOWLCQbjEJPaWZ4AbXwmuGLdz4NOPUrxLE1wk35f5j1/GY55NZHFpkvTYDgXg6HdYV
7iZvVNSBdBmyTkTErBMXWHgGT1gfojO894XTRPgSP/dqac6N1y+xZXoB1ItMyt04koqKUpUScbaU
dVCmMBilDtv587cPHfAi0F/LW+D8C7O/zGWxaRfnRB4TXYnAfJVXDQrqku32BtZOjRFwIkqUcOXT
Tjvt02gtk8NzvRzMn0ReD9FK/1BI+1AKqmgLQswz/7rRVYReO44pFwArhY7n2UQDj161CGOBFGW9
PgQ68MttxIvLAZA0Q/vCV+cSTWGsdh1/ZUwW4vD+ejt5X5BPWyHJyYn3Ce5ZqvqCMAxUZ40zrW5S
xkdf+gQBt4cuixq3Zl5lU2/wmXS5ei5JlAdLUFZmtkluoK0/MC04zIPqs8qPlWTrtxHHnTh0fvq/
s1KKBnQBYTvFOPm1GRZpRxs1Vf/uZh/PLNRO5V5gR3Cr/dmSM49RiBUNXhdF268k9K4Nc02RlRH7
jtXXZBWHTmciwa1t/2EJG5akyf3CqPCW6f5WoDmWJk+n1UX1ok4ZgpqA1RkCgX8apWyZ/W6cNXoh
nv5pisjhme1TPRsWQ8ALJmRJBPdj/FtgPZklq7S0AwuXDmux6pYRvbQuNgsj3dLMLlV0WAXxaR7x
dDs7ZJkn3p0uyX8OgHrsg5YyUe9FzPlQuxymavUc8J7gqJLBkeV4Bij2RXlnJCh7mFTdbSZQxwHU
jvfOSZr64Uh5gJi6dgipK9uSpKM41Yhkesyoyfuf9JthvH5LaOyZKIGF+2d7C48Itx6NkytFxGEa
GeVVWiBTfQ265RS7tLSl1N6jE6o3fzv9DjoCePpMMG/XyVuIvWPtJozdzl9VJDJLEYDlxJFoKYdC
8PMwfGAC+hwKNywtQpfr28dMfMNguHI9V9py70YMA0QtI9P7QxfxH5uns/NfI7nNNma/BdbkUfL+
qEKyR9ndFutPKlqh3bROCSjEd4g79RbaftgJbpoWqyVV4CtCHlOnpH0OXftQ8+pox8YYXac/O7SX
2ta42fZNIYNwb5D8jUFlq6/cIABcGrSfCuzIykG9d/IHV9Mg8v5Klywz8xozJItXjcu6YksaxU18
6hbNUejrwC5+faYIt2YH+MAhhVHIArWkxzac7s2UqUJ4s2ZufhCf8jsDRBM3gQRFlqRUqxYMLpEK
CB4mJsjUwLaHiRCAQl0WjK+5kn3PTb+vEbr1HoGwnJaqUY9gEh9qKVT2euQBMk/tdq3aS46f+JpO
6XvSjhXNmYXQ/DJkEnh1cRnFdja3MmxuSu1cCyV4lhQbo5y5Jw6Qrju4PJwbktlOZt2NWf6Paw7o
XTWkPcthbN2BszCzPS0WodbwUK2rH4NmjPDByGuoOJlmCBMEsGXF+J4ma32+M5SYiUbPHTUJp/a8
UaEsVts0NgduYN+qhVtEWuNhHI6SUNJX1MkW/PTKZeeFPDNvd6fCHxiBXrR9r6T/XBmzE7BNpta2
iYscA93rIfzCZtSr85fxmDPOboVMmMsJcg3GSPIXFlxftsghRcqJv/Kc+37R2YMfXI9t4Mn16wjS
KXgurVwUBGYxJ9MsynAenNJ3iTZYaCggIO+ldo6VAOvrpfhlsCPoTaAKmmJp0HeiOrg8tuJRxZxA
elOoNH706eHM24jJu7uGE289+NkpC5IDkVaUbZUSXxlm+2uZjEGN4jU4koXINLXxXDT0I/tVatk0
mtFDvN92odB27yYXhM9Y7C4B8znHCdVZw4Ys1Ft/ZKJ5SfOUSvurN71pQ2p4jsTwGHcE1s4/Y03E
aKIfrzRaYbtHseg571EwS+5RvuKuDzJRXVpmkBBvnuwoMSo2EXsXQnseqHLzg6wlj2S1EKO/XKTY
cvfdd1pSzQyDB8XTWomN5Z0HQn27+krKaqLoxrck1wLVkA/QO1Ogx9HSSeumKwejAYSbhwRiLD3E
UHaoG+ce8zkbADaCG1wQJbbJh1EZllY119/AOSmVawZo3F2fN9doDfCQ0UPngX9LfDHU80uTahFK
PyGVODAaeZYo6cbVEhlsyRtoTJOLd1d6BPgkJecwfmg3w02a2w2YjW5LO3SYrLzES4LyIEPzC1Ax
NGgj7GdQ15Tt9TpOaL69PtEIPEnEgQEtljsLigqe5o8dL0g52gVXM1OwLNcAWfb9hTl5PrOia2p4
mAQOydKORF8+rLYVCzoL4WLC+24FfAxs13SzyiZo8c7jBdmX1xGBUpN8crmWLQra6Q2CvKQ4Co01
p/hXGx0pEexnIMp37/lBy+n09DwRPa5aJX6R4wNoIFOqSLISWR76Q+kyWjeMooWqx7mwIIIwNoHA
PrArWS5LTjuSEd6OsEjgG3EDbrWi+EkWItQGALmwW+u5OirFDQ5s7dmi6IvU7Oye1tGVmacxWBRK
5cUSUV9znsGBw+yxqfFAcGjntl2mcIhyiPNbkoXp2hvqnT3Hgro+ZsOBQRpdSegwE47KimsiReZc
qZWLIslMAv7zdfo9qjWcTOfXo7PSHLT5uTyR/zY5XFp0cYedB3XrgWM5wwGVQbzUWm1fOLYuOF7L
E9LIBdhOPg42FdrygVMA+gluWObs7IdbRJAYDGpJ2aDpVW5kkdox27vwnw6TibFSVZCcipwDJ2E+
rGxbWVxEMeCP+nlCP0z+noVKE9/lC+iH6KmgVh0RwWzciaJdT6RQcwhAyc9rtBCDgnWkAAh4diGg
8VTt2VuP1d4sFbeRQWXXCa5Mrv+tqEe4m6L4c6zDeQxLVj7X1nrNioGNkjwQD7v/iunTu1V23YaZ
2qdoBTMuEshe1i1yxvP8427Si/+Vc4Sl6YT0ifL9Nn63EVy2yu0WzEhIIt2DApfCdKGMgpAKMIFQ
+5hmRDUttrpY7l2EUyLw5WhWd/S+X7xGWDBXoEKvqUaR+lfV6q4GIX3fAUeuHKDIDpWA108zubwo
P8/AvQVm4rJoQ5SW+m0uR57tzSTrIDC2KGdajnvF1efiXZT9hxQhRKWbOnFRUF2gAR39C+qROe93
YNj6btYHv5mtEfnygvaxzw/nieHvGm6scvOLWu2Tf/9sHTJxXlZq2Kv9Tl/9CsGLOdN+NxCxtU33
UYb1t3sA9F0keszCfBqX8pWKDQUV5tF9hFYd47cXvm8JcEFb5T6gYIbSymPI/0h9kjiP5JfVW1ip
mUO6fGPYDU277DQ1Sb365bv2yhZ8nPL/mOkbYIP1NtIiQe9U9XoBqE+8bnFodfy7JDNarbOqeKSp
5dXu4Uihsk5CS0msmA9xQqyoA3GuSrl+i+NWK1LYJ50jXlgp4E1+PmCwUfM98bTpZl/CovQMevIH
VXNbhAWVf++Rkcp5StcU2bZ9GMcBLC7xY+rtz1PMAS5Typp4KscNtsM6wtV1DZuUazNrHLEvI5OP
dQTQWvCZ9JvbGVTyrEhea9lD8ITASMAr0r5USGGo0UXc/kxwND6liwE47/dodkd6+slQhe/krEF5
vCn1ADk+s6HsvKzC5d668cEfR/9BuPGNbMekSR5hNx38O4QXE5UhJfXYTcYzcDiJafFXaDm9375o
834aB9un5plNJU/Zph+bN/YdaVRCSQRFR19g6ER1XVelPC+lTJP+uU0WUrKtgPUbbZKP8+dG6q+T
oZqqz2Sr9z5bQioonmtEWDydd2z+9wyOmTEVLIFLAIi+ZoWHdqh2JQ1sdy3LpU9rGEXliZf0ghtS
akDUfxnI4o9Pi86oA6pw20Ar+NKmMpnTcx+OybVj5yLRW4OuC8kzMrqyN3cnAmlxNkJckV/IlJE8
7e6Aqjb7EHYVttjeqpVPYMrhX9MMjLLoq1km9cgC3zZdCWbQbFpqQUnPd2V2YTTOyjO8PAuFGWR6
4BuwiJJO+TiA7cK/evzM8h8J8AAorY0AWtR2Rqkx14Ya2ehhG66bhAoID2URvbUZ36/yayiajoo1
nUXebBpEWRIzFaIR4/QX0vUZC/GC9ZKyjDRL/M1lltys1HCkqR8DYGqfrIlRwXreOEXboPaJfDQU
D2NYBccWMW0OuEqyD4xvbmr9CDUVRKnw1vwewjy/1MLZxbWFMXUIHpz/zc6wRonlKERQ0xtUECI3
kSr+LYxRGr9fphbBPbfa9rWOzyYztWP4cPVV6dGGW+SgeE1uugVN0RpFNT1O+CnP8R2h/SrWTYQ+
t9kgW12tcGb3dN6SzeExe0AOf2qqYo+Mp+Qn+MyeMD52eLIo7g+JMgedCt5x3XTcbe/FPRiViTv5
0dWElvu653/Uz0E//zQKfQBGH2N8hpb3eHkZZ9+LkEY8jXD4cJD51tuEgyOuf/nYxLdA9F3VJM8h
Y89KdqUOxdSd2006itF8sxkSEiWfxsxc7ui9v+uiYXCa4uPgIENECGWwBZTdzn/0ov8VsSDaxF0V
ecUUXRG2kjJynNn89d1PgNuPMkn0Hcwa7iM6r/HVHMpGR4oxFMiSLdrUOGnbrBFq+zPjztWsC4lb
g8jmcbP90iOSalMiHK5mbQwvYQCxcxffMmWKNPsJJUeXALRU4jpxilhOQ876TLTLIemqQ5ZCIBlw
RVE2NMqiduHCBBOG++Dj1tX9mCw1SQ+oE+Q+V8LNTyi6Ob6CQ4ccuwupKHV5uE1vjW9E/QzF5FgP
PeyExAE/2kJuJTz5BKw/3sS9EiBF98DUe08loNtU9+dcIQyx+64BR2etEJvpUR5VK3WT1WhGpEkC
X2NKoGjS4WJE9MHg8tnBpgazmaGiZjYIQVsALnMaJZvQR0zZBMMP10QQh+GwqONxWqZ8jynhF4UF
TwbULSiweIRgf2bpoitbi/q4TNY3zYVe7/mD4tqmjMtvK53XShIi7kQAvBok8EzXWz0hIvajK/jy
6H12EGwWATFtqoP86fpqqiAiTNmPURpjD2vXdQNO2wiu6mll8ZHfbG7Tm93JUyJBow1YdFlAzUcJ
HbgoV+hrDrqm5RQqLbm9Tjn2pKm0s6GbkEhsmeWvnj59LRVI5RsUFyS2BL0mPmwDAuaeDTkTtTeI
jN/klBXyxdDZDKZRmPaCPjLAspebOzGjUYoNE+WXdnoy75aune20TiOHHzkYWcfOATh04Anlt2+G
SCkbZU8RWYzENctHvkupOZvzp22kQFxrrTr9MNTo/z2RtKAuKkUYAsgsoxxMdGEFQQB58AbP5DoA
AMm/HZvWwL/bwIjgI2Qd554roCJi41o1XPdPjaF+Id/32ZF0Y7KOCWbyB8h9KLuEgVJPYwCtxpbA
Cl0+iioHyo3vsRlcY/hsg4E/URodtHaNood2WCOs20TEtAAHI5GlrAgtfdnoQaOTmUW0696ySTbC
wz9gNA5yau46dtjofqweXzZC+7yTZmvZMkmjDnB/VShNMyON7glse1jo/3pK8GQJx66maT+ffw/k
OmKsBlPNXyG4GJW9rEcxEl3ga21JBOrN+s8uKQF2j/34aKSC8nzND6lS+ZoeVUBoz95Ff4oH6qlK
nODERLTR5S7AI7UJQM8HCoR+zUxk3YaZNqdnPChIZMf8xP3nTDaVmo+kO9xJWacKNOw87hSfpuvc
CMpe6rgYdjwwzLS9t7tScY5dMCWDjBeJIzEtEwSbaKm19q58kOComOBqQyjtZwxfjljzYA/t6iWF
o3Rf6VmkJDK4kA9uVn9v8rIms3eD1MD3m846/T339RIgUqEu2sIYZFH2mKMwffJWN7kPWx8ewOTe
lfV0DOwblAyO5s2bULCH4l1Gahfk3BFOqOTYUgiErKAp73c7IgbEQbcpxSBXYLWLh6iBjSxAxUrO
FIYPGcxuk6gLumgX5PkQmNFnVxXGJmuFJuanaKOGi5lAPnY5vofT/yodMe/yNBo7zchiBUxll1QI
PgfSo9XIUPm8a59OvCJA69x3COqtTl8QAiiqR5xdyHLUorT2UnmOlafh6RCcX/1bvVr51AQywcGA
O2TxZF0tLgMpeOyp2MZl8DqbQqZeoquptggKQ68cPI1i6bGdR/yK/DFdjdNQ2glsiucVzOht60tJ
rrQJ1U59fzkeDJfP9kqq/+3zsUypBvSqhzSWWpn8gR3M11wop9DcUh2Hh68fr++yP5tf9fKE7xE/
lw87YAb3GmSRvLIJkf8nyWPxAkhaILElmTf+NWcZD6r1GbXtehXI+mOD35+ulcykTZbmt+QCIdjb
0/oJcglKRO10RKyk1U+OHrUstm/IgoG74abRvYCW8qHy89XyI12qgVssZVLG0icIU2A/B4mivDp7
c+zab/RYy0pNvIihycFCSXUOWlqFIkmfpEspFwPyFI2bA1ArBVfmgpvQnEed4FB5QcOa1+TP1kjz
05BqcsRZASPPBBV9WIvev7hJ4g8okyXTqXuOfO39gj/db0Lg5aPsHum/H1YMW83wtS5LRnuleCqd
hK8vUojYjN8fIw4XZSsYOCwHj9xr6G+aJwOS2nKQ+0/VTkpJ+qGgc7wk2FTKHSld/2756moRmqaE
gkQINJVyywSFEus85AoBXzB0rdIwyYMOAC779cOsNI3/eosnQnKI53iunbnB6mRx6PTmeyStzEEX
F5qljEIP9fulTpy533ZHkG+s/IvgjTmhIQRgcnLxBElViVDk/Hj4TC/xcpqHh2uy41s+gy08kn4t
YzVCFW+r+mIADzLaEvxLI7wwvGKpKGh6rk/d6Y596XqXEqwv/ylsmWiTGVVNVz5VkI3wRM67lR3C
qA/ip62gSorkI2xXMNQ2jVQ+0qmS8gYp2ESOuYSQjvbE85NuA3om2G20xJi8AS8buiomC92ochi5
LxmF59n+cfPEOd4rV3oDqZYVhE9Q610JBrNBCjfwlwPOwhPLWpUZuPI88RUSuQtzhXQERPW4qh0i
GAzDyO8AND/ozNsh9+Rjmwhy67NFzXDq0OdjX2UcvT67If1LFbPZ3scjV5mm5ORLaIVuhREW00g2
AD3Db9Qx6ZSWMoooEgdly98LejgD6Oh9Rdw8x5isIbPjVHiElDUKCpXP98FTJ69CKgp5QJmqHDI1
1pLMi49b6gVfmofe7C6yZm2YRHE5eU8OcoJa1/lGAfAO8dmXpROtpZsrY6DpHViDq4UsInv/zUqY
X7PkSHo62CfLyR4P66r9Xq+jsLd4EcJBRghL/QENmoKhbFvORQtKVRLjwzWCYol6/4fg+4d2LWUG
4p1BuvAlZ8xUaM8NXKCCn2y0AANZXBrMldRIr/1RizutQF8TSFIB6n5f2gvyvLVkOW14D5DuJ5iS
cNZZilZB4iZfrGW7xM9BZJV5qu6sqvzSG42s0wmU92/RvmCFu99oy+nvwqgImY8gcyhVu9krf0hp
3fO1oxazerylzOQLneRl1lglU3uI+odoYTnznW1bI2qJQFO+c/OtNaMc9S0dzLFMHYQLja37UYVJ
Yx96IxPGxAYsChauQTklsuqmxI+/BGWN9JNPYLspITU9/sHf+d77+nv47Yy77urkGO5fp896ClMr
NTbDOnIJAtyxSFF8/fudnX9loQvgsZkjJ8VD1UG8yOxyDdApEjQrSHhiMLmHJgEHyDIK8Huiog4F
AjF8QLK+uBAM3t6F4WVfsyNIR1Tg0DJUeGGtkv/s4VXGqmACMOJUuuOW1z8oRdq3PiIwmS4cZLiE
BakRRsz2Z9tbU3vR2/C5/IZTWH18KBpCZVaJKFytO8gn4x8roTDs0ueFt4u85A3RGKK98gUMAJzr
cwWF8bqemEH0uXrkL+jaH4XvenLnQPsinpgDumW7v5+Ni+Hc5TEKiDvJVUE0E/QBYN0T4pMYLsEf
3dEPgkRR+7Ior5HEhc7ixDf3xNiUNpl+V/bXFUcLVSHesg3VRTcIccWRHqQqpRcQ0L+mGZK7Ua2q
8QObMaceNdd2PsZIKr8ryuY+xCZexxZxvDxZbJPLXrAgz04y0aYqrie0J2+9Vj3K8BLSnEWoc1Z5
DGf+CkcCj34fKIQJjV6+8kymTgIt5jNBPKnJQqlWEIPoZ4AnjBD0i0IjYmlHZnyxA6vVa6JORqO3
C3RQFTAqQaj7lckT8M+gcn9Chq/YqaF+dyy+KCnDDOLX330rCsL8zM5ybYjZQqgVTK3BWf3X0gxr
F0NzqdfBqcWVgad1sLcSiDo+Ac4W/ytXEhpwj4eqpKXaY0wN51KRqdQDIPvhFzieB2FzkTxU2kK4
79/6xqg7LBI1oqYLFh/H3pCKv7jUCsifT+noGOqQDGnRh92bWfrE3LqLgeJGB8/e4yro2ipZt6eP
vuGkrGswH16efl/oddpDIeWNGc6MQnHa8k7Dk+ot69Sc9KknY8UYaBActMqGj2xuXxml1NMNjLI4
jdhDTw4wlTwFhCUnP9tQ31/wUxaWUu6dJ7aovR5OYniv/CTZYDppCHS/94Xeo3cZRspFMzq/QEPH
aQuTtvqAKnZ5jX1+ufjeqSNLhGBmtoYSawzvs2Gem63YpHuB8xmXaNlJ7u/eolumCA7koIRIpP68
eefksAi3TQ6Eiiln1VZByTxoeWhTZ2Nx1FFb9AYOpR6DJa0a+1A3cEPUJNWKSP8iJ4sUHm8GuTE6
ub8u4E9oBouOA+iJyfGlpq0CK0oT9nhnrzPcNyfsvzv8D4buGeKf4PxExLkDusu7nPvwsWLffAPE
k3h6tA2tUkKsgqyUT6OK3ffK+1dQ3bkxRVIZ//gms459sGY+CGbj/wqDfRCMJCouOd1JwEY/odHk
WnNoojmnfVOKQSSu7Pq9fzbzbsTaSgvs/Zbu37uoNnN6p++Q48WcDOcCrp2zNcG5vy9i9VKOLSmf
/qpXb2RaTO+Q32nMBfJKSe53r5bsDlgPwhIS/FF3FYKTiSN+4vxJRUCgtkuejMo3t/3xvUvH+OUX
+SAy89UP2S483EFkCw+e6QzuNyJpZwLzauM/lWSUHCaZp8d8BfDvjteE46yAJqm53zZSx0bZVBSw
/jYnCsyjgyIByvzf+mUMr9rnFjLIQ0ut2R8r4Ac+YdFHJ2C0zSmAFgUmTHrch/bzYINLG+WON91K
PULQeHrZbK8/F0mh+hdk663fDbavqZsvr0H46R9x/T3Lz6LR0etQB5V13nYbC+Z4lNyCogqSH/Yn
1UKGfEmRm0f61OVYZYnZxhPZOp9mt9INs1NgQL5X9uQVzWBjFK/D/9IdeMhRh70BIcI+vf81xYys
AD2VTAWCxt2uEFWJMYkuAXeliRGU3aeU0eYN+t6m+kBp+WGGqbkX0Lq0c6owx+vBwydH/561UKO+
qRojzUh+GcAIPmif3sQ9lSeY5NTA8UnbHr99Bkd2Lxo80y4yfwVe7oufvaFy/Xrn0W+i+VKhV5Co
ti4eP47+xxY6mxFMZgI3nBbNKK+8yfLSH1aFJLb+mrbcodtpVzusMJd2WBQT2k1Ew3mSHHs55eAK
3xbkePN9Jd3aLo9u0FILTRb2GJemtERTsD4Xj+jff0mIMITNLLX+0Zk3OgVeU87tcRZ2tXxDgAi8
gHVDLeUWk9WcJ664Qy2lfNXl3uU9SVmM904jeFw9PP7fux7suKC5gmlnsvJbzJraNmSA+3em0+XX
+o/Xe+J3E7kCFbS9IWoCYM7iJWDQ+iiVNx3NKZei+oW+S6MLhxzThSw51BKDdq+LX+x6Vx9XdasC
F5kXz8Hnv/ZhNETWiWWFy/ZGZsZcrFd4zNofcoJOwU/UIE7u0EBEon+rP36/ECpKnP3juxIzLIBT
np++1NqL6czzxsZ+igbdlrqkG0vJ+EuG6gtbnhVyygRAg3jhI/RGa+Wk7pjHIqzkK0DC9WTZ1+5e
huyTTvUIHHWg1obYnQSKY2vLIdbSka4AOMKbZuChQr+06rJSC4EIAQUXh9PB+NrOLY13g4+YLfRL
4gRCgKf3PoQIHE0ELDaJ76YQooNRWRpoEht42qjFdOcfNeKdoCuMV1C5hr6QnxL84hEa1FxgurJO
8LJPf/Pim0HbeGRVhZDbEFjHujsW6Smot3ZVVa1J7p6KR3I7wbB4QSolWbnC/SyJ7Ff746lsWWdz
LQdwzPjOezTdaGuy8wJGkG7+rb/ffCXvEutkoetVVgyplzmKg3hbtKietR6Q14uZYFSpdGPa/zTu
JVNuO8HlR3VEA1FTV2UVMmmi+i6X89d+KRw3PiXYYNiuvQkzjjRpGH8mdvxU3lVtsADoCItv5sfw
1XT8dB8yrdUydp3+4mT8BdJ1XgfL/S3yLubnI83D+4/lj8P7xOfA/Qsj0OINVqMWmELj0h+8hJUj
i5WnUQNgOv7Po6Xh6Uf3gQplLbEAWVNFzMFF5g3xzPBvtNInm2j5GvOZkLhAyXH8yufY+KQvg3Mv
vxnjYVsjxvZh7P0xmSEfRwtu5Sc6L1H2HvLTzMmIdncGgaLpjQM98vyh19k7ABhLU9dbfyYAbeOc
LqYgbzKrlNZqdiV2uTTbFYtDDgJGQShEbsfwgV32x1Pu1SaCVYvHb6uczhc+hANpEGiDlIN+VNWE
uioebgrO1rpl9MQG7hJKsG8PsDY5+xyoutHdNjUOa/PNDvH5/hztqZIy5wvFhrzBTArGGn1XPrBM
tdH1Xl/lN5xiuOzLdOmucYUj+JlKK4Q29aVmMD5rdUz3NMKYSaXl5TwyOaWI2bWLDjRbXH3Kl+VF
9I9Ko2alE2zYGHtGFiRVrksW8HbZzPjx08fjez9JGUG2PCuq2lKivTs4jc3lYQ8DabKdzAYWt/lj
SP6giMGPDHSVnCDWeVTjThTPHgjMH6lZmrJ07bqWLoQVrGWPbfZZagONepM4cEYUrhMgmo+psZWd
2M/CN8yYQeKwJp99LkIisEld3+JmeKFH50Dmfv3WCl9lln/7vLzXML9YnZ97A4OKb8y4n04XwGgP
Y1QrVtByKp3iizI5uoCipvikc/zFlKfOzM6D1JcL7p2kUEVoWUlnEUr4Zz/NZrX/WE+VUu7LVD8Z
pARKGR2RT0pNqXrSM+65BHXeDfvX18y68VG6tY4R7YjW86iQZOA2XPNpN0Z9PZ+ajvd4HyY9mdRe
QgdZpGAs4sW4LNZ+m70rLhKeJI/nVIKJ2PZ2WaQtWGSqbcXmFlQWe1C7rjz9ZbpOzu6utLoSOjpV
/V0dXZc5g9onEen35J5iHKCesrmTxAlU50TuV/E+FtPETYGOgZA28hPmdpzkReEt9iy1HYXhq00R
mwwTEykk/19t/cXA6P9MaEnqbsvphmmFE+BP0PjYczW6j5pAib95l8OyvN0AxBLGkBzzkzRVShjE
xwJvg4VojHm72ebadL8tCNhvN08rne4TTJkR/XVwW7mFJS9KhpSi/WxTYdrf+Wj3agU/bLhPeEZF
9wKzd4uD1oVjK0BuIvvzVkZT4P7sXVFa+4PR7itrqccw8Hh2T4ki1dwvkgQaKjsoC6dSwz7lqLYI
1j2nQzzsPXyj6T/LinuAqzkMaGC0EOcxS3JdcCTyzwlY3XvXxkb5jgyX/xyf90bOcbdKf1PEFE7S
I+fNMvEoiXPgHokI2gC6ypTv4XKSye5ary0qXSVxykrrfPHAuVxsgeYMrRmC9UkpiNYkdzroibJV
cm5Y7gD5A1+xS7iwPxmqL0CbtGtykh9No4A1f9bpOVCthX11KtfAjjB4xj2JKcbXa9+4LMCzLSrx
PDeRmMCo+r7IdOT1BhQhimSNxYaZNowrXwo8Ly4GqiB+8jxNN553ulQWoXULH0rS5/Ixo8YIbRtU
mxGbMoWga9HLCctN/C5FZHbnqTERsjUFeNUIOk+dJtv4cCfXJvA+wUuLBZ58Wk07P5Fink5PTSpx
MvzW1SrNCK9hnWALlR3alkadtBYjo3drecg5//81IuqUVHDilZA/zgMubB41AEKYCupN02Uc3FY/
whvMQFTgie43VjcSHgw7DEy/bZkqLG7ysJf9XW9o93HglbDCHv3Ysf2zWv3OODHNOOX4ig4FZPJd
F1mhB17YALEkR2lbFqnyWjU6lUE858IBosECn7R2XUKgUrrZ9XFzz9b2Bs3/TOQXmffLSB+hQKNe
OGiCZagufB9j/X8r20WSO8HhdMMyyxps0wPbIO/6VHAC6TZx6Uk6mgsjL+6JicI4X6SnRm1sYAxY
4MUpQDs5uUk1gyaIPKgCPkuLKJlGjG45cllWcmwi2R+ndiZYhVLB2QhtVaT/CX6IY/uE+mftjfZg
WDOxQqjzoXXQGVtdGuFazhC6AKVzZjurLDPorg3tp1ZB8cAxH33SOWQCDwF5DmONvu3xenjJ/378
3wLaXW2py2qF9jAzm75d6j2j6mn6Ad3Ycgo3ReOmZSt8z4OeaqqEvhv1KOYCIOrpeJrBR6YbLJhl
T+UvUtDtdhbmLjcU9BnKt39PQdqPGJ7fpqLi8s4evu1L5chX3TzQDDTPYOyu37dV34+3gKZDv2u0
u2qqgqG49x1cVNk3fEuslWcTmlhPN9thvM25d2uDicfcFm6CA66X8aJZfNWE29NxLa57chILy0XT
LkN+rda+C1YgqrzEvh9IRLAPzcDgV2byDP3MspnVZnEmFDNCFjPaBoSPaO2GRLrooQpLIYAM8VWE
m9IGshC/CWt6rTJRu05hTuiXmO9/mLiW32YRisTRcQasYepzF5KvfSKQXgz5l1rgmB4kSacDJ04t
KhXGXQU60xlJzMWuw2Chv04M2LOaN0jeB7bQhrYDlQyhURyqyMqPcyyPLohrJgVbfDb8SeYHH3Sj
QqhcUDEuzR1dTsZqjKp3zoemgdf1ZyzT2CBfUzPKU5PDf3njusVmX9kxB7wmWFQod0Wj4AOaLwzR
Rdb9716eU1oHIe/xqTo/JTo2dydZy1UAneDGe9KsrZ1Bo8rg44FQKrU92UVg3Nawod32dHBzdm7e
Ci26wWYw+uepizog33sKeahTFZVrd8IqZltdZ5Hk8YT+tYogFjgoo1fBGaZlSFGBub5qUbBrHZ2U
ijvdlEY9KrPhqkZjy6dnyaN1dBpCXI+XXq+0I7uPUz4EOa/dx9w2IBiWf6ZgXlWuOPgDJdU3o6Z1
To5v4ztwlLJ66+6IdX5TXVFveSUUrfVgWZnpsrkeidlZEWdZhrkSOGrScKZbBSVYyd6w5OaCVO29
gVrQQYHtUkGSCR8Qi+0Mi4gsU57AGOdd+6L9hoaG5WyMMYPAF0YAuvrD8xf6ku0mnytQKdNezCNu
GJ0QT2X+1f4hLcQFSoh6BdF51BQh5jQo1F8VcJaA2nHv3YAa92rrtOVOFSE76z8W7V6ua9j6eFZ5
7eGrUtJtVvorTfMREF+VwIBtXaXCnrelTUfssDsS3I4bRLqkFSKu7DlfrrgSwMVYLIDv08KNMvr2
OJEpdxAylRcV+AV5jTvnUIYPI/nVkLKYKR2iZBPGLTFBa4SFajMdUShD1DRMBY7/+gkHgf+Pua1/
xq769MfYZk9+uWIy1mzK5WYrMbV4WKD2AJTJt0+Cb2OvSP736hgjEIlvSPdQ6B35E6V2BdpA8hVb
dcvCxCCg6MKsHL8raaXWGovzSjD8YuEqVIpQvTZOZQGlPggxKs1Xs1Wbzg6iIkWuFaJQY/pv7qcI
HGIkJ2B1xDr5mYALSuFCEShkE7I33ATWjhpYhsfu461W4GhuW4ffnn5w7pqGdWbIP3RYvDBXFXKL
X4NP6k7We5Xy1pLVaL7Hfp/dBlPQQYeSiGqlc7IeEzcv0T/NZVFYyHItyZ0qYTICPNOWDlwKNgXn
wqjpJrb/L5AnIhH6ByA+kcCXFysYCJbvViUWCrMGiroxxnY7UItIzRlGexZoIsZGJV5WRv4S3dlO
3hkA1xIRpVNuVlVRwyQH+Chy7GNDItdp6CBiYcUwlBO01pQ4wUkPtFH5QW3a6nomAELQ3AlaCgBD
nFulaaiwSjgmNpjo6K50YqFwVoNmtjxwbYZDSXDEMm/mLTDbjdmnF+X++v+aRYieufuC28Rr2nRd
CBsU8vBr/jBhWlfhPd2M0xtS4QXsGfG3uvFpzceEKAEQltYqKMTN21IBgxJx0l4zC0OJd7deA9iQ
zdXEv1Ij4zgFYadVa7e/uoUW9Bs+ipKTOANb63p9ukzKeE7UODubJ8bYV74Az3BbKt3gE991Ynl6
wAjnefq3bftkd1s4etAxysCKVG8q+PMI9PYEFbpqNBvrLnlagBxCL8EyA/usZQTaI9VmuA+uYwRe
3cValsBsMKMyrYj9frzKSs5JmSrX5Wsg5mj/Je8bgec/IfQplIIfwVjqv3NlQMi+noiE+h/I86cv
ZCEZEkEnND3QbtaD0Zq/oDpLiM4nitt3S0ikjYizupKSrV8CKEh8PFoANGD6t6DS47x8ll6K6Yqt
KC7bjWb5v6cpdOuSHkY0xOVA2S6K1tIQfqsM08XLwumvIsFa5H/2oNR7yb5wzc0l16fV6E0F+VAF
2Z/UlGnAS8ml7qFHXwjMRl2oMEeWC+iCaZJpscHvivz7/MAx4x9o2ULiktV9Na11HCjkNSRssLkp
V7IFInDLvXez0l82NmYLO39CqbtONLCywAebRI+HWScZBzrC75yLGxljUFMQFH9KlyOYGFBxLJ1o
1I4lSwMuALJqZ+A5kz996oRwBLeydSNfyBn6picTL4qWYSvLoDDMM2vFp3JYwxwWTteCJfKxQha/
Hu0yvDpSGecPTyX7ecFDu/XjuR29y9Set27sDQXQceiL2/w/eLGyqHUfoNNiFU2g+KLMlwACfaiz
WQg7xS7DXQYIuNB0cfP9gI4iv8m346Mp1dm/lXz4faakLTVN6CzWobsp4yadM9lFR9lt/C6zLwNs
75Z7HNzeXoijNdUuoQuXm8hvcnxsZ4z/9UL+8Dn59MKbg+4vVQC1rbiVdpDJtZ+d3a8CocN62M4Y
lGEd5x31JjJ82Y51iLf70GqCq39NgwFwoU04acAi0/nx29BDSAEwJtnmKw9GgvhD++WhEt1+7l2p
IHsRQ2jqu8qxmEoWgGBhDWP00l3YbDCNAAqD4OlfmwjTHXpVnGYM6aUr1i+L8tEpIhfRStzKvace
Axzxuf9XuUPVSjYpNxzhQaVWlc41I+E61+44Lq2hMj6wOu7uq1ZV7a2IVR09BIMipuD84WQKZqKK
MzsPsGVFviCYWGw5/xMJGQOJO9IxDWd7im1ex/j9G6Y2lwKq3SfLbte987TkRDPO05Z9YVE9Y6O2
UamgWsPbvsd1RnUrdwAGK+gVr3j2y/OuR58e5/X7ij3uV19x8MCbFnVGWM5l+b6cSpGJsNHnx5Ft
+fC/ztIdCK6o6CLscWLAXEijgIMLtgA44d/ly/7th8x9kxH7y7Z/ymUCMODYU+rvllzei3xTdLBY
bQCR04BdULScnMZjAWTsk1KnrCaNOHaZkH5T1Ro1NsN3Lx7OksayvRbY8DVBB9OWkcH7C0Loo2Bk
2DcNvn62yGcmnrAuVO/fdLLGM08hid+2ThE9HN4oYt6T+vAddXeqbY6aOlNbn3n0dUCBcCVTIkBN
JQmQpvyzyDwaWYHWe0auL1KAE1t/JI/i0sqAc4N7DXGN59bvcEAkB4qn4AY0UuX5NIWr7AXnv9pE
DRFEASN87QnnCZFvlbjWWTeyUgfTpeJQftns6ldwVSpEgSWgqn2C9+TPnwgcNmJ4CFb8o89nFUPz
zDSWzpKl7g4UBCJP8S2HpUXasEUNUqSf+VBQC4CS4Sn+zGmHpoFfpULWxJQvIryIIk7AUkLc8oAw
FnEUofoA/hMw+xbJQmjSpZwhkQW08ILiw+QomtYykOOpga/Rv9uZx+4NcKm//ZDnJy9sDOXxFu/8
6hTV40qU1fMQmw4CIZ5CrEP92Hc4wOZBIkYjhWlbaW//GDh7y58B/PuDsxWK7bQOplVdJ4Mc7lE+
KRYkL8YDZxpcsIz/P8gmywjvq2ZStWzsb/X1E0Gn0pJvbdFni0uG1SoJwMeiXpJYaal/iA/d1xid
oUTVUmiRKDNrfx9qICHATU1oiMb0GGEymkE5+BZ/kZt5MUcIFQOHEOwsNwNIGxsUiAfh3WyPyTvU
86+ztfUWZzUu69mHMJhvqNyx2rdaPBpdwJ61Jl23MF15KkvUaPGQa2gjm/akSTOvKLNDwMNER+8Q
jxnzsqBbDw8/P81yneZn2QeRtakmFLL15EVmVt3raK7JXUfUbzh+/1uNNlRHZW5KMm57YePzvp3D
cT/J/Ea0ShROSdTHf+OSYYlTMW8TgSd5avct/WOfZ7Lc8/fyyGMdnfbGjsLBD3ogX7OaPkBL35GA
78XKcPmPurBEnmdAmZxctejU+5WvzdVxqKJzJlBbUhz+VUMAYFsI8quYa9UMWVCsywH/1b921Kw3
6cMey2ruunnquIZSFOt0X0YQL0YrhpGxQMIsypxonkS39ePWIN+SncY+vg5OxLZkqz8a2AVvfQKJ
vmoN1IZYVTtX1zI38Cu0GGIm5q7NTEANdJ0kgigaGSrN34qAwPCGkczxrgG35RBtSePZWpnxI7hp
gUxANbPJeP1pSpf9qh1wTeXs4R08ai+CQ23sEXxVI6S+aBnaPV1EFy7oTBb79wyT3IzTWwc5qi53
j4GI68wjcf0YI7ndL6Jt6+5Lyi20elGXfWq6ktTj6twjQHbIvXo6bo65jHAkHvqnR409hEqrgWKx
ZZK5WsrKIESg7rGEGctHiwKvEevIQKoKUHaiXVXn63DdlklI5ju65YMz/Mo1/OAxSywS8t3I/chz
vfQqWSTHy7oiK55zUum1ZrBOFc7//MW1Ky+aCMHNjk8B2oI/f+vrBLmw+1dlBundRPMsM2Y7gglh
/MmFpuE78/DGi4j++U9EKzni1PMs3itgzgsmPuOKLOb4RJHNyqw8xj6UMt+teh4m/9Eei/MhOoNt
owtYBN0Nr84Q1JbVaGkoJS1gbvr8Fi84cFXgqkcVBxA36XP463RjnypXJuJiAmCf8lxnWufTU/hA
gD2i/VgDsaxgRqSNsZlxX4UJtsExTB2oPxkbTarbF+6hNJBfxUXBa0jzu2eAD2nS65CU7XR8pOOe
0WiWlAjFwYeNPENjJUEwV6P2mmNCUCEUtZGqMiChGYoKqYoPCyjXY19XZP8PCLpfm0YhZx7eiXh4
/0zEWLw1kdSv810eRCokyGEiKk4xoTUV2iTNyzqapKyCLX9K5QmPScKcRf28imJg5cL83DjsFRB4
zb4WZCalMRSl2J/6NUVlvxfwidSfXLWXzgEjhyxDRB8/3c+7g38w3aNb72m2uj5GLBNMLvvBRHN+
AYofA+i8rNeCbWPtOaUqTlPZUk2BBm0AxbLfWKdempTLUMERsVO0TytZdIl6otzAO8gvMH3YwLTi
zaH6Z//lfK2yrdvzaNnhzYrLAjsCKySuq+UDo8gHhfm3Zzu2y28ImdjQd33vJoFExYjnm8DwjU0P
vDahU7b5VU2ZHpyS30vUbvEPld/NjBdfaIb3RBJOJwYe6X3I51CFph2M3BrmEpQQ81uZspxViNar
hxUjp9kcDCI687l4OfVuyXVQILL+E8VkNyGWzHdkuhlshUp26WEAApG7V81zxiBb54k/cGtkoB1i
AV0n6PfTxq4qZXlrLKYvY6tFiC01oySGYVlINU7uSZd2eC9uPOPHO98GQPq8SGPodx1Y6RSjk8x/
Ew7XwGwUySIhc366c1kHquaiPy9qGWJeHQsYV5e7pAkMmxcA7pgZCBGjMU0HIYUWVB4nxgVuhb5o
1/IUPp2aTCvZTJFg1UYo4uTAKb2tuf1YhxZlAOyZdF2PhYX/ar1WBOYVci7R07sSNioKAhyAskGg
DQOSPIT0o7zVEEXOY9URwvbdvib6YvUC7Tcp5svAb2kKFdGKcKUFBS8rGENH6hPIRE3sdxg8dREM
dc+KY4UUyc7hKrZQWbug9y9YoI/Pj6I6tOYAClL6UhCrH88SJdwLR68peVfHVSsNDwsgPneaczmF
rhBq84Gx21H/bnGYbnmevQh3S7W1vZCh0tnsrkFz2pSdwno2UnTz7a553tSCtVJ0FFn3VvxLEJq+
AbrQ7KIR1BIY9mqZHFkW/mVVGBDBJZBzqeD61hwip3I+RtnQo7S9QgcLR2RVjuAl8IV4PUl9wlml
QgpiG8wCVYbPnXyxrRKHdTnOnf/qxFdZURPG36H5c/EBzG5BzOgahliIrsZ/XiG9JLzF5I98nP9v
dnGLlWN/FhVLoCFJY5eqM5xSxBlyGnMS7nNXun+ExuUz7fy+XwDP+4/+wobyAZ0eofwdy0XkTuzi
lhy5JDtJg4y8r7qSwshuIC5zAGwpC95TAinjBdWyuMLCX05Y4OxEH/TbP9CrbIe1aJAoaBQNeU70
meByqmA2AR8bUAvW0gdEMobnnvxZApYupdvpC603LFgFlng7uBYNsN0nv87tC36uZ/1O1tgQ35oT
o83pRD0LrRN/WYrwVjESVM3hls2ONup2XYuwLm87QixhEj/Odp4sJe9m9tEeg1kesVGt/XVdtNuj
hzcQLIUSp3pRJ+BZU8IuEhNEi2zehmSX/NBwM+kSaWJoLsnM1M6ZHXEk1VhZzjmHtWfAcAnQqQ5M
cNHXmCQe7ebhYKgXhaaclA5/4heEOo4kgEMf92QWvkEIY3aAGWFeL8B5cz3ZPkYlkcJvtO0flqrX
2QpjGaDkp3FmFBTuuz1vm3dEAs7FFw7GIF7iUqrRrM3TeYYc6w9lgw+n1Tc5lIBcw5aWDRUfcvrs
faBduiwqiOU0TZYZWk7tbNfkMgARzH/BU/kMgScDQQ8wL/2uVwrVxhsaqtnShCb5bOg55bcgeHQX
eiMScLYUMMV+W1BHk3BWFuxcgNWmU/lIcO9LQWrzstZu2bDln1XaKdCwgOSsJVnhderQLmXklxp1
S5WXNLfxsg7kkrspZ9TwqVW7CFXO9hidoqRzW3mpxR3LbEb8xk6J/p9Twsq+J7UHYS0eIlDXTQ/a
tjg1IxUqW6fgUTXJyOl8QMynTKjy0STgVGOyaFR6DZp1B0t/y1tYNsJsXKEpMmKR7R8H+w79QOFK
TqjLQfJbFgXgPBv+QQOEIWMkQhyaVarJFq4DSkD2ya62vTnpHIiNmjU+nDJjo7cswkTcVPqpAjRX
eeU0juEu1M69CjIvMDXtssMi8VB9YNWqUAkBF5yQLGE0MOwpE0oRa2oULZUjg+hLGRbb4xLxbjd6
1XN/ai0kLqc34C8aC5y4HCd9vK/3c0B3RFXL1GS0yFx1Wx7RSlx47XebYL2Bk26DiMf7HUqaG2Tx
Ie1cbNNm/ryTG/OVTU6AcGjicuD212YtUbOXX9xBsGtyCEB+jaGhc0NbIBTW22DbjKvD+OMha/LA
gdNKUt3C1jMj+kH0vk+Tw73X8J55PVI0RmFdfT4ytj3mKKsLP/166JTl3PuWhmetHgRO1OgHUhzg
MUsuzHd418aOLYLLdpCVkf0JTU4KO8LfpCtP9qkDP2OcBLyeB9FOW4idaVNl9yTAzGrcP0cO9YYp
y3flaIwq57QJwiH1nAE77pi7WIoLcTLjkdNANJMfBF2+ekLsC2FpgoK1gis4YTjItWa3MgTwUlAn
ZjXiTRDin93XHpmyaTBw0OiEmmaZxBCLgl3830Lehvj3C2r7fVSPanFQu99zG14Yh+uj2jy3xA7S
1YUGmBNEXKEg2sNK64z8JpI+KzEp73p6fiY9KS6dYEu8P+KIhJVqn926X+7s+DTW2vXFWXDYfh9l
GMeXvXa6tdSC9BBRYA2GPm5hoik0DR83tLw3+rWW6XZTe9wZCXDvOULm5eBJLEm6N5KdUSOH7/Xy
FaeegQiBJuk8FOKxpohSWqd1ogQJWK3UOXB6WzIVdSF1PhThnCEaZLw65srJ2Q5TKEFJ8BTlnvC1
mVIlfXZkVxGzf/vOGXHAGpJfxKmAs7S4XfpVotyf2kbKKUICyuXqltTh+Q1LSOGtxC/H6ETFkLRS
PxNnPu4DqK7QIaRtZhOK1wybJCEC1mHdQqUrAWEGrKXWWqRRMuTZKj4br1YJk3+tEyXMojOs/nhp
2ACdP5Rsyf2xuhs9h6pvX8NDrrEAcH0wM+OXJVX9JMmrbriiu9e9EU4Bj3X5zkK5dmqI90pVRTmH
gbGEy5XJQqJbGniUMh2b11m3HH+WxXxr8MRbx61BejTd9LLDZPq2ZAYJ5uRHeImjWjQMJZBFFzIN
/tt7uYTB8cXBBUjWbO6C/vXiCrz27wCEis1io4zpuh5A/MP35uPQqyOhweNm0Kfjk2GE8EMLqpBX
D07kxY5/JVv0bNJngWT9bsBsxj8ALye6lxrb3fG9ZA7H7vhrhZ5qUM53s9rW2YssDbLenl/pH1gP
BHv4lOKStDbwO+SfQvnEoW/tLc1yW6IT9T/WMrSUYhveOI5y/rO1E1DD+9ndvwofyJ6TicFxOf2o
V0j7sItG1323dLwQtx1H5KBG8V+1VNg60HdwE0cAnmoF233lA3c3+UDrBHGIaF2qyd115BiMNhAM
7BLMPbEd8L0nCILkynwV4gno1WnNW5X/Aq7RKDSu3B8f0Wxtkv+BHEH9KSogw0IOs2KmTvas3tEx
+IBJ7fdCe5bNJ1UFbrNlBIEQ5tEvO1LzguZQWYq+x9q2SmwLn1tXf8NgZb7Bjezi4WU6dse6FgRJ
6aF/+fSuPmYM6BqXDVhNn0QQ7onQdBoKkMRWx5HzJn5xAHtgNTWDDCPpOK109D4oQTSS/ZW9L43n
t1GbuvnpT92a1FOta4T1Wsm/2ufljKzn+66HXxiDGV4RUdFYQw02WipTt4ryN9N2m6MbvLhRY8iC
PLnZDqYGOR0VZZ3pIN06ysjcGbi2HiJNS4QCXzssQ40wL5LS6P6/yhy5cISl/PKzRMXbFLYySW2l
LVLbWcIN7nrpLg0lAAnyNrUywzmDba4HY+Zud7++tYi56CjvAgKRUREVqDbx5c5oanamRDs4uxJT
5mHfPa9bt3ZuSgKrkM04q2BZwwXHNxVMbUNMzumkZqie/JAZxtLo98dsKXjxcMfnI+K45HKKfgXl
AobjpTjAgJm2Paueqj0fvXWFCHNtz2948nka69XW4WVmlZ3p5CG4vP8v/Ku4MLUsvJV/wdXU7baQ
mUL8WpDXkbD8VUMnhbpja1q0V1nLNYRk/wgUvjQaEZvIGPI/AqA7DdTmxb0YB3C7/3EzuP6V1YzQ
tgH5xk01YLDBEFyPD6H09SHCoYzcJpKZQRgJcgb2cixrBL6/jOzAi9ju7gjNFa1XTm8HeCSPfhmW
ovJWcqQ81YPeoH0kil9K/uEYLL1kWxpWM/8p6Z92QaFfzhqsScFZMHOKHch7MAwWrtso8PKQi7j5
lX3MvFvFg7iD6jBtAZhWBm2XEZMtjnOIfvW0XpmrjQ6oB5CSynFNf2Cl/44fHcws8hfxoRDhPoiw
02CMCje41tDOzxI4yfnAga8vC9ORVJChucScUGn0qZTFEJg2uRpfpa2/6yo2n5iJ5NTqvffU5456
9oMPaBu2DLA7QkT7v7pQqoH5DMU8hyou/ZiM0JLAM9oQKxfdodXRs1oxrd757yTdQ5kiVPPOxU4v
Ot5oNzlWAVX+Sr6T7oIVVu3sP0of/jx1HZcSGra3cpyoQg6Po1pSMIm18ukvbM7ctRIuQUtsxx8J
8LO1rWmT2cj0AmyJ+3WdrjE2nAL/EcUdV2TF53nGgtDW5TBoecgwm++g6gMO3uXhW21IBdip3VAn
SHF/ZKeQi99r0y6HylNT7qczPNJDUkaGSa9aoNLA2YhOu6GtjurFn1ekKVEjoL3FyFf3+PFo8GAr
ZYkRI9+RhPH500OXEORjzKKHSJ7PfioUOoZRzDxuq2hjCcqggGlhggZZvXkbuCAdxuXtNt6SP79t
dtpXjncErQVXI999ZRpWvyJ6lq8nFKh6UfASqYwUqkTv6RJKhxSGc6CLsmVLM6IFBU15oskmQQuD
JfTo/fH9cWAvbgV1fUSnVsbVBQQnWDjlpmWUm+rkPWIWNQ3FNHu6qNVqGMGGpKUfjEc9flaVhnZA
zeQpdxCIuEn/yubn8E9+0dGK6/WDnCJOcUUy1xP7IkJx/Tlb8zz4c6pcChLsKOVkpPP6xa29Dw2Y
Hg20DSUwMQP0SDvjMaeYEaXxM3yvB+GoTz1iKaSNrGlLPJPVr1dYc/07IC/Ser2MHaBsgPTBCt34
kfKnVfbEXlrcpbGeh44+drkKf46g1PwAY6GhA4OiA9/kxd2s1/mt3t69Lvv9vmKDm7CV+9ETdTPR
J+CfvLsHVm68UCNgCFMl7CZZeRgijXUJNMs/Z/poR5tIlu8GHAfY4OZo9uMQ7w8X6rnnOhzRiiVf
vAHFpQlnZbseh/j/Uyqq4Likduf15j5ySZJHBxIcNgegEddOY/ezXfFlk3oJ8j4SjF5XT2glaDJi
vfNAjEcjz1wazBTg2kUbhth+b59Wsvv0Huf+MMmIM7W2zq/oQoCFXrKViaYLQNFmc33uoZLgyZqZ
llcv0HDmYq3CLC5hhCscHfqc5yL3qM8iq720pa/n43MA3MYqqOuKwoYFLHT2ml++04VLgIDb/Xzt
8pK/pgzwGQBQDGUfvjMbh+iZz5LfFLC8aAoFdhG87iANcQLCIWJ/vJ+f4TSngyfZ/0CMnEbhOxoX
V+frsx9gWYxFCEe4No0Td37IsgWJxUqNTz7x8xzJGvvvJ7VQxaGySbpFBLhjxaORa/fFvseVJXmd
/ydRBUYXdc5mgpxRpOgSooE4Zk0qYTQuYPgfmJcSZqoSj+rU475spJCO+NyJY1b9TqaMWDqpbdIK
+e4E66tBhGrxKN4R65xEz7I/5zXHFJYj3KFqQ+KsRqKfDqf5trQcuFRyLrwUWtpP00Syz3cfJ5NA
aqNHFAEGScJ3rwVPStLc3PqCNAkjMFytmFHCDj6kYJBBmIFDu6dhw+yyVlI7ANKfssIC4d07NMi5
IIE2lFPkhGqISpO4qBQgDeN1x7daTujPMCeIzKYr01nTCSPQzuJdWDLOlVjTYABI45NliijV0DK3
pCvZydJlHND93bp+5SlVSJPMb6VQ+RZRwH808+Ho1StXF8qEk6ZVrk7Wyz66Ea02kWOZfxFPzI46
xv/LvwOysiF/nuSj2KLcM3SBtBXWTZZdlmw8ZoYzJLG/kcOyN/1nPYn5r4Ox5iYfbcFJxxNLaBVe
KgazqRzaCQVHoVs1Ti1l3VWfuFCeVOea+4UB2PxervFaTe2bvJgPdrPzvidtCJy8WQhRI2rTCZ0D
xHCd4YsWd+1iXCwhPqxtLdKodVzQjAN4P54xk/5+C4W8RNeEBOT7ssilWqK9f5qufWc9nWE34ZF1
heMO384TxHLVi4XH6O+PdxOxJ+TXKA+VWTHoHBZYOtw1bqUdIfN+qvaLuputwMiVXg3cXHsuXkZf
UYgJsXwQoRgNk2TI9Ngab+0VElBPW79T2zcoZwNHWKtmD7Wwn2olqHFjAaBb5pXJUR7c+Z2Xreog
Y1FamZVwOnMSnku61B5YKSCk39qaOEo/Wz/1yxVb4+qM3ilTIXFye1TJNZd1QMJSBSgmX4sptk9u
h5dy4rZiypU2BVaREpvov+lrQC/Ks+4EaoGvA6DFPBDbRAhpOQCgfgsZ1Yo0cBFVR31BVoJq6tPX
QBt20mOE7s8pZV8BBNdDV9iEsHm4C1MKPrapRqZlw74l345ttNxU7A4JvqXiBiwDpeGJAMyojytM
uFnRzkWfNSnsoQ+2ZDN1Ve5qhdbk16CpbTI40hR9MvjJKSBO7aHr2z8DK/MS5LXf5MiHE0oecDI5
pM8It6ydgN4qKOd5kXzfSs3wCcONoW6PuIAHl2Qtn0X84bWA5TVs/vGpShD+WEaojS/8lF7Hdak7
Sf90dGBEV49Vi75SX19OOMphJUwsLDt9MTbzZf+XfWjEGThJIz+6IeboluasX+6LdNFsCyjKtIgc
+nCL1+7szBTl+dz9eD8rjtTLxQSM1JonI4yvq+FN1OXSb6wCrYmorw+bPf5o3NTFcPC7pFkgpLqo
KbIyjZpb44Hq3piPIR1j9h4X78DvePsy7HdiA2gn7o0bR4UxQN8Vn+xbjKxsV40fakYFjBDyl8Pa
52mzyHrCceWzCKGnCzv3xud09O0351ODnMPuMvQCRhWdlfFmlDqCAt5Olsijs/QFua8F9zkG1yma
Q/pZ5JOZFyQmxJg+cTP4zCl+6ImdOUa5YbzZw0Qx5LkZEhaguMPnhnesNf1Z5Kz5Yru2COH7yjtS
uioqjz7lmRATI2UCcE/0WI5MHWtnL2bbrTOcdHsAvY0rBsn8+ECc3Zs60/T1b/XzL82NdEnAHUX7
smUbdHg5kaX7iTLne3L+HpYZtMu6TcfD7ae/Lu12fwjApFTraLGMPjeJad72Esnc8C186RAJaeAl
1+FVyx8zdprSZNj7aNBn7do4v4hWZBgX+Yr/HeInvK/ezEElPR7J25HsN7SDDdyUDQMwypY3YNgG
Y6ZTyVXhUe6kCQEWWRcfI7Y8u0TMh6zjRP59RvSBmpAR+7PTnm8M61vh04QEMzJ7mTyHBxGjisPK
MoteDN0eIrPWvo5VEecyBaRhIml41e0gSkAXBYakDWQEBwvFb68+3vqQpvr3kzfusbVzWB/ezn7i
nVUMNdqMRDJjMLfrvFDDaKmTf3sTHghAZ1rYYuo3h9rPqF0MWNdA5CkGHdPMDqcmZ5wnuDwoLPo3
Fo/jb2SzNSi3ohfQbmUbcLRNy0VR1kDiJtmrxfAzYvx4PYvIlum1s3pvYfRPkowPtLKrohVNkyGm
c4HPHJ5Z9qGJh8xKbhPHxY6bE6iJiyMV7fM7tkqs2laUupNWoBSmi0ZnecPPjkbWrH68X9gG0uQt
F7M6f0hB2zBvJBB9CxSIBJ8jQ4/9C50+3X3Oc2JCjCjhoyKdF1l8rzGbWj1Oe+qTYsudrO3WH/sv
l5B+lIOdnYtoyO2iGqhMEvcsOma0sacvKnnr55gYqIQZhU1HAHijlFjkmOJDufHYA6ZENFy/9Tyk
dQN7By3EG7mS4SggHJ2mbDnaj2IuUEgsv+tGhAH7K5wpgp+5qbiIOVU9umTCV/Qz3zBe6iquo7fc
sy0yoT9Q8Q4zbukPzgwxIhuubDZgKDae0sALdr9lfTTQAkyPFA04phM9+al0h3moEk8srNnwD/g5
82haU7fxxe92V9e7E/kASTwYMq/PJwtaUHMI9x5ISykffOoC8GGS8s2oYtwXrnOmQlxp07savCz+
+J+HvbjwSNFaNPQgAwUNfLKDPV2mOqen2UAPP270W2ot6KvgK9RoqXwhiJ2g0GfguNlWlD42I41n
V/obUyG8whyl+S2KZ8io2xswgrdtM4R3AaHnCxadjr1Xm2rFlrTPfcPxmM1iGBKxzNzoXGWMIsj4
FFadgVSDbekRGkWsmaO3QJFYUN0VhruRxfpvmnf2CAgh+2pwvycaJ5yKzNr3a2oydP6lgANBGo+e
mFT+4W15WWeN7SRam0GdTJnSEoM8tqI3VKKmq09kZASNOL0V3Gr3EZzttLs763cOJnnM4pVf4yZp
UfYER+djzhYYNDEIpo7fx/1+GoQxpcUnAU4tDO6599XjSjtCaCkChhLkKn7/t+XDYfc0AuWFBG9x
9lSLGHSY7aeImM01A8D7REnBzozQ2u2+JT/WMJeUqDFKlaNltb9MUVqwlPK4SdPv1VdjB/83lUiW
nYBEzP9IZX3g/cxJwwOcV9lvETcQQS3VooPAb6U5FfkHjJSjLhzdG8cYEE/hLkz9ofgZnLzhITGn
qrjHD2C8Isn8CT0d5x9qZw6+VUjs8MFRS04Z9HMnpPkJKrUObZj1KFbcW3yd4wioYvhQOdAIzzSO
5dMcL5JXOR5/sqmyQ7s38/gZ3J6HAliRiSClvwSd7iGW/K+S1ZDQoBs3GncWDU6ZqO07GhgNTQDD
1SxM8e+9UT7N/9mMsG47qFyZ/CJtbv+HkKCEsm2ONkKuffkoiiPlMz2TMxRaCIqEQMpZ3QyBIQ3v
poKFUx4oTX4AuBcxvenopKUwL5Rv4G+zoH0Ka23MqDATQhauSBPS4SLHGmKyFFZUvuw73GRzoHKt
mdDBLAyUAgBFtiMTvNJxyrcaCbVFQfKD7IdKf/UNr7oabp9YgRdE5Lw1tjQJxq08PnSWo1sEMoqT
GnYGgZYb+EhI4pvS8agGJS5dIeQ+SuSUMuEylt+Do4EE1CST4t+7HctK/FUuBcEykk3EAc/eWXlf
eCM1T4j+NWGVlkCgRZNG5pj0d5/ow3nee8tUohy4yn1PgsH3RT2bE68wu1TBRzluxJCwalM4mBKr
H0Bg+YVDjgdS/zsjyPQMm7v5hEluF0kKOUMpn9E1N2JifAXlOKdIi5oL5dL3xgbBEBEq313wHr/2
55RMIxSv1vdunwRUVvgT5oAn7iH4fRDX6C2NLud0iptBst05iw2VLLXP5r+/T5AGqc23S95RMk3g
3RkyEGGeYtxmGJbvGsL5GJ2rrKokoqLwz1oBnrY6Ynr9zG/Mh2YdPmJNsnpUkjCuSzEj35I1t4N1
5dnVdmeHSBFRdmoDomA8NMligo3GG784BJGGjz265+GUdTO/OxjTQnPEbcud93VR34D1CvWXdOdM
BCTDQ7DgDuTyi5zfWb72cJblARXJoNGP5eJxZmQ8zh2MKYa28LowjMC6+dRKkvqL5iBYsHlNC1TM
SU72YKMyV6C3dnBBLiXIUL07BNPuAfeooYuFlQRO0oi9RtoU5QV7AECAVq4P2lGWdWJU4ExZ6767
1NrElUImLd7kVk9wpqpHzmY1cSJ33pD42pU4clM3FJ1v/+qFngIdYX8eZZ3vr2z6gXCKDMfk6rkj
sHpeRhXfk529JQ6GPiRuQpTfJWuEnZ0HbWBpyYOnkMA7KGTgdAzUpIquVdQUnZjbrhwF52kuiqUi
NRv4QQZCvzTymebXIXQqwKAASZJouSuc1BbKv58Mgh2j7a6sbE67WCK0JFRlYoF0eiXzZ+CC2Rge
8fBWy2MDwCqxGJNhGDeg5bgj5vy3i1gtS9x3vgrQLefEcpw6QOa90NeTem0G45VjkPjBDr+g888z
qFSSyestr6BzBQt1l8ZEaxWol3pU1XSyZQjrSlDUIM24Z/UtBn8E9LvllwqN/ChSLA0rBXcXFEWh
WAI2hr5Q4iqabM5HqhTwuNmaGe2nQhhVO+fmQO4YxYebf2QsgOOHGZ4jVoOJML5dSg+9RC9cfxdJ
Ojy4UalzTX3j/99T2co/ulEFUxCwRbCAAJ46xadhIOfbt2Z1gDKSfSggkx/mMELPPmPXxEB6Yooo
ZH6YzCPED9DGJlT3XH6LIAiAzMjEikwIuiHoI+NHBEcpIc2Vxd986WgTjnxJHjF/R/EOv667f93r
GJ1gBPevxSBo+Vc9L+HtUeJ6BNVvNYL7y71yXFqCoGeRc3HCs+tT+FqP7BE3riVbVGf41LxOy5Ha
+mdE9YYp2edkkMF7Lv3lHwUmm20oaRJuCYeK3ul4xdoSMYo6NoethSAR/klk7K7E5VWgEoFHdLvv
s8mazvmMahj4kH38IVbfdEsUmM40wLb2r/6vO5+s/3UkSkIsj08X/RExMOY0YeELO0SuGk55goZc
1oollbcpe7caBUWDv50KeypbqC793Dk8tCKIWVIkrgcDU1tcE6hMvt/n3cBLaScx7AZOSDOXoW55
bcj6Y59HHZu/3ffKkPhzZ2Xy2Ja4QRerrrKzJn6qfH9+hOwQvLThdbUi1+F4Ov+T5hQJq3RkaIpt
RWzaMrKVxG6iUDdWXAAi56s6xm2TNKzqOscKFE7NAltRPqGkn+CNDztvaWRAoYKFiZlr5H/cNwMy
DXOfgDfNSktGxcgs8bpsz9BQrXU9h9OthpUyrgB6SSZxIW+MM0wxyVFkePgN2lgBD2Je13kFjWrY
YaHkX9tnuwBmhlZ0WSe3whmWSFRImNaIsDFPEVNOtQOKAjJHb01W/wglbDUl2th1t7aK/yd5JVvB
k5D9SlHzaLHm8jKaP0RG93Av0bO7ctr4e/tXkqgmyi3By1FgnwZU3MY0EudgZmXipWz0AChTBu+g
Or0cws4/QMAWf7Jpq0l+ughvW/tk37xAikRleZFWp/SBo5mCo7mvJe8c7oGMwk27iZR+3l7R7d88
FDgDd6XJbGy7f7OfIn0GZV+sUyaN8J3NS5lzcP3n37Jop7W2ka813fbIlWUof4gj5xTJKVXQVfnA
6mVEY22GwdDEX3Vzu5ad5tCC6YlO+qsa7hJDuxl2MEvtNdHRY4bt4+k26yVP0t72BfJjPcQQeUfB
s1a49WYF9EVQ595DtXYmcTXjLoPMlh0JUpqa3fR0Nk7/zvTdCYbXPY7U21d2spLV6vNUp2WY8rXE
1ZTEriTXzSNSFFTC5C6qb/brgCYD+Dt+OdkJoi5zXcxy16t2gjKAAw5nyRBvVSZtGj2b5pQ4KLxi
u5nWVrxn88V077WUnq+eSpJ9ON466UwAmCqM3+P9M6YSsxCa80DbleHePS0kMh0F4NLqVrO4TpRE
COg3CVFvNYu8D4R4nUbhX9N981KvSpjfuqJvnr7Q2e2QrDPeIHBhDYkFiWYZZqkMb4H+LAdI7BdY
Pzubafo+J4lOCmjGWOhFtHs7v7QCTTpy3PfiHWC2LME6s95CFr+1jxnFoZlZzupfqu/m/h7vDWfP
0DXYUti4RS2XWFwFJXwfsWikkud+/lxoCui7SvqtlfokG5clDAFAlMe5RfZ57FE8u1DD5E14z1RZ
ZhmJyJJkvdVnbensG+ykvl7AWeGqXCdzLSPmRwXx82B3Fzz9iuIQCxviR6ZFANtCZsNiqNAdiH/I
5Ja1ww+5eNWRGFHUxJTn7a3KJ5Oq3EicDOjjpIwzlyrRtIf0sKKLUYCaLG3s8UUB2kfZXTOpiEta
UFz/W/3sWCTPOQcrGmKZ97130HkSO0aX3PgfrLt9gt72gDghnCNBjKtg1Rq4k7F05lPKGNZ8mQtk
vRytNESSe1aB1gLC2WYWSnBYyHYmysEvFuF7xZqt0cYgFdJpJeaQ0lXqPdRF5M2EILYi1u+cDXTt
j7DdX86wZNLoZrV9KR00/tym2/qqD2GYP8THTYpWW3296rwzxSu2FWERNw3+s51hwUGfqxPmfHbn
xz/i3POT7c+cPHRE6CopoC5019vQvINRjXATavVDP/oTNP+wlR4juIWkCTzv6uBYcQJDpFrJ4CAt
L0tjaVqkeNe6OmsbCNkt+jOYl7i0BzFTM6vk0H3H0N4fqPf3Ohaivpi3/HA2lCNDeMsbnL5dotgg
YWy3FnqwbHfcXVv+HGHpU3qw3oasveYD2zpFEZXSXPAen8tQjAfAkO1D6WWSY5I62xrZ6rWm5wVf
t0Vpfs31o2GNRKGMmb638o/NN3/vOsicgSDtscVM4d616rhtkvGVja1f3YSDYWID97NLjo/bddC/
xOrhuMDaQMfYvq1DXS2vfMJvrDokjpZRCMCtOsd/aJEJAGln3SVhwvvL05tpn7zcK2HwwRXRdO9j
m2cm5a0oHFW00GVvGbhA7Og/JWzSbDEwWQm9D6YaJEGAD5x2QQada3BXCvnIcqh1okS57zTVER3r
Owe+ZCcWXOczr1OkdmryY+7mwVn5il9DM5HSzbHpEEO0kmf8HC5iLqYn3aVTPnjE9t91DuWe8MP8
sA+jEiNUjj1Sl+WFAuSntUxHEQO6KxprU1qHVz8kQvmpAbp/YKsMKixnJgvCyKdWMuX2ZNoJpXiZ
ZWi5tz99LuCiyfuItAZBvEeO3c1i6TuB1KQcSCbVlOUPRkwE1g3AjLUPv/Es79d5LoEog4ybHkL/
MUvXOmetugJWWxdAVlN7/R5j5/I/vES0wqBWznPRv7kZjxpH0zaVVhQytfsQIFCN0r9VUULe5QIq
WekzZedmGRBh5XbDECj9ei6c6Cy0fppk1a1rGFfcct0ZdbUK2Oz8j1vpqAPCa9naT47lHAQkO2Jp
u9Kc9K49Qeje6yhuFVGTulMn17iIKmeBj/I7xaDPPIQjhHWTbVNsQrz/iVDiZ0H6k5n43LPukohv
k8krUFL9rDQCpt0iSPsTR4nsC7/ETeYLTWX3AiZ4Dc0qQ+uXbx/UIJuylkiBC6XLH8ll+KlhRpxU
5fEOxt88nxvHS6ipYeXh59uUIzg0qoding6g7SjbvVagdGgNk7MGFDg3UtVb7eUuZVcS/RuKkN+M
22T52XiaPpJNnDio7tFF/xF8QU3aDfPhKD3HllE8L1mA8LUmxbPgoO9Hv3JDjG6mFclYsNWKtYUn
DAeAd8QvkpT8D88ipPg3wX4tXb4piahZT6APYyzgSb0uOgipfrbfVO3By7HxTHFi38QGK0Xs9QN+
bbJH7yGBHY/ouRLYA4l1Vbp/yFKs28KELy/odlo7kwWZSxOFSlzvT6V5hTTZjhDSR75th6kYm33F
Sg3+0/IKOMmOLzETIz0UhEYAoQBRWWMPvFmVjGQWqHX/412mJqVZ2xsEQ5piCwk9UZSk3bKe1hlo
3SGpwT4mkTfPDpKCAZlr7dRRmL8XV+IW1dXYiLEtSDicAsT09bJYwY+FpDEE8hFI9wtIrgH3RRI8
bHfDl4exeZTDb1bQ+pfog26iXkGS9y0bbxNvIOX/LNNt6X37JLkeW/RhNU5fiOpeDw8fOky0MYUV
hjIPho3bOxAefcbnxRVXlPJNkA8Hv0hIkYg+yJ+GgiUn2DPIbZz5m9Rs5CR/MqEDWkC19w9VLkdy
oCJ8qHYV1fZBL6jgIh+ZVeZIouLooLEEp+iugE7JV9Jea0qYVL3WXOUJXnszh2NZFGJpvAjJkg7h
doYSMR2l0cxUBkhB7IMyoEkZdtDH/6fQFFzZLQSi2gkrQhU+n/HH0dQwH55TztwLdwu6T4dY6wWi
Ry/NXoza8KpM6uQiu1eM4fbBJPwFrh1qK6hVE9JARMxa5Fact2+mhZinYDKt7vssP2leV0Lqslgw
ttoJHg+VJjbnZqmdHO+s27i/vK7B8jXpAs3N6j1LJMNNCVapjUD/+Q51/XV+NipTBt6wRpWDjxSJ
eFH/xXNRN3nYEOCpSVmCwwmtEo9xAvVRQnpWlr/30h+MIHmvre6/yCAOzmXZWBjly/YpgBinK49v
5wn8TrkwnVw/SFU1X/uytxLS5D1g99j3zHASLaWy5XStlL5N0hFsUciKvPXCk2BrJUGTTwQFF1nb
mGS0yoBYsoqZ2uQCIMLsCSvmLKIVUyX/JxVWvjHHBsbK1SWT+yDovPWb8jvceL1hcvGuoIlvD42u
1k0bg/eLtlpLf5UvMhs6pTnyI2+TiYJsVbaOYn/6vT2SuLTXA01BpWJpMH6OJxo3VneT5hk7IKTF
x3n+ke8MsGuy7yh470LxxRPMOUvZIU3k/143BBdz3t0DD+KYgeE7qZLSIamnWH/IDg8MrmIYXuFT
q5S40eYHnSYewC5u0TyffVcJxt+ENqSNVx0XMWwwZ2xyQ/rXrnFkj5oiTiTP9nKUoYrE7g3h9KGg
hFEgUyWYsmM3GKGL2ywP6JwMIPkRQy5AZvzvRLfI154YDZkUFHGqNce0O1f4y2IUpr3PlV2sxQUm
WCQ7O8R/AUrHGM/zbzwNCI8bdfIt8mnrVHecy14sUwVuNzyHSgW8PKoqLdMlvoWpqjjxjK2Av0hK
hzKw8DfcRExdJ0v0pUBmvmbTsQYlqm/9CppN8e2KOOjsEVqBMAywsxsrbNUp9/ZkxvDaxkJ98Yun
sqYYwOwa5aAGMr+zT+MO/0ODTTtI+RYDKpSQgqnzjXK8fR0UyRYYn+9qc3mw23bI/76mReruiKAo
XMgqeDFwMx3nxVUcpfyIrT6kJO3a3Oa094qI2HxAw3DyDLnmYkn3Ahh+RxEgRfjdn6zh1/6v7sZ/
0bGcghuEn0hjT42NMFAi/ZlS+o8naxJM8uafuZlI9spxfOeM54X4RwP38uVdjkYpHlJtNEBPgsRs
X1FVD01ZgDHh0jtYrvHraQc4j6Jf3TwXVgj5cnYp5nawfMV1vVq9ZBsyHSJGSdC9QAWJwfM1k6Kn
DhAcZ189TsDHmz7PyYDFufTmoFEzabH1Wh+8emDoiav04htRIEfA8qaZ7zNxJGMMo8dKEIOzKQN4
wFspV74Xv/PvK5hVDMVZiJG5xrtfgfv1pCL0w9TLc5UaAL2g/YdhIvXBlBWupcWRh4HJuA9kOiwd
mXfb1INE26UGCR0q1LWLwMEfJUSpPKEFqNuUXI2mhrgqRNU9KcAY+Uhv/O9z8FSJ2l5sj9GpxOXg
p10Rt5XGwXMMBgDs6/RhMTdH2LBz3BZLSP/8IxjdfGUcJrwY7pTnfrZpFf8++uQ23mfhuEuC95hK
BdOHSkIbdTZyk/EQLbe04kThcyTWmo4m5uw3PgpIapkhsJGa8/3mDNJ0v16JkpgZQsDZUtMKwdEp
T/7Rgva5j7VkgPMk6Ep1u0oJKImSJZxGrslOBmgdM9k5GrCIW5JtvVGsNxgSB58YxiNObH30d9tw
1YBzamXNavO/TTOaeHvHYIIvQHfpTLGKo35xUTLpriyIUGlelKuSBRXNFDbUoW9c5xR2+wVQjzwA
pCSEzlrV7lIbqleSLPWqyrg1IgmFnvDpvRZxa8Qv1os1eO2iQfn4zRQgCzXfjAc+72QlpB2jSdJo
bPwW4lQZqG2DrR4F4SF2OgKc61sTJqcgZK2MM6hld2w5YbsDUjb80ERPIXbS5GCm/XH8ovErY+gh
QYDIfJc3E+3GFc2ZkRBu7IifgXhBsU0pTq/8EJPlfhHL9HI4RXbkHYeSgs0AGfv3YcCLWzT1aS7n
IinUKIuNC3U3CV+HKIz+IkQG9lzm2m6aJKbtbLx5toDg63E96OP2QFdPt5frT7l4d+ayKttaUejs
3qnkpBc8VHIuSY9P2yY8u2Ubdb3nfsb2GVl+MOdIt1Ev5iY2n1ObUscgqRtgyu9QKE00Wo2O3oKo
+Sem1njDQW9l+WnFHcWnvKVgR90DWp8zToACc17SPujM+RNNWB59uFambry4+hoGxSB1os4uHBI7
nJnTOeHGQD/DvhIo6Qa3DK49K7qfoE/SnAd4OrwbG2v9GDLWdoaK6JfDa/v0pVT+ot1seLgZDajl
lvx8TpjpxA860GSWMEYgO9ruBwTf2w67OItYwnLI7JkvCUYEJa+hhdhsTPsQ820IaHmbtvNP2RIe
YxxzJg8qcX74vGnmD+kvhjwQOI3oxYCSRuKwxBCZUAwUJ4fLQ77zvTloBy0Xt1Bxat+rwEgC8L3/
Xp6+u4MPkmnJaQFY403CmPq95orfi4FN3Borp+IbmLyLTPpAir6Zhr1f1j5VB5KH+/NKrETlVDh7
b+4cA+N2uQM85t+rkgyoAdoPRKI8vO+F9qh4dk/3mjsZcKabS/fmATX6w267BsQEaKqp4enYaHJc
1FX1vZZqb8yxHWh44B5NOSH2Gb3xz7pXkAEVPHOo+eVhZAAODJHdUfN/p8dQcS8/3+Cilw/MVJDV
TPHE8rEF+a+5Hqd/zxEcLqmmxYSX1l1fwYr2mCc3Szk6V3CGhIW7WsBbPubMQ8zbXwdMlnAXfOWn
9RtDYKg+/t4sH1/Cgf9klddxbuhEIFhrm+4xdUswBHYT+ue1F0K5Bic9TyX/o8+HpH0W6A7rHrx2
ljXJNTOzbbM1E5Th/NhSB9oTjcAlyvc3vr/bGn+8p1MivcCBQRWfSOKQkCWlDn55oh5B8o70pE84
gTvkABPqGYtoXfb9wCftplsb98PMJy4fOiFC3+69qj5/07qTiPMlb6Xr+Yy4lFsZ007MRfqbqVa4
HBe25BSvDe0Eca8NKISkT76sc++KNY+Zw+kOUqyLdgQiEnST5V4HkBx66W8ww8bJ+hQebxCX1Tns
/uWPZAKf8MCTL7Hu10k2kM4b5hdwzakJOP0clqpramdY6UTS6y/ZktNvEt7jChuHN/BvzzJ/+iMW
5MDAEerOri9J4YZ9l8EISwqR33Cm3QkrlcggOKrFa0bV8QUP4pP3bN/iR+4NPRleL6F0ovbAhVm3
6C+7rj9s9YXLUfyZwp1t3qiyHkj8k86Utz7ZITEGARgd8UsHvBLM6MzrKF9aAFQXCp0npsf2fXIK
lx2ujwlvIO3oG3ddsLQMPaGH5ssYh8D9n6y94x144veB5ZUiphYNEFSyWdJmNa2sAJ/EzdHGU6Lb
i5J6sxC2vLQTyExKFqdgiBjbsuuXn34/TvGJNMk7SssrCXBKRkOd7tAT5JFSlFzao/HrfxM6ZZG3
XE+Z/VhXMkhWiH1BIVjjZTMt2CK0hPO+4VqH3d90MoGM7oUZAy0TswjuGRI61hcIby5GgGFotRqX
4/d2kYGX/Lcn8pUnh/2y25WVN53Lub1OjmLGF3P0pln5eIlZstNC793+/c4j2sBbMVwHOKVH6x+I
sxqru05HZrOFUITWPXJ86BsmHAtysgrDYkmG+73+lvGKDi9ORI2qLUKSClytiwiaLS4nAFfNmmhD
Z70+5yC3rGaA/PUHP4595HnS3LIGPzW2dWNeSwjjcNN9nOmni5DkJYltT5bmJLaXAI/pB06Ozh1O
kQPE+ZrnnoKa1p5QLoLfWwWnxS92Il9R5X9BX4ZEFBKtgfxd2kRitlNaxSYBC9FyRAvE2QzUOqw9
13fd94TvxFvcZSbeREFtlaP8DojbCfaBwYcPi5k3+thvD3kgf6E9yIgBWvoa8gY6rD8Vcm4MjChc
o+r4p2cm/jqR2mx/nFE3u4YGLEHab33OFRTqx7cL/DeX4SyzuUJDgP0XK/7n6wx4X05yYfyVzvmo
cEX1VuXPk8JHgbtea4GQPEtp/XGmOTxaWpG8zZPFk8qDeADVXdQ0AOQpHSYcIoHp9C7hhM3jhb4M
8Y4OvuqCsOYH8bdXgGeeTbMrQxpgVeYGCzZF7JTJHzKJWJkWJR33pabPAwY6GBFnieeHYoJvaMGl
5swjrKixvU3E3dsM7ZGNEzNZakezCoT5TTulwPn2tSP/m4ibAiJQXM0hgmcV1Dvwf2f4FXlVUKBF
Th6lZSPslhNB/fk9JuMYqk3ZZodGBH0wHq5uI/ejsO+y8s9sikVz9Bu1Uhj1lDLJSm6BoDrS/HSH
eKjjo9GtihLoyPwauQ9P/FNp9U2jgNMH8rlMrq2+xDgmQ3Zwxgf6o6GfPxGTClkJmghGDA22X8hy
V6OIBLC6L0NBrBA/f8V3z+IOq89q5kwoOGep9ie6FxNQ//MKiIi5X+bDn0o2IoxvXlFvRCMQRzf2
ZxxEvTp+CHn53HeR/vFL1z9jbeQW/Qj6c8nL+SgEm77YHEXLSmQLKO5g1FatsNQe9w8/lQ+2AGdf
TvcwRpOI3R/VX7zjmvXRCDRDJYVajpa0l2otckDU1ALFDye3LS51S9eXIl2qH8GmswepUAwHkXcX
u3rE11iN8QafDmzvE+HNCYY2CcNI6u0EBPOfKsyW5OyqPUpbnv8QwFwig9VDNHzFS30/PrYVpR78
6LU262N4+tLcSL9Rx6s5IHULBaKbrvx7Itm1euGKpa3I6ZXRdslYg7WgcjQzPCQvQ6DH2Op5WPOY
1KmW4oJZI1h7vLVGZSALUUbiQ47b4cOPaCPVU9/tGCgytbYUuy+Y9OmeBUjFvSLzwG+yN9dspY3w
/x5IcaFRToTPWWkt67i3SMgNNwIJ0gzEULK24KtfHYoBzRQMDHrgRsY6K5flgNIeJ4rtnjH9HpTG
xD/MtxkqxQl7X/ockjC5PMIn1bq9pNFHfQtxCI0Ch6wsMZV/TcWHNiwtQBaJiEShp1R1nV1Oplzw
KQYaqQgrW7zQ/OkQImKBwPR8hsWo1oE2SuqX+NT/VkZSCs7rXNjQ/BbEJ/1NaIakgZOGu4LM5Pba
7fBS1QZt8CAiiSFo3yugyvBvWAtvvt2AX366ihJSYg9lJvWDJAjXsnAhT3+xiMaEzJIQw2FTbsAL
EUAES24WBY1NeOr8D0npDGTZVXkwYNplkk+kmN0umLtKu+SchtWBiBLie9Wl/SvicnHojWPEQj5y
UTgWOxyBtwuik3+Ai+Q13GcdgP8ookbhnPD5mb9niOVlhuz8rupxpSciuohrMqV3+vsD9jBciZ/G
wux15Ksm0eOd3gX+0TQSIP1a/L9Kex0YWLacbeBd7xxORjBJs1p+LMnEvps4Yy2S9VlTVGtsDSWL
0XWrtjzieCauptMlu4WZCK0qgEaLXB0/5mlCos3Z6EsWqagaqaMwffTiTgrvYAgGdihUalakLvrF
Eujm7ggaMQgWOfwhsr43TBWn19I25wSgp+h3Tz1i2qHzPTPWcu55PLKIxkrMGt9YnDaESKjdM/N8
P/EHmZ217lCLT25cAG+uVVFyOGSUyaQNNcSxu0qjt9C4LjBj//dILFmFxyEczQLzeeV3ik15ZeBQ
Drt6we2wUlZRSb3FblpABHFGP/Zwy9dkFo7o3wwzKKRaugkxZjbzS2Jx+SWqgqAdqo1CBIaI/5bM
NHBIMp/NdImE0BIFLXjt/5oOCOvv952V981/UXlk56v6Y19wmnpRFJ9RQnjALC/twe5lFDxMo7ps
+AjiwFUbBMlvbJS3gvnHHBwe1LDB++QcOfyGNB6SbRP2aKARRW73mUSmEOVCfKwehaZBTyeBOhiu
izPIGGeV5TeQML8lxbexC7xK8lRiz5MNQ8nYFQUF2VF5OQMKuvaX+v0u3OSM0QIWAYQf5ow/PfRz
T5Ta2KPY60EdyMriURnrpZ+mhOqsHuLHSRuY3UIXhefYA/ckY+kFnbOn6fX8PCH9q/rAbG6p8OCN
XRpncmnd4lgYomlXwXzFXu/Usi4YGG396kz1VOLUhTw2+tWjE+GY91N5XvaNvb196wGLkDLm1RwB
bub6rrzLWLK9RyaJsIBTMFf2b/+24L/eXzSqNC+n1pQgxsQI5mK1ioeQjxge05KqrqHAlEwdStqT
jpGQtD1U9qCYPENLYmQ/fmv12Iyr3jrIDbb/U0BVOWIzArCAtVJP6AGY88WZc+NTB71ZprUL5AiW
vbwouxrvYx9pd8u22MhCwdoiMh6fjQedB4U6I5nCuv9SOG3qZCqjc0OPeloDUYp4l2PUiMNqU09y
UeeqrX+cy3u8b0kditk1LkLbC0zxZGln0zNdufKxwsQT1RmkHknyIOhll4evqOeoFF0pZvIUTVaX
WxRLfchkgsAQE3CzcS4rmXQGqDZR5Fi7jI5QZLz9j4bX+kfrsYggGb43Z95X4DUD1gDYKj/0kCCB
enuPRo7MfCugbYit4Y8aKSwsp/BXn20i8G/FblLuYJWJysySU0THwNAfyr6rDcC35Ds1rnWYGFSv
7SDfWduyGDAMn1IKRT92jE1fayFvQxHehdwe7y2+miXwXNUP0gewK+k9Xck/BhuvFJEkbv92TpA5
NeDd5hVje2PjL7TpKhCUHhyh5SR/bRCqLlgvKOgF9enarmXjMUQtf0zLAm8Ie7a7Bp6aEIhe7VM4
1Nb8nKYjfMKzOXlOroaP4Iec1H2f3X9rhEeLreN0PeukbBJ+unsvaFDAZlOBnrv+YGFxFBrPdDyq
JOiulGbuULgC+pxGLDA9Qzyq/x5dLya3YRuG/lqNEfHmVn3Cag2FU0qW88Pyy6RgYmJl7uR6eT9V
39JOuLXCPN+rQtcDrLjdcoSPhNLC3AIi7pB+iceKW25KkFS3FCeirQewBpNyn70lGpqru+vxqg2z
/N8h0zjt+RhPA+UOdpJ10oR7UpK7DorrVtYrQxgn7uyuhjZMLVAkJDMcdnAF6jJhn+bPYdb0EkBn
BInYTCQSuyySVo7l+QVOvZaMFDf3lPjbWBXEmdwXISO6QrMjt/w0LmzgaCDjdHZ9X+jMMlZpjYhM
AkdJIEzdUHZoMbyc/9PXQxHeZBfogGuEFH8pt6QNo4GVGQyDISNQReqOoZ17QIAxqcYgcdCR3lr7
UOrZNQk3IFYXRX/KYPwD+wRpjnHTfiPapEg22t+wHkDU/aOO2fOP2+ieCFHgB0+2nbPpaEnSg1VF
cJTXM57hn/5XjAI5JEq3P3p1BVvvfyo07ifjVQmcoJmwWfM+Vi66eJ7uCWrSBmrdSR+9Wfevyv5e
LgkaIkHoPP4djqWZtmz8FOecRYTYAP+ulgj1+F03pZQQdJyRdxEr7z0ITWDyX1vle/lABexqlmbY
KU3OpXEMCObsepnoD96WHGF9QSOhQ0XvxNW8+nlBhGj3QuBbvZ1Ki3qduZrjx+3Lptab6XKPV+DQ
e36zOeFDGfIVx8rD/yWwMzpEgHOTA3Y3FtE3wPh5PJwoxbTP+7/LxVLsdUugTmbQC4TlOahhZul3
OuEMI0vaof1UfrYNSIh26euW356mCMlGDMuLqGKDFaQFo1IX2oHt0FsxiOXzUgirrbl2WWMfvqKU
HZMUis1dfRDoOsLweRRqs+7PUXJSDi2+7N0GH4sGzVLbBR4TGX3wcCgUay5k4s/dhv1U4ctd08WG
HYfa0uUwq1t+tbut+lwZBT+rRTwdTR6xWgbAm3qPANsuHDIdm6D4kZDsxJD3zHz6cfWSFYQJzc/u
qwBEbN3Ae+Mxq2WYrP0eXG9CjhwHgDvKyKnub9m02cSPGgYNiKyv2suwtCtZyzxUx86u9TEsWNLN
Ja+4q1jztBnsiOzOn0RbYrfJrHt1zHvzebzkzBo/6sqisCWFo0Jba+z2d1lNk7bYCdZ8IOciCNYi
f9cW9Xl7GMu4Sm/pi0NpB8MkI0rtgsWRyavx0QSMPEh4a4g4qdccPPfAdcXiZpkwKD7FbRoiFnuj
eNSy6qIr0jQqlRqYwAhiKdzIx4YwxB+J1WRe84gKWOP2ZlKPJfwtsgseQPtwlJAPThM8fWIu2y7s
RJ6RC9B9tCaeOGkY7oKW7jkOPPO6mC17axNkbymTRIYSoV3g8ZrqIBOZ3T9CqCsOgTyHL3GJuyhl
dX6wjv/8uJFM0JHc2XH+Uaz4ge5aWsEkDIckJm+zmWQBLW61P+/Q+2RbMe5TotIbywwCvXSLqsja
OJMpImXPerme3V8J8nVY+SwE+/7/rIjuxIkAtBuTSVAH8MbCajfvyP48CNdIVn7pvH7GjiJyhBYD
tRNqV4CN3zHctXpWwvWcMEaH4jm0cZBRrUyLgOwRmrwEOOHUOAe+adOQuOSjD1fwRoOLObW1pMpt
Ilqo5bFjqdCeVGHBI6T7piJlNyBrRX6kEf454qONOqLeMQtD4dM8x5D+/h4SpXXNKJXGiQq+AhvT
MR3NkqJvo4fum1/dxO7qHDGBQmaah08wHna2oe9peE4TV1ig3CJdk+IX+1ivEvyz3k4EuJEl4CB7
KNuPnC7l4F84SwK1e79IFratwlW8bcXNBnz7gw9vOS8ieq5pAqsvDiaEbwup3EvJC/jjLUuSd97U
x5YbTm6KD/jLNi72HhHdC+wF43WRP01THZ1TvYXIQc7BnX+rrlLz/nbjIJrg0TH2CrfB47YYalqf
hyrK4J+9y624MpBxjsmtkkktJIqajvRZaR7p1LLoZnHieUT9dYa2xfc0jODqTn2KRydBP10IDlKv
x9NEoQxXJFpqYnF3gBG/mRCav+mg0U6oYW6v3ixzBlR+TJ8hzaJfnpBhuO7+YXLRS9FBKnIARr/i
hg2FrXXA1i52HPRQ8jeyrAsY0zgBoMSgWYoScON++4RBwGsyAkbZGjt13ZJMKGsvwllby+mWXlzv
xbYeEUdNVPRNaMAUDkWSe0p7xwG4vh3n7+vwkC14xGtjOGJvKDcT6yjtw7U7it3mP8dZHnHe6HIx
kNbiEkyRZuL7cuuK6FvPCkI7Jaz8InEXUNy5wIE+JBjSftVTlhZeKDUVvWOWEwdLhoxrWj921UqP
72zaJdGYM3N8RU/C3gi24+3PzO0Ot13WOTasw1Em2MZPP2O1wK4xUv5nufLkYyAJVJK3S2IfZwOD
EMYnOkWibGVQKCCbv1Dd7mW2VffGHszuqvZQv7Pp5ootHhLuiCpIkf85ZlUS+O3BerWfLOwbPEOe
BtKFYV8S9SJ0mBfh8mVYUSbaXW7SB3QlPoMjGhbArUWA1GBdEd1VdTvW1JgI3cVTsFNXxoCO4fbr
9WoXsW+dpzupz1abi04INZqKCodEchr9wQwQ0rJVSPdOtyFdtI1hBKDUOixG4fZb3VYU66vvHIJ8
LfQWS8YsASOg1nbmPA46a+SzZ2SmVByD9g5OJzxpng9f8oYUZIrQYdXS2tXEPv6uKiwAOoLgeoh2
CvKMiZtfVQLnpEDBC0p/XLz2aTuxvU0FuYaXSus7Cznuxe5YwDO36FDHm5SoqzLJj6Cc6fh+lH8T
NMHVntk4xFKEXGNQS+uIsdHYJmE6vvPogGo9UWfxMRca36H7AnI/jlDPvcYsakHSmV2IGPQuS/Hv
yA+MPSw+EyHSgYkgT6WAaaZNAnkTxb1RK++wIRa5jXtApoFf2nLd0RXy+n/YHaB1NGaP1vrfWB8p
cXbkHrcSCuFFVEqvkKwzwP5hBckUPUFT/stq1G+7LS1EcAHlrsdsz7sODNv4mRnFShym5Y66pfZz
OIWPgO3oM/+ER26C4n1+oH+eAthNn59AUCXc8WSAX5SILg8ST2g3IaSyxe/hCTzvo12M7cxIaU2k
aMinmy1I9XFzm251Aebrm2dcIQhvZKXWrP8ch0wnwMk8auG2P+CDtU4KIONfSujieLtxcRouZZ0q
5fBeSwoHtkdrVn5jiYztshiaTJMkTAmAQ12+3pMmhduLcCuqLVI/lOzQlZm+HroYxlXa6AoCfCOR
+lQXyt2ZFdmwYbyqu0yA2FPdV6+DswpzWTo0OkpXmllp+tRPBsCSbf/zk6QmQ3SWc9AiJjmM53Wq
2QLZv/9zCwgBo6JJIRyVyciRLEK6RzBj7uqEp4kXEIZC3ClNKEGYAd2R7JzaBoTVpablPQkKn5oS
AOklw3whovFOK9P14PXjOf2CWb8OUaZ+8fSPtL+0j+x6FFQ9W9HvDS5hhOzoG2aYAxcE4sWXy9NU
yYipxY1+Hd/P3MgiEZd4PV3rY1pi4r7V4qLFJ3VDA5eTxhGAin1+hdwfuy7O7KBOlhF3CThSTCmf
LPPZpKUVdiJQtwfzxM9oMyP4zYbNN8KUCZ1hex1Gr5ij2eQuKrJTvPYPmEUJ2wXpAnyfdly46mBy
ofK8Jqjhznemo1KvILOv3uwyNmUnexW/E423y+bYcUchHJSgLLQRI24qsjSUguDacvFYPZgt+lBE
pnpTNx7fjaYWIQELW0XOvKZQEcw3VYMojJmJpCXek+8lQCNCxbDqO4VhHaDdxk0W7OkWs9L5YBVf
Ek32L9LEEMDGz1PbhVdwPQ/X+s++LayLbcX8bwi8VIjBztuI3cHE6+cDxGBfj1wF38swIJHsy7y9
hZr8cxHlIRQ2TziSuWKkb/cO76OI2/qEb5h98FYWtJTeavSypq6FUZdIAwUlk6q+r4cIqPxf6VcO
Irq/EBa/YzVR9Mw0VUy7x56jng7ClRr1MUA/Mx/5ss/3ciTZOrIavA2BnyFf5ILcomzKQBUbmIaO
FXNxZFPrOFWnnN4N4X+NLssP4XRbffnjquVh35dvG1NQlEbjc5/WMq6723CS3zZBTCQJlAKZj0m2
IjCrCNUKn5ISHdzNHSEzTisg6/5dRIXbZiHvDRUnmksmVWa852eTCDk1KBDQ4dUs+sES6DN8/07G
HZIyxEFbfAKq4LrtINTYKz2BIL/vTO7uIlhlQVoYBARDYEjNizn/z+gEWsgT/8SOiEoBM1N8Zb0H
quaki84FR6xOlrRlz++aaA+SSD9JDRu4iZXO3Og6ZxTNAvzR6aUs6lFz8OranhvSybd8YLbjpXX2
B1GOZlOsAzMxTwT7AQlYmYJRLoOheXufuERCNALoK+KcKINdZGN7YAyeu9qmrcSYTmmOP3mlnWX2
KcDUCkQjh4hiSU70KJGSpnDdkcWh8dEPVFCzGtuDB7bhapzA/0iyCzsJKFVFLM/TUMjGWKedqFYN
vvksQTkBdof/XxyLmGxoN9j3gmTTb70BItT2w+GZLocD0wZCHijX62RcJ1wBIGKr2qvgFgu5Pea4
eBCT+HYlddDrGptIOKFz31FrbrTjOJ2B8rmEmIaSJfxSL8zI+9xW5gA6nUuQGtcmnq7HhT3r1mwa
VVjKhJRkT0msK+MlUQLs0GphNpgDplhb87Tv6bMdY87X6KpHaVt//x7BZxpd3rekPR9xFtUbTkpi
u6safe7MHt1VjUAJ8p6kPDEmR3xzIP56WvP+xfBWGw/gR5ISSOdaUl5db4gzOqtfnKtkdLtweulh
lzqeFWsizByF3IKJvVSkMBqXi++bpQ94sll9lG3/LpiKe2YA2E6f25DhspkyMkBYHDHNkV+PtmaJ
A5P0Jsx4YLWd/p/uOd/s6vq24PJmRHosjR17vPbm7p4n9xVWqR/rcu8C631DPuO5ZkypVrLHF/6M
Alg9ncF7QxsHdHNpM766wYA9NIVud0w/f1gYVjwM+11Q1pVKO0erzDb6Pr1qYXZHtsSM3yyNnQ2m
C/g4ptHJ2GlUzgAA/XAZBi2ubzO6LASYFM2qNBz0fc13/E9rXH5kA61f5meoXcXEYB4Jo7gT6NuF
M5ppyEOOc8QcukSf9rB4m6BrF3LzF9cqKrMs6VHK4gBo8rDyanTe2z5ZOixFwoHbud/x7EaxDk6S
KGTULumN0kCVqNwsnEi949atB7QQ9RfDiIwfAnQyAC5yFNbcn9h3zMCRgek0q607fJBeq3qc4vd+
RU7QdNt4eVAdAixjVwmRmAW30rkrK94e7zFUGgFvovLFEi0ZoytHHmYbyvId7LroD8+fyxb/DcYR
zomhrR0mrUn+WJ/dCJH6OLqZDqyG0YM3seEph2EB18cWBlXuLkYzrvVRtTakC4DEGFanhdpRj6zW
g2LFJ21b0TQrZ2xf0BBqlrFlnmAqnFkHApzO7bC7az4g5yMG5uuct6zBP7EhVFo62M9xpl2uQyB7
16heWRnjNOrl4xrEZ1AMEKAl1686bRJnxt4qJIOtiFGqqwDJ9SbY1ANqLqYJ7CavdfMWkBEPzj1E
7/CtRWcMu1gJ2uhb4BXnIIFFyShJ9DFN4iGUxvppFnwlzrgAfZ8Y8FmONj5tFJqw2j1TCLy8FDIA
UH9ec5R1KrEMXgrS39c+tuRhBJGqpAYfgdzpgDB+HfqdFRQA/GTEqSS2bfZ5kyz9LKZdrcU/Liqy
tKr5z2/Ds0Db551d5c89v9tDKEXcBUG32pRGP/p9WO1zHACJf9JyFXzkiWc76CRROSdZa0nMrNZn
vRB/NzjwFsSHbRRaAraHXhkrne1+t7e0HH1aFsiJzaDeQT7EsUZMmr7K1Si6FXpPtXeDpIq22C79
uR1PmZro9ueieVodmxbxBqcsxvNYKeZrB7aJB/LSknXEwgAkZ3ZBFja1BBLP2jDW5DQKKOB90DMC
BZJrAoZ2BtdZVNuejGie8xiHY7C9+I4HOyEAniY+vYEkle2y985+B1LDaS/TldQYsDNMTsJ/ryr0
+09AyjF/mDT1fnzAEFUMUoW5KVzODKlp8I6gVfuPZRKgJo9Y4eRhy3JgDZNiuleB81OBAgTDqUBE
TfLkaRPBivYSIxRd2qjxs+T7oBToI3cncG5DRkUycl+B+jMvUYA1VU3MYE9ncX/ZOzNhbec3bael
i4GbueDG1lu5ajAPnCg9RgBE3D8QwNGINHBtzRx1c/XioC/xmPoR8UtxLyDJbivRxcU9WPdBS9NO
r/NFh5FJ64p80BZilh8+HL+GtSZrsuTfigNHpd/l4asUz2pWpwVW/WlX4j6w7A4DZHm8txLMNHMO
nKJaoq3HTvMF+fCMibsKtPjBtFIFA770nAWV8A+Y3bPs3+QoMWeWlKYNyVa4gIlY74lEfkeF4QCn
ItY7Qv77HTZ7xznZzl/77szEOHcMfTj1i/UFSJyG48guexOxrPEYeFCgBN9uupCteXeDcBv9+rYd
XJ5BpXIezFEI5iYnEb8YpobrTNFa0tWkY1nznjqpg9qBY9AQlCpCn39yYz+NtyF6QqlEy835FE4p
vUmGxCwNwTUVTU9NwtbwWz7DXzjAs9k64Hfr03m0ZWGDO8z3YDxJcl7BN5EDDT79aYhn4+Cp7TYS
ZIaRw4aCXidN6KUPkU7H+YGBaCSR4iAa3qf2u0GXueI0xksCIAWqv18FolpjhlV/xhW5a8YBMvZf
24LGmSQLjHzc7MRNvLziSNIx9MiIFwvCKeyoEv3faVSoumIvdyILOQQMFk/FNeRYUuKwIuX1hdOc
xfV4dBHMIrth38peQfn3FsMqcqOmjSZYQ6LzCObv1TG++upZ/iknoKneQ+MmdAwgi6Y8yKAZAbRx
MH+rc6baC6lgFTYIw+7ACFctT/OBj53u3xQNhuY6E/yZVTDgZKkc62ZNOqDSy0q7IrTGcc7u6g47
cV8GlkIcoKFxnyekfD+fd1fGk7nktOHg4gYpr1yJ2nh5Bp/V7LV1z1GPcWx7KuevVaXI93Mcn0GM
xQCObZssGR6iravvgod7jBkH3JfiqUuq25IFq56CF392W71kS4HTa6MtKTvcXe2QQS1XNKAzaydd
vMNqBWnQmlHRBBTwWV79PBOxUKzN8RL3tVIWoRXzi4SFRmVx5cml4IgiTARUlmblVleyIUsaGst6
G1mHlKFUJ9oeNz5si2SQlrkZRhyNtcia2RvtWOQIEYKBraYd6gnxxcRPIDVa9QtJPuJIga+y8XgX
GdAm/ol2VcSxea4ITiX1+iKAcuoOBtSBmUCYuozD1U9UQEIYL6UylKMxNEh+yKijyXEeGmp6MRC6
RukuiAurq2gV9AaH8LIn05SVJRNDre/9NWehsPGScfBSM4wEe7j3/d5MRvTfgAOr2+q0DtZ3EmDG
UO0Gjf5MD2PgFicR0aVXB0Km8hO3FHGVW/hd6QOHQMzSfO3+Wbf4IecX/u0rSy9d0z1iILzMdxTN
7oLquG+9IFFOD6/FzCox1ce2trTAROUP5yJ2HK6u6eq+3uiqyfknwDZmeEhxnndRssgTYdMKZD6D
rZd2il81Bu3pS7wNK2gh1mXV8Sn5vYFVUs69Z/k8vuzgUWtIN1BOyp93jZR7Hf+yt0sShCSQh6kK
T9+u3aOge3tWcnh28BeZzzYGBfEDsUd9GD1JRAaocVkyLWU2QU60Mj1t1TEr2K/netb/Xx86f/G2
CPBAHlsnlEmHxdqSCHTtIzECp+UfBPm8gcwU7k5sHsR0DWWHM3VHk98SBYUDxUhmHGTvs7RBA56p
DdmhpqYX3bF6t3H9rybp3XT0H4haCeFVoLO0p/6+uGpzzY+ciuta/s87WHPjTHb+pUGr6N+D/9rx
WE2mqvEpaWJ66PIcNwtOfNcd0n0NP8FCtzdczLoGmV4BvWEBcUXyz0X4xbnqGoBXv4E4NjW0iK0E
aSEv1LCZMkcsWsD8L8F8T+NsbH5L+nmXsigjaU72i9rpDP+zzs0JT4pO/H88IpYsEd15vLwq6LON
5++1tY2jHQfE7qA+U9Wp7Dy8y0JjsMmbQtcWckLtTjNNFivnQTgaTeI5duKyaPPQLW6g7Y788b95
D238xrA4gAHWSDAIUJjRAk8xLyFU8Fsc3odwEPojf4e/P5NXkJtWHtvn43FQa7QUxFR+tOUf7p/c
cEDuMFkzYYvvvnAdGxrvxhcYhzYm6/72ZjfktCgm5AvVfjn6YnJwyFrc5MraohmGBlWJ2/LwCCZ6
DzddI2yGlUBZA5zqSW7FKVXYYoeH6nZ6cvQNzQ+tWfHEhhP3b0OKrx8U2zpCzGJraXdJLUXliRwU
9ZkDQf6pE8hcf51RjQysUxrVF6pn6y0lU8z+TAPOCgiw8WbfLYLqVHXKI5di2Aq6JCgQW2Wkvicd
jb9m+dgDpRLqQ1cQsoq4nKs1uYnk4stBQeQOuSACdq1hJ3/ljBhdYqogKuq+JE0pVrzBOFLfRseI
tfFPiMGjjqQZt/UAz3mo/x1ncPAoXm3PuJteOZ7U/6yFTYlXu0T8mGzwEyOwZAasFntvAi719SkJ
XAy5+WH85GgtnBOkmH//sQ7hD19hBuU9draftCiawvQgYOvbT7KyX/P/0Ag93lDMxf7gjmOHyTsl
FTetqf1Mf+mD6WC9dDgEEerKszVDty/MLm/Vje5NjCUZq2TEK5ve962PWFaJ3CRqYvZwqiVL6sNd
Twjm275bNsFN7MP2tux1oYGuOe6PSuR/S+51u4wDGCeMcpBiK5VlAdHJzj7pLnxkZ8k/yUn/la7J
asTcF2u209LiijmkUVlYK/tPDM8R9Dpea89yeXyc9daSfeFnVXmJR2RjZPLTAFSzVD9dydLpw4ZM
UQ51hx8g4moaMqFRxo/RhW/t92UwvIA18/HcR/bQl6QglV3mVHKHWSGMxJvURKQ9m5pw+3uhEUpf
kh6oeGlGuDzP001BymplyfzG/+OG+Uw3knkpwuHKXgOYr3gNHvwslj1iSdYhqILn2TgqJRb5Muz3
Xjv4pIQ/r/VJgr1Q3nmqKDOZkhBLyTm8yY6IOvZA4DqCK7mWyEu2NCY3MFG6ku6xokADEoWbGixF
xglXleC8W/JcQr7EANMeovHFvvdBjgQ++G4TUp0V+1J1hAt/jCDd4xkaeupbkiRM4iZPV6ZEHkTZ
QN8I1pTLIqaPYlNsDICHV3vbHpk7AtUcIy5SAjNuhUcvMr+Jh2+nAI1BcCHFNo68nWFsJ7SE+JUt
rtMNQMYV+gsFz87dGoLVBjSqkj3O9slLK/AkOsiE/BhfKuTJlGIYa0il9Vmj+LkPOblh/gb2gMoV
hhM5A5MV8IxMszyO/wIwY4/m1IM4u/YwgPqMJ7UJ9wktAaBcEqe/IMtclT3d1ysYg76jk4wH6NcC
21e6WlbJJwXmswu3OY1w9eYKMvSeTqiLsdw7k111eUMyyJdiezeBq3O7TD9BX7kJrVIxw21WWiUv
Cut9DyjFoN3cVdCSHwaIBK1jWCyVco1ACm3tdhod8A8kGsh8B0qt/OfjpH7x3TT0shhTYtuoesrP
/35HuQ+dYbu9fvbti8hoA5V+ovFPZd/G99JN9RL1ckmbkAJTVhCH9IiX4Kupekbin7Ns2+4ZmNro
qI5f5bTOemXEYf+8H8dd55LweRY+IBeBeViQW0UJt+gq9pfIZiwBS3RFsoiUQdjrm8Fb5pLlJZun
1hV/xHqGA3sr8I75hnJ2C7nau/ZPsuPga9DCZ4JSkW+z96a4C5CV9fXOAvfiOzVxCJurRGXYDjXO
FDtoGqdvglDLnAnb5ylccDILCrK5whg2CPC4HqCMSUfRO45Au6KW/PIquGkD2aM0Cuorhf4JcDRz
ccgS7B/1wFa1/iI0+IvDvRnNnwpbso7o8X6zYhRjsZhA9XeHkM3Ay2FzbWVrQwzsHPhuU2vyqJWQ
ZKKxj1S7G8V4SDrRjKESBepInnFHQBkX5vXna2SHZ4+OxXA7oiBjBtMyKN8ixU7MJmaAL+Bhzp5p
RobbGQnvK9WtF+mZjOSwY+tI1uNfv3zwn2IYkEFYqeVATk4P/VtCVs08Riaa2PkagJRjsc3+xQkk
x8i5IKB4L3Zm5puaD9QebvRvnnXoGtd6O4qJ9MnZFZSeKp1tRZDnHkpianLhk/EqcNvjq6TO3AiQ
Gf/0C9jyMt/E0teRx5ou3nfhwbHR7LJy7q8F+lLHeoQbxLNpVlLvA5zT4kAtjiOrw+DyFdfQNgC+
fHHQ4we2ooZerU807e37Zzd/R2i/Yd1RRYMQCvVSWGlYoePcE3UWbaESYhRokfOfNBO6Vk1CLslw
ugOBJBCUuJEF2KPAMzt5ge6gjy4YXuikYZaNcbURQKDftQL4ypYPCTXkp07Xaf5d89JBIak4mz3F
EcGyv+3CPqxOaQEly23bEClnPuTBt+4IDLROHmY550RJXknMSjonu6K5QmCwzxFmwdpRBhTgBAK2
uRGInre5M+bW98EtUZl/KFyeyl2C7+zIiKtur5nbd5zT9qMw5DhLpRi6WiSuheBroYCoc4OjGy7+
wIE5AHvQKbjlue9UEZ5t5GaiXZQvOWiJ1e9OB9S1aPwOk6WYPYTDSDkSdcEPIZxluTkqdZYTC2Vp
mOYVJMevFWISuicPFfUlvYRSThAa3sDLcCCahHfl0k4Duv8BwLWi9sCmTdzZe7dyW+diMfdoIfrD
oBbS+oDuMIcGFiZLiVb6N8bBAoNpBGJOeYtnUFrPOfCvNSk2H2P1ALYJRafTw/p0kSEA66LYRDJ1
eEejHm6Ed/R/IGV0XoMXh1K0hWB3J7r+FJc6SVHrXpzDceGAO49/SnLJlvvAb5eBUmtUb30gQSi8
xq6a9iziyx9UaRtnr+EsT9R4OvxJAwWiWkIW94J03t7oSAo55BFjHNuz+JmrlYyZFoj/S8d4F8zF
2YVT7BrZPMtGak+SSugZ2LizHXFyty3liG0uefuk2MvdXvZQS+kbONZ4wnIcWtFpe5tkV0hI3Bf6
Y14rTRB1uZwb7H+pO9Yak59UOXhA9DqoXtRwm25m2QnzUkPQeHyywZqfeHXeQM/V2mPQDHJvN2Pw
Yn2pq5J8QziI6/ldpBR/gUX6m0l8IGL7h1n4r3VN7Mz9jmgJjjTrnNueAvnLVM9shc1EqvSQr145
TlpXaI8rm0/r9JcgK8SALMarLKpWNQoKsEvGv3ngt9gtC1r5ul/exubhOa/i+gxkbivAQnzE3+7c
fxv6HhY9U3rqra7zhasz/r9/BGx48zwVvGw4XvwDZaLfg7g50zJj8ExQsOowPYKfQZ+WSJNjklU+
i7LBUa22FEyKgUxiLYGyYLTf4cnxc+7RvLYYejfLJztzO8PKln8QD9XSLcqqyFmf6d5eu+3yULXt
hN4lM+Sg6Q6w3XhLOEF4urLMD/nGIXHl0CzVE4e1bwwLbuSH26V4vZRNSY2J6oo6C2v+zDlclgl/
qDnResmvRDvPIspiQR5ZIMXMQ007bX0bOJ5VdjQVtYbQumDsJmMxLUwrWky8FCLuHnjw/RVY4+iL
y0edvcNZ0ZNvw9BzUiYtvaoPjro8ba1vvmnXgeYgeqionypeFeCNBbKVsWsJ0JpxzG8OquuVxfL/
YmFHF0SpktTDoTtSVh5YIj4cGS1UPYLjIWs8fIlaRtC9FTivnmJAZ/UhRmRlNgznI095/FIU+0MH
o13VyWJFL5sue0xEnyVqdw+h0om8z8cn6Kitt162qlGGVNJiNNrOxOv9NbIS+57ncqF2ckPu7boW
C4QmQ5kPreCMG5/emWBjVKK/DYILnPnKKCKGkkkdtumiEdj5I4mDKYo7H943W3GEaiaqsyM8eUE3
cS5u3Oj8DwJIgvqDuVzvw7hyNo1f6DmJOcXUmuIPFMtUun4K7EQPAREdT3K0tEv1gfT2JYFdIlrn
qmIUBSGD/vAh8Z7YvLKT8o58sWdRkAoZHJ5uPvojaMjmUArm/mNFW84ZhZzSly+vK217oKM6pqXb
MjB1gILWMZMv5lAgS+VdSxAv7lgdJM5AYE3Quas03plZCx6uVQujwgnrWynLg39lLly4J9hRO0eb
YGCt2IOK7b4b5LKDyrvm+ksI7EZnheT3s0uvSllghdEXpTJdn1yWKVVCRGS5Cq3TI27X7kd0ptMm
d8QIszz0mmzuAZZGuej9Bl3b6MSH+uDplRDLxQkVsBVs4EhxmX4CO/pxWG73jJ0DIllvXP5vP6yT
y8oTEvLIXA89A0W67a3NL2DuFzUxGv+fny8Zp52q6Xf7Tbj1f0wmnAHiK3eSdP8pSdLqPGOMq1Qy
23i0PxhAUdjUpbQltVKyISzTD1anXmts4UOzu+1KXd9Kte6FLJ2D844qDVO8y6tMzfnNRiDxS1qp
wwCoIlSDOy6Kk24IMkW9lxWGAlkFu4ZxxCyprMes7QnlpbsvZ5ywDZMcxCtJaZ3rNzqiG1rUEnLB
ogP30Tnd3wE1tt0V2I8SRpxLYJrc243gSwtXoMY2a/SteBThSst4zMdTixlLbX6C7hBGJbOilgkR
wpsHNEABICMUE1Ys36+LepQMIuzRP/KugrI6ppoAsw6LhFTcIYyVC0jDvBv26rBNXOa4xaMQuMuY
mzwujYtICZqUIbPpzbkkKmlMWX8mXXR0JQ/aeh7zfAcpo6u282zPyL8hQeieCG+4nDN1dTQqCBnh
B+6c8lRsBH1NSN8Xm1CwsQ8fJg0p/xotRG4u/6KCzxz2gFrUHljZUDCbU3F7Gbv99MyydwvAwTUS
liHCC6W3WmsvNRfxPl50E8WJ1dLDiY7TvosNmo0YKzH12RMabGNl3PIixGFZeZZ03Z7lRr2WqIVP
xYJ2eHnFtAZG9480R5/po7/W3cIxHzRP6Srs09iF+kzBUKPysEYHTo3+BfY1mv77uUrxbdshoZkA
c2l8r+09oTkyV03Sna0w/LQ1G+SGKFLshQLnY2y3ejSYQKBGXWJ49HkehQa3tON5LdrMsHGHwbtI
mELLe2Xz10Z2lEVJI6hk5DNFWZWQsEhrVOFi4HENG3Ghtuw4ct063OFQ1r+vhee++vFgahs09Qae
1eFpOPYZci4s8GiR5/kJN/D1PbG5wl1rnWrqZmvzZ4GFEifp6Y7SyZ9VUtGpDI8gaFWqY5qmgtJb
ROlp9Jt6sDTfRLYh/hQ2dCbZcVCRNUjIw4lYEKr0JWYYUu9i2d2e8RsPVhpNimELyfxo9uNvF7wa
bgLk/7yRSg5pOTQAE77/851k86F72Bx3Dr2CKYCcF8QGU1IJBRMCZdyi3ZJLjdvJYvFtMOcjVVIs
s1K2wbzPd0PhZ1bBpMt1Tlg/A/pvm3ujCXPa7lxZkrxK7qs4t3gGzM+e+iI4q7M6Bouymv3ostXE
l/1TQClQ5aQiU/IKR+2vV+dN/a2xPW9kmayCsTbgTx8x350mQqUb68E0YVWjt3lUx8hNXw+OA/MI
oKXHoIZUXgQhJDbHWE7Ztpx1X58PvRMIiWf2/Q/4kwZm/1Uc8nq0iexVeUrFe7totGk51MqNfuDf
Yu+Liu81OARmWI+CXI5sGmcPC1FkJmUI6iVXD2es+wNGjf/6N4wONQbAbWQ7Qyz2KTHPr8uh9l8z
azL36veLqbvIw850/6VPJZket2hIGorP/AwgTrsD8E/ms/thHS11FIJdHRjS3XsOPy7/N2lSA56x
3aVdht7jKOR31s7yvhw5gWA2UgebY7OR0D9CbfLbZRiBDY6TYkIngUHP31cafD4tunkmNLtZQJUZ
u3V11+tpG12hYY1zm/YOtDjIe0rAoo97LmXfEHOueE2tpYJVyeCEK1raJJqaf/+fZaw/NeMj4XmV
4jVkZ5o3QOenQnj+BLVDaGrCFrwYyFawQf8k4KkrwNaGr/0jM58VBxir7Qp/sQtYlsRXN9RVk3Em
KBluwUSkQndcCWCikl3lEUfu7ZAIDzOE84/yQw/92y/QlbAsbN95eayJ5pOUW7ssbcrUO9ki/0t5
YF5YIQO/0gjyHRO8sZHdCCskr8Kd5YFvFa0Lt4UARtoKc2zsHPlSJR3fYN1Q1SyOV6KkRFbXMTTy
Nfx+e8n3pHuE0ScDK0Q6NOLzQGYcuOPPPc0YGvfczUICunxU5Flnk649ti7DwTTaL+p5GSMdZqRJ
iSJcpRsjz1QJGUoOBRekKWGZ46goBcG/p4ubG8BjaLv0m+0GunFqR+JFwFDjUQ4JSlLxaeUvYVEF
QApwnFs6g8u/BLtzRW4mYnbp8HTtyMPSIAUmkCFlIACRCrDl8H9nb+H2NN3Oq6OVtbjDHFByWRXH
/l/p4nz3Dy4wOx4usFvZxD92QPBt2bQck3/i3bC3+TQWc6r0DO0V2TdghzAYOw1chkdumgh/yHtv
tocpu0n+pAw74AmNOcOC+0MJ50Uj5WEmGb+rkVkJCyVNiQoIfA6xdgOMJzG9mB9PYI/GkFQ7Fs1Z
oPVSN0BS3w7um2ZnDhrXpENxSkBCiIpV7M/NFYlX/jNgpP3Ohj17+uyafPHlRxtAXs+Pgywseinq
HRt7C+JaeYzb9r3MkUZzwQXoPcjq3SnxZbmGUeFJ6pQ69jJ78w9aa+nYniech908je9CBJDJ0kqd
grV24yPJ5uX/Hc9vSOA4WaM2AStmgJyGuwvilUJAp+vobfx/hjQamH3aM6ImRtpufu55wjlZ9d/N
jgxfMBQpzVuOkCqPtXKk7I7h7u+undZt/+AMRCzV8mYWtp2dTDvxQfDLVVppPkO5fNZU9YJ4nafW
2weohDAUO/Du5JIqu5Rb8FA+bxUTHF6xrxPFhbuhBztMV67KFLtQmj5pCQo9kYYzYV+GCk97nvRj
cOGeCMBoIN63hOuDBaDysdyqb9HeABFLzoyC+VteGJITgDxceyPmrixjTMgWtvXbK9MdtugkSQp+
2suwSgpowqSt/B2m0jalU8ml0BJ0dzhqda0SjTN8qNKf6CjHaRSVLuDbV0gVcDbmuuy46uudLy5q
XaRqpmUG0Up0XIdTwlhBKQhRdoyXEeadmmYL5stZJrswcQwLgqb23fyg+Pr1a6cX1TNFQyBp0LBt
SYVuVrSHFnt4HkVcDBmskRYwMFXwbh4ewHiObsm5ifCUg8+Vs+pe2Jiu9E+etjrxcUqw2W1kknwZ
Y7RBO8sM18CK+Resp8q7R14ig67GvDILt6K1d9i9DS3Vvx7HE6YOK2O2+efrIgc+TAj3Ww2dh41C
lLW4Dhr0dLwA1nEGj/CUmYrG8m+waWoo6ZfV4gYqFls8qjpTXW+AJbKDLoI4Dv34LuHRBs43ID1O
lIMt/sjKJ8z+jUzJzyBXEh2/+S5PChfg0wevCP1zSLvXW/1Gv1ynyQmKiytPBmAycL0nCyx99JKC
wBp4CBCPvbHrmF5ZivU59uG8bGJBy/Ggdbd0Sb9uoO8jtbKBWSTJ6r3Rg74DfGthMZZp4abuZokf
42cg0+EkcUMbPhJJsT1cPFrzYgSFWC5eD3wVykDt7twQqxyIjCSA+l2nDBf7rG/pmrJoQGGYtc/M
8C/eTlkRC4O+lxDTBgndiMbPEauYmNdj3Bs8G4KTYgVnpUNkHoyvRhOV4I59gmgM6ZUFVi+JLAMm
6keR35U3E5yXiYla9XLbsl6mjzVc6QAeLvxNM8I1DUcIifYTSnTmrb3Sx1YoZYMyUHSfx9/hYwLZ
s9rBiENFUNgyIo4sFLMuC15AdaI6juNy++BWxNhxhT7D/IR4OOwe7KaRFNOW9nHZlUivmFxrhHQD
WZKHwF2yFarDkAuM+7eZzVkp0rNJ4BqkM4T/UTwG63uLdKKaGqR/qw2XIu8+9iRomwvmP4IwYw7w
28xPnTC25KN2AL4BoKNLjsovZJU+NwKsvq+K3GKVNFcQYrcyay3V1vpN7gNXXJ8cEATy+rXXA7x8
20H2HSqZ8/BtmjMb8GweOX4UkyTZ2KOWZ29CF66I0JYcfYKaJDspbpX0Y4OsL2Z+JAL5T5JV9KQb
/49ypSOahW0nXBgl7fVajl2t9/1+P6696NDAqTkF5kcBLPPWLwW93E+wEmzEKZ457SLJ/0c7zxVz
/2FgxPhigRsUQwJhA6hzUdoSXausVjzdPrNpr5/wsGh3KwQS/0/WB1FnrRGwm1PMC7YK19BFKDa2
JQB0fEPUDlQADXauglu37LE+8rNmNuX/g7pDNgUmcZQjYJumdHmbjkJYSvae56cQi92Jc2zXUsg1
nI8x+AkL+Jx/Gl8MiWWSFF1LhxQxmW7xzAfBksCQwHVi7aZwLnUKHuOomTjaXfow47MBq2ENVSF/
jodLN5zxGXe9yaM07suJzIIoj5U6ChwSLdRe7SJDifziO0wkuE9t0TfM6H+meAkprPG9U7ZZV5gY
k+ThnhYlIVISsTHoRRx0xiESI+AZ228PD1RccWERzFGlSZLrEmco+BMFdcGgZKN6/4Ad0ZXRp693
BdXO38nFRfI67YbUtrrJ+FeX2+RGesVRWjX8krpIVSWWGnqfZ3mTutCbniJCrkEqe3q0fAUm/Soy
4rM6TfnSTN0OnGFyPmGmcdgz+PM0PxOwdw8IOkIJQ7kIsHObZI6MaUrA7K1xc+vvy9TXmSyTe3Vq
/RgvKYbBhKtNkKzV2nS/KERD7hAqTCpIycH+yGCV49xEpq7ubSpXse+2Ma+/NT5qspSCmkJ12zUu
teAD7sWtvbBZv8fkpkTh1Cgu9+34rGQ9B6/TYvuAQlRbz7APLvJe7JRAe7cjO5hOwldpHWtUwA6E
UWW64I/n8NaH6CNbwSXOzvcZyWeGhhEQsoNzlU5tCiMZX/3B4JNggcK/ADfzEvFjvASI89Jljyjv
13QfyPr63kga4vpsZ94+apcQ2G6kfVnOx98PBXuYfKgnNbIZEPbG9os8BVROpk2JU7Gl9x8EM5v8
L5itJhZ4ab0p+lbW/1b84Atz0zTuwKoNfkCxjenwIQK+BnPrBl9MlVptXhQRR1yodAhpAFOuM1p6
2gT0MQqPNMoYJ+APQIHEUAjwgaylOk8YJC65l3caR8unL5AP0GGA1fSUlr1j5rDoX9H/dBHBQrly
BcasvUpiVeqg3gl6rw2e9fzHQVAG1X0Qkk+rY64o+f+DeaEDdyOI5foxPvpN/RUAFbWfhClcDaOs
aJXTYx1hqV0Do1v7zD9jvFCDYWVlCqTonhGWjqQ+NTohKwEON39d536pyEWz7tDJjjokY+abhesV
Ejcmr78kheDsXOs9SyDXsLaV9px7e4E2E81WMgsTS5BRb2KXLvAiqXc+8WoNcWSa3n6RX3w=
`protect end_protected


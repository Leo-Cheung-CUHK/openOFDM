

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
R80NnScBgIZD14acGTeYZyZzlDoMDRJH97QvrM1z3/BPxjYOI5xO+RmLRE3ogivikKxeQqDB3hYo
CtT6MXJE8w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pzFf5UkhQCihEthT9/vXIu9qyyEco3ugn72RSG7p68vod9TXq7nS9azLrnGkzXHs3PQFBkq+3+ZG
PNN41vDN58/lK8pIjiAlp2V0xXr8ZRf/QoS3nU9pnZ3CEwxt9CGwUMks2MBnm+VSjWWRxbkUaTxZ
+kjzVWvQpUuyFFsOEs8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xDcafb3KrEW7vk1Eyiww/9CKbzlKF9C0uKrVBz5bHy5+6GMNsnwfCSkgxU14+VriR3jhdDN7viwB
M3a2pKPouTEOz066rknyw5X/sQ4hniBD3iUl4NQWkHTGym3kv31ZUeZYdl5ODPvzfUJOWUvkAXp/
gf4rtgV5FBbGm8qJS4jxuFSsv4rhcb7t+cae5sULvX9h7Uh0lEoAlNX3YmEW0fWj4bhIgTdzT2gk
C1ytdGU/UAnitwmujc/k+32KWV0i/o3dHRhIc31iawLLSmuBJYefDEaLG6KE8nGHeuho45Se0dhe
7kIaZp4SW1wGf7C0xxqwh1cgZ7+6eWgYBqVY1g==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OrzITnToGC+ryHZVkpDHCj6CgE4vEVrPZ7Z829783FsE2zjugDCdpipuFZ7ikbeX4Bc52TEJ4mFm
0OxylPcCXPIE74pJ186gBXkmldW4bGFMhTmUHJ94bRAsyJjr329fm+j77y2NmfbHMVOsljahWWK4
OMppytgOrZcnsnsORsbXvvikZALiCB2t+Qc4RdHc3/98o+DDvRf+gwTZNX0GMOitJmVVvqxqw6No
K3aHL26WS+5291/TUz7aF7ySSp+k84h+0omwPrcy0Xc3URWaoYbqLrWiEi22RgQYitI1tEsa+afh
tv3h9WNr+65gWTbdbwWyOz1NeXJSaNV/mc+/Lg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
riYGAyaVfIXieMgcJVFsucQ9kUNBkyzgx5CLlDibSmqSJjCaDvK63ymwoZpsGDT9Rugub8H1Y8xX
XUpLlzZGCXrlWs6NgjXfNxVpLlkmz7GswYkQ6KhUkZhRuPh0HrpJPt1ne+1pTM6fzi5LXsyTv6sn
TisWpJPdsnmBDHgM6jupb4Iv3OG7/q/NPck9K59oFLN+AyKeQ/8pEy2j7xpMiFTRlE1OTJj2mjHF
yWQWyURMafr1KK5t9Wu7YuocfKiTo0f6okHNafEo/nNpObW1D/liUJlS5GVguNNbnFjSuun9SM4T
MXhUoU0rVPqSkeCGnTpMMYK0MY5IwmbyZXn/fQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HyAIbEI1uxEAA90t6+VWFTmyUje1JDZQZoMv6A5VyFWA8tJ80b/Pwhc93aHby8xZos0WjlEANrxF
3hJ/l8XJYMVZWlVytBIRAZYGbhnMBOGo/5sjE6O2Ap0308iwfA50rb1ZITdKRqNiW+PlWkaGC+3R
QMUfNUa7cSm841V7mmc=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GUEL70ZQ78wO25wq2V+5JNZcUKzj485nYHAlIxulC+dFYZ1T3bS7X0juNGn/cdIyRbeWgA5z1viA
KyiSR064Z0BmWFsIYHfLEP1CENE6B/DkEgUM//4pBnGxH0CUe8wWHQBcyJQAxQHemECYQ5/QfTqT
96OTv0jwZ8yRjX1vKXS1qZKREGwNAsV3Kgrd9M5oaNz3PuISlyOOLoxPx9Qvu0Z0QYAzZbksLAI6
oekHTbR7CXs/P7+GCnbyf0lD6RFUyKASz8PAAvPi/+knG0A5BGQv9W8rEQ1GlCyJMbWqS7UMYIM5
Aany0Gd6zUtHqzCJMTpR0Gv6o8IS9bMCD8CICQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 125824)
`protect data_block
Va+mEYC1J7Xfs1eMBxJQx+vDVjiHrCZAfyNdSOhbSjfRTsOUfy1BFtYEwiOa05CI7x6z2O3XB1hL
PUX+3vEcYRDwUW0v52Ft1Q+qVwY3nQGHwmNTHP8pr9XNGIGr1an0x76KzztMyA8lcCDFBubTBWPm
4AhhQ5xICxIiP6pI1zR7tYZoOryMDuf9s4afAATvW4Qg0k+9KVmihDS45A4LpJZRfeW1n8Em6GcU
Y4b4LdZ7LdcaLBKyOxOskIG04f3NZ6mGcvQ4t/hvaTC/+4+df42mWUamwgVmawp+NKCIMqF/5G6X
7mtYrzkZQ1x9YExZn/n7fdXtWqJZQR8b4GehEZLXONH3LvrS04kvT45WnNL+cd7NDCjhMca9Vh3J
42zx05hYABup+tpTHelIg/dDokbrdXD96Vl6aTAzpoiibNKYVeJi+HBe4CE/L0ZNxyzmlg90gJJe
NYTh7S0gmvMfySaJQejNxjwq1kyeHS+MxiMV2ZOzxjPagc8pF2hIpWmjfD8V8B+kOUwSUxlZUisV
Lzld3vPX0V+g1rM9Wx9IfkzF5KLBuxaetBibZIb5w9FCdFe1X+w4jarT8JNs59VTfqkutyLyHHcC
XxgPqlAclgoWu+f9uN2xsRIV9KNOqwB/HLB6OrFOj7kbW2FXe5BecMzGQ5qAZeKevL8du3QuVxUt
HoWy++myBdQk05kxaio3eBjHQv8TpniBEwpzYEH0oe4ayE4h2wCeuANmyDRxk82du8yBV+xa6jmQ
LQBPsK9Y+YMf4JpjVAKXDWTYZJzZFdbYIkfgNUUrHpm88syXgzATBDuMlqX+bTW8qr7xiqr+E6yn
yObOEGcn7RFIjEhUF1LNZdjkviLC6DADRMR93knVoJ92CSCaq8/Vi3U4h0UK1t8xSS7IoQpcZn9P
9vprUiOusCf4HYb5MPLxjHaEMOKKEC9WkuqqAaTtX3QIBy8At3ET2TcEk4WtyOVvUNFNENuYcCpY
RN6CTDi12FWOhG90Sx1CLpeF3v9unKnwj/BBdlC97Et2Fz0Ay4YoaeVTzl80zTI30uMS1JRSo+2C
Q3eBDIC3Ii8jjzyHaN/XjXml09RuCkx0BSofnns770SDyxNZ0+kJKSI3D8o3Fqd36U0K0GFD03eR
QGAr0UiSXBrZViCUIC/IN1t6Ucr51lonOZet0toE/cX75+RdQF4gfcZ60xnM88WFUhkVLXDa7nbF
eRxRXRLgIiL/mcMSB2k6+7pPlFLz5P+x5B1JSg51HKZOuhlinXthGktxvKzaqaq16huuSbeNkINk
SYd4pT3jogdN4q9QXwt4P0IMYjk8fHZY+5y8kUC0PwglEGQnyYpOZuCOK4SbsmwFXBWN8+s3G/2E
YziM4CzDmWIDmnD5c+PDe3YQYfaUB8QkSULN7xjhj2bTPlOlgStKKf38Ha98yONPN3a1iOyXKavh
lhdni7+OAj8SpDPBSDWU/HNwouDPa4Taapib+6SO2lNEKhiWJ81cwwvY0qdJpy1Lg2+DmgDtIx0/
JMJJbMLmwvBXO185Z9CbYNHMAzeRmENbDlTaHtRgvVg7gFgeRwPfJQmWHxSUCzpSUSkFvxNSNcnm
JYSDm/m8Nnh56GAuxhfXCgGDuHCtrsxyAURx+ISOnReBvAnxwhww6DgrMpiea20VGrcKtM3/E2E2
0JmyA4FYk13iSu+0JHlxiJhWhp4eTD6Sl7RYq/T8szEo6sh+hYpn0jd2+zVOkREyLgT1Bqoxe9oU
RTa+/FZvNZMo3t91Q3pZaP0Hpop9+jRVVUvqxuoVtXdd22KIvoyW8v5oyDE8pJtI84CRy8RS8FqV
X5zFuG7GVRtyZo68/kU2A0CxjEzUCGcmF6t0/JmX0pyp/yql0wnigIWfS3OtP/l+3hGYgegXUuWd
+Mp6mCET4ggwVhZ4Ky3RDw9q0zJY0OtA5xbRqMqG9xDb13rPuL6AUuZmpurWzP59Qz6yemiCyaSd
ck3qdmhjmEJAwIBsHzz8dXsl6/X80hFZdVl3M5QBNUFyzPrDoJIYHnWO0OSoLD72SQ2weU9hx3SC
j0/9siZZAL5TxrnBa5WnAsK6S/EMxNi0oZxOwBKksuxUHhPjuX7ZrpzJ87o4qSg8JdICq56Pw4wK
Z+cbx+RF62hATL3b1S2UrzhYz522WOIjk+7h8HIubbbA7PE/4ACTuP/lcZfT99OJkmKClih/P1mr
shlzZz9PGTaT4x1EnSe6of0tUFPAFgW7JkGerLdpoV2aA/YDXzWIaT7GIU2w6IARS7HsWPKc/wlO
aRiInDglDqZXKoK6hkTnjhnLofqDePO+JhteJuDIiHlfKyOXMpmzCaeQog9RheWNOpwCmemMnv9F
Rv82lrn1gJ343Purwj5373t47Tm0QXIFtrUIbAFxfjrH4Wj/clD8nKj15D+vobR2NXPqvCe1h0lb
1fQqbr+E4qdYFEvGiXhy+8eL4C2yeyAjXSu5xsVS8KoyJFE/QmRU72RGwYZrtYyxkUOt1zc3izMR
xk8RXErqZjlZtc68BbgnMQXvZ9rYXkSGQFieHq879uiCGbDFvMDVI167dxngbCiCjJunPfiBOtWT
5szGD6MeOCRRCdefKM+CabsBY4GW4tESNXXCKmMnPJeK40b0XwzwQIlSChTe8QzYllqfU7hVpaSB
404BNtiZeNQXXQ2Y4xOZtijCYlM/EIMB+xmrXuOLoQXly/99N0Ybt91NHx5bXNwsJIw0S1ERtYET
YkGFzaMJneNLTAW+H28hOUWMYP4R1Ggqo6QARFHNh8CE1aVSrE5aHieUymQblisNrjkPve/sLwiG
kx/a42tUvfmr75wdjMSXWCfMjJzjKaefaRWtNflBiEGvJFihyn58FtVpBgznm+fUA6jpaaMF9J2F
L2wYpOB+P3HRHkFgM6gYu9LjZdFfLFGOfUoYL+2Ok30nrLJkdXEyGVn28HTf5rvS7VQ6IapmE2K7
ewv2b4eXU/vCsQ8YC2zHR1p66P0dAr8iklcz7FKV6wnElrTzERcXwU8qP13P4vbpmBk/ZCVjK5Dk
WvtQBn7ad3sFlL9zZ1Y0xINm7hZlP+oqpuXuDMm/blT5EkgFPTrd8CmNYh5uurox6MNIc4h4496Z
HCViBJjl00/2QsUWIO+3dxk/fUD+0UpcYrou7+kbgcaI5cMN82mexMmrczLRZYrVTNv4Tm84wIYe
o1iCCNBAMob75Zn+luRe4xvGFKAre+atCS2mxuSQx7S6ar6QGKvVFWE8bPydmrLlY9gAIAc1r4Ji
vZaqryyLVlTIScYLedqqkQIPK9CKnxq2hyxSGXc0988U8c0RNfr3np03wVZjfOkHjMBejazmDzeF
GTGIkcJ4921/jLegkRWsNP6d8D3FN7mPXhtZh/KjZe2LBH5jvQIR9WnPi/o+YCRU0uiJaqtjxVZP
funcBotYwd4fKnVnht10mdt5HjQ7fmXrZQvqrDBqYSXaBBJPHGNfiZL/khna57wIAesP32sLLjTW
IuAlRDe/NJXJ50naoeoIXExOm0Iq/nOSdY1YrhPXboLJpcMdBY90jUsGCkJwypivTM4472ma+jrq
uwh0NtrIOOy7cCCvILOoehA0QaEJ79citLFYN2w/ES7YxrwYFre6iWSTNlPDy2oaWZ6oIZ5FwrOI
TAO2OsFX/mG6UK/ikeXtcRxOnZoF/4Y3f6adPUj+IUky0Qlkh1iLa2b6tdXL6eWvwA5AeA3PGzwi
5ACsp18G77x08O6RZw9e40xCkZcUw0pzI5Y7246ncFh7MhCQCeJuUxfQGg/P07Bul52yH7dV0KMF
8xROGTvE4BbhUOjypRtKUkBmnaeaxP0KrnsKEitrJ2L79+tbalC2z18+gojy3mnEA4CMS9JzsaEA
wda+vEppB/wPeC3X3G26gQqU0sCvg6M1Hq8PBHaq+k+0V8QlXfaiZX/DvntrVqJPGq4KQpfB+kWD
k7rzZjTLuSr2MnlSKkwrSrkxd9ioRQ3mWHBA5jXaY7yjvrIMVIVxTWK+1s20T/9Nw/68F6Uw3cuS
JF3f6wB8P4hedP7coMHWwbQIcsNV3INKgJMWJCdmsBM4n9JVKYwygDoQkNwFFRnFzcgGqTpgwJYc
rH7wEJa/4NhPwyK9dwkfL1YPsTnJ4c7XE6l4la/P64ixebO1XWV83mTQm0GtYdkEWNagpz1BKTxQ
N0bA1zpF5OUTUPSszhTuOi/RHi7wOGabry6hMcsmAyAJTNKEu41EWDu9snDB7fT3lvR3nZGzVr3Z
ZDtEA6DRuFmR6Sw1NYu6Zw/OWIaY/hjCIc8cPeWBiNUZ34nWguveqG466RwniqRlWXT5j+EE/aIv
8dg+HNUkiZXrhJ7yIKZyi1N2ulGHrhzLL3emxtxW0lhn5cnM5VaSIoec66X2n5rELxws/Vbh/ETX
HeyrCoJNoYU7reV6rCExpJ0GoHRpB0qnq45Lhrr54K2NZhALQiyokVF/E1SGcQtP9Y+ISciScLKH
N9dcqUgMbryuincQX9j1D4TVFon1IDqNnLzEMOJGIZfcP7a1arHlUstSR1gTyfXMfIbBKsX5Gt82
zFvjpQBlML4lI4XeVEX5ynYI/ffbMDxS7mbvbuxyHVsn41JeDqtbUi84sES7brsILjpvi+ucq4TP
sG7rrutjkEYlvwYMHUO6n/KHvaKOWD2Anb+xtpfpUWXRG1njfLEBuvMMitgffYxY+1AYyVz7KMPx
ZV0L85/o8CrIlw2XWcRIYeVhmQl/6V5xJbuDl0FqwtWPtgGN8M7q9itrub5WR0jPTXXTQysOmSMp
kFtDDDTXbPe+WPjf13g7f4oz5/tQ0vAup/aKD1CLyy+ROj3gyoSy7G5AmIPoolmMteVnUOrjZiTn
3Bx0ufLouFIlYwFN8aLEokT5mVb35KGKkDyXDBXdxJehuoBYuu9Nl8pHd1i88srzLCWQOy0bR7qj
3s9Ly4GaO1nnDhjuxDtRXg/9evD+oXCbykyHOja+JrylygvI/6UbCW7j65hA+ZBdLbmZ/BCoSInj
xCz8oQ6yQLVSUqsy1nKhUpwtFZPsLSO5fZ/f1Vy8bxhWfXmum6mfvg59CQaUkBhO7fsFi6rU6PJn
CZEf11608X6WDNT3sC1z/itnxEkvAXV3e1QxCEqQABDEZhJdT8T4IUVfzEinzyd9+Yx/3NeJeNdF
Kzu60aMCGF2TrBbj9RGSx6b5DjduNaY7dQswSXX5sFPzFWaq+flTjmbpZshj96NaauSDpsaXDCpX
0xGqOUNoOcLqpjtivkbD+fmAYOVxPfxasybeplWPUnE7RUPz6XEhmjK+pZXKQBf7QQBe/WKKFhOU
1nFG3vT1bpfZ2/QAOxvnS+cj637Vf388RH/FjEKrgah4SAqMHMyZBXrJXH2pclFyzsKfI+vXT1BG
NkWwBCqzaeeOXYeRPt8dJ5Bb60OUwOj24oMiHGc98NwYfyqTNnJDvXFT+MNTn/Nus2Sa/BvCKQzw
wa7iTe7xNTx9JgQgMGaOVZ/rNIv3oYUpJPk78cQhONaKCcfRI86Qn4ykwSwvif+YtcfA5hixc9Q8
YgZyENWo2fkMwpIxKmIzyynLt0jqC+WBZEhSj0JBGhqyfMP8/oIRqUgE9F7nGbU6v/1+4CwEZ+CZ
bvrUamGT6cs49ZDJtA6qmYsVJB7VB9dDwqwQL2Ia9bCiVkxzhd1AisUt0Xeatxlsq3/81xwB21o0
k9QZyl1XsydV6tFbCE0oCVXxwqt7u12rrOzkp7bvTV6WmGRBQVsiOr82HswUS01CVg43sv2ar85H
OxQ8NpMpB7EmnGG9fAEu/x8laJD0I7u5G5aQihLJLFsghIiNj0VsL2hk7DWC5MMh/NQAqZjqsJUp
SWrvur6hCGXl5TDe4cGPD/TO17sZVpW/hS3k4ZCEsZWcDc30+dGsd1AVPAscRNUR/I2+NPXs+5TK
zKiVNK5XjknxpPWV4+qsK7T64gK3AW8p/4+x0n0mBU2jA5abSW0D+/zr4aesBTao4xB3uK9c2jes
XGsfNxsJ+Scuc9m8H8Dwrar0JR5BwStQc660LSdTR1HDRxr3X2VFsiBDS3FSvccW5QZ7XwyINIRi
bOs+wxoA/a1xFOfnlJKsVs7dOyy+PbgXse3zZohhWv9FUrSnDAILkuATiO39SyikjyWuWr2BHKmf
pEq3xYvtJuOVZzciYIwHGTrlpJUzNkWFA79gzzz/akj4XPN8q4edtH6SHKAOCwg1HnsKmOpE4a7d
Mvcj+9rkjQrsEr9d+hx018Dyrk5931tXvHDdHnl9o+3aKeUzU1/2zgyILvRyhZ/GHXHm5pGo4vIm
DUVVstmcoJIUkvOpGH3IZ3RTP24cREHiT7rPLw9uPZLH16c+qOrsgFrRg4SF6m4c1+AMKqaOXk4Z
joANV+Z+zS6z/SIwb1DSWOY23WMO3LZsxyy8lHUwWcFuMgeEtjuA2p5EHbk1CvittsJ8tv5weCbh
O6doopxgt58qUzWUc5G274TxPGZoqOTv83R/rNWwukgNHvbn/wZp29fXWIXsJHiidALvY2eB5UwC
lcpYkUVbeK3BJjEWh6mC4PfnxQ+J16eByLBglyS/ifX+uAHKxolsn4DZ1bOnMSHVKZapA9kUFuxJ
quvLiD932FShdesfHiJm9PIXluWC7nYBOSel8JRePDhv3yT+DtlHSZXPUGE9fUQSFh4a5/uwAcWS
99Sh01OqA7nsiZ4NlCha7D867VIuJfM7uoNflj/BYzCbCfLpg2snaGFk7LnG7wzQR8AGMT0+1Ctv
g/Olptbe3t/Jc/xjCo54atgvt1l+5Pvh/q3JBTAerQZwRtvkw2phYd5hruk5Lh5ROyWbq6Q4QEsM
HxEgYfP02xdkrZOQqQbFzD2aEGpWb+RrwkT6yd40YMiJEcMjw33PtThBw+NTp/zL5+Zk4/s+4D0p
dV864bsRs7MT/OR1v4o1t4WETv1I7WQHwd44xzg7072qJkNfbwSKBSqHnnxjScSqI4Hg1e/jcVlL
6bTqhfIlfsLV2PnE4jFhJE3Lkk/HFHIx9KIiLmGjwTqNrvDYjtKPxlHmhjImwL9kIzljsA1tjcvi
yI0pQrho4RMe4XvZXDUnOG6HJafXkG5qY0t4JIY8q/rfpsh6dVii/tYeJ22TQTfhFPnnveAN8Hqd
2scb6d8jA735oa6eRbYDtyDLUzIImfDLWr8IeOMX5Dt1T1vwSqbGL5msM5lNgSPQAAJdldPgqHkz
3Q1x4VviagPF+RCpxg4yzcyXZHGHcw1QBiVgD23G94LFcD58lwQ3DDtTAAEmtCmftZmuEuTQC+7d
3/nenBNFDvhlUrkfleFCAVyMQVhK86JbBW3wqx5lptMsNItJ+s8piifEQqC/9KnTIc8Eh6M+H9FR
Bz/SNC0YTY0EfKEL+ofhZaIeeR+FvGbb94UhDsXJCOC2NWjLH8SpnVr2Vz5G9Yoshe2dkm43fZ2I
FYIuEbWBtmW5dfVXY7db7sC+4diiVrRjsQSdD+7G13Ub9CMOVXlMiS6uhio5HJrv0UIYlR6/8t+o
xyQH0NCgtqigruDLMD8r5K4yEV6aMILye4PdKjFJZhDtIWfQiYuRKBVXD2JbhS70fVL0KSsbmd/7
RJOIgwxkPf1GIr/k8CNCbj0CwIcmuizLjG9deDSwL+3LRu/L3OcrgIvtQBC0HCVjmeRh6NzlReNu
tTcw30wt+MkbB+9ofOECQSxlwNSRU1HZSKNiTIlF9CkXM2HXkEubu3luox19o7OfSyteKB+0qf3q
uD0peKXfnY9uZLaQdCfwaulKGlMBxDq/1yPtn04oZJb0gtCGn378hxpOp6+DkKVyo9TSHrjzNJY9
8M5s9Ybal+Bn13Ba80R4j+he9F/rPhhAhAhKiR9u+/KtRRsjO2AddHjPfw37hGsKnp646Qljun3i
5kIvjfywHxUt4x1oP0m5Zw3avbZzhvzHwd0zV4guWQ6u8utkuTXF48QBvbfA8sdco4MqxWJPGpDO
O+HafYsjruoRVDWCk3fiXRjFfxYknBTK91eHCrskZXWzb4RUREYV72j6BW9nrwEF+xIbmbuVvIk0
rpmepXHAKxogyW1LcB0FOJkZMRsew7CDckOG8mFpurD8Ox/pfoXMtB6Lp2ITVYXpEW4n8hfinKRL
tELjb6w7f+m9aNkfIQlkXE3tnyUt1TpXE/fbhoXYl391EJIVe6OKPqzlajalTj5leI+Xim7Bsg4R
+XspEQnEiO1kQZDHB23ZPQjK+bfJtniu2z7tGQwt5m949J4/wUzhxY7nuJ/8RNz8fo+t01wo8pn3
55M39feTySek5w3fdr6aCFp3K+0e5gRQloyTDP/UHlr2JGmHGKbbVPNqjHu+jZlp4KOcD0Xg6xYm
Dfm7PsGqvGGS1ooBFsZPQuorgoWsWhGuTRVZYV2h4YwFJc6+WBfBIJ57PkbJTdoQIikWDV5ZNAE3
y3zbMunVo+76W9/qZH55HGrZtvb0+Ye3Z267Pq+eJI7/EtJ+MT9PMkYbX/SxCUFdUZ5+B2vX/Met
mPipvsEKPJDZzLf+AbTnbxpwhXqYi3H0DEznxEzkyYFd1Z7pHjD4XVlA36bTemlkEADx8ye7vF+B
9SLo9fQWtrBUJY3AAsQFrQ/VNOl4rLfQ9ufWdbdcHKaB4qHy3n3pcWTNQVaCKXMYyZEQFuUOYbcj
ir4vyiOgDTlZYVVfDwo+FS7KtKNsoVVoHvi7xjfYYhq563SI9ULlLA1So8muFhtCiXj69vTn26V/
LIbyefm4FKLb81Xz8mGV/kaN82PUMJdNWsLdYHXOA5Z76PVpLVy1K814XvoxbVYCrx5Q0yGBcWHh
I0kP9YSJa65H1cCC3eeFPWEOMScwIWHIO+NIU7jsD1AEdmKjwhYs5ijqIuZgbc0JtaII3QjTPCUJ
vNpEwuKVD5n7dDbnb/3Nj7zYxSrIiUjlcPrrTa4zAUDe+6qpoVniUs32Guzf+dFH4IYZ5WfaoY6X
yHFI5pq6RbJUiDvoGBuff4aGZmnbVGuD2I2RfcNjaxAhjuwA5nx7y+qJydNuWMZd6DEJLBO3YpLq
SpUILHeCGggjLrNTwJXmAFhMcRkQlIENvAs6EE6b+8UXaMUa9d4OPSAxEwUh3VN6Eajnt5TZu7PK
tDGrnxo0XUQevFbi7XStWb8wBmaxVFa+z+HuSKfiwbtxm1IR/YtxwSFc/5eAiP72ve2VtqhqJnDR
GgqkKaVRF4NJCSh7K91eV521abf7FrsBAcjZAvZU0JsXIqGNvzDsbfGuhXvztSieH56WDyjrBTaf
NCFeBrekoL7iAdJg3cpGrQf49VFs6+PGQZIqUsPb4zUszDGW2bMothpVQMvOlNsxbwINyMMOjJhN
CmrNSSCxX4efG22fMHMRue4xWgevKB9iMWU05i1glbXt+vPN7I9IaMeGO+M18TImTxZOV3qJ/8xV
nRsQFUSt4ADVdjyd8/dOid/avcgCSDPR0p6a6UdZNyM3nNnmOEdM6NEW2AtLeTWG7rQOenQfjlqD
LbIhVCHG+Xa4qifZR4rgHHvNaCXiREPyUI5wsDBRHxMPr25cwelbT9wcfVXANOCcNldVrfZTwPvb
BySaKmOqb1+8D34HiHTY/dt7vDXrb+fy7pfspK1+6AA1cTZLr1E3pj1EbKSSKDRoBTUWR3bj3dc8
Kyap2AmZn3RFrwqysSbGsJxFwjfAj65Q1fVugEpb8N3Ynom32vaRbbeMjV0bBz7anm01MtPon1mE
DmCgHnkVgSVcSXXwmeFBbYsthOerK8Z9vzuau5wehpTd7LYevWJbE0b8mmdnh5BjOW8pZFv1K5ph
NzMleRH+YXj0an6gU4/ruME2UqDycCGA5MroPdC/EW4tUD1v+ofyOqzROlxi+3m5O+kRIilxukBV
kA29JqoYKtPDPYCDVsDk/2UwDJE9iZBN7hpzkdKjnstTRNRA4yYcjyvM128RnIJ7ua6b+YjBgqqD
Dv9kCJi05aRhiu6lvGV96GzWi1I7e6CAwhRVOKgV6GM/lPwWP7OXhr6lZlA9bNW6gXG4RUrjPgSW
iyOfbm+N192UU5rKq9Dvo2yQWmPHUza9SwShOo09nXFpKvprEKZ8GOAo4yh2Ld1oRdPvdc2OpdOW
1GG2fze1FGFtSqNitk5Nnw0exhug4axw+MajKk649fgUTeMfy0bNHdeYBIGTxEezVYznjIZkYW7D
0ANj5GKY+L/k/sz2f4nUZtravpCk83SUGRklBW66k8sYBDHn6zPyHShKBaYFxd8wRUB8unRNXuLZ
iJ+smNpV08ok2GZ1M5i4elTgKIGLVII2FbDeruPEhX8k7G6TIPX0SPbI5bZ/WvRKRrJrPmUXSDlD
hnI5lfAHuXGq5kecj7iv745VEC9VTx2IYmGGAkeDqefMh5Y+KvuHSgxKjLnKy/Xldogvm9lwtq0d
M20jreWAA/rjKhJ4mu8vEvBfnRoEBW69gUrNEDRXaDWpVnKDzkpoR3Xb+gb/p2EkVysE/ZNy+qwt
Ofu1lxWKtI5c0bLAfqdHsjq23Gzu6ysYNtGgsTTA1ntVG7paToKW1vXBB/iq9AJUdFkCZN8K0RLf
vAv+9Ya9SMb5o5leKPtxB463LhHz1vUYZZdsZjEJH4YcECaapaNy76WhB9GQTg0cy2FVJ1CsTjku
sfyB4ImPxQupUohE0S3mn+S/kpWw1OqEqYsWkwlxDwrPZ34vPpCVZuavDwrII5K01uLVApgUWS75
WoavpN5FjRz4UDYa7YCJlIEMXeSQ7H26b8ETM2YpeoUfraGPyRQKIj9YutZ8sdfSGXrZvp2rZMVy
LD0b3Tt7gc6HFUsickt5LhplxHWR0jcnu04/RmfXMnaWbHivXaFJ3xPKY+KC4iOF2oel0LfyMuh4
mBguXa7JaEvQlqc+l4EV16O4JTE9VW/qd3HHQqoYacj6Et7Co8DIt2Duwy3xKajF1HXVo3Hz9UDr
1ahSU0r2ZtQgfjYO034S2jcfABm3h8dSExX10dnRReXSJbbhDzchf5quHKbqkgfO8wZJqxGrEz+9
1IT2SK0lXrl3z03iLrlyZOkXKV28EmTUeglSCpTLFg4On1IQSSJWQxr/Ufv30ZRzLDoqAiNzrCfR
2jTm9SPCfQBKkAXPm8HSm5rEAJxT7lf8wecKP9YwRxVdS0wXSZ8ztRZiTv9hlzAUtLG0DG3DsQEz
A976+sKrFMFUSiGtn2w1oN5p6maWJT2GV96v9dGQcq0QW7YzrSQ7zHsxCsAMSEMDT1mSn/VnjN7G
CRtGPKgBdr2BVMyUNmv3/wzzhgzn+ryxKRX0e6PsyMnl7W/WJt9FD7qH6aDtFtNg0sWXfDeJbErJ
yEU0FvqCE0kVG7hugRl0krtf2jTnsHGsckfVPbvpQoiTjgADtNiHvobKrTpABpmEBKnAFyLQznyR
bo0EfN645OkvcdLFfG/4bUiBJYfiSZcJEqSAyW2b7xArlXLQ+AGAqUU2Jtst25IzuQa8znglirhZ
Q/CZxDJj3Uc/ARLJZdvwYEWGm+2Iqq3kD5fUC4WEaMPcIclE4AzP8fsF+FusybeEIh50CnWRfXkD
ZM5JotvQ8ahS9hlNCXZJoGvN2vgTL3qg+v54QUGiF9DRibhUmn9jJWkKJSkfedGLzPTVWuhiTx54
onFdUJ9ilDAiTHy04prCo81oWWDqDGpN5Lfek9HH32BQ++jbpvtqomvQnYbNnfdOnaAnr8Q6wl6l
tD1ov6XFtSpqtZwoqgv82CkaWWGfJIPME325zV/7WNjuF6FTPyHJvpplUhGVQh0E7VCeJUZkKlrS
92iQ9QNXC119v3nA8BZ7sNA4otaBI2Io/TwRK/HU8zdzR+XUnjmGEuhKnDR/5F7JijJw3eAf/cA9
jb43nI1/5v+WbeqE/FKmhVv7ezDl9Vcc/AXfq4C2NZY79zy+9Bui/r2vrqRxtzGKgCun7iFeeVFo
9ogs2wJvKDyU3jo3+/I01KL6Zmf4uiSz/A3XhX0wlHSaUkQ3jpUc1PZgOgwjc2hknrk3rJHryZG5
knL13BR7/qM9dEy54qRfRh3TuF2alEoY35ojVokgMpl0OzuBRU6BADjQQzFxuKDRjEY+0mQatBT0
Kcw5gnkka6VavIwYA6cQgMgcDBxWco8nWo9wA1+PQu0eJMCzeTbvzGaxAf/rGGkC8K+MmBEfT2fv
RYBmEQvbJKmNvXtFEbY627CGtt7kxPJbSZ0TsrDl9FGftUaLN9ogTBmgbAOC7QKNF+Db5yhUjY3K
IdxqbElxUgAnLjllXqq8ewKgkQAHjfIR1cMJHbsHKEFOlptwe+T1sTpus4F37GTMvJ3SCqsuDcA5
uG+KJpWCzxjE1GJWgsCM6jjxnXAgcaBJYsOW6RZwtY/z4IzR3U0MMaMbYXSZdyOqUjLwz9tyEKkU
yE7z110v+fFG8GRVfFsqsV4D0584KJ9LqXORRTRkBi6NJcrVu4pBxy2lyOUsEVzHK8XfUJGIQq6z
U9OEmpLdfPnMMr96C4BOtuV/xBk7+wTtm2fxOVJHZC5lm+pp9gwbqItAhuLaWxRFl3+grCsHyRYw
geQCAZmnZeugQE++SLOgMiJDXKe0ImqWbfyCZOlGP5SWzrMiH+eHEAmqz2EzZnwEbtnZA/9j7zle
7Rpdveg+kdXpBwt5+u9i07GcyrbsgFz+nzVlVZPfrsGPTZmBTe1oOcEOqPcaP0ljjaZLwNLZr/ZH
eM6A2KfKaAfaIwkCduNhQD679lzIXRCHVl93UfNd+8OKEqY048aujtxXwwDUfaW8Lmg78G0SL+7z
HqW2KxSG/Zz8SbQcg11Pv8oj5u7BtJWKcrSN6XPF7K2jcaQ9Pjqj9FQiFQOSpoD5yIhwl0PhI3JI
N6+EbxsFuqyn0Zb8JtrtsMdaf9fNUm4DOtlg+yNoLxrAFntpmYwCrm9STF5qLUl1iMTAgXIxgCfT
hsCbbe1O/RxVOiQNCP/aLT/pTxR74fWDFj55kFKg/MhH98hkWbf3wLY+bfqK/aQefDu7ocJDlNI5
1SifPycegNzJPxapWjTGSBhx+sOZ8tS7ooLOqbLBoG57xRa2WbJdGzmDBvmXOuWUyCP7z4HJcVW/
OgGRkNZDTH2WCr0QHJkGSPhoTytijybtZROXOXlJV/PI7hAsYgBrotCIey7B5hssUGhnF9/h1lqq
K0J7IxVNzN8b8Ay47TYcB+YzG+i+SYiZ3GzRwJuGLEmbUbdTnaCWzogEkHivyzlpfQwvCX+DjYNC
YzZQrU2Vupdi6AZBa9fXCUYPe2+CX2f2ErkVBYd4cm9ucPj781EaRENrD7GBCi2juUJlmylzBJSh
cnzxH0qyvVCp9Gi5tYLMXWJvmX+gI6LlWXGRPmn9H2wRPfina1e3NMmhdb56hw5ePev3K1Bia0/l
9okgD9GTRcBYkht2b0+jUAiphP1MVK6m9Ti6pOWy3LJ407Xck/oo7nWfqcdwQHbWZmH+pRVZra37
+vLyPcqyW0ylx0bj3Z5QdJ7BD1zjf9DbQJxBjy9iIQKb0apYIClcZJcA3pkh4LgJISvorL82D6wi
O5XKE0++WyDhQl40ULH7NElTefFjhYPs5Cr/pXi7Khv/Gntpcy504f9y14s1griRqklUt+YJhClN
gAmPTtyHlPqXNAkqHhlpv8KtZiybBNHJ3ewSoZtBftSFYo5cPRfKg6NsU5eF8WGpMuwS+9itbhkp
MLF0QiCBgGR2DGwugocZaE9TAClmHffuTSLnC9AAN6gXcVw1yiODavEzOeCh0jIriqa5zPUY8uCM
b+j6D+blpFAMAN/8oUxqwWOdx7gcVNZCoMZu92nO6/l34kh9FEVZmDLGyR+7II4weh2U3wr6TMf8
8LlRMv09a6NP7zrUsQP4spD+w6ukgiBLBwOvlBwc3WUgLKavRq5+UCr07qag2zVsBNMT/IAa/O0C
rkD/MH0uZy6cNSEJLsUfOdQDOWrnXR6mPoFhPf64RmVhT8a0hqKLl9us4hmu6cQQFZuotFU2XM4v
PsIsY8HkLGJlshdZ0JLAWKupA9VXrf45W59ebTYuHQYRZ+HwLgvBkY945AyEVE9zEmBSofxGzXMq
riPy848Bxmj6nRwCppKaj19devgFTVZ63eMHT2oVsh/vOEt+k2/ZPVpmsGgLeYUanpuMYh2Lj4R0
9AuIruEPWnNH6cswlLbjDKe4FhP4XpqCLV7kxyW0s97faqy1xcPwJWnCAxqEWK2H6vZGT0hREj6v
qEu78vjIYgFF5mha1M91oyeOXL8dLXlAw67E9zvADU82JaLq2zeTZots68ZCM9E0Wk1SiNpzOveM
dW+YtVY4+8DsLbJlkirTaYQ5AtayPt+VZBkqvvp0NzpeIBb09KiZvjmvl9zA9AV6PkXBEjRULCHf
/TScoZyyBImANHu0Iog8A17iszzsPtuaK7QfIfTTQMW9MPA63dwn1AVCLbZHMTeCMt7TlEq7+s+u
tWelcZm5kSlG/J7/GNLr+qbCwx4tBIt1xxH0GqwBwhY6vvV03UFPqfUIeYQA2x1IABTc/8oSoo4Q
gg6wDiav6LS/7AABLeglAohoe0X68aMyyvsSst9XW+8h4ACN43OXTVZryHwJBNw4Ki50SuOEVXRV
xgbUCHXLb2tQqppCAuDsYeQYvwuGhwT7/VKz3zGZ8hOJiisaXnuK2/PGu8TGxGiZoJK0/dFj3n6o
K4aIpgAnEZ6PitAt7kk9KGhfv+9jMimSnG+VU9axLHTl3Gslo9+M09UPrYorZXQNjsY+Pw2QJkRA
l/SS7eGSpggogD75Z/ky2jZMsQ/VnAqHl5H2RtyDfO1TL0XaY43O3AUK67Xyqz+3sPMVOlMgGBEu
Tm0TG30mZwKQz6jyqD9G2zopuJHLqZ9hksIzVmZ6hWlgfVcaqRb3rzC4UDpSqIt76pw0cVKqo30U
aXj0NwyldbsdXanIX1KbOci+qdf95RzNgl0Jxjv4M9OvPKfY5WNh+IOPLRSuoV49g+ccjtbSnRLk
H0ibj+pTAyJFQP1kBI8oXdLMiTWo7BYu3jusii2uMLt6r33Y6T69Kl/PfuLZX/Gi358cAl7+UIyy
pJ9Q3I3/bZg1TgS//r7DxpADy2+i0NXZ4h7175aKaxDX3eFkc7d1Sm4Wu6l1Wr1YcZaUol4igNk2
34Ax5g8OwaDP7JHzqVB+mjFc9hvaHOYeM/wQ+qkAj65laBp21X7DExvtIi2zOrbkfQzwXWgZO16A
O6fADkLqduV5NTutr8PDrh1ks/s2GUxusntNpzZFZq4XnLllCeqcXw0viUtlvRIU7SCgFeBD1OJJ
B3MPcxlSfSFT4IVF+tcl8xN69hQYkdm6HMoDTgdhFEtIgzp/NhLVXRMnHSH/fSd5vKYXIJhadRYI
4dDd12gb5ckojmS8DxU+79lnfmFgZMfzolQREUSHSVnzqhkCPSuKOqVT7Z2UCTRBdOf4m7WmKgj5
nbBbW1FviU07Um8/OYFk7kSEutQr8RjR6T95THgL2uABV9N96jVZDxMIVcWQb1+8xlTwdmPF7DOF
VsCdIvKtD8k5EWyNW2nML/r3nZC/pKSnQSZD5/0apKVp25DabtiIIvtWBPN3Kn7kdHhlgN1r6gHt
fHIZrMXB8yUiGlKID024ikAHcuueZpEX8jjFAmMy8S873YO3kcsnxJLuC4U0tDGbY8TGvufd5cmr
01sHOGuetmGkBYosLKMO63/FmwQFd8HiwLVrfOaZZslvupAsLTmdOAiUWoeo1552DKSS/VpvRA87
nZnd+u/OXyTnI9w4TW1E+RwiFvTO1riAL9xvQ/RfuokDBzoZnlnwnt6O6vnGSH3JfIpTT8Tl6z+Z
IP/9X/G8r21e9WIe09cEN3K8/aS/Vv2svlW4EJEKnZYfigQ2R/szzl/8dkBwVGC6TfNsqSureESD
SwYa5SxkiNQZqSbFt6RjQod0Xg1ElwEG/4x9y8HN1pnTNwQGfTk6m8DFb1eUGJXtiF3t4U2oibtO
ySMecJo1D2Txsn8+BhhNNWeAIbgDOfkQ8UosqSSeZ2td+vm2WUdEKwuaGrbcS6v3mZHHreC69IkD
LdDlc5lBd6rQU0II1Avq2JiOx7FoRGLb2eoJxnED9PLw3iJq5OWLeuOItHbbf3LkS8B9EWJmKRx4
qslvWkghG48JgnTpBLmMNP/6seWXAs6gbPv0PovHvQkQjAkghR6NyYHq2RH/myCR5ea/lGuF9Sh+
DxqYp2QkZJnhY7x3Ly0saaGgWnuexFrjsetQ8XDq6fsu0zhoMfJOux6an/3ch79pg9CdTLfvPvVf
yTp/jhaimdURQvrOOeJsDC8jb1Y99rwDJQXS75udzNIQs6eDpOgyE6mCjdO12EFw2yeql9ucJUE3
FarpmDyg5Wf6tujIObPQP9LHR72T+/7Eg/726/BJls6Ghs8ADnrjN34byWcbDavmdwY6cerFGgB9
1A7y4onM0XiepAtgYdcxdxzto7nS2o+NBYuhT08fhS2P7FoMgWquS6sKVlDTAW00FEOcymqCGLIu
0fnr7VEfv7UkKYXgRh216gnJGeo2xPPKlMWNKeYvBLzSPT6L8rmnuBQaTbaacIqE5xrdzTd8DqGD
QYjHeWXYHONePaAp7UbDwjHd/7lClnodOWHjMHBmYgO02B+7K5SUlvTztNmUMqbrgNX5NW6+/BZ2
xa4kifoJSaB0fkVu23OzbCQL60HSGM6V9HvIfvxYmHJsCDKKIt6qEn1hA36BC+lD98g0tg7nTJuD
RPNKPZuQoRrQiwbyZaTsQDyYJfWCbov4UdrPC14Fm/Swz6TJ9I1ZFtHpix9a3bObKFU40lP2yC23
03kBsLsHCKRRDTDbnnjRq6hpNAb9zr7gXG+po1bEiM9B26x4RFEAFEFIo3+1yoN8MGBKDohAoNbQ
oHqwRrf1Bv0wddKlFTnhIko65/y+Eq2rUk7SJz7uARgR4qGXSr7lrHPeAseXxBkOCdjS6SXOXYYZ
goS9ZZThNbv37VS2C+KRLe41zucIcPpeCJgudrBuzEUkUvKVlMXDZRDyx6xeQTEf0sbag2Dv4FoX
cQkua7xPCJElA9N5+Fae8CbKKpdFzBD7tLIG9mNsJ0q4Pt6sZauHV6cajPhDxyoTtSlGXe0tsB9h
2vYKcVs6j3yvFxc2f4HP49AjuytHdsJ+SgGhyqXlriuvBHSUUdr59Ut5W4crO+QT1bZOR5myiTAS
ae9PjystwlqHdXJe6+TUyGDbd7ovlxe6OOJ/s4lWmLvew1fHyfVq1etHVMYVYy1cGDr3vFZd9Xln
RUnElv1dRhTOrf5G2As5X4iHotlZZu0KhWVDYEIFGsKC/8BvZs0rodIM03VqZGWMahMz95yt42Vv
UlfiVz+7CpyaXjjmiuC0orLFQ0trINjK34qLZspUo3vN4sJ968F3fzGc0jJsc48Z7tBjPLTYkNA4
DA1O406Y8hvCYgfWH8MeLH1msRxvdATzoUY72ZJMdSHMWDttouPms6X1bkX3yNBmThb66xdZrfra
axoL6I9tXITgu9mJk3wiVfWuQImPasRDySNlttdepkCbQB0p4nLUz4xKKEjI/Ns8f8j7sylznhJ5
bkv0ygVPkiXP3gI3mZRZXSSdDof+h08KeMtKVinjf1cDPKtCQrhGEykFTqIxb6v1niiKdbp11Jl3
24CGg0ZWAv9ZGU0irH1d0WJTX9P3p+XfPKl4bXevdKdz5zKOyXxTg45mr5d0QS4CySeqYWx1YACo
CDY0bVzgK8WplbdUtMTvDQr9Z9vyCi0Vx2IrGEyqa58xKLBhDDQpRjYGymkAMrz/IB0hMp9Esqab
ebH2lpcgJBOFFD/04oaYrVkgr9U1rRZoUn8hg5H+5/6wZq/9zIWKAuthvR4ymmg4EyRfR6zp7yQn
BFP/N8xtFNgQOhXn7QiTqVP+xRgy/4lfW9TWjP5DgucCL8/PA1nWFfWv4U3WDkI4jaxrSEUrMiDv
iXKigYXodHQPYHGuwxRCQEFX7hpGNJyRCrnUyz+kyqgM9j+MWYrzANvUo8lhJfWYoaZcnFklOTVa
xHm8PIMTxvCjQksZeEH7TUsY6QvAlbj3Gx/JtnBTKlCOFMm2LXki94g2gPrXUngtiLw/ZQawD2+9
Yoee2TzmnWYoPSGjL6jLRrHnae6jVaAsZVZgjaBLMj5wSIUR3s8hLepI5Q4ST0qmv65XoIT3T36v
QCQpI8HnqZzXUfVf5dkh7lMz1Jlo/IH+0JZRJkH2RknrC7T/Q7gnjjUmCOG/8MlZdQDrfYqTMWMZ
x8F2DfBdcZ5saCR7e5pYi9FKCXLDstxGOw7SO401+IrKF3GuG9QSOnqFtIN5nyfh6WPxyMlVqqb7
L+iKGU7Ccwh2j+2U+C0tz3h+Dx0U22TP4LOTuY0xQPUlGzZfTlQMRHpLHbO96eVB4A3pm0vlE8AY
YckYxzaDb29H8Xw6UGulgt0frRIcEcfO3dx0lrTi7DJa/efYF9/ucoaf9of04kVTzjm5dK6vbJi2
0XXGYJmPD+v2sQ4/CWWVkD0XiGbp5lQEg5dW8MAETHvsevHmfXkMIKU1lKNokPcmoescq80JRw+4
YkPIbXed/pQtUQT0VsHa5/q1fcADT+/NOfu3e0Xaadqy5BVlxjJDDR+6vDv8RIkvyy/9uo+oSpeZ
EGIDJYnxanJ6FDfcyXqp9ZA0Fn0r8yRx1yCG2lBTXaO38+9Si39wCt9j2KK4+dkOST/40p5EVmAL
JdMhfCHGUIGCSnE+kegtyczamPkIuzFUP/LqX57UPQkkkXDA4vNXYke+DSVcd8XTBJKUdNo2wyHq
G281qk4Kj2PGbBrLxOYTflnaH8o7HAlakVEzUq3xVay1mmSiOycqTvaIWXgeja79MLUGEH82UOQ0
uVAvA1D4JvL2cPxiEqgtRBtLwfp9KcIT/eA3bd9gEemNvzOnuzXyj+6Uo2R9JiWKUJ0U7FrIM98W
gSzAqZNapB0ngeectWn37TD3n9PTzJIGCAM7LuNW09u42Z45fTKXjOVRTtCi4NVuIU6WaCO6M/ni
EcYXUSZPgGZ/w1sM4b3mIpRUTVwuwO9w9+8gvZXov0l4f9ObvAsmcK1HZ3cBSFO9C87OOjUMkuE3
ZEX6Pgk5yOYagQvKxDDZNOOqI65tJTy23SGgxOxvyMK+m48uNB56uqRhpXzhl2Spx2WFwmetGMKS
n14ub34m6ESkaBHMHTlvTKUcP2gJJ/B+hZDLORrEWOdP/ajyyIjB3vyr2CrwmeiDxH6OQCLf3xps
HokpNS2ynjgT08mxwKIWXzm8GspBwr58qi+mIdNkv8vHVH/nrqbqX91LmaJS2mZH21/UKf4lw4vM
UM92wziyn+L4euE7Dhzs3ZW1jPWZL3XsdfOIwd0QC1sfBNMTU4ErHmsSyVzgr8KsiSYHs3+rTxwf
x0sos7IfEovih1o27md3XLcyJh7hDHw5KhxRP0sZlo5X4G8ZjGhV/da8c3l5vBRgU3zdvuAa4KRY
5cmHx8HhPhhGUB0oY2RKBcIUpeXigEuUEKNDMlyFPShml8ehobD5fPNJdw1XTMpUIWBbQpZnSQtN
k43QaCQtmjwn44qa1f/RR7/fPixPNiF6FiOxDAOByDMxApiRNPvoakDgrOm9L9Au50mBp0bRBSTP
ebYSSL9oqN9ig0OrXm0Nn3BFslDIyDrkuX5lvZUlBw37rraR2UTfDBNKKyPjkpO+1URQjyqHHc0y
9Kh4uqS9P+dc3+ONPgsNeFTuUgoAZ+pgjgmAyOHHt3udNeCdVtuST1vP6LTjeDzNBjCl2vzNwKep
8j3i3xrbMmMtnXuOqmcSGCv+r1ZRmaC4bFX6HAaEl84iRrES+YdKQyC4SPNykpn6SB0bHTEetzTH
Re6W4e9HXlQ3yd+m/daOda2U41cf6/+01TSQJSdhpE2H5e2T1VYqq/P7mTUyaSgIjtTpILKMhtB/
Y7TqJ/RwkBy0t0Vt5FWsGuvqtGDx+6Crp/gKI07hBDp9D8g9TF7IB4eczR2yd5vwZ5KEYsmmJ7Hp
lf20UAXupSsqtt0GQlmAYr49Xg3yUevVzJCXJef4tXaJKHjvMSaB9WONutOcKU3ubb06u593y5i1
Cn+z26wa4DQHp3k9vALjxF38zt7C42hQ7okiWoY8XEMxyo+15j2PZM/CF1jIQrTJHU/KP/0tDkqz
vukbRLM2ezFyjmJNCQaYIhJ4EFpX5BKXvr1K7k1ANiXeOzNjP4Zh5FYC/9ZEbIrYfEWdk0DyOWCR
lF+ODoocjodgO2h9W6d+HaSc741dEgmeHPxB8Owl7Szu8jytk2qClGyG4Dx77zxtBBRXUt0f749a
X2mR50dJOC2hncUqoZ13MjvXKH2Z8xrpXqGb9UK/AvB9OqwRxPDDorjBaALxdXRsO9XUIkK84Luf
Y4zZWglBp7pAlPH+X+hvFfZqyuk/EYUz0jmrtByoEF/NUQU8eOUGw09usGLBNzqQIRIvRiGILVgn
9LxBGVmpjJ4Ye5qVKGSCTdKSmlQq99mnJAHbtIF/mr4VbqGHjM3SgtEkTtTg+h68kSlrCf103AsA
Y7Rb8zolUO6RL2tAt9s2oRHr1JoMivt5rQ64xyncpT73a32bZTjkMKraQyq8Fo1s1vDYX+Fpv9Aa
5JIgxD7M/AYW0Rrwk5r6pnCYs7ZgFW/kAW0dYW1ZkJoCmbuqoZnjJBJnjVllDwJKojr0465xNbmF
YaLEqHpiHVf1twl9NLCuUfDomhEaaMCIE7vPIPD8bsjVxb1hz6wEAJ650tXhmUcpCrPkgukrHeo3
krc9pX/rS1fwTS+Qq4D/ilfhTlrIqVvLZh1F2dkONqbCQzJVvay+gS4QABfzxPGQ9kPLR5DkduWB
RHPjX4kJ/gMoFr1V/Th3eYzOqsaxEf3Iy9hwg3yQTcp2W8ij9hTNtQqgTqTQFXXwrtWSZSGUK8Pa
z+pCUoPioJRvglDsLhx2ejPFydZpwxu4YEmUnqWAdbYKQeQCvORgSa2kZbdakv98r2XVfBWQGOs0
QL9eLg5Jw/xz/zUvMmoeKA2XfqgBPy348aJcB/8TkXv5pdjO3VVu9uFBZ+B9pnI5Tp1Jpgnm1k3f
4I6DBd7WZNIJ126slpRZv4j7NWQYcEXKHRysKx0MpwObBW0b9eQvGh7+OWnV0oHBJcT6FDAzxEAj
Wge9TKbsy01nxTU/pSjbxEy+0Uszg6t+4PlHjocppDJPs8Fw8xR894MzMK9CCYnvJbaUsFt6hJOX
4LcXZ9PFXHWM/jE9Di/x2L6OtrshawVb1momyLIH6pfd6MsRy66AYh5+JS9vIH6VNIcYSmTVC6y+
A9QdTFzcPl/ksyseKesPGYsnJh/+5BdSrylfCJ4EB64+bpmwlH+SqfGXzQxOW8M69D/QHj3S3A/f
ZW7FSaQExeZ6f2OIwNYTEduBn3600xo22IyUDUnG0JS/I4wkOnMoxp1j19a+TEaQDelTgGp8GOLl
528PaEWJ8EZTdZW2WhaSe0G9bGG7qLe/slsdX6kdyM3PhAyYQz9vo9jJFPY0k7GhYqL0Hl8xsy0t
0tBLjCUZ+Cabb1sPViMHaCHIfJc9OSG2mMvffRVhrO9enNmWSHaLzBrFxHAg9Me5Eps9uGL4u5oi
87xjcBmDs7dcYpwpahEleBuwxeDJAsQtRqoEDkNEcq6+9ZGHWK3P5NvuDXWPX1mEGafVtWFelbda
uGTYQb4KBDqmAB3aAqI1UYYUbvzjWor+s7OMuV9fAVeX7IWB8yZ0Quvrxrmj9EoKmjroKxh+3ttg
yZ1xOmpq9dCbLZFoZiT2VcL7wUBFk/hS1z64OpzCCDJUdQy0xgV/VOGkPuUlRnO8XdmUQCuzeNkY
VpWleOAyxr3YC8Ulyc7qgFh5MXrElsOdjgax4G6+o1UrDrPXK/uQdzziHkL/wreWovC2yZonV//o
Tfa0Pxh8YLc9Y2unYaeQ7WcD7Qa5p2GiUbiUis54/4qYHYK2eHrka0YCe9t2yY0NOYlMv6xWS8hf
6UkM8Y5mRfBLAQIXRbgCpy/ACxHmSwuQVEomH18PMzvLB7tenjDSMFTmi4PJCcN6Y7LfEDu2v0Uk
81HDhdDFxAgpWbEESDDtwk0tbhZkx8h7R7GNRxobjT+QHydRM24ytFvBKNx07EdgcoqgpA6EsoWI
LyV2Qu1qsemiYM+aMkwHsLAdAujw87+kQ6dV4/ouKbPsws1efiCLhFrmu6xgTYfaja/B16xoY+Z3
/Ctzel/80oHwS71kNHr8LKhcdxVBalSxdDEepDRzto+x9rfjriykFnry/a06w6N1mB1eikuJXQFN
CvesPs0JInLvs3Pyl3EFFuvuXLbKYTW8Gt5u0z8XyMLCRH6o5RQD5OKS9+HFyvSpZjLLyYREynSo
Ku0xtvJcJzYO5n61rONV9rBmurXa7phtVkAMKy/suW/a0t3Vysejdk8DnRu4m9ayZjJWiEHE2YjP
BnBSdn+QiVyl/8pi0fpsNT3I+KCwrFZ58jTwUZswge7piPb1EU1XFHru2LNuuTATiIEt4X2ziwkQ
NZWg0aWugn8hzgERPn5u+EXs3OMThWFfKWZr2s7Wb8coRbpEddTSvlq+8Mpz9BDdvHJyb7RxIT4X
EI+oaHdiOxztcwGFhHYQM2oyl4c9A9lKHuvJTVOwO69HStZ7ARrAesU4eg9GHxEERWeimGRaop8Z
irBGCAjUXw1GrA4BI0hHQPzWA7DEVfzrcdZwUbfWstPLJyBhMi7fAMqlRweVj0wf9jrPgiX1V1P/
f5T7F52qUy8q1a+QbgclvC8ANN+GvQZCdzcXvOpAJUAcGYwvEKW9W7WXrWQaeqAC7TiUG92HOPae
dYdPqaHY6JmBjUodhp4p82Oe+T7kS/xsQdjE6nkwl/5kuqDDKjmiFQukQr3hG8fX2s1viNyN9xQj
jnB8G3oTFGgNsEKCfZGtBRvaongcVdkC6cIu9yf6U17X8uv9YJht9Qb+9wtW33MMnlr5bl7s+uRY
p6WDHQOijVVbIGAYj3G4zvabjR8KvVe9uD0gS/WsNC7UvnrJgVtec2ZjOqZqBXrCKzaBlRwbtJY3
ggxjqPfCpbJPaIlF/PZQFZDhTFBUg2v5IJiUhjhnuMaAeaDvb1Z4U3gZE9lVBqGXMs32zpAmU7RF
Siv9BsxeqBVmWS571gNMmsbInOMH46pyGfBOmDo3OG0JQsHo9bfDeftD2BGm47yW1kReqy9pOs55
wYKjyAVfgepXE+1NQFbddszD8c+QdIdA21UIiptprG5OlLHqstZeb4geJSEZ8qPkcDDUxn0c1wZA
4+771U4xbBv36YVS2js+JfUDVNvA1D0whZokWuV/mZuKKNnEtz/9VPSDmbwGO8IMoGmYFJG4ShER
zjnDjRpUEqqXuSt6dCnKNbbiHBQNOrOIO4yyE3xMjdI7TlX5Ifx4rses+dSoj3tS/yDrlc62QFwi
XJtvSF0QDtpg6f1yPBcY+4zlnxtnLf088WdRQ3Ppr0OxaO2vBgACN5s+Nl7ejE8MljRPuYlV4qhh
vPwXvJCFpo2mDSj/AgN/UterDkI/Gq8uRxwrYm/4VhZlGZunsYyTsXNVj6/78ABVQjmkTSqugGh9
tMRUGnI7JFmBq1weY1llr4xCEYcdkjrbN5WCnCzDs0MSLlrE1/nZ4f1V0sR3SC2s9A/9z0EMTwav
QQLnnWKm8zj9XxUPeDACmM/Hs7R42aGNepIWiLVkkdRI/6MOFHdR8GmMQNSdrFTUa0MKHqUe7J39
dlz2qX/ixTmigN0esmRwRcuDp8DIjBtL249tfkrBKRXSY31VMEkOqyjzdKqNZVwAN6G6eO62J3oz
tV9QYOhVlY7ApaWfVOWxpWL+K4cxGPxK+L+zqYNtuVu6yPolHt78kYBuUM7kaf9T1KwEK8aIPDlh
7byhCYHPhCdVQke1B7MHgUknzS3d9Cr7Y8cDx/CdalZsrx/x2zzjDApdhG8GPvGXmGimyAqP8zyy
Wt6q3c7jUk9DN4KF6zegkzWSL9wgPX1zrrqcK6O0TtXNSlzScPhZ7FQAsNsVp2e1Xzn5xNF4Ltn8
OkbZJx2DxqV0RvDY7lhZpA+4inDaYR2bVsPORByAFMPCgIszh6JPR4JMr5eC65w5RswocjbEH6CI
YF4TgrQpmQlkKJ7TIvsrKb7uxJcY4XWa1nAyibFAg6dMkgnva/K4dhy42SEMNQksH2dX68tHNFsc
ijiPTs2D3/napm4dzmnQvGBqaziIB+B+IHJ7qUUN6vaYOriox/546Ce2adkH7enEynn/Ne95joaL
DoYOJvzbU6hjP5ZVUV/ADJyDXi4zoIe2/gTsinRLiSguSLARsWtVu3VHS/p94rBVByIknBOqtckR
euzYEVZMke3xzBdBjS7s4KFAjjwn9MlszAvhFPbBwpjaU4x6qNTUGOb1+ZVsBHl2Q4cbdNJniKDL
6Aj3zpvDoXd79O33n7vRbQKwljQ7lwSyvMIm/4xSk1C176jN50Ln35ulIwlhamDleeMTC7p6KgsU
AqmiAYn6xkItvdzM74YtS7ZgqJRUQw7NR9F/DlephRXNcVnavx+FJW5EGUHEizaU3oGy5tgCM68Y
XFkpQvkm6N8BnrrBDgf2c8CMMOTRcwx/BJp0NHdOogMd+H+Co+A+eFRxvaJEjFo/X0pikOfjkM7y
aqNVwyLHNTs820b8xdrnh5JpBy6QspX41TQoSc7+KLjWlSR7mvRuJr6zaD6gUJT7NfEr45vHROGK
P88xssoi+Llzo4TFrvYfMpzsBOxKHxqZp90nXn6X4QDbJLXBqrPLkoHJwE7HBO2bQ2g58g2LkYYk
W/RkSS1ELYWri2FhMdBT5cvteV9J+OPiOXX2Uos8bHVMq2I9nYvT/Vab/lqAA2XwpDzY+cqRpo0L
YQfUZlY08Ibkjmdr7YMbYHOA89rsHGQyI1VcyjXCuKgYA+eaHGkjJx02QAGi8iokQb9uUkqGULcL
R9qpUicokWwFVDbVOiIGimj5hqeZhprGcAhNyrIDSnlLwBjkpg6kUOOnnZR89d0EV/cABc45OUZE
H3DR/QO/K0ppVoGLpfFl8tAuuJ1w7RU4puTHZi7sYtzWpSCE/98UYNXuMza4IUyycmmYn1TUwzVS
CtVUo9DFZE25VfkgGwBdUOchDRLGre/+CgsTVGHSv0ODdVqUMtYlUDXZRZ9reOXyro8vlbBqughG
nFtREj5eveyWl9CdmIVj6q56t2MJtkhxMFBjR3SgevAInQaQ6plNHonrZn9s8SpSdYMfffku8U7W
rQdTRN8xzyAwwI2iryS9Anz+N9HnGqX1FiCeaBbOya6sZgfHktjST2+UQkTeIWqSOXxHKiM6QNmM
nC7mh+pCnGFF3r7BBTuPMEANebnTEj5sz5euaK8wsxVSaWf8bXbpO3ylzX9dbq8LsfIbVDGS105g
Jr0N2HzV1U+mi8wAGSsdJ8gJbYo9yzSyH05hd64p9027sa46802q782La68ZYB+i9JW21XujOJQn
YQL7Skvel9RnF7PGKDd1FIjAZrZkx4FffdF67mlvsZK2dA6oh/aAiZftrZq9lCWMX6ch6QbtiPrF
cXG1Io5WMWoIiCT0+TzOusp8oJoxa8m2liPBThh7bLOnCC1CtVCDOj82+Isdl8k5ZGMk4shdXDOX
2/LkopXkSN15Bd3KLEUl+a+8uu9VZP9qzl1EkUSmG2jwCMZHccchA/pc6gTX2V5U8L/xXyZQ9scp
JdsB9WxblCfZM3eUqUjaTwSe/fBRwbmAQK9D7ap6hcsFD+NGNxm4E2VdoEO+oo9Uw1bpk1Dyi+c0
sAKPOz+rn5h38xcyPPbW/aLIGGHatyAYyGi7FS0j4Tcs53cQx0WKUftU0LsQbUSAszNODds9ClbQ
6w7HYnrbCB/xWbt0vWPfS4tfaNiAR7ZDbVqiihqZ6KQma5lHBxMqwhS3GbzkTWY+JdniXjYCkvOk
f15vXm4XVBh8374dWiPzxAomOALetF9XWoXdWDdV3+B2cf/imnS+eWNarCyBvvnLG+u3BUlxeeXA
I5ZdkiIotGjKMO4aMS/PSY32M4dDBiFbmx3mQa3KZLqmv7P9nliPUYxp+AEimtw6fo+mRDcEWN+x
PyODOJvRVmh8u3MxuqSdeeRbjLGXuPyNDv689QuxsVcqoLL9U9bd3lBwzBDvGqErz5gEmhhClnKY
tP+rExZBrOTUch6BoqbshCks4ogfQ8WK7h4Rp0qjt06y9yn3wmWxbcFLt3GwwGPuLsSZBhww1OLy
OzeUF3uyk/PvIen4D0tMkw4ZMDmAGfFPIOYAdbNUUg660TuXzQurcw8ecQ1ud3+YtXlmWxnHx8c1
Xe8ZBN/wTOyeTclYXut6Hd7YXacNMxV6phWXIab3riHiYoMWhd3Ryzvdl4SMadf7YD+7ts+TsMA3
5y+7U7HackPnYdWfM3E8sQ67GhGVPhHqCff12bxl3a/OEz6YZx2Shxm1sm6hQHAKt2xoEmJUjA5b
S25csNZ/FxsBB6Fnu44tWn0Dk4O/Eapn2qfxBRLVGuIA0YR7vNHTLDtokbiuXPwZ6kEyaM3wb92H
QC8GP/XU0bPuWXyQ1jGjg2DMCZ0mwb9dqzlAPmFuAeQLEw6/HoSfRGwTUWqglXX/w84LgUGrS5Dy
VCkAVWV6lj5ukqFrN3sZTR7rHzy/8XJu71he/TU4Cw4ce3Lapyd/CT8XeoA/q8sm33qcgq1hdT75
cJeNrT/0UZHQW7TAzWw/tRujbf28e8DCk9mjjdTYzFcO6Gm6g8ql7IHH8cg6aCxgGxNaHQ3Pc/eL
t9Q1FFh9Idu2E7fRan8RGeAcbfZoah2ylnMlJWkb9Iq5hya1YvkBVfxgjoAjka52CiPhLk1OyGGF
5WrTST6J0QUqk2w40G+iB4G4/Wvd2WKTwA8tEAFEz4MuJE8qlzCXyZhMheAlUDGt7aSZD2hgU1cb
87AbPnKityk90mO9rgnNLsPpIhXKbWqSZf97JIokrP1G/dkH85/xeM22ZlHg2ki4yDTnN6uHLuG2
6ilqTdSoxDWBZ02ON1++LG3+UYPLEH36FSzKwn/EIUtSAEx0ZTVBMs4f5Dxhk2gIKUM4tCGcLxXJ
fgmFIvIVx9GYqRGsGAoux+KpO9eYztHtTDb0NTeVrF2KpWgLbXCADqIP9fuub3FwZHrvRQ6B6enI
cntyPnE7Io6zlXdnpkD95kv2N235FPfHfXPpBRuM1eoMW2gcFUTw8AGBRVn++iKLOnwNT+jguUpW
XxkSkKnDCY6Eoq2Jdcm20jA8/0/FEzYLy8VZ0d+FyR1DxSBeSViG1nHrYkm8o8yLwblncdMrHbZV
bshud5Os0atWmtmwjwwh9Tc8VXLHqOiYi5sc4Jk/tShXyNBI/kwEuX8JnHzwbMCyqCo8HIsPSRL5
+XC0/cSneu1F9gUeZ7+/ARNRhpn4dm3sIPW+tyGB6kmYBpNN3eaHYu4w1WelitKr1xYNDx8Tcqk/
ceA5QjFXDx3Rkv5LB0pyOQmQN8bTGoaGx1EgLxDt9vRPhpORVfYVDqWeVdow2pEXKYrObyjwqzQv
ojGivMzFpfOuMRIzoEkLXPPryJj/ryes3qr4M5LwicZKoqDTqUnCvR1niiXZW0qVvXNXRq83Bnqr
UH1id6MUdKG53Ma2fH2U9RMhh0EK9GC3AQiU2npTfaM7CgVoOw5dwVmplGiJjOP0iTa7CZNltr59
rTW2HbPVxROd58hOVVNmRZG0LSRXCwT9cGHakeiBgnsLeVh04uAYfHmE+jLdPs/lqR3UVUKmtfOP
2grVlwM0sb150Pmv361NWKNNVxr7oNKqwp/0GCbWUuF36B14XjY3t+vcvLPceO4rFVng/Zi8zHuz
f6/H/lBnovWGll2Lwg1MCUS1CGH5+AL+KNP6D8BJzMBykUvNcTCV3sXAWqfVp9QupkNK/WjlTf/0
qdnes0rZFP8dgf4GVlGmV9Gc9/Qi0m+SyMZgGpcuU1XafcENvU4jXP77kiIrgLMQnybD06KUnXt9
GyC+qDtwzdDyHa72FEoJqE3x5FBd97VSjyBHmX09DZdqrqcvWiYEyZIYJ7FDJgi5AnuMLPO4jYjO
tpx5UceDzIgvI0ChVytsVlJLpVT/byHer/gdVtTDPeTL6aIDVeF/9qc+BYkMkwMCREFQ+ULqpV/A
ngaqwwRcGOSoHJX9uuUKyIMIz59UA5HX6AYDvZdCqBf2AHNRFm/Ml/na9gT47khqM97q353ywRB7
iSWZsHuUxMm4DTH+mcMXYpoVipQnD1Y9FTXv1T9dFDV3BzfsZbks0RNsLZT22eJT6WnzXTaouJKL
6+4gpTBznZaBopW7XK27V0Qe7UrZURdNX19lw5cLKToKS1nh/EO/+QhlGHM2aOQ1Sukt57euhnU2
zASy4ndz6pIgl1ROJWK8zRVTpsIgIYI7SO7Npwkpuw+M5fEFXR3jPBZOaPeThk9ELtONG5le+Bbx
JGfivkt99PTPeDF0mJ32fJeAjIr0dwJsTDaMIHk0LlgPBvc7GDAd/gVqOke7Nvcoy3n4fM3epU2c
3cgxI3g4Z7Qyn2l6tV13j0DGwPLo0iB15TDbacjFY5SnSr8aFC+F5913JLW6ewHtNTsFDu3r57mT
YmRlwPdbKdVBnLlThn2wMHg/kF7K+cn46uWNPC0bXV5NRT4HoqB6QKSCZLfkFXjEiqXJcGEIztDv
nHJDOPRnKTYECFYRNnOEq2Tm4bsUw/YY5ZGLDAit89UcUArv1EW71UVorR4fFIzILuIDUGOBbcgO
/T/FkVjTfo9++o22S8EyedEqEApfyWK8+iCFfRZW4X5LaKbRcJxpeAFA0vMzZ3vV8s+qwzdYVbo/
HGQrKEhGfwZJ8S/v4+bYxPoqcflZWn/aOkMxsbLsGlIHehIrVVkCZL2ph5U+TBpEzZOKstIHTtHq
1zMhxbMDw7yZE086TgkCI/A+ABUC5qdjE0/MP2sDIkeg2JZJDSWzrbnMuqp0RakcXYVjNQCJcWb/
HzQjwewHwRV1mv767htkHMnTlYw+doM086FYL6OAE+nR/CQfxw14ief5xPhaPLnzeFTBL3FbwtTT
VPpI4QekbMyeAo8cRVlV7PdJQSV2/37nY/5ohsXuVm9QzmUv/zV1hQYUqFolVAgvWDfu5EbMS7is
Kwj0Bs3Pj4BrBCcKM9FCLCXv1Ee2Bl5oWsb/DK5vp7wGAAqi2jp67LGuD5eQn6NCaGv0Z101psZ4
wkesmPMCX00xRQGD2pIDM2B9iE+RiP2lQtAA7BExrAeb6Tp2v9S2z77cGQYeLky07SXJjtjP+u6F
uh2za/Di6Kyw3ziLwPkIJlpKVjl7XBSkBi5NNwwWq+yrfBhAjKzthdmVt+uozlFTBPP/AcDFeSQ7
f4xPUTYUMDjX3FYxqKbSVU+i1sQVo1yDBHbimTUI25gxypzTITP0c8Er+jTS7L2SSPkJrjsxMyM5
AZ5kMXlaEOhnqe3tRmgWcIVMG84cG8NhtrtRbxYOOtlQCmPZZJN7ujKikI0la0B+4EG9FCjyQbEA
RAlAr6fBEOUSZ6atNcFmyHerOIj2Ld6MXjmxJDOLsbfSEf0Mx1vcKh9ATwZTTob/O/TmYVTE1Jwv
T4aM4ykR8fzFIGHNTtdct7C7ouXZP37LIemAWncyVUqCka1l3Fi2l2G6+2WGjTmX2jgy0vca2EhB
xLU5UN2ord25NRxBgxG6r7ssf5g24nWngdQMmPuqhhCn9W/pPoal3GrEskdDI7JrR5+Zp4060XYa
TPv15rcfgQv/tC0m9qsv8X4Em3p2/D3KXMAcIST55eDtBEmGBZEqbh8nFrTT5VTfPT49hT+q0Rsz
d40LUtn5T6c0FxyseB16PlxUlJ+6DmRBzMzaAU9cXcKiDXuknX7lPNr+PqrPheJD7gecwIBScusk
Rowo7BE6vxYZL1Kym1u8qGjxd5pkhfuQLNDQGgBaZbhD1HwEnyw4XTredJn2SgoarGODcwWwtLzj
4Cf+SujsUJ/4tieHEVDoPPQ9VBwCiRKHEyKOcmrOxyUZ9k/XMgIs/yrAHyVt3E68pWJVRqwd2oWY
1PLiIuE7gIyEpAwvI9jsVPFiLk1T5FXLn4wM4ToYe2q0dIZziowaGsVV/oLSfsj1Z0IGuMq1sPxn
WY8P9VCSwS1YaLbsSCKBqMtsD7yOIuP9gXX7NxwcBeLNvVhD5TZ681F+fjTFszEQE2RZKr0x9Qzo
r+UDNZ8gRW1Vw27ce+17TKVwKY6goE/HaHYaSOJvTQUQAKKX1GHJMNV2p/RYi48DI/kJnPiAjTUJ
4JgKpbNxGdenWPwIgRrcnKmq2tUUgPmE8vgjGOVpB/qse0y3ulabNLIj5wqjP9IgxKZ3i4U9nrZW
LZ4hjey3d+7fAXY2RS/Z91WCkyQ7ukEl4TxeNNM/yuXyZhBim6jFGiA6s6N6oSR7Wg6+/+Kimb+D
0Btunz6mgPwSTNxOy/nLaOvDZAI5yr3PSDctFydSG3g27oYmrvC2Zwct0kh7NVWLL2pLkdZU1dTn
6M7+9hYnwp/DhqjKe3nXL+YEZoSp6fogyeeLFkcSztTAwJN+5+DYQn4YoxpP57fgCr+u2c3er2Wt
Ii3owIK8iPxyNBRPv3OqZWe7g904p28VEfkd0iR4aJIn2U1T+vDNtJC5edoYQXuopxoCBQikgyoJ
yrL3YinHWGAwqNfXM5+4fiGLiLEUzu08bXtQeMdy2Uc6e8tc8qt+i5iOJC1EHVxUcDc9MCNK+oFI
5Ba2FYhLuiEnm/6XeiYjw2woDX221oIiStMZTMR7XcrrL80OO6UrZXxhTYfOZQKMy5nCBkijc19E
mXcOWjsmRQVyV+NVsk9GiaZmAc6BhUfb4kW1WHAqWOdaN7zE1VIydkVGPIUKk0skS5Fniq2H9qB2
qvOcQYnN6aHcApdV/rtiD3nNy1qpsVTL/b8pN9XYIq9lXtn4Re9wPLp9s5MIo/3P2NOJS3CTNLpi
dUN6GBp8TzJkg34lCjhptyq4H7DIM//UO23cXMsJAOtyS7aet6kBn0TmZxlVKiZxxP6hJnh5gYns
nX58sPusuh2rkelCo6kwHIy4pqp78NlpdxTV5GSLLz5BjSKKxhRsn8XD9sN9eiX10y3gpK00+rie
CecWY0bhmWesSOjyZ0xbA71KOIIZ7Y2JCXrBAZxom50WrK0qO7ATny0n3WPHopH9WgwoeWfJDo1z
pa57g6qUZhdpLzXiZcJy+tx2iWQt/OTLuojIE+XrGlpf8IQgwizjJi4qSAPBIsur3mdMnh5JuflY
1mZXhi8gDj9cpsutD3AZ5srsqw2HJIh+LNxEaoE9IA4Fr0rrItIc3qQFC+ocPovul6qbuQzPExNZ
QtA4a+D2KdhGzXSUDj1oLqhYKiGTTHQyZWmZ+XaDCMl9FqN57n8kOrmWSOllG3EVNcs/N2c64EUt
fk2n0Jwl1IXDkcL2bWaihvTXFRMzBNQ6vT27mWW1vu10GYAKX9Qk3CybIZZXe7yeZxzzmG04+J36
FW/Nz2aexW9EOtKlelwr5TLaoi/Mrrk3KLqpQHPFnRsLXW9cgkK2eYMf0K5yoKHNeABgcd042K8h
Vs+j74YxlgjB9x1oN8YzM96fCyYBDNjguvfeVdlMCmMM/Y5wTNjrvKDcId48D9M7912rfPlZa7VB
o79Q8vGO34Rhv4y7jlnb2VZze2IMppTThAnzplv9SQuy4E8B7MtN/yelFfn+42JrChA2lRR9oEYN
MqHhSWqm7XKNGIyDqlWHKMm0Td563JI4gmha9W0pjgHtQqZMzHW0lEFKnQ1e5IxX3UYxqSVGK0AK
IISrJeGGhE4itPZJVbiaIJHNDmYzDOe3vAmDFxP6+f9cOWKoZ1Vd2/wiCBhqqT9P5cg/ZXCdQVHR
sa6PIHDpS/97KqSF3k4MUhIXcsCUbVaTvAK1/RzRf91rkiud7eVz5AzL2BTdvY6klsq1SXEdGAC/
kV6yYxn+E8OErxzGHcpbr4h3sL+TlV6dUmc+KzKRa2vPSBoIrwfzFD06Qbhu0Zqiw6/O83SF+3Vh
uH/xUg0XVNe2SsF6eEZuSJ8UrHHCraD989TxFgQW6q/feRPfKIJzTVtd+d9DEMzEiFv1mhVoiUJv
iwjQSxkewgdaXI2fuuW9DIFdsM2hMmAZxkbDZbQ9yfdLoutG68VImmDLdbY/TKzVPIGMzY2h+r+G
ju5vav7AjcEiqndco5cHMPSmVyVYvEsMAJfGiGQUukijAvgHLjLRM46kKpN5TRnaFhH6JegqS+LG
PA3+qyFg0YR3cFlNWpaE+nGgb7H1WUrsH2FjmysMVLyNEBPEgESiWsZ+AIX53BuvX5ZJJiyoko3W
q7AD1qH9+1kdFjhKbdLbS14zBp3C+zRsLB7sHwGVuloOOMRV45diwpbBgZCdFKzbUgVc6DWm/PZW
I8laX6OHD8tjfAsxnxcwWCWvAjqw7/z+2UmuIfufCboFPcDKawitWENjcH/kMYb4rnMdGP5BTjty
OYCAOdEjgMTl3ZGFBOumPAlHkQDioASYpQ/0W1k0HjkslfqzYWa9bdiAC88gl22Y+8z2ic3om88w
UPZa8B4V1RMUK52mbi61NKP/H1mocAz986UHNmBRv0QC/eGS2spIHOMplGaoxWjIiw03U3zwVr3Y
xIQYMDjUOuSXYB8CrKYI5F+Ga7pRxTD/sX6a9PDPGx8PMiaHjBstMU7UTwx79vd6FGlsaiZy1cby
4wA8o4ReuKffMxdEY+h6EoIna5g18sxP+TPh0XBJokBijmR0fBhdauFX1doqAe2tWDo6+lgBQz87
SEGzBJO/mGAO+pAEt/p2d9rUAN3FbH3bsQv13pYSBGavN3jJy3XRbBEEqfCJ99T3LbD41NsgjCPd
ow8DyQeg1rVsMzMOVGzXqfNVrXF/PBkgw8jr7VO4JwTX9ZLDeDtaTjqEdljMhpYVdAXUCUOFMq8y
S4FGrveQyWRYS+4ODopX8GVBT9TwjZEQjjXwfpeeI0pXUBtT+wSS5j/hpI0nIFqzwTZLf1xIcpvb
fbolrjclceXIJ07bzc4HCOo7fTLp0dODvGqxYrGNnSxOw2SBO65oWd6t+UAQMAKYKTLNrvqdtE7u
8StLkl7q7nH0S94+yRDA6GjrLSqIE8tzfH0dNrPzqiiLfCaEAXxdRRj32iAc7Rwopd0VBYu+UCrf
u2Qvo1nV5fWdMzIOx5StA41NIZ5CjhM3Q7EjmUKPwdNcgyrM+JXfaJKp3Q3lacQHqRQISkSw7a5x
bLo9cKYk0cHF5IVFa7IPN/NVozG8l5wZCHDs13iNz7ESswckwjbIUBp0onT/MBZq0enAS0qh6Jfg
DdTfh8TCv5NZaF5CIN/oHfzm3Mv2DG2l0GO31nTN9lEIxpof0GwsgajYbKeQ5owuhWkYRNfZOyJP
va8/JI6S0pGHbuOBCmDRiIfI4sxsyZv25uAr2gMF0vEyLF6TEyJdBbq9TPQ+8S2I7hvGH9e7uzTj
s0/6KdwKXjzgzIHc6dZ/h9Qj4FzEZ+fgwl4aiBJW298npRQmSlqhUp8mS55W6/MJVBcspMPuS51y
UDYl2/TcDPcXK/SmWmgoRWHzInvjqvl+0JIVOgm72o5gaBPZAGdmSph+8sMlyUnEsMXP+KtWIp5a
KzZRoI9EAcE/bg5MKXdoKpcMq9f9qaVNh29tcZZ09cPaSoacweSor++HSWH1yqcDqJ7C8DCZn6zp
GZEvoopxXSg3QSnwgfKXtz1fDjefgsssFtu4DklRGdu8gVs0+5U6UOYW6Iwb5pjjM6qdpiMhsP8C
WHmbGGn4vS8AEAC12Vv56kwq1jhdbU6Hg7GPT2DkpGWuFZTwWu2OcaejDimlsCh69daCTxnMfWjt
pEWf6avyHIbEroKe7O3xeZU7evI5ALJg5ZDnu+YgRiibXMrujacMKLZ+JPvBSYJp1YrjqKzLbKzR
kJ2oRZyZC3WMXJbiPbZ17vI4ykkMWRKMVnekkWJgpLBeQ49Kq9YGv/VgYzVeKU6Uq6f0rJ9zfLzw
7yXUp9VJT/zvD0Ujl8UzWIJawDeRyKLcViU+NwyOdX8trVSDqvYHbibf1ogJePcTZ+wEyQJlrPcQ
Gy/yWwjwJ20BeMbllasuv96J0ZgbOB2jdkUmStbrnL4bWb3N84GG04zPeEQ97y0ZY/VjnGp4D1tf
gAiXa9sgFTiE6jWt2sn/hQfbgJGZPZ3bHj7K36PQ0yjTHOfYoqNxJ70J5OldNgqH9DzpJyzgZAhY
FJDjA7TYwqF2aiLv/CZHO957KyQcXCZ7QVSNl1Wqi7BMCVk+LSmhjzrIIPn8X+1t8d5N9n2hhCEX
WJb2tc2LeiPMcVC1JWYyB8Zi8AdHjxQitoD8CmmeuNXsJQH9IouK3tRXv4Lrn2h0nPwUkTBuE8oa
19ib2llGSvOloQ8nIdipoUpCvYryWIB8hiwu++Ekv8XQlVgtvRa/QyuhlszXsvw0LPG2bQJL3HwP
53MvYNwdbwgcqdT1i2ES3Fcz+lWIqaUaTLLpfTVdNayB5LENxTY2YBa3H8HeZrcipvtncJkKcDe9
1D6+hTcvqA+iIyxC3Ic5VOs+T91BX0OGEH2XuMeM1Din1QRmu8K2Qwl5p6nPuF0RJg1WYvxeqqyP
As0y7Ccc5BOMkk26BGMjOmZqvjx1n6xt6NqueuQCfrozAUPpNHMbSbqHth+3oOiHR0GQR3N++EB8
BPiErGK5z46D2G6QZes8UmOA3ICRySg3VFQLDduLobUn7t9bvvKaqjkSRypSxj4by6DstBdbC3YF
V0oMx3bCM760rHnKfMx7Y4ZFDUUnAUVea/2dpaexSFRH2cJHI5GE3wvjezJipYdLPM5veNMvBjOG
kp4/VlO9K/JpRBC8CNEqyRhlg5cM4gfBDZzZ5SleSUfC6YkGIHtclKV+4XjSE2S9R6XeybkcPG2H
kvwp+W8Na38u+jiKEUWLL0bD6PzB6s6FeWtUalSY/245eKpoT/xTsVTDS0QJZ8aOZwVjlk2bv8jn
3yS0EY2dwdxehoQdzTcO77FD6YZrWTi2vE03V2zZDrZcvq1NkuL/6IWOeQyecZKDlWvBvaQqBem2
/0NinU6lzjuQruuJnFDJlxmjV5ajylKcIWOtD2rUZaec3LDFAbc/BToVLo4x1pNfDE2AbHdR6VgN
bs+1WIRAEBFehm3uGJfmRTmS3xm8hSJcQq0yGrI+CFmN0S2LpSqSRPqy0dnef3O5TkyvkWw7kOQ/
due1UiafJ8JzY2j+obk/cBQ1O70tm4vxZUWFMX74iRlUv3y8//K9WQWL7cyxul3jG6KVEoSwW0Rn
wXiM+Do8ZYEoRO17hIBxAAuecZ2rg16xgq3mQh9YVX65WQpp72t+R+4dU8Ahk4ViZf8gMk5hBohW
nTxfpTSm+VOIXE/onP9TrKeDvNgL0A4d/WYGazrEw0uEuZJRfjTy1xKNIWxvzQv0hZFbFEA9yanX
DJLRs4LB3s8t+7KEsAZSF5B7waOHftddFvGkGpnesbkjtSu8EJdFgj4EWOoFLZ489mOi+vUGppev
hsqdA5Gt6hyaGPPm1NCABNDfJ/J3D4fuYWIyDodQxzQ/gv1NzY/bsa14Xb46BYzzemawJZye1RZ0
VvU/AhzPbbQ8ESHqonClnESXeKZVB1Nzv0aI9Xj2WeKtj6s6rXEKZuiNzH9gz21V0ouxpEe98IjC
OqofLsUHwq8ABnDhZmoQKLdyPrl8b8wRaKaJYh6uwSxUJfYLGWorUqONzDLgyfjOyH0/HPTdYoMI
zy2f+P2D0tA5ZZvNqsczkMzYbV4Ah5Fmhqe2qYlNwmKtYGxD6EExNQzl1QI+rjRGCnrDSFKQ+uf/
1hamCkO9KqQlDSBrKFqgy1J5v8JLpznubWOG+TKhi2Ss4efnRc5gJ4ugqrtWRAIZhod+FXBku9n9
hmi086b5v9UqnnJaB/ZTJ18hLNZU30amEvLrwGfo7clOcB7diE7aiAB022datdkyBYV/tbXq3xiW
4DzR7RKeMgfSI+C1HKoLPvBoIu2zFJPasS3GI6LNF4IwbtJNF+3MUnguLfrAK1cvaIFEkk7vNQxU
mdamiJd3v4dGBb+/sE/uOgLQ+Pn8pX7IQj81kzDvy8n8UQTySat1qP6qx4yvnLksxJtbAEvXXVu7
OhCzKAkUBhvDShWze1oZyUc7i7x4BcA7MCNoNMLZ4nt0dTe95ae6HpNnXfO/jTOF9KEYIFohvrJb
rRY9WPK+LcIo9jXc7RJvmTBni7GuCDYx/AT2hDN5P87OM2GUqclBlT2nNH5i1souAK1kQ+KKOEHq
gfF9suA79iVd8PpLXe3J0eIhl6ShNZXCfKXTybYbAdvej00NkQ4lJivhKe2+nDZFDufC1X5mbSRv
CnZNIG0cN36hFTuoBeetfxWzI1ejNhAPQMu1+KJLugUPhLyqnvMGolUfZZahu3Owljk+S5etmbDf
OVq1HEU5ybtWPb8N8lGGw0kK6Iykc575bv3ebdprNViucAshmCIl/alHc2rrNdgpGyUGcuklc2Z1
OdeYGFmxX6FeL6Oq0LMuU5L/gGtTHhM06mk5HJEpqSMuyJMbaMiiKZPt7ZfiIcknZsykTeCOpafB
h2RVed5OZuGC6Jttd/yI41yWv+hyMj++QI8J5TJn6kK2iGzu6pVGxNy594pBAGSLS27pzmxw4r7f
MIa1YfYSwnXWsGEzd66csUPaVGvDTrG8NnuLnvDOVRCrPWkNqgIVJibNlt2DYrFM7TTUd1fIEkl3
dJfSEqzaYVd/1WxheqjZ1fit2nzM0cwUvgiCAaJv5CqsHlGolkpsCAuLBBS2o/30XzbPdno64QAT
QHHXIkLNwEjrSjudPxSBgzCozidXeeLT8JNbzH6+QCW/iAQ7JPWkohxNMhT+JgQd7x2DVH4ayv5C
ebGugkSfR8Yt9lDl8eItcqjMwupJ2XA0GoYTcdyBMK68itwxr+odJVQmmOtySYP7fLC4E2n6cGIK
fVB8zzUhFb1HJY6g0trStHZXFUEFm1Ahq02rVBvRri/rWRcRzVjxhffIWJON8AW2oxDGjsX3DvFM
rkG7twgIS67bS2kJe2nrQtDPohi6EuolcX4C7Sxnro0N8NklqVEkBAKqyBcWWJs3XTQBSpPi/RMd
ZGrLAManYnfpqj8xptuDuVcp2fGSx3CxfzFLSrVaOkrWkdG8aywNNtuHEJJbWy9zdQSFW+xzVdMo
2wsGB0YGFU9mjzYLlxSZjhTpv9xyH4w0lr6vjaXLVOujSwXf1epv426pMETfFbPTu0NBQS0UZQ0S
dOPn1WrqOzPkmwCWKY2UZvCF8WyCpP4D7odBamyHRjkmDyUaFXIl/NJKGG5peofR4Z6lMd6ogMU9
IaUPLc9e57y1BRp9wKZbGP4FBYYOlQjS+lVt6FUF2nijQytjrlHs+kNdcmeFPG+cFm4HJUzsHewQ
L0mKBCD/R4bnl6s3bqEbQ7b03sF40m6wiqzKHLf2Ckr2cEVkqXQWez4pEZi8SCI5+xj0/LMIjt2z
E+0mSHmKtDQ6M5BmO1QFayo8K4ZFPxirwzFEw9lX8NryM8o9D1f4U3xGrNHti7k6uzyfL1uZtfTS
3J4BwXag7KF8E4raqIYg66NT9IQfBzfGXHBrasqPJecUzI7UnveWu5NcLzoW8ps3XR+ec3yigGIo
kDhRc8+xILa7ZhjRNKzdoahC6wA2ImUGTrFKgSdedZ2O0WxZCTVS7KVPmFIFsKf5/Sx52YQ0Mckx
hfqbzkSAIgGgtbdSW0SsEOQonnwWZEzDZ4fPQUZ0FM0ODTnXJsDFSwIw6ltd0panm2xboJQXBlML
sUito5n7hbmRJvDxm51do4IMShpzwf6t81PNbfUFio58tT4HTuOUiTVJetFFpFQqYaRqCqLoukpy
2nD1fNMYglP7uZ2KkWslQ61m+z1jd0KEYubiKiUqmfKF6QdVY2Ajy03NV4Qg5DbU7J9ZJM79+yLf
Jl+2AXVhld1yCN8+9ZTmvWdPLNSPcGj8zMbkreYETe6BMM/527yxu6TTFOkCGENm1Jgn9GzLtqak
Z3sRkKUbHZ0NoAAihsy4d9+DGKaZNX20/QQolh+KkSk/9S82M4i3Pm4xlqCugOnC5PImshgz+7G+
ZPHNxNqxJCeHn7UPmF1P5yZGyCbQIqArt0bSVUzdYxD4i4/YQXb8/1+Pk5Z0OV7tKPkrK97c8NNR
SL+ng3POyKuoIbJTqdBSK/ESGsJ3cXzhDm3OJpq0mBKMlo4HjhjqAmiANGwJ7txZQnvobb18Zg1m
1eX9T39wDzBO+NdJ9Y6kAzwQMGaKlFjrYagctnd40m51C5pb+ey5DH+Eex1fUOmKENUyBUkfgu+F
8CTPf/HSYUoGF79yPhFw5GQOM0wR6n19JBckgRXZGwgz15cRZx1bXKrpGuuTxSlVhKAnlhIrmT1L
MDrCCFks/l1a55fGppADAMx1qKKkAA3yuPEvPOO7bB+IQIxVeVIEqolkuuKjjNYGx/pwzL+stM5B
lMmfp6WprxziMWwQvdWLJVQ7tqSUiiQ3JNHAcyQ25PtCcV0OzOts61nUJMRGDF2nZGfVRJU1La36
M8QMxanVkaZBNTq+u6j11z0kiHz+afSDMUcWl2BgQYNIt/wPyxhcQ4gTqRzFsoVWsZRSN2EqfoLj
aObflJo1k7yvfevQ0dre9TEs4HSv9OhulbIKd+XYQx2/YWZY2DxiFo6uVUCZwH9eNq5nX9+9mBEu
cBBpoQG5GoF80Ks1/kWUTRTxd9fhL7vKNczTXUDRIVT3hzWWliV1yC9szQ4sQlmioP8AugMpS3hu
zPCOsy9jA6b5XDXaSvWNukZxLxeFWOKY3cpMTGQKTBVrzCCNULiJ6hDbtAqMmZHpw7LYNKqloH4c
eFzGyhN1gAn9bT3CZjsuinfWmZO0OvXOcQzd8v5pTv8G6W3IFr1KsHRVc0PDD3OT/Tgr7EqspyPa
WlkGUmJIJejIC9SL4GN1HCYjiQAkVsGTRRSis2eBLU2a+T5/JKoUQtRYLkg4HgCK8vYivNtV5u78
RM8LaKrrDuK1IfpOk9636J570EuRo0i1yXpqQn9SuocyUKDUgAmeSQ1OaSHsUXEc0lZJJ8XNYb3/
4JEOymnrOGf4hvZ+AuZF0c1BKkkSgVYH+QVDbGIoILG0INbVkmBVku0hoZSFnHPsSTDTIh7GV99m
1qpdBkBQ2Ccn354nodBBGFM8h9uhuYUx+hJenvAg/Qhd2nJDhQEiLD23Zia/0A45hSndk0QiPQ/6
hb1C9L+yLlY1rs7tsvcGz7fMaAQ3ayPaAUFKC9ELaVnOUKH2Zn7ZWjkSwgjw5JhDutJpin/3v2b1
djxoSndi4v/swtJ0P45FA8YDUUJ0iLMiqADjX3PF4kCJGdI+4hNiKKHWsa+xWLNyExmm4AZ+IPME
aqTfiZTFJEsSIJu01/Gy4Yz60mfht5VSjrY0XtTBMaQ2VSAxpA7InIKQQxz7kRg97QoDY+D8kE55
IQI8m90sOEAeyPSsV/rwSrafENV0wQSuV6x61j1EUkd8FsdGJDlHUAKaaztRTtZcpqVCql4PBuuz
cGDKlcMLhFJn3GbY5Rnx07bpBCNv9yLVmBLKhE6vnXvLyIF2FTE5raBTMyUCzYQxYvfeNFXSWo7N
XFvlfdYyLjYWkk+aeIPbd7EycH4LyzhM5+cvnAeMoHDUNL994YnQFQeMRJgaV7NFJfdLnfRN+g2W
9PSl5LULERmtGxwPlWZeyrfLHYx8+3q3tjAfxoLp+nF3EMpe9JSrby0B+rREmRmXl4sfK1Ccyd+H
iiC9iT+sR0QDgm1qE6K5FSP/0YYoBJ5rlMWq3t4eraaFITuN/QBucybts1u5jsedQEvSzQk8RISE
Ip71D404pE3SEOWlM8Fh2xk9hnD2ao/RWkaYG3+Xdvzrt0FvNYugvg16r1CLWzbCw1KA28ZS+Bkx
M43xbWOrG2ixrs66DLCwLpDyp4niZRdHy0OQLO4Jhu8ovO1zPfOY6hv53ODVPSmqtz1bzFzwIfHU
vxjtHzSoIuF6GMoojZrWGp4J8DKgsihQC7/m+c6Q9YI+lyBJD8zJDZVp2pMqoyijufwR2X2Z4NyP
NGCoqcMyWV1fAsKw1JW7LRnC5uLXReUTa6oILRuQoDGB7TdyIQPO5tHYWAfX8Wi9vEyCEwn0UX4P
103raDEYVBYAkWCh0snfj8Tib6QICzx/KvQ9uN3D2H2rYxN9JlQv2Lct7j0Jird/BLqSzNUq7DK7
zqC9MaMbadICzEa07uxIKK4fAp3DY/kwha2MdP+wK4Akl9VIDQK3fP3YpIhZvKd6+ydAO59lcsm6
ZB1kD87ldgIoD8SziY8+o4MShdudLj98VkBY/gd36WZ535fJXmU+kHsJLUSrcSrV798wyx5NHZEB
hfH+rs+W0TlooMt3Nb16sJ+EH0/j/Z3Id6AplB/2cpujOwS8CV6cKjqZhD9SEGcSA0dkNLt3pw9O
aN5vQquYVIHrhxr/xi0SU/lTEWMnvssxNiOPGudJk+rKamYoTC/pPmINIKtiKDr26cTyTMmOF2Y8
OWFCvFnGdb27STtoO1Ob4/nwN5wUjhKnGnJEx/c0Jylk0YXo6Aq+KD0gws2o7ZcoVC0mRe/kzC5f
Jf5WrNXBr93G+6atmEDJKwdWmWGPEfKi1HoTeZg5KTLz8yjtuW2ozG+DLS5so6Xj5f6T9Oys6vlb
X7gE43QtPnzch3VqrNIgB59aM/Qu8UKtHjd1UHzknW5H+yI3FYohUuWF473mBd0ItPsoifBYjCgj
BifbePKoBuaML5UXu7/w9gS4qBVLIPagrNWeLgMIrucSgcX8ee5C/hda76N0RGA8xn/JbFq7TYgl
bbmCmTXDCS90/r4F1v9EaTFqvpC0ajAyFj6RAtMvCdFlBCfowVMwCLU8aHSOyY3Swbmg9xpwpRuo
kMjwdunU8egZUBidTCC3NofyX42F5n1tbfr5XoC73V+7ozUIIX1GqahKcSXbIt+2x2Y3cmK4r2cF
AtmPGroeOyF/UYNI2SxIAn2j/+Pg93tab2A5pu4sI4bQLylIf4zZb783V1mZ/CZy7oknSL1QlIqp
ytVpBAwtBdkMGf12E6Uh9ug1woBU0p4PFXIGI0SjM4ZDa1+XoVauJUHO/IUjac7Av1FgqccVYEax
0x7vbG+LLSUegaK6S+/hYaWSZiBXTn/2d+TisJuZHpKoQ95GobyAd6UZcF6VwQdtOt1gSwF5OrhL
3R5ZbTVPGi6uNCZ53wLCrASlRbAXWxX+VlzEQqFujJqgpyMuIjrY/Cu0ZlZugfyCnfp3nwsvWM3J
bhpLUMLbsA/puj6F4ueKTMjslxzKY7LWWePbj9fcmFdNwx8ZGxVjgqPQYCqFknX5pMqeslH07/nj
KQ/c+QCuu6CsJ7Odnpqt1Y1K6FZnPkOOA/+yvqJcjcJgP6b6dtuOczbJtSOaVktAGv112NIWslzi
4iX3rh8wFUb90xauxlQhJrCzsrpBtHkgtN/Tnl7hL+laMepH9Vb9btZuLNkueWwktqhaN3QGZGL+
WYk+5jKki3BCsL1Yw3tgk1Jt5dDXBrcRTo5Z6fi/jyn1pP9BLAR/F7pqKHeP4YGF6MPTnpXkGSch
vhl5pXEgp9FXPTo0AlSUhJQz/sWoD6pjnyMmnQPTPs8jN2/rLxkY4kMwnnRg4r5VmSl6FGvQkgDm
LlU6CxmjyDCqdeWfxde4cFxer1yfU2hGbgsM7Je1pCOL6EktnaJLPsyNaSRecxHkmpXy3MXfamHO
LzIBST5w/vIMP6fta4txIVZ7D0NtvEDT784RGgYpOJAYKkjlExJMMowGFwZ23gWAUZSk64kKo2WE
+Y0pMarEcL+OUil/HtOEnEE1NjtV7414LMke23cqsgD3jbe1GS1DDJ9k8g61bS/YZhw4M3N4kC78
KrvXvBPWgpce7QLWJQ41lIZVi5Cr4eo4ossAppCgzfalLLFT5nd/NJx4bsEIEuaNDFQI+6uH3jJ8
OUEiTU1A4LE1JX57+6lGvZgxrpjWsOecSdwsS/dws7GJv0r6/OKcc23BJaZS/zihb9YhEcXwFJtw
8J3w2+EcomTGa2dpu79wbsY9Mwi7fPfb03abqqOxf8LuM41JcXyLmqWAXF7Q59sLnwsjFpm/38/o
22oPgQwdevezGX1j2RVdi6DVUzy5aiYsTJD2R31UHuZx7WxV4AhMOtkZKxUeaXd34fb5sO/tCDuK
2LTjPt49IYWqsLsq4iat/TSJB8X+VIt7vm4cpeRZhwt5dwRlhcKSVXSRPsfpBT49KVvlrI4X9R4u
0qymuJjdhreI4gbUa4QCyIUEkwTkscAiCPojTDMcBWKa9iLub+2NXn8olJ+RBDsyx86Dj6dzq4Ga
pgNf9PFU+vbzBmvz2TLRgqQN1CZ7vPkm1eCbfYNeIiwkTX1FCjjCOrIG2onV+NNCkJqOGfgD5lSz
3KZgWWn9SoscwIXO3r+kPwrcTAm+j76BCc60yg/Su/SsJ9iNCHPjBpr4vHQtl+sw1DbCPtEU44G5
Q8287uM+hNKunxxbsn/WP9oRwlXPEmY2LLbceKRK1nQGPcfAxhEPn/6S9+dRVlr2682W2k3G5C08
n/zeoPNE/WL/RHAdvAFKQTvnYkmP3IfyItwZ80QtieBhI1bkOnXUVc4gwNq1XXBlU+onxkbYt6oN
VxbySw9ShnNe5j/rFFcTtLBzSrl6OiI9uo91rsLSGyn8hG+0epibJpx22+EpCrtn3/tEHjgohw1g
3gV17SfOVa0Yv8TARhtiuZcq1pgZBwM+OA4TkLtZDStF20F6avJRVl8Yz0keRBDy2d/1cSm6ln3c
4sfQCw768AuY/S14ls2CJ+aZKt80etkBGFhh5f8eqwnXnqwnlk9IOyf8tI9DByWEYM9cK54cTlfD
/P0fgyg9ujdqiwUy8YbYRRgfPZ3SDAgzkaq8Gq3Wl0Beg5FrKhfSgk4cs4w3XfNeyhSUdB8Vvdmt
G/CSmuEwPkKJsfpH3HsVw1Z6yNUrSf5CylJ3Q1PQxur8+PULpvzFCD/Hnp6PvZetJaM34s2iuMRQ
aAF+9aIWfqIJkXC8Z8Fa6+k1mAhnQpCb/Ja3fZe7fJLRZf+g59DV2HwxwAS15BFCKrV3hkYhag3e
hG8T3xlFcI7lkUBj4o4+mnxwMHtYzl4bfQZvkaDRRluCKkrlCDQOBzLJFWg9wCfPYtTSg4CZ5CMt
O85P2kwfvIDiAYqR79iAun51zO/ynASYfr2z2AXA95KcdIzmqa7QJWvpKPTCkFdftlXyW+ST5bv9
xcOlC/rVgnLvbowNZi0Vv48Nfj6aHYkHR/G7xmWoPftWOOktFxyw+6aOxw9An5wUG36VSvD6ozlA
vjhfl5iu6Z5H0qZ9wJ3tmNdyUFgnYUs+tY1lARa3leTEsj9bZsL6zN8QSancuzM7DbWqsKctjMlo
RYqBnWWQLKkLWkCRgP797jI5L2raQjwqbZ24+XPc8vY/NfP3wyxkgRdp9RDB/VnZZnA906KhhHbN
Zl6s1otN9J6/E912Dv9S2mllaS3tENZauwvP0xNC9pAdFH0EBtwLtE462v1efOL2x1XJmcH4yrg4
R9LmFywGma9toP5n29PTsjU3Y9iib8yfoyCAOa+aaeHHbjRqh03MUGXZgRg/sd7oZcCvOnqnG1wS
/IsEEEnbvo/Qo43jvMOHntrhDBZhQqUTz/Ed0oxpbdAGlNz2YWlkzoVXi/UY+7ksLepKgFVb9eYx
HKfuSGWqAVx9mj4BvTU0Dp4eEFIitNqRYLlHWGcxiSUM9zM92ywj3+c+skbJO66G/MfjgxoysslC
JJjGFWfzQ7jRUQN3IOmsome4JEz3HsdP4Pm0DYAg65mpSoelnG4i4biVaDoz3Vp+HwJZxJV40slv
KOf4Gph2NQ8xxa0iFHmr4stbb9Vm8jZNmnmSWgC8aQgDF17q43vzXmjD/gHROBsa9JSUg6DGLw41
ZdkSXDwpZVoQpWhxhHBGRLcXo6wsYD8XaLmI1CWyQz0JrqpO/jZtalrGpOVmYu1ItJb0GC6VQZ8R
hIjvb17N8jN9a3QKx+g1FeHOpEb1V11fnpqbpc/EtFv5yZtrsAGzkk0PfMtJH7iyIbNk7mPD9zPD
pnF1f1PuNuysHPOXMvsw42Tghp6WpHfjtpjQJjQasz2UJDsfO85pwqi1SkXJWPt1VHeeVM0iPmlj
2TM5jPIkkZTtHgzkY74LcfhUjwIW35sjrwQF4MPUXK0BhbLMhYNbC4eZK8fcWNccQ6kd8ym5U5nF
1+T0uUBr69hTVcUdOQNYlDqr59oUnCOeAx7hOsH9oQ7NCXpsxaknyFvw/jpPxjNFzA7JKuqt5Z7L
GmuG+cF6nm4IqiUen06dYm3Zq0XJcxsP7M3YAboIko0O3H8mgKms8OP3n/c5ThZgD3s49MvDXO2v
/yTor1a9ln4pJLYuwwv275pEEH2l1LgbXs9CiiL/b2nGM57YSlAaI5VOj978v50oJz6hscNnrDWU
tw7Q1U5zJDBuz+rXq3DFIVC34y60Ryvwb3h2d8+pwBmngl3ZkUyDImooMPuuHraIFeh/WRLJTI6n
7P/MTDqdNEYL8H4ORIpV7TnM3wxLyKWlvXr75E2jIfza+bFWZEbzy+gJy6Zg1pGXNfXBAhP5MEEP
v8rsS9cUeCH+5ZOPymME7FcGTsLzlvmA2r8bxk6se62AATA1wwiW9kJjbfMxCLkWprbRkd2OEAM6
6hLy0zue3rHcfY8nU+bblBpylcwGkB6foggfTKIWflGaHRJbJaBKs8bVM0XSGp0RhVNhVygKbA8+
jshajV28o5OM62fE5i/LVV460zb6U3F8y+kh4T3E4/Ldkeh+Whji5STtVVnon5HJ9J0T+m5iYorO
tHRNQAxcqSQfDoAe+/K4kqh/EHRtb1zkAVqYkFS2SgLoTsuvYmXSKcPlA8z0WtpfGOoEvk6m8wwt
e0p92cLUE1s8KGHsHV4sq2TvR5IpkF3ZKoaortKEN59Y0rS05qktSZrey6PRulZasoQYPdU+HX9k
tmzI1WJnjbRxBJqdHnhIkAGoXcU4Pv1kkFehTFiek5vuWLBdAHufIF7y2zDp5P1LiHUh6TL17HRf
kEtEkvxgcriw+C0KVpNGlXRyvafTNFPvMPRnadOKBI1rrDksKiE+rM9wmVS0t4ayXqJPDvbCvXZl
fkRBqmz4ZWgHFAXZFgGKHwibomh2R+UBS8WlujrBuR+ueZ6A3frflD7+PSYdbIAWHFlNGLRGLgmz
WTSMw0KRs5U9CLsxKDTvK2hCgp8D9OwYf/ZfP/sWf4JHFcxmRN4HjlTeP5BZpRmM8h7yLPur+xJR
dfNz7ic5KtqQI/RstQ/h5e+bTAgGTt8ncz0OmEYvXWlb54xgrvvF9i6TkF6V4qEcnVTSClZJvTtJ
YR6kE8CLxcZQejTguyAjZ02UGyPqZ6LChQRn3D2je9RhlwHXSO6pSXr8jmjLrkglyDDa7rXVecg8
f0dWafJ/peZvcc77R5BtVCqFl2mzkSCDPqlzQK+a9FdA/UWhH7Dl1nnZFIhnbfrYNWKRzXW8+A9+
DgEpPWaMeD32jSS09HdNwvlRjx/pzhiFkNwXLNX+ZWrNzsFes4gIOVckeicHyODIpXf6zZjbJ5t5
1weHypsRr4pF6rLIh3g6jnFH5GVxm/IQXEYDiuMxfEBoGru0h3jHBol1s2Ijrg1LcIj90RpTlcZa
Scf2QvRUWqRbHOjoIsYDH9xO3qdBY8zx/0fa695P+54SqOrQGn3AjVxaCyDf3oFamOe9FSk+m1L3
kt+pjyncvzABSJLUaCskWn6ke5DeoI9nn1FBC8kv4Q31AEjrlWkMZwPfwYuKOwSxTFJ++7wEl2ni
UKiL3qa1fGTbOXgj7DhTBSR6NdAFhcG7lCTLBMOLrsnWdL631VJjaKHD4Gt5yHs9Q62lY9WB8Z6h
3PDbzi1/+YS2lpyzGp4FoDGjRqEPHFisOP5DE4MozLg5boxi13at4TWYxNaXWa3ySX7Ey0IV6cV0
iukFn++Kz31CZfxq5QT5dl/FckfNwbkmn20D5b49DyfbJwH3t0kHxggDkBxBsCVeknZAmuYTnehY
+bOQVpRmOOQMHbmo1oW24Ve2bYlJE/hfQX3N9dRGB5DwWuPln930vh+3h8XQXMCSCAZ1UeVJXCrg
eyGqsvzT7xTO5r8z59VNsutKNxTjY7nlbS6+eVUy+pCoCeDVv38fmCVeqm1AKVB46n83+QwU618m
ZfFn27b5nAXA8a2IyHTb/XnJarubSKC38O3L4QI0e9rGq71S+KCLYFnIB/abl4bADykrAaCRTaRh
Mka/MoxPXzzyCNYALpFIrqVoX14MrfvNJUW+K+LadC5b85LMax9ja3CMLX4P+QJblb74ZokzVSFo
Yw+AiKY9tO/gisacQjlk66LA1uqoqgLJXaU9K9bkv5dyRofZOFMRve/sFgsQ/KnH7AY8aIuNVFzf
kurFisnNE01FHP6nrDugmAKIw6s4Gpdkrd1MUAKZNhrCCBGx/dTXdVA3HIk86lWoKfvvi9L+Yj8v
vit09Sekr/sdEqiokaciEsxrecvyvlGuD+g1R3dDAs98k6jAvfnGU+gUW2mY+kYfpSJeA38vtUIS
ga1okQjBL6xXa6GuBQ83fq8BfZfTA3ExzVtusA/4IeJsFK818V180rpGw2MtKddxYalDoGDZfB5w
hxg7LyCDv7nysjxaz4A+S01z392lcUIrVnISDiSEglWiIoBlUohBrwUcvXeF6W3W6G2MWMlCU06E
X98BBo5YMwoRqnnO/CRBh4OFV+LVVcHtBxjxGUyjtrmRA2G0ddJNgUwW/GNVvXJ9cr+b4zWbBmX6
b33sYXXYZZkqA9qcFC5jkfCxMNUtGDWtpPpWnHxeWg+OW0sICfTU9N/fVvFR/ErcF7gtzxJQO1z4
Q6nKX8K7doFOLEKCEESBVussfYJR3sEKH9OOlpxhm4qfvqnmYR5JOmaYfHBy0p/rvJrOCUYUT3QE
EGa4ew5NKjgzlGKPWGijPE/qsC7l+8UeyDrSMX1gWz3pRAjSvIwdVXcMcyJfHIf7qT2beZns8og9
RGDvqoUqIY4B01CYQR8aQGxbJfysJ0pbe+Vl6/2pzwfzfs7/3gBbVBaoYpNt5iYLQiQ8lrsYDaV8
3NT0iTSVcx+jcV/ImIH6NP6sHqpr0VCe8ZN9Jv8XELzyhhzIAOrJ/UjKZNOqDaXihy1uH7kG6NnR
3dpRJGTy1lTHACjptVdarIhOdQe6BLSyj2+kN1BAVTWnLjbLGtYW2+raKGms7GDCqRjzhecvnyV1
FFjdibIO/i8mEBg0kI7nsLdZJjeqrKhWRr/3eiOOOzFaVl6FfmbYKsV/b8Qqk0jQGEV3dhsvJ9yx
1LMG0UkDYeCOhIFjdsgyeA7QbWSEOCZ3dRRZ+RRFMmiKoFkBWufR6myZsf9P8M04+ZpvAFE/5xJl
n3YfHBxNTgrWLEtO1sC+ZEZpsky1rWA3oBb+FELbRB5iijsJXuUYpSjaXh/uELEFQFOrGoN4Bh58
3d6583bRwwrIShVaYfYBEE9qa5sOnfERfF9G7wZhWvvfSUMnd6CFcivBr8fWh6eT9dwXtAhWYZPH
/Idvo/eq2eeY5gYld5T1N0kuG7m7GPm7pyNiuQ0Ytz4TX7//RLkhuhRcjst/Zedb3H3XDmtMiI0b
GaAcRUsM7Ns+Ff1zgJfeA6JgMAEz6KJOiPe1HZLtkcB6ncxJUpc+Rups6oFlONwYvNKNy8r1gwjd
g6v70q9ejMJ9X78ide5qh2zn63yQQQNDmZSG0y5HVsx+V1A4dD8T3Z061zjIlu9gXQk/r2iIL/hs
SvzEByrwAyuUayJnbcVmsN9JU8NsCKI2GJ/n1xqi+CmFqlXVP29LykOh9Oxn68RfolDnQU8V3SnQ
JLVbmSYu0nqWNmaC8f4cio7SxUZBJwnBmUsD7okXpIy1vyWCJ1/t38f04OwPiAdzgNeJHh0KLycl
7OGBkajEa7iEzJ973/fxCIeqQRlr/Fuw8AoA/d1T2jKZXC4Px1JSeb3VSxezQEC5dVrJ+AgfIW7i
yyS+lR16PpWAfK8Mas8CxuGD0d7v0REXxRfSL1QwCYmNFxV5WHAQAVp2qwMJxzZdJ09A61AZdPqb
MWbph5vuGcaQQ+vqfTmmIBk6F0262rfT/NPZmv2r/EXVyC/bgCAFdh2RiUvMGObrUOB7uKu0ytKM
FGFRAelw6COZJIKOsjam1KGzfXobHL3ODkQOrtZCbQjlbkUrR09CY74O3Te0GG1SJynvcu3Iyglz
tZPe1IYSOAb7BVrg2oeUIuP5VI7llf4HYlAwHyVxy5c18dP2N+gMUzMnnpqG6WeHDvqaJArrM3TL
4ptib/mFOZ5d4EV0VySGc0DShmZMBVS50rVLMs+X9bZ/Owo+ABmCsO6ybPRybqyUu3G9SNf0uCZI
0k1GYw9WOPKr88dMzpZHmZRGPUcbd20/QYGAp3X2Gw/C/rajx8bUDTYacSpqS1CZXx3Y0zRfgMMJ
x22PYBVyrlpy4di1LVdkzUyEEK3GkE3sCyFE7EfDSaZPbyo11zzj3WstdOkS5oQZggRAd1gm4QZY
M2B0+vfIzcEWzgnA2OyXkt7liC6FgmL00noJq4q6KxG6B6JW8ZZjR0TCVA4bz4WZDpnjER9V6i9e
tRY/4yr7nuP6WzWetnNTKwoMqrLSbAaiAobijXQuJMTiK4Nv7Bvl22jOggIBIOynbSiXQcU42jT8
JMvqVYMxDHqSy4ThDW5qz63f/AZ2qKN4VumraxBv8r5AzP1rE39cA6qpYHOg4gcXtX6dUmKJ6EPG
tp7HGLNv2qLhIC35aqvuJGmQzRf04OCETOVJnlF3bQ0HamK2IR+/rKAFYiBpiEAdnEqH7O+1H2rS
mKjvzfSBBY0o08ilzGQn8OhBEC6vSkzwg3Pem5MrUOc5i39H7hdhxIDh75WEGXVqvtryOx6EwQz1
695i6ZYrOTlgA8ixg/8sueh5Jz0SL9DsW2EcK4CS4IVSwl6+Si708jU8QFWomWrFNmr43vRonb8S
tCVAnQXMzXC2E44e7ah4XhP5pX6e6/IyswZEjWUUowBAzl9trIwwx9XNfFAIdY7OsRGJ94BwcMLK
+kMILZ4ToVXCMxmo1vNsYiuX+Id6kL9i6uLdyFjiXMMF/s1kcNiDRAGTwZ9+EiEdc14DCgSkphfo
JbkpmzkE+ES9EdjxPjW1H6kH2S6z0RM7DlcgkdLMTsH01300qWO/Q5Ha6A13xuViKMtyBtcgd4+S
7/OEj4adeo3AzMekABcRA9n37UbMva9XNczwO9djR5Yr3Y0mkVzhac4WF3QxrQdF+ddEonQ55RGC
aDau7JHgZKXGh8a7bW/PCTaCaFkImy3CTZ4BjKdcCBoH6ghQ/rli6OPeE1CDJnN/dFPnaA+kgGD5
RS6N38YE/QkxrZl0PuaQwY9OrIPXAqWeASRY5cuDncLqK8RbXMwTfDMNCgEOeQp7WzgvAVRngsyo
p3ifAP/CWwHQ6tMRdCuVJgvTNUFGCt4QvOsO9+FIqVpZPKxoxFrv6BammqGSBp4kZ5K7Q1urmjyK
rQnaHxZzpigcVr6EE4NIOo1Do3Ns4t0t7sMiMQtt0q5SIz4oNmox9gaoONumF+LDNZQVujAtqPim
LcrsVo+UBDugmsvdTrTFr8JgxOKCsB6jt0KE04c1gcNFYU2dHFRUckTxEc6Yp74oF6AZ83z4hwEJ
1bqskEv01ihbFPDRaVlo2VPfPLALIrwoHwFybp0nN3K1U7idLaN7OXwS1OTHkVq0aVZhbzHh7JeW
r2gyw4ZXe1fRO0CyJwQmHTIketbO27j2/5ehGHexLtywVQtYA1rxcqWTC+7QrOY8ozQc4ZT+pNnI
UB0OmNJZB3NUbG9zG6Ek4Wy/LksyNLBoxQTr5YKyjheFw40buYvQw8LffOc4ZMl24BaRGwLoWWRZ
HSPobBjMVzg2FRZfnqBRryQ6BJe8hYcKIyYc6OVwvJgSQhUUp9Diafmb6ty6WF1Oo0P+/JPYrvD7
/x1QG4U/AP4Ur5+2Be++rY7EE5wYoKVTNfbo+eg29TDL76pvCDFkNC2L/spNF7vYSZZLKmMoqM8z
8tLnrqMs9PVbkF00Mj6LoJlYnmPbp3DDEwREgYjP+GpXrAJktGkcKfEwRI/fc1EHub4hvtxpdw7x
yF639KSv2QQoqdJFIpm/jjPWzeRLKVj/0DDPjC7/pk4aCRWOCvu+P+nHq3oTmLGaqVzc0JtBVO7x
a6oz88XYiq1zXPB4EqC1XkXPNBJKZ8TsN2UCNjsRhoj7kpqz6RgEAlvdeIx/4OWZlhb8s5yVshCV
jHNa8hQ/X43dfsEgFDJWyfiOzoeRzdt7iW/dR5VY18fs9ZNrtrO2qdj82JGOAodyKw4jmVOzLlF/
HaO55rn5awESylYfNJuuBTvY2Rko6QdKyyVDw7p4FjerCkSkPYlEUwIbTT5aez5h+E7KnjDOOrmN
wmvPfuBisR4TaJOE+B6X+D48teHByR3BHTNBUa91tbFwQtmsxIrP2nRr2sHUFsyiVQQuWvbCoy1I
algAjHnytymXZUKHuZeAWjyKUOXpF3Mj0gBuYf99ZeGVfLiMl7Ykg5XwP3nUizIzQxAC+uIRppNt
lHRdRw9nTHhgnRnkJPWuqcIhkL1MRwoSZx+SNWXhOLLkWDJFUr1lH8McokvPzbnoyjuUv6VKsXgv
ocvR3cR6BtQcWVExnEp3bu5kSnU28povovjoIoguUGlZvxfgUmDZxAP5nLklepjXU5qyjWsgOMb6
jHwJbt7wTocjN6Gs5UwbDiYDyH9yCCUK7PqnMuZdzG173b+sP0XrXFI5o6AqrE5A+ky6nPBnfoqj
NexeF8SUMr6EOK0aC7uESq2Kn9AkCoYRequdf8AFtOjJEpwiV9msYOI15l55mWOip2Yj8WMnwvQG
We6O5np2OtGbwA5GutMhxqzvZ/4my+dURoWW3gMyX+Z+C++fDqNUnOFew5L3zvn3+tUxda+NSeED
EJEThMJiuhzLuLZE2yqMt4lRnFgoroUXOEMS2U4cHd18CiOitW0Seb4thaier+bQTwEG0y2pqA6q
nCFszLJH12/P6p+/NLkzrZxx+hI0qbXW7X+hYatLhkyvQJEXR2y6LXsZAjovQ4cbQFewh14gEzZx
/Wdi5N4NhMq7NhuEjlvM3fd719ngRE7MAbMp2GGMZ33TLOqksB7UVeexVgMf1dcETX05EZvrErj4
WsZ/lhbe4oWLv9BvD/NhtUhewJe4zZzTwYu5LiqgVRvsUYrCvvdKaX7z2JknGYLuwfqZPj5V6huV
wNArdfuR49xRVSX/6PX+ORKUzx5sH7eDa4KcN0UeRU9d45vI+M6psi0DXJf4DsulbsGcAkqojOvt
VzZEl1qSilqBcIs/12SqzHEtYJie8RBvJ2gtenQyOJGinmFkkpksk6LoDd9eJ+74yCaQvJHeQ0+E
DR35BYiyhPBmG2s+z1eGUaZdeaYhZy9UVQRuLwlgxanzwQ0NDo/vcld8fJSF4nup6vav7h277Hva
O8DXb9SWKRWawifcSS28Y/4EYpRwnqYVFCBwzdQ66/HLMNv9svMEMlMhdLTdg5LHPUoh0yp37qAN
d0eWGr53PuG+fyGXdsTxVjsPJho1r+zzqoi4JT+hFzI7mJwEH472dT2ZVSHdvQo/w05OFhTHKwNd
sMwZNdQeFroLdYJ8KyheZ5yHRrskaBBB0bQVW2RpY+sdqWhZzUknRRP3mAc/kpOeEvy7PnwT0uIn
GC03OFGuQPLHzxTEjV0cViWRQNyntD0AliGirVplW5zhhCKZof9Xgj4YkzLV9BJYmuHHMKSEQLfC
DFaRRQmG8YuLijH1zLEvW+HrpYJDv9On7/1gWTAZdWttCKduzQ0ES1W2Nr7UjCsP8bwwcytJpQo/
hhDY1nwQ7rzc4wb/tiWI5TwAEPCzPifvNhkkehg34B7FMzWeTc7CltzWVKv1Vlj0KOe7JCQ7SfGo
rso0VC+Fm7S2ae8u8H4hBDv6GzufZ/jWf/D+dJys7ymQvHfoyMqrtIgNt+qiDSmOLJxy50tBM/QT
xmRWR1kOT3sw2yjPVLY8T2mGsmGKRIJkBqbGrS/FNzYdCBrvvrCuuvIxxrtSQXjjKmtiR5lxDrfj
S6E+qaIzhOmYQTcSTmA3rAU9Vq4TIkLhBq22XVudqrQ7mo2NuEOUrMid9Ku+9fepRz9nDjXHBrMF
rFe+4Ia8xqTvTx2JRxSZJqCRtXNjQERXMptgOWANGyDSstsPXOp/iOMV1UBjzAM9NgKJXkwtoG4e
9G2lYnN75EYWADfkXj0NMEBk7snrBL96WDsnaEwRHGHnWMl9FCoxq67Lz0OeyUBXMCbKzaxXk9DK
Vs2pY4XdPK+cUHjcC6ZK7xtnaTnPv8djZNrfbszKnNdSx/pwPyNc/VHUoA/wnPA/JHCMynM4BU5J
N5xwSWg9MoHSIrHVh0ofn6GnfjS2Buucb5fUQIJeuqNC9Z3A+lhpbr5FCfpAuinW0tStXDxq6vKm
uY21t02i9fjj87rO2MdzoqC3CYt9tAwiilgZRP5YYVbCMMzL0gXw4qLfFniz8JkQYYk+7MOhF+E0
NO/vimHaBRP9xfXdqkiH5f8mh9QQYoaNG4xULWHO1A3sUDS5UznWe224053UHi14OTVRB3sJFbOr
TiHGtpMAygd2b1A4cgkywjfFmu6Q1yaB4yKc0tAy9vvXxZSIJmm90/mf8I6IIkDayTcR8BQgJGYl
Be6nvjD7rKIT3T87M+d1PUrckk/VmbTeft9erLisThmkUKz4GdVvFBGQJCT3lGmq9NopiLwfkFDK
Ps0HNHs97yFyMZSyvSWhZYbz0PhPYLAk+/92e0iBq9+cxDU8A2Mdr9x0Hbq0s9SSzlC3XK0QlQg/
DDrx8rVL6I191A9Y17q3EXEtR3yiLzx+sxw4yiGEdgPSQVcbmMC4O6qq3x6lu2aksj9XSCoC9OQ+
gYECgxVkHKYz70flx6UuYKP6O7qtoyeKDdXawLTa6cKjaZm6pPEFaqQVzCh3YwJ6R4Qm61LW1r2C
1TI0Ub56FU2H/yZEfpGX6UlMlcHtiJcXuaUqQMzexjpCfkAD5SdnYPVk/if/B9yz7s3nMRZobi5e
EAfR4/Ey3oF2ymeKev/X1QX9Jo2zVenwfajkGfU+A3k75STYnmehCKbNp3sMehxHqkVL5EXO37b3
/+Dn+ZRxQKNvo0oKGN4rT8u2MNjql3OoLYcENkZWmfBuA937cq5KivBrKhca3VdFF6dnmX6LPsOt
mtNajUx7uObw5L0YtYpnL8sBunso+yETqORdfN/HIFQYQUfGcDTjpc4Yii15TRULv0aXRrqEXgOV
tdIIIQZqxTseeBsn1WoPDefS8AOVXbQHnhp1DO/C+WhnoeKLrDO8e9Gpq1RRiO3tVCGXCmqlk5ks
CV4DtT/FdDk2khg9qqCAL6hWHOyzx18fLK7nPDsMrynbbY0MZG5Qfz+vbl2Ifli0qA8x5qeKBpoL
Sx7P0lVOdKRTFi3eDPslR5CUg4JGYTAkEd189bUn+u7liLGZ1k44y+STVHXfv2WggMh4FstJTMwc
XCQxp+t1NWfvpM+ULZYc0m+BwF3ejv43BQKq/9zhItgVOcjDTrsvwACThgUoceZFmyv90WbZwy+g
GjifmUNXWwuWEOgFSbvKKp6SGnM7V4Fa/Lq4ikMRNoL+t/CaZCJLbh0P+HeA3URQBnIKoLzZGkHP
Rw66XrRKCPWzPrJg6J84jgr8W0Dzi4PGV0qM/RJY1e/MiAj+G3iN0FPNE6TJsLMJab4CWJPrp2uw
attnf/5wMD7KN+RJieWt2oyuqOLugCUKuEMqHYAu5BYthKsH7Kx+jzpQvjR3ObqELN/v+KxwB3o5
Gh72DoiXpaeECMxPxbuDvDzooJ3UOIqhXn+8NOjMuLbWlnT1zXmJHQnJjn/zmOCzSOE35tpJ8PXg
rw9fCHALhzu5Ude1WBnVESmp7Kx2aS0c/zMJ05bTMRF33lp2qOVu2vmI60vsRRGotjT1KLrX+NgX
vBKBZu9iOV5oeFEY000DuF6RyTEHST/VcuhNLAz+L4khXarYULikRpag5hvRK5URH7UofO0zrqJs
3S3f6FxFMgiP51/j5ObSKiZFnRR3RLI5r5OvjKQvnvTHpNSiXElrjeWaslpxrVhCriLtrQU6beB1
SkuNjohv9616pWFWCAymmUWi05LhiLw4gyCgexnKcXRSc+aWIAER2253Lwy9fOWoDvezb9uWJFY0
O/N4F7MSx0JuOYXpAYxmMpSh3EmTvakC9qZCbDbLJ+58EpOI69nLWXt6u1Th6TQacVrWLv7csxrS
y+qGjoxnrFti2F2Eofwz90pPqaY2/9BEBIkDcKA/spuSX3Y/oWJyK3T4+/rb5s4h2auAE3Ahc3Im
yX5xCfG1DerV4X8da+VklPD3fZOnWRfzzjnZHaeLLztaiMIv+4Fr54dJqQtum8uhM8Rrf50COu3R
9X0zv/ipha3jsN55HSGcv08i5O7XlxFj4wXXdX5ScEiLrQ7///4KFo85zt3rpxV8DvRKxdOuN553
e/rbscOuroe2Dltt4j0e0hHy8lmNYOKEz5bRazk5awCkiN37IiHwFIjuNJds+CIbTx1Yo8Fb6B72
q9H3Kj222GKHkjZgLwwp/dN7iorb80wbL4HMLXs6IbQdaREFybhtJwsiXRbTkWkSDpQFjZMrNenx
1TtxXS/X8VbIILlkNtuRouEE61WUHgBnhcvSPE1Vj+Oj4AjBXt4RbYuPloLVaH3MUd53Pj8jmfCs
D7vMFvnpImWN2C4dZVWHTMUC6Y2TNI5Tmr3pt0V4T8l0qTv70dhEYRR0bKz+6YcyuULI6bU8QPCb
7VB2bak5uXJPCX3A3KzElHGeqkGuAhMouMLfSEeZ1PuPDLUdiIrHTOod9XVDKYDctT6uez4aaQZK
mIHxc4KeEBdx+8na4AD0piISDBY5t54JNlRFJjMRunXm4po38II13uXMW3M5PSjmxj35YLr737+z
FVm3q/Z+TVQYD90gM6Ip053BdfskN5JKPLTDZdWDMP+63glQPKhXpYOtfnSxNg80Sk7EF/+gr/tI
6d/ibcU/JeI8oeriwu+Ugxy8sLf+bBePrxyh/NC9ugA6xVuOSS+01MXGRqgfgVD1ONh6e0GN/09N
DR6YLo/6oBPcnBqQ5ZgR3MOMQNe+JV/bQ2bqKCFXGrHChYzV6HeUVcLNF9irnXj2prJAI+FHolPN
eVoQWSVw98SA5mQsS4M56tyrTSkweHY13EYp0kjYNzdX28/umfZ5cAScHz6334xJIaAO8IB+ksDt
JGhfoCi9rKwJxLJXz2Uce3vwvkkT393Iybw/Sihu0K9QxmKJ30yLu/rwhAhwJEE57AKKW/53PxRC
2PICizGh/OAahjtJENmdv02QxVeBFatj2y4ufG6ECL8ay10MgFJK457CP1u3zdLLxhvUfWnD0ckg
bt1kOHmVxF0QP9WMXHvtCnnxsJEPUJhpq0B3u6286tx53VtdFxCjz1Ude0QsNg/RSgBtc3BxHxJs
Q7I8+pEUwQWBnKDIBIq8aAkV0ERr37iOUTrbBZyMe4BHndx5EH9QJJyeBCJo8/JITpuAG5FismVS
Dsnn0QkRTwULWuvCro9mbCQ9tIvXxSwdJ3N+IuDwajhUoE9BtNbsQrRV38la7+2lUajQ2MGEK0OV
F4Twzk/hanSLAZ/iPZOqAEKIxiGp5zP6cNCb0BzaR80doi6gCdiUItY0n/SK7dxmDCGy7Eh46X2k
emq/O7DIkCLK2H9dzHJmLLw9QvnTCPeasjAAuNRVKBg91tzBZbRRw4XuU/MaLDC6PSIM4Hn7xyaS
WHzaeQ7p/fZ/D9gOdWyVYKiYAPa/P5mUR/aJ6XTKfCXEhwPMrqogFi4+S1LeAqBE0IN6GKmmrIHX
DxJummbiivz3Ci5zF6gfyFHXH+iWy1PVMEtsT8r8Iv1/wldtBU48Oz883MXsLiAlv0/ic2WQj8Em
nlUqd7sS+GOl/Kk8s6eLUdx4yPYRts2xU+45PG+jOfKkxIwF3X4T6BpZmwUEmK370bY5y2uDnICb
QAIz65vQOzuCEZYftVjlJcLF3wFC1u0MCkx6YkTVRI4XflZU7k/P6F0fHg0eqBfiqrViGwMZt0IV
lsVIBa6StpYRrOGuQvegebW+qOwvcBIB8bQKPrDnWnZmLcTU1XVM83FGy/qp5UpjBtwJ4U/aVz+S
b2f+nfg34goI+fkNF5taC0wpaKsHASnvM6sLfI1yPNI++8Y3AlCA3fCOkxXGDd5huJleQqGJg0zr
K5TuPDnPsSUOZeGqJ9x7rGAGFLDXjmwlMMEIupA1oaLxMzhcOXptR8FtyXbCsxK911a4iXiXpzJW
CkcGZOu/W6gcIHfzCVRjnsg9Asb3EExcBNA2y0AugZ8xKjXKwKS2PvfZgGulc7aR9SJLfgBoB8zu
JW3PtiyNAnlnMz+vYd5acgDLACwM3Nevabe36zqyCPBS7Se3nZRS+NnGGvtE8iDlvpsersE38Xpp
lK7UJi6DTVIAdgbsVXqimcGbfRHvvi4hGyY9sZeEWq4Zksv4tR+CVHM3N0psvxPdD3qW5TOeQzaO
FQ0YEBclGAve+o7abTDXz1eQyBx3Z3LhRjRJQr2iACeKngxYMYTebpPxLyHYGFg3nPu5gZBuU9Bn
j++YnIOm5DcloIHw3xUpgjdecV7pQlx00ckY4g1CuN26XjMH6pZa+3gPOOv/5ib1DMIPVn0dG1JQ
Cpnn+/E0ycny8SslEem8cJdYRJnRVccJ7TSpWV+UcSg3YML3/ymnCG1zWQGGZGzLBb1USClbqjqi
s80dOGDZSCt9VCE4N/CeM9nk13rdRJGnWCQTIL7WPMFSHsJ6zdqO8mPamuf8wn6h8cIZom9bS2Z5
gBVVlDaCX3DbjaNePawEykBmrwGuJ8ucBgcgvkdgWmtwHO/WDp5/qJX0BbIiv3n3nWMAsC7zxgqC
ti81F8IbX2Ykkw+t6fFqbMMFXQp7t9yfbAmpkJF0jKpE0R2XhvWIPAi6kMpwD9YbCP/P9pjlk6IE
XOGP0TZFPNQXpoTjOKvnLpqDeqMTrSk+jR6Rt1oHcYJPpMFB0A+bLl7X18sNN6GnG0KY24cOWc0b
TTLp75y0NFbj+0Xdr8mWaOJvr59EA37QvgVlJh3L9xfIr+5EI4oSU7ks+/SOPMWVRfjYDQbDH+sJ
ZaExe3jQNWf3etjAe11YNrIqdhoiNACIY4NUS75FD5TVp+AQDXOzEl9GCkvdldsay0U3H541X9h4
aaypXSpJ9fneI/Y5pOqVUfS2Oms1sLYbRzhOt1kk0pLI71sdW5XNHP2Adm/9PXJESOgdQchFdK0h
Fxf7DM6oF4yaCyocJ+ekB9K9DkVUbK4lOhGWC/8ywFjNe3DHsNIGkk9q+e7dvsP93r+Y+z5oRk7B
/9XFYDZ8K1A5m1K0s8jBQkbdFpHneX7JIoZx3+915DuJmySzS+AKNVGQTG3oQDkOaT0k4IaDlRK/
XIeNI6YLBYCOaoHs7BQ+5rHODbsEYnqWaAjl08jVPCdtxsryXQ0qeH0oX+BT6n1s3xnWGCJZncs6
7RNDlhaLXIOfScpiAx5zhHrRxN4ODQyiD7DcNh2GctEmdY6fdPZ3qsU0BOby+cjFaiOrM9POjDiJ
qkWJ6Ul3Vq8fhfKBhDPYBCIOSvgug/jGWMqjKgJJFW/4OuxtfeusVmLp59va4BFK9JoDvm9m+ulB
S3lEmZo6UxxgmKetf1Pkm3OQjv/RHQCHYdLoOJu4DdPVvTdGayVRcJS0Ivy8LreAMESFYj82ECT2
FvUpjkCqZvxM0HlZ+jPpQpm5Ab/ECN33zhX33Vm1KSWDaWC2IhzwlILKzMzkmaLyQOn5sECoGNwP
IHFL6XsN70ZhUYhlZ9YXHHMZWsjqEE4OLBxph5NNXLm7+ytuBtET/KvZsBy6rRiI16277pAiuXIH
PYS/L/YPYfZWQyFD7J/NIwiqC0sP8U+42ONS0QzvVeM4BvloFe31WxkCSifwEoNrV1Fgp4sQuazj
TPUSYA0SUCpf+GHfPCVmzbEwg0RmyTQUiG89848Hp/v7LVSEaF5LGGAsJzZ8hRryJVT64qt8aJmt
WUpvi2d7wqNWI33YaDGvrByWLyDWYv9vJ+dPFZNRuzpDCGpO5zdOxA/szwVCFede7xLD0qc+vZdI
phbW5vfmfTyM48UZyZnxSY1WWcSxwKqsqI8hUdh+cuT4e8n3y/vt/SNgwWLOMW61xL/CAGMuuJAv
ak8UryvUkRmNzm/YGHg5X/p8XgcwSKneBbF86dQHZWb08ntNw2DCRfubgSEEbRAojQuJr79b0Mbh
9bMl9wkrVoZsh14BNTK5ZhCOXZgF/dAj/ol879wxgqgb9EcxhbpcqKEIaPNPyTP1oF8NvvbleRuF
/hpvnmFWULrSz3pOvQ5u3O59jlHiLw957hXDMNkvloWOLFoHPvFlrzHrkd1TvDDbzbtc/iJIc4iD
wPhzTLSIG/GRB6Qv7Yve+8vkQGp+/zkzs5BJik27MWUean/q1XiYh7DEUoT+VjEj9qEc8ZGU3xwJ
mWXr2uo07h0cqyVX3XdFuE0sqpNTmW6IdaZ5aZZ94rRUIAqb4JjoZHqrsp0pG4Yzj6rITo2HLy3h
h24RLLtoTAYwywQxrb0kjokWxGcuZAUu6JEBdvMyMxE8Rwc8VdYPQRkchSE7tJ2BJfuLQ5S81p8C
plyzOzfSUdUat73dLUINZDjgfJEa7GXs1awznzTYuCpygrPxkwUKxFNs5dfOSdM/jaaTg/m4ceOm
QphSTzRfJyThufqPkId+g1hs6sK5kTfY3Bmelj+rGL1kOQLxPJfjXYGi5+8a6fZYOoe3I8EQibRZ
4Pg4tkepjgdLSIt2yi5JPCXe+huhFo582/v9lqWZWJnrjhPZ8UZb4DoW1hJb8AC+FMwSN3C9srOa
e3kPff1miYJP5nFSavrvYCHJcNNrGm4lJgyVQLWo+UlfHofyDK0W/OAXnSnPuPfA7hx1Hth+L3g4
aeXm1QfWb+IPk5yBVygNCHdGmYwFRYOvp1iROlv2BUNBOaHC0Stbd7y0QQbCduw8zNZ7CLoilXhc
sUqzE6VvXI7OUVKR6WS3ijaxNyi4szkcuG1qfn5kalzZ3HuQc6mqgDsJoaPDPvKqNxKRtf5fxqbk
jChcro9MO51cSW2W786EXp6C1EIFgFQ8VOM5/isgc10jgIOFI2QqA03HzSfZB7Valj1qiyWfMCKt
LubhH8ZULQLpDoCglm1kuAuCXXxY8ArEzvf+iJ7YXdsuiSV3fP3gYd+DQlGbEnRFrFpnb+no+kAv
PvMiZBdlTzYH0JbDs97sRaSzX5qVb8zS5mcxpE7CJ1rlxa1U3SFTE2CvBEne5VpZK1XJ1f0J3p9T
ilKaDHrOZxDtmYIyC1u71kWoenKtYyllPg92uj7bzP3KEAbluKptvYT+VarUgPYPZsugvWHKUfl2
wTJvb5zeMR23ZSkecJCZIpSrSH/lG9nDXqTCSRhmFqIgPHbBtLIi/XC4sKkNorSfHIRVb/rDoSvs
NXbdJHdNAxr1KNryIjosj9kvQq4nk3cN2ywOxj4B4qLNLytwtPjYmI8opcF4fSAX44zpSbZOoM4D
qwmWcMLAB8GmMbhboNaUQ0nkr66+iZquIycZrEs17EgSGNnPeFpeZm7iShzuAyZH4Ei3+gq50/Ax
EPj9vva+znoQS6nD2UMgsvdcpMroz5vYJtEy2cxtZ7zL3LeP5Ozgk4Pmqx6PBfX7tNGk8zehbIrs
gjSWb6rhd6EtQvbfAVXD14dRgTsN9FtfaL6WJSrWKu62hKUdhnnS8DJYzaV4/QlVYaRKjX20KgLM
aElvwlpzouLdmV1ppcQmiSUkSTdy1joY9TC2c7JE3ixbPWH3Qb/Wd2tpYec0WKoc7kEsdCu6Z+gl
4WdJUc+bDmeZPiEEFocH2FraWAMTUGJMX2WlL3Hojj2OAF56HH2rOJs21IGBfKXGWxHLg7DI5bui
3Qvz5NkkClVGbit/SN+pscBM87vo+D4hqG7jK6APT6jsTbwTcH0CDMewiWh0iFpMGLjASDchaWVZ
sNo65MCYB3FMN5a9V44aaIcbsdB5YrulgfK1ALEBFKoduApQt3u+zShc9ozLcmRMLzZreQxM47Nq
BLGfeCtPyhoQnRWBNHSZEeXPY/IiC5A1CG66ueYuZo0IvVRYWgkbHLWITKfAKboagJxWYlTN+xIm
VSqud4YD33Bvdl2hlzn1Nt9J7IbY1fzI3SPvKnA0OOt41YOPUUahlHFqw+nsKZZX4vAO4nx3Muju
4TxosCPmXA2MlkAxnKExOXiv8cWoJEbCgX/zNO+40XNSsej5dRAxPZyMceeslVHnrWJ0h257CGAg
GwRMhG9vq9WMNLert5CuTpdOwka/zHWECJJrgJjKl5gMSIJVeq4aj7Srom2gItLSx5W2fmw1RAaG
iWMYUfB+WgkegdluO65r4hkkXrZf03AMwuIIXsgkyCsIoYsHxjAk2H0NcVTVPNBikWM5wvbRUPu7
NBcIDPEsCv0q3Ei0Ea7zkTtwk6wskoQipOh98FJWJCoxK4cyPTWc+jPEq0KR+1eF5BfVMX9yx8eG
p9noIXmKxKOqQhErEv0SB6cPM2Xj+imdDbI/C1U1MfkBmqAwDLAYeO6idMwK+BMkGXVtf5z9BukW
dycuvV7oc2nF/9PbASUY0z0B93z2ERzbRjUYOSECFX8i1+dO2yAYuzSWz9KBrO06nBScgqaOpAr9
ErM56jgFdEu3CQcowk7ih1YxB8dYfLXsvAo5zVOXf2QC38lapNg9dp47HngChNaXItTq2A4Cx9pw
iLWmE5HudDNtoVuGHZ4ar+uuk5ERWS8AsdeLGkHj1IHoCMuvA7rnMic2CFQype+RT9QaSR/Gdejc
Y+bwma+XZWYr/ncHZx6KcLZWt3m71GnebacsoYvkDUTRwXvC3QhipVSCXuAQ6PNO6N2JeElESiQ+
m13mC9EB/wpbS+RKjK1K6TghF4DSmVCA018K3Oi81Vd7XDlUw6IeZufbBqen/t7sEQV5D8MBOadA
VN/LBB6g2LR4pd80lUgbiD5ax7Ct4+KJEZaVSUEFt82q6p708UsvPpxLUorsOTFaTaoIFC2II8MA
r3o8YhIrm4Rr+bkQq42W5QSVGglZ2J6EMlLqayZFlWPJoyHLaLPStE82A+G7zJxdBlx86ttJf6Vx
9XbrV9T4LJiKcwTp8K41d1gxA+TqfNffKOlgLl5fDGQKb/HEvPPAhWtvu+ei7BnazNwm26t2ITf/
DIKZQapFR/IfV0ZCDEemoz+eHi9/i7DK2/KTufKzq7e4yz584rhz3RXiw0NkqE+9V9BRObs7s3KR
C+F+DcixMFqqqHxVgrVmkb3d4CUKewcGYEwe3da+MmFhyFIfwARoWgz88JjnlREllhL6EbQFTnrH
Ccs0E3YYnHPKJJWTtw0OIIXRuWn3ZTHdkZB3wvbVS+tTs1QsPwUrUyjDxoMucEqwp1Kcl2//d7gI
KtV3gh3FixVLli8E/qLVRge3+H0ojyA/er2jlQyFxj9iw4WijHnu8sqcmlK1SCMFKi7LtCYskW3r
tivC79fIlTj00c/SBFkr1FcBApTib/eocwMFPztMJMUw6vuGzGci0+KoJwjU+/A2rYiTNF5e0qbG
KVsXW69uKL7IVKTMUmSpILu2XBEGv/X8qkh2YQRZ4k9E6mqsRKumAhT/nDcTczOnzq1ZQG67S2My
kuaUb8ZJkxfus5ruAclCn8sQMgLBD5Dd7FXzqyK5QnPjc1y/7zgJf0BfG856PmtF+pUyz5fp+4Vp
SL8f8sJTcFJleBELgu5L2/+Z/96OV3XFQLTRGDOV60i01JYnV5UBH/RIY1DMhS5hHeNxaW1LrIjL
US3BVgpbIxR9iIww2rozN8MSqfbBdDUXpUiRhi4habN3iR3U39/LCFXV+bKFb/Fv/Dbi7f+X+Dxt
l8bxeHOMIEGjBQY1C66C4SDMWUeXHtkK1zL21ifAV7/BKyzuoyfOBKgFFEkqGVSiqQAQBo9kDlJP
pYK1hR/rFSMtSCHg4+PlpKXZP6/i0Yno0kt27kgOKmyFRRhZWKzWL+mB4kT3CBJbBxtjYIwLyRWh
WE8K9EQohC7g0VxrGZONYFhMsspm8Jm11IC4JaaLGHstOvLvPcDph2l6IRwX4KCALUMZb0ORXaxw
7ixomuaI4b+SpgltvfeL1lF6IPb8M3hqovMukxLc2iVSr67mAF+F6ztV63qC6hepFl2LP6uoToH8
qAxt2ROnw0WhUaa0olFCd0D3hpFRcyqjsnkWsM2YfEuS02IuclppU8mb/o/92qsg/KvXt1BI3fYU
dqTqERx8poR6LD3AawhvG6AMHMT5T54/tKbHYIgp54TIHH9TSM9wT+dNMZ1CdS9qdl3cZsX4Vefs
a9JdzYPJdJqlfz8b3JoyJS7T4PuYrv8upeyclB1jvHx3KhxzFRodGkV0D+lXhw/JW+1SUzQuHT0W
rxcwBXo9ZI6txhilGN2HStaH2WQWApQSNdUAOMCYi8LJA+kHJAiJNT0tlJ3LiYEvx0eE9ws674FV
aAVdBBqX5oakIFQruu0N22SKfk5Pu8PlKbGYEp604Ax4thgerV7i8bmDL4ZaqWrOjyhARHkVadbP
9DwXYbC+Fm2RWN6Fkk8TN7ZlbY88G+RUluVHfiOZP3qxG8/Od0KZNe0ZDXtR4cSTD0H7/WETi3ZC
/Xa6aQehedrFG98WT/TyyQsxSTfDOtCd683f881gcoCypfYll+rlJCz1lBlmG25R0P3YCG0x0nvi
2TjJfVpk86mHKRofEHY4IVQ7XLtaw9TTeLqwMnBDzo0wG9Dx5TmRgeYzQiUBTTaWwC5IE+LnNxeu
POVrYZB4tyc83doCj6d5smp5OteEL0+ZO3uQzG8CWqX43fSrMqVVc/PgRSmwAVoNDB0j3y26ypW7
IBaIG1zislOhjpWwV62rBPnJeK+KDGtCBOYnB0+5jXXgKWqQnVmmTfvjpZyXppIicTjGLVPsLaHN
Azhlnga/AMoev2nrbQFLxyeg9uQmZh3Q+DmB4gsalxsd7h8ng5EVkXncscL8awBzH2UdC+SSPHGt
29JP4U1tpfqmQOLhEysd2xBZZYIgoORRvB39PnIQ1q4aABmVAfL2hgJdJFiwkcOw1D92ZqADnope
Nwi4VS2oeLaiHeHCYgpRE9PmqO4gLTRaBMtBuYFn2lawOUJ7MGDbzVeSx8yipsfGB6jzSzlWUVni
QTMHKWv6h5Do41tuFogDsSOuVYhGLLcMkRvVz6yJgs+CwxXoykZlJ0/vnkR8cJSyK3y/Q1kJ1pbK
FaSS8hBuRsjmrZqaFph3EYfIR04ksjFv4Ir6gAlRIXvXXgDTvs1WZtmQ6dMqoNlmAQrzAZCAyoU0
fAe8iSVRm8AnbdnKNIngFmVJwySLx8WY7ejqLA05pwAygQmF8NQ6LGUxGT9qc+rtZ6ASGKdUzDTr
ohrX9tg5qo48kkxf+CMGaMOl/jpt5TVxMgwEXRHbfm2LlVD6vpdJOMN1m681p6AOr+rzwY16Lecz
KBncEx1WOFRweBJv3KySDYCLD5B63BpbEqnKkNbTUfi/zKyhzgo7yxG+5J2Q2L5VbujWPtanDMXp
CUR/dzASm9M2tQvshWHeAxXZ6JBB7l+R0ZXIkm4RPkiSS4M00d8C5UvFtCXdt3l78dRBRFNVrntw
CD1RVeqBwNDrvwJ/3fSRp+wWeclJ6Dt0p+OE8ZzMsGLskR3vgzGQBA+XpYzCD6G9ZoyTeaW+xNDG
ryXUW+iQgpErpzAdJ/urs6dnCm6n8SF9G0wD8LlKwY6/LzfojgKBEnwATACYsU51kHSgaAYgcphz
/Y1WeNMuJQFyKReRTwgiSm/ijZrE0qHOHXrrDVKRs7jbIMi77HSUil5evzftd1T5j6SuGQ6/J1P1
n9qlhY3LaEaQKDbVgsatAiB4XCsn7sdUgSub/kT52mRVPR6WowI9wPt8s7Pm0eyg9Zltau/W/QVx
ti/t7V+USicD7LJL+7ykOYZC0qmNRlqkS1s+F7BqSCUNDCWbW/irPPUUZPJPxihtg0CBcUE4GBD8
UOV+gp/NhPkxmFBbkVRiEmcrB0qbJ8panJ2jYYb2yf5KDq1LV+26RfWxjMG5N+k5l/aMZoJfSbjN
VsnbSTDJw3ORZ8VhbjfJbCqikdoEBV9LI6w5ITGVDr2k+Lp/saWHOL9x8PT2QqqGrcN5Vr+MXUuD
Jj52ZJG/aW84OT7K/wXtBzv6LIgGO6mZZWlYzaWAwDm+EVVL/0UF2zzhruhlpdgz/2nRRdG2hHwo
PkT26wd1LdcmZgQiC1m0GX8FaqCc1zozOe6N3eUjxhGaMnqrFCNN58qlQf7RslipL4dQ8RUPUdw+
ZevRJfpHckIxhS3mXzm3hGATmBlKCNeRRyba8ynnMCXzmcf5jYntuAm+DrTCK1yoJBln+Qdkw/ev
PSTV8+yLLXUQ5F0grvF4xgKoL26wC3dpAouYYOWww3TmcNfoQCFjCcYsaP+r6Yi/aBl1m2uj5u59
FOUduDxEfns1O9ZmybZJQ92xSWtCY2SmFui5F+oWiBoyMh5MVUXRt4BuWV8IHOODQbcmt1FsWGyB
cd3bYmpQCxpZrvUdJxkBjo2AvrAPCGQr3qewbwtSHXpgXz3rAECAAGf7s38Lgqo5gGdVmNs1jacQ
9qd1fftDrTo4l5shZKr7OJz7R3KSKN1/I4qiNtLk4+5cPPJK8kByQ3++KElZw6GmEP9UgdUr/hpi
nkDNi6ViVe5mkJxlnh5gVgP1nnHT7NX5lz0y4HMaxkCwlzvGo2NPmP8UwW8dBADRcY0c1g1Qc1tU
PMSbJhepmJftcqHKPzKZx14KaYwi7O/0VvuMwTay57wB3rrU6dTqqK6UckVZVaqw79Ds9P/jiZgd
IB/A9KyC5ZR0S4Dr5mzAr3UpCGiSqBioC8pVvsR6OvAspLCT3V5P1GZ5kZjUUk6xxIykc1nPM6O4
I4tpxM7Hq8ir63RkomAjmVbKOwcjQwQOG+b6oHOpV1mWboRbkFhc03TSE38KZc9RKJq//ZBqGQa7
xsA4Aq7oEWdi1CEDxcjR6/0TVFnNIgByj6HE5TTgFPwlePZS/FvUMZ0C0jVcYXF4KhjVBZWkZeww
LB7ay3fmqSyG2sr6WEAYAbS6M2heNysXAHucVVuIaepEmrn1lSXuLtZ9bDeOthZE+Sz/Brq74DF2
uTdX3CI2O5B3p+CEIiOFQwrSkxQbV2zQ91N/K2yQimX+LQzgM3dpe/MAdIcUNZTB6x5ijxgyg2fE
eDmDJHpTG06bjGiKVNiyL1NRgeRW4AZuC1zT7LemESVfCgSaesjlT2X87MfNmksrlRCovHHwL4KL
5kpwaqCaz+TujZg/pzeqcrc1aN3ArmHtBfkPyuo3YvWL31Ubi7SiP3T9h7y4SZcqLKIEhe9EfjQn
ju4GN/y182CXFE5z9rGBD3C+a4NYl0yNtY72+W/McaKxnaKDD5hx3Kd7PP/ZpauH3GNBqFhlZsFf
g7sg1AX7r+s8kZV9HuhyUVd4Cdh/zU9Ms0w/S9bWK9lsFRqCOgTSF9IUo1mzXI2RlLCcDejTV43w
ftzSaMhKc0Duf8hqm0+bgRA1D41rYLjBvnVLMAkZ9Aw7ITyOVCNhnp3hF/V8R7yM7ITJxs3+fkJk
W6cfbaX0AGNiXrji6upeiQrk3qFr+dk+6IIyXDqkfQKeOPwgcKU3GzmQwIqskepOjIabOxsOzw0g
DZ1FSq9P8ZIkNOpxzD8WIa6+V59/Ylnkn9AsZ3vX1vvjO8E5eY/zosghf1izdXoFPL8vitx963eF
trKyWMSNBFT9h7lxJK7wZhsGMfWQHEdHeJclPuGC24+tarnRfRqBflAOQ2c4aVHhtT+DoG/nC9CA
wQZIv4qzNmJ0h/YGxTDnBT6RCQhFJh9yZbUM8iLbMB+NA1QrMgTmZX1ZXTUkVRrPDNS+UImKH878
CybPbCwHjty5t2sVg3x69Mq8XJgn+K/UQebwUSjeQIiRG3aS4VUayRm82EZMlfD92ZGQajZa2/kE
9yjz87UuB7hXst0AWzoWTfdKLuJJMjvHP2BouhKOhHxR/qTHSXvgGuSzGvBFDmY8TkivYGETKBGB
nMzY5yjtUfG3IZsjTTSmbZX3ThG8AX/K6f0fXeXYt5qJZe/tU6PcrsdLo8CkwUo2YKQN0VAUaUdk
VUjDAqx2+25T80MSpGCL4FVO7SrdPJ1xcwhgB/2XYwA5MX2woJeosSmiWQnrMIg7fC18ZoKXLTAC
/zH5g6JckIo0y8LZHBkTsU5iLH8j0/RbXv4v1TJSVDtYiXdNtJerCVCEVTNiIoEGIwaEc5SPtVrc
ZJU/tH580l9ASUv2QP3GdFm8uU5J5LYgbanvAZ3YHtVk8IFYWd9crcEKSGFIMdt1uKpnXWvBC2W6
A/aoCXc5vOBiYYcYpXQUo2bLPAHJtC0GxLfDlYq1ojkfAxwmqTbWLdU3NEpSMSBBQyaZrtCvrQyH
CoG3ftB//WEAdS072XRiNZUHaVtzwD79ksoCbuFH+bQTneUTsV5KL/Yg7lSZ6ZqacED4Of50JysS
/BBCT+m1dq0mHmnM8w08yRI+IzXbDC342WcM63nLyyKqmGROH6tOsMYPG1x5i8yr8Vgm8LHnt8d7
OrMOao9LylPqbjohWFiTy1QSuqMV0sfzx4dy/7oDPuxfVFWKVlIG7PmFHwXhh4cI38GNHYsdZphA
8iYl9BAaARBc2n+/2e5xegZOrAxcbZP7f6Oeb7iBtyLsRcktIYV1dgYvC989oxpLwoEXI3gjKwYK
lZNVGhwQZQ5wN5yh6vfKBs8bAZQt2LiBYkDtnzRFf1FYsNpL5N48Zw5QzXaE4X3fUdqxeOuot+a8
dIJIEFNvxjVYDc6ka2f0PsPMDQUqS6mnm6sXQFFDVMx601uKAtP6DXsHe0tjleytAvHYBoz/wYge
n5Riz85steSI9BTYkiQewL2BiIZo0HER9aEWYM/Eq+rartKrOgwkVmhwjMJkURNs0tErcbDrIIr6
XAnm3DJNibrIy3eOQtJ6AJ4M9DcNOp0xphpe/SzFtbvDYQI963kG9AkusLfHf7hQm9XUr74FERsh
rcJqGheMtqwbvLmIPX0FnIf2rHxzwaSjJKtGaIcnTJwoZZea5k26Jp5QOJXMC+mM8T2b7oNVidYh
o+gJW/32o6q2goNqCwkYfrjW6a8JGL4Ob+1Fy1LXkUbh2t6J67rLVqvGSJ2H1PLHhK48CVDtCdYR
e+03+TMw78wDQCyXWLxxLMn74nVMOemPixWU81gxUUi5uQ7wjZUbSIrcEFh831AEaaTeaECYZFlK
SNFy0X5MIDwLpAQ9MK1JAIKqzc7GzwbbQXh45IGQbmuvvd11l2kO22hY4guBvqqljtPQ73+bax+b
IjUL94KaTnElt0tmotnZObjef3Ah/Cp75d71LZN7CbrXlsv64bzfL0x39z8mpvrsP/sWyx+BpS8X
3PsEnthzCWi1XfqLl4cOM5dCEDlw40d3OLtuAsDRYUFHO160ZFtZYuCORy0cwRoNdurLyMqUty5G
pPHXiQF0NJZcJTG2pzTw6UIDNfyOl1KWo7I+gNHq4C6pMu/dIHtRxhTL41v4cj9dXHqSbrIyHytE
6ZqVbXWc8niBIWotAsJvIpaC7UEfrpyuj8044WKiQz8TXsT3TpZTkQx6f60dFrJgYFdlU4Tt26AU
X+Dqv8mATcPnuNxvtKq0C2SS2JZ2UJbKCIlZfx3FYa7pCndfxjY5cvVA3mu1sD7y17j5ARBsmree
T6UB30yj950jmi+1d6xthI6xi5ol11zyHG/lAzEr6rrPBUCiuTirwZJdFlyh9bA2AuYb2f7U662o
6bpkueBaj+II7csCezak+rtmn6qvStUvYrxT720+r5wBD+VbPmC4jj6hYW/lKySvp7OwMbyFwpRa
eiRuytfJ1PTLMyV2XkutmwUVCdhEW90m5kM+YgZD2WFIInuuKwtb5jFdNtgD9+6NJgP7RKNM2daH
8ZSngTI1shBfRh4nM/m6xHcJnX5DRCFzyIUfxUsfwUJL6+nXVVUFiJWhkq7+wnCPStK+osSyxhAH
WeNGNZqRhKZQm+P7KoXTWfikpn2UcLJHXiW4AB/1YDxfLA9tk8EreIO8YUE7DBiSsMdA4puQnlyt
sIOFUhDcA4I8OeTxTT//uoKGbqC9fqz53uSC/+HxCBb6c/LlYztDvlew7cLBgZX7V518l5fxjWcj
bgqZOf5K1zgnq6G7Wn8MkZKyQkC+yIoJyBJoyyGU61POBCDY9jgF/cX7/dSvtZHZBaTaEDfZm2bR
pQgoiwONJ9AdUHAuAZ1p70qwYHBrkGYBlSivfGXgrD6UNyUCasMJIVe20T+CP+GPb5qkae96b2py
C9wXN92++uDO/EgTKOeyAmoDO963ZecHnwOo2Nbxh658Zyw+4rdk8Jl40kd6Iv1B3OezjWpbpQHF
8KBPBVSKkOMIvUXV9j4RA/YVTOvZq2Wfeet4D0tYs7dhTDRNSthKShN5qBNg38U6dPhUIq9CZ/ea
EnXmEsCnUt1ZGGvH1SaTPMY6H28RJsrBly4jaDKQ02gIpBcpLSByf/SnerDsvfkq1FhyMZ4f/r/X
G9uevyG0cjXStAMEZTG5H1SMxWU0UN8+/qVKUmzuGX6G96rfBrxGkdGB/K0m6tIchihJ0A+ZJhF0
WUzaQCZdc8nORHcB6rymlKHsE6PcBnGF7qYhZfVhSbcnzUNoIpP4fC5fUEUSfDKgMoBiTb3n2EZc
hfs6CgPnNuMGNgOb5apfzuxBI8WW6/joevN5q3BGjn7kC6yRFf0lZOI+cRV4rBCE2+vgUiDVIR6u
rWrWwPwXEQUc/w8cwly11xr1LCGigNMOAu/oAyRShcNDzDcy8o3JFBmHH60xDvDBESsEbo2dhvIe
yzqnY5Yy7purxhA2KtY3CtC9Fp/fYKn04ow1/4RwwpoW+LwLNdQy/4edtGViepZLGdLuZlhityua
cq5Mfahnvq8DPTtLZ6zoJ35SC4u52AKdi/T/69hnwuapu09lUiKXORtFtI6pgTETTmGKpP1h35SK
Nk8lb7z7dERylZdMseQ25QJdnJSlsw6c+y4LAQa0PB76aRxrXQG3JA+QY/7Q13LXy2ljp91kX2SJ
BAHkblgDfxrAItKJovcCzLH4NxWaVfSh0qiDP1BaApAjgUf4UUTP0542XLtVt24zQIJHn63V9NI/
6/tyQcf//ePcCBDuIsCcBlA4OkIHfF1Jf9wyNzJ52zxrULjTUEUP+YonY2u6VGw/m9o1X1ZioWzf
V358vZE8NvMwe6OjXr6d8V1j/tY1JMYcRHsfxgfeRpZKAVN/mpy2QmnTbVuDwxj1C5d3sz0Pjhtd
LWFjJuY+XV5UEaY+pijV6CQVQ5qvk3RheL9xKUPX4zIX+ZeNuMu/4mN6B3+IIS5F6FR7LqLrfRi6
k19k+cR6iygGc6lO2NOQEhs40m9URatoKnxA4sI7ivwiTebUBAsLix8OncoJpDULnzAdb50W9UaD
DEDuCwolZxUNLQiurz7/xRzdGPlWY2FCztpqf8k41oE+pIbv1hk8/3CtMdtauoupVYnxNjpKMQyv
yhNNmEu9gtiSgHxWyenxvZjbt6GYy38e0tsqT1ZAiEYB0k1qEqVdxZ7jV2+TeZbrfOBrTHqdBRMe
yOeVds/W1/0bfnCqz1sA+UcvQ0D7MLcgIHDx02qi4qpfW3jtlpZ7t4rD0mQd/+sMFH2RiO9XRyyD
yUqAXsbO6zxSDHqmHdKaGYibt54Ozp9HjzzLhL6d/5FdBQb4i3/XUvOTfs9pOqq8fbt1s9OQ8CO+
vuSVj/+JwEUEr2+tb4hRp19jYmScRcTyneAJtPDe9gOI4TjUM/NTlXuRLdmA6viXg3O9zVX2qR99
6p1r8/3pNFvjRPaOo2aZp1lHlaBpfv1TI/OeU+yjPk3HufkBAJKYe6wrLw9zMGm/F32TbrSw7C9Y
BjEnefaY9D++rAJJrgjaJ0hK5VM7XRcXS9L9eGyrGJs3C3Ea7hbijkUb2HFvzUgUfN5sYLpX4hq3
ZCWvB5hw0getZyNrRU9edx1mQKc0pBuSoyUUl9qBgYXlJtowhN1I2vNdNE9B8AnEYjfiNgmI0IbD
qd7Kdl7AmjtUTffL/WEvZkBcvTaPEG5l1HHkU7gRdSIXpWE/KW6C4ng17wP3KIUiRBnCuzC2Urcz
h5ouT7GCEDe8YD1uQb14oDCHXBdIBz24l7Njl5tzk5nliJ9BWbv8audg3IQfODtm8qlyhILwhINK
VxuJHCdIP/FQE1ubdp+ej5NUJFUehg/mVWhjc15jyok88SfpXruN2OPR//sVU2NET9KDj8dVTwNk
I/E/AlZShe4UzM3t1Rvv+3CWzo6dewNXDIjuKE6vAxZatvxalpDhf6nauxzLlrQOxDBnFJC+3uyB
ArogOYesxajKsoJzqpsEi4LQk7uDjyTnJ8pUD/DWcrS7j0ABkEmiUYeDs6nPWWUTSW1paQeA8wRf
YlnE3KXO3NfjdS9qQIrfQ8Y6l2kjqypjkIAEMDNFHROmRcmOmLIOMjDADMhIl0QhPoHHgpsoRwGF
A12CEVB3ytbmAQ4IarRCYdesJQ8Aem6ZW1HiJyNwg1jtocPrnHt6N8qWvnER1yZgs7UN76zwjtMO
BgUnBJ6E8cjsB880K83Cm6hN1QmnKL2gItTP5B9GUPsfgSGbQ6RVY//W7aFHs5csZ8TSug3cZSnc
jsxZ03AtCWoX/1Db2j30wa9bCkg5DyPAA3/qyqyjaHps+08gNw2iZ67uJdGXp5WM8cSevjYhmq+J
UCTew4cOGunNwwh1bDOngk7WqsSXabI5vap5nDaaohfS8gnGbeFANVzYMo8cZrmT/CnBOIGHce2u
jE19e36eW7J87Bi5b5Xa5EYZ6FizQx6VRORz3XoSC1+rL88shmhk5bRmRO/P5FGjZx8HmiDxBPmI
mmeQ5fKCSm3ZULeHCEiOMcRaZdYMbHWSXY3qLQb8Ej1AgOo0z6iWxwVmiTlf4K8urdH0d12VT17q
WTGtJbOcuK7uAnadt7tg477pxgXQfTvOq1qTM/usGKkDNF4/ntjbNNOV4jI12UVFakK/ZK+9Yr8H
4aZEb4+UGghaVFtzGZvtLIrrCQWE+a7GV3rwIBp0W+q591k1y8zxuFGPhIPSOuURKVDY06A1bxFk
LidQjozO1+EGXEMj20SH7Ys4f/qxeVF2mWxrEl1juC9pxU5SQ5W747GaUl5FWruqM6QB4GjX6SxP
dOX4ckW5UPeP1gXTOTtGKwM9GRLivPpY+SkvsBOGnYcUSyEst1m5MVoiQtfiMJmhtTr/yXKM/ApW
jHFFg2SnlD3mlZR7rTqOnZCyGlYlwAL+FwMn8vUjsT/8vaGoB4d4i7FRseVFSJL9872DwHh2MSlk
gnPaQjkEyZo6p9h8du2BQptaLLnoHnWunG0JcKe/RLmo9RR6e+V5gl08whoP+yPWKXXYCYmsc3s/
ixMIuuGnYm4S5VZp9gnk+9s+EA483CUM7R21sJOMaZP/ALRXsjLe/wbvdQYKEuCIjI5q7gywYbPU
ym/5xnVanb9b23/e+kDIZAPt+TYo8W7KVBR36DrjtNyPYgSCfvjbqXCFKYVzfNnC+C5iZYmMIro/
4MZi1kSAXapRH9jahLJPJUexqj2AM2UYwoaFhI08ucZTL8h2DzpPZ5+3rTUebbg8bcMZI3qYCXs1
mWMVRvXE1MA4kqgr4//bFJVBA4rooEH+SXdwS3YZDqiV5eRJaQP6kU+bD44BaVFFLnmNFYBB91JF
TMp88xTHesIYCq1VFOv7nQPVj2PErdWHu6/6F/pVf7k7q2z0rMTDtKWTnOyJ4zRUBmbswb4ObNeT
1/ExHz61mfs2KsLOtMbS5GwfVcslNhO2OVJ2FMiXQLeOgV3p60PaYlxandsefwPO+LGSYn6wvIw+
D74HJbHrP8NGhDTGqAjZl2aU3pEexEkz8erL+eX3SLsyc++lRzCJGK1zZ8TAoL02N4YMfzivr9tk
cFERCxI8nNavp2+V1gq/cje35BLEjRc9C2MPndsfL6WX6uWnUEkWdwZNSYYSZtJDMuLuT3pWRwqZ
4h/oJPJs+a3w3lpRkABuvW558PLbIix15pw4uVRzz64xNV+DX74uvlLAclz0LmiKPFXpAkKPyV4n
avDBJ5dcLK3F08pt6Lca/RbOpZmOHq2a0Da60JhyX3MhloL4pSw8BCfwN8EG5Su16tivlMus2mLJ
qtxt2cC1GmmQT6cm8LWxfoli9ehnxo/DijLOjvb+EhWDBpkpkq2vHd7iHfsWYG1o9PbsWHRV9b/D
ltaz4yUsMBIp9AooAyedFuRyLC+qBRwfU2uJ1nGhEuWtJ+HkntI24AWdQ+IUeQucB+91m3OhnkZT
VJuUyptm0PLPOTxzgK6DB6mA9bNOf2+opA1sVFVdotXBrc1UAkCzub2bFcTPsPUc9LipPI0FFBG2
VEKtCuuPofClavIE1ePTPAhHD+qC6f6cR5IyO7okQbzYBLoanTJMrhYGXmbfrkMfKiP6Lq5kTQiY
vfuybE+ZDSa72msOsP0Di/Amdbz458SmkR2fnIdrAnuirQAQhPXbgWQNxOUue94gCzaRigbgaSI7
IyOnNNvZsH1abwCgBizcIQsZlWMF4JNaEFT6eLx71hpAqDUdUHxwZYtR9WWrMLDhQiZ3uYc1vewE
FdRMQw7mp0nrzmHjMtNmfBHYHgBtENtEl4ApFn2KJYXwVrAk25MHFZOaP0RuJkc+AOAaRMug404e
GPPJg7J2+oMegW43kXihPMmrGQIvfVq0aG7Z1XwoyKTse7ZBCyzqm1LW0i8v+D8ZkQZnnNppMOqK
0BEC1nZSPdZiKbLGyIFN/HZkuwCOOzgYj7BM5GuomnZm3PjKuwLpGqN7gEKgCiuXMC5j5IfW0+Ef
HfDp/E7Il/gfMS9OTq0o9ZFHJezJQmXxRrksBpZRHEDc5oo0c1/qNUFb10FgYgbtwinOI6BhOhkg
azzIbGH+GdwiPal1pdJHwP9G200ugyhBAa/dPaqC+fOH3zIJCA2Kvvv15JR6zYBBUayi3iyUOJPT
pQmwparDVUJWEhrWcCVKdvIladDjXuaEDhax2AA2/Y/Kl93OTiBsjtZqxzKgwOv3+LPqyWZpA2T1
L4Cg8uWtlRq8X0KYSJm4vTWEkY2r3gTq3nNW3cWYUk4vEXV7GD0QFA34ghV/u7EqdiSWp8hjSkDU
+t+XxKzxkEC25BVOKfONlo0YPB2wkXZYymC/g7u6WI6DaE5makzWJrGHIEXNS1zyRJ5CHKZtay1l
yWX9XgDAcNTJ2BjBGC/AyQeRGMgz8CrTMVfM0KSvXCgBaq8cNZpEuHzvT56nVSPjq+pxtQ/Dhl46
9XgzoSFORclXpLm1uXhaWk1EnztP/YHPAu2AGnEjvTjNHccKK4UPeFvzJFLycqW831r7QD6fXYjI
ZOAeiYfwv/pRIlJ6fHbJMfb6RybvDpHUpXVR7f7zmD7WRga21q/T4rN6cun4ROiVEyehOG8nVnwi
gyIsseIEa4zPXaS2NWziqoXvv8XaCfTPecaQjgfNLiBL72NhuQalb0dmH3vjpB5sSx/qcn7uS6WP
FtnuFUDsRL1tOpxWqwUFyVYvjU+B8dXe4HRWmE35Sx3PmIcC2LfhJRFv8GBsuY0eUWDf+EdpkexM
h9WE0y95cdDrwvy+8N88BeGJzlqUla2Pq2UvsnGAgKC24RXPvV8aQQqNYBPTKrC+4EdG/fv04aOH
sO4xOfFmP7O5t6aS5SLynn/GULdAfSv9fY/W/BtazknZGPbQdMSgLiR1GY6LpXSyqaOuojuMqQEz
cGd904VWN6AUfHc7p9CiPcjADYT9icN9vxgR3EZsz9yrkk/Ft+h1QZBd2au7eEmj4MyYu2JVXK8j
L8XeNQ3ARisOVuFZMmEm0fEIAO/5+iFwoF/9DsSLeEmHKZSPINknab4kSE9tDEpZxEXLTz4V4TCb
Qw7ju9lK6NlOTjlt/v7fu0nLrnoxRDCuahw5ghlXXdMfD+5lqQq+zyMB8WIF7cGH7kG0g+umGfza
bBujjSDjcDzjnNdCiLjf24yUqTUJ0KNde2EXWDCa7DyMczfJ13ZNY2dGzpU/8mkKANyIEYOnKyTS
QsyIP/U5lh4hTtC1usldmMzlec/hUB9T3EjuByjvYGgk0t4xIjBTJAVG9oGf3v2XmVA2R+Lt1cH9
b+McJ6AK0ZprqCLljc9h6pwTjzk2XRNOWjR3RfBGEPF7CqZnjIZusEkc2UGYTRdqNFVSv9pdeyDt
+RVj5r0J1oyCLN5FZvHBJEg70gR4BqhkEn0qw5yNBUaQD/plgist/XpEOEYAQ+L7eyBV9+2BOAos
X9bOgJW81gkBp+kWnpZERXJ0ZDndHHeJti5nxXDJnBcZylAiDjkJO09ckUn/ihniNkUifdUk7tsl
SgV9kTKratI8XQkCrCLZhPqsJRtDkwwXit7dRXu/AhI/Z2CbCa8bYpNkBv+zQGDDl8LfDWOMMV7M
nQ6nI5wJVWR0fwQnVpknFYoTq/aZSXKdnQ4KSrOYbZT9QNFcmqrUl61toTD0OL7w/u0dqh3XdYR4
Cc3xqS5sb3XOQafqxjTgyVugdTpeakY21e33pEfd0U2RMw0DpyAEvZ/2nxYhEoP5wjNtESPxy8QN
kBWo59rFa6DSzPNiCAaimnPA7jBdq4/9+cvCKWNRHN4I7bdURrXv13voHCS660AbkMofHl0AXcoZ
UzqqmDMXn6Kyn6O7dpmo/+BdOkyi42KrmUZanZPO3MK3dOxDnhVWMk2iLsYgvWsw1KGFS+itJ3nT
EdTPzedsp5FhQTcz7cB8bIbw9mEVeUj4OnFN1V2fOr1TO9ld0VAEhx5ZDcekgcg0U4tpj9Whrk30
F2B3LKZ7R/4pqr84okFZ6Tw5hbQEhCWS4oycbVvG86WLSjiNUS7If+Nl9mH0VF546PWsOM32NEy/
I8YA3ROhOVKpTtA5GID6VnzD8VvB0RGN1nHgeTEtLHwAyux01TFxAhWuyrRj885U0d5akO1p5R3G
QdPgDWNc2eCt1gkS6PWmLOHDqyWWIaoWXQ6z2l/ZlHmL/qPOAX5F1ZCF+engMaiq7sZ+ZkXLn9We
2i2fjk+uPlQzBO1WCaAnBsPh44tCPdtZkyebREwgLY5ozpNjuTmtzfc/sCT142u3setzUbCjrE5z
JExjk1XufDsr+g+gDkjRCDPRLYY2HLs8yX3asdJa8mtfTl7Q3m+FZnQ4gZivAkvrG9BvHty797hI
CqsC6Iknt8qTqzgX9a0STxRBDM1Y8fjJCUXiN5xNZljxdiOTEVdG/m3XnIAXkFNxpVZYDsqtuDwA
u3f4yPiQ0OaBT0LX0fi9pU8yFuWcIp1Yg1kgzNG9jJNvvofbyLnXAdJPnI4D1rdWPX/Y/bTIni3F
OQ3K5nXJjLgTUQHosZZpqL3qnwBwaD95a0i1bbRqTZ9XqdLYYU5JlVU4CblImirSewhOUj9RCX9Q
yXF6fiaF6OzfdAhE3Vt7a8hfoAYLgnWNjd4wgANxQWQE55bEqnZlnSW6m+I9NDM0cRUAr7WA7qrJ
M2q5F1O7bvHKHZzO05RG01WKC0z8p28NRHZkYOw/nos5UOwT2QZMyY4U97cDDCi4ZDfoC6Ftvxxw
fq0kVvmQO9YTDm1cjBCc42zVa+mqNkAeUsu+vhLtQA78F7lfiwhl+cOV05V8D5ctmYrksjRjRMxN
6lyHXyEXimPhnry3IjVhG3/dfcMBFs16HcldDuBFtTPJR/NdK1aAliqGvba1PKnD4Yn8KE2RdJZB
wHIjkq7fwcejIXSpWdUzD+8X0tO2rFawh3Tqv7+LkPzX+ziJdJlodqHiKhu7InYBqL1O8qNM+UeV
4HPa+5CrdRxhKz3gG3EqdqFaVbbv9FzfH1qrawt4hYvUbM8emw2Gg4EF4GlOjkkkER1y7mjOJXu3
b8LQw0RFvLeeFwBhPQoTKZmbv+glgxRC/XHGh92EmkDROUnHCAaf8VLtRz7KIGs9a5LVdR67Qj7B
4uVrLhapHvj92AnR8H73TZ1GzrhygdnkcdNvrGE1hnf0oQc5MaB/Hy6Lyv0XGlKgqIwTUuyIz9Un
gPgPW79f4S6GeaqdgePpaAy1jgbEVO0aaH6VP+odDzsyisUZIzM0Wm74ZghcwhHkXuD2hTtBSRUE
RwjbwzsWPGndbQOUi0cSNOu49V4PuIBtva2AjkZLOgTjmiqqoCmNqbzZi/79GL7oJCSJXnRBI71Y
av4iYr/LiyXIpIRTBLbUYel5X16UDn0oC3ii0GX69Ma8Wd/Rby3ucoB8uALqZj5bKDdhNTMtv1D4
Gfq4IPMyeGtaBJKcU9mJspB+52pNuHGOZj2a4WQxmxlxCvlPSH4d4jzjmXPQCdQQcZCT2fRN5R7C
Et+XBZK+9xUBJSFMDLuJc1ouJ9hxB1nq5BeqsSJcLFMpyPTzr/LhO2CKyzgLKJw2pW//P/C3SQA7
yXT/LQDSGOKh9inMr/+OzHR5AthP/QSkeFSQ+k1v6mL9BhYtlrpiF42NLb3yKA+JImnvwcu0Sl67
AfFdaupp+khgwcKkKWq9R+8yR6rUQogQQXi36w5mHm2iPwi6/0+HnJS7SpwEgII9D42NvH/GgRPF
STii92PssqfnXC4Ro8rsdFwpUtE0LAfptaXrN47IdDdCXppDM4RbPB6MLPN9AJivA2K5f7ueu/XA
r62mSQc+45xlWUaH2Ox6ykJ6AgxwhDHUcUJsqu317lJ82/aZ7Rz8Wui0xIJFUaoPws0mwKHzWC3e
TbKffoUuXmttsKGQ4r7fggzkjI6Ne0upOE/f8BoIt5Aaiy9MBCzui6B+yj1tAuyQcqPa2djUOxKa
gf9VoZDdyI4YaPJ9Ou2/fJeT9XnybG1de0JcS3MWvFq97Fkmve/05gVFnz0KOk7VPvweq4N6Ob0U
CKRtm+ESxyTqNd4IvNXTOrL218urEHkz78owB7xYJf2SYkjIv6CSNi1oTaGG2RhHUSFJqEEaNmve
6WKOGcEaNM1WhNfMpOqccpP8W+koZK2UOWSyNeDnRGztCx55Y7jrV5oZcPnrTtdwPtzesH5lRxue
in3ooKfhKhn83Tvp9MQDE6HZ3R7OD4SfqjH1kvG0Sg/VWGsz7/zjTFJtII5huNzh/l9SRDIv0D5R
FBa9xJbfpk1lDH0LN6Ebx7gNOuutnpuWjgKxkewc10M9tylnnLGU+qYh9QeNcpEqtYg7ulWEIc8W
j9awYaeVX33jlqdBpOYgeYQeL1RYn0DlvRJ10oW2TtCkVwDPiAX1AlO9jA6jZee0YseJKiVhahEX
nc/VTXeS4UXC+g9QLKFX7lmWPzrkyimU63a3iKwIGMHTNOT5f+I3I6CewjDG3bWYwFPCDJ0ne1r2
98b9/mMKf2QjyA/UDV8oohSUTylcxpxYCm8J19ICmFy02BudI0T8nxzx5LUEkXbvHMcC+RkgmBz9
d8O6nXQWUB9vhe9Vyuaovdt2fphOf368DNT3MuzM2QwzKERFtc1uBQ2sw2uv7oFpWF6LydIvfq7M
sOJfP9xah/wuP6p29O+SqGcRaItYgzImocKanpAcDLtyvlUcvpDJkmf3H48Uhiaa0V/AhKy5Rx/V
xoTcoE35I/QpHFzyfjGYHfHOjU7ah3hOkEX1dhSSKHMt5AhgBe7GbN1NTGLBc77ShMl+jjXMZEK0
w3EiIicKPcUQrOo4oIc3KYeF0gtW+mFef2/GB8/zUlhfDcAhPeAbUKVK63EyJVK8I3hROymZIGyz
3782M82yiITrcK2cEaOA8yW5NnvhJHaVFgcAE1bp60N+cIDtSA75JOAty90KkIs8pH3C3mS9u0gQ
AHGlKucD8gOgPZktvIjYXiPAaMYJj2k9+jrBLxWmZ2QxGUyg41ym0c/+uZfNoQ47yqIEoI90UND1
ywIflqPriv2UxQL1eSo6lCsbcJeULpqpf5S6WK5TcJ7LFMKs6KXzJt51p0xMCgNZGmw95Uw8pTWQ
4GYcnbffqfVDZV4iV3sk7G7MyUkXpr5k9cx6rTp+dhCIbNOgAiLsuThcLtH4NITkFsNCFE85lYbb
j65Sx96H5kSWqLRHrWZ4u0/W34ciry6PFfNk1kK9rx2WHDggpDH/o6UvCD6Zb8YT0SS7qaMBaGbp
p7yHLVEcg83zVD3DCvR9f1SwQJXQFdfVWjdzuj6FR+Rtge5p3flynMD1ejUprSgkp80rWWKEyqr6
cLrJNbspi4LKmz3qRWNYC1EBgs/Gx1vbK6sUSnqxUVY7regJAKirUVUJQ4c4YY6bsVtppAI7hVBJ
j45mzBzS7TuZSpsjWOfJVSTOe1xme9PywLbBsqvfcYajlzAYSRy0++3ViO+qnA+pG2s0yLFA0Ygy
eNcDFZO/YrFKThtndbc1p6XnS+K1kmI62y1cYoh4Kz7+FGmyhr/3XjXDTPQTv19Vz05sEaEzlNbh
Ae1Vkg5tw9xOc9MXS7owARc+d4dyAqtffgomOcQGg2S/RmIOD/Fyq8XwM2diFPY2kLsXlHHYypdZ
3uuLi1HMuIBRzf5SS9Eutv/GTU26Bbzd7+UhOpN5r1fgUc+p0edCjJOzo/j+25HP5GNb/w6Jk1td
8eoP9YNcqF7lYsRsUYORFQCnPQPU7NYrQOf9VPiat+tR60oYLnArlb5wTO83FMngShnCri7TrKs2
pBxnTit50cdWPyfSv0mjLkxJFMMOBvOlU1fPt+3XuIkO3tB+sn34HcJ+LWnoDSlHJ5+91Q+bcsbE
smwCAAQGl83bUQhLMM3DXX90ZFYOMsjt3dzosFV3oeQ/TB2et7aHrABWd4AILKNKs+28yW/YutFn
Ni0krbaKYye5B72baZqn/5VyaItgZL4nRa7ME0yXNy5KS8l4RuRgm+mzVoAgnFPBYYtjz8PPPcAp
Mmvx2w6ZcJMZa5dLlD7irCiPXQOOxjA3CrARE0SnvM4f/Jd+U/74bTh8AQNTi+zSDlw6++Rgh3Bn
eeLci39v8ZfiOkeA2fFo+FgcqKpw88P5I9n0BzGGHaot4w/6tEIBZCSsfez+W4F0Hyp5BZfeAwpG
n6AFK9FK8tV5i8c1n84EwXgqTJiHIowsOC4lLXam8Ouu9OxliZTGyWVSi1x4bgCoJUlSX28Bzcg/
13E4VsrjGkkwQLVHcfIzPUsovuRigJx3KLE6O2mosZC8lzjsTKT2MDLFOVwEtklaclC6wF46rj/D
Aczuzj5rTwxd46IN8qtMhjQYV3PNZaRPGbNFIxeVtcWz5qWR1W2S0gg8FiPyB+/Y6sksBi62G1kW
+VZtyzU2sZVs6YLDftgLNSdP5epvkBORxORoLmn/CSKRxF9duRFJy6XXvppgsbMzjnjS3QsOdXyu
ZeVoNlnaZ0trOJisrtqKE4Tb0qLxGwVLHKiYcS/fHyjj3GHsUvpM9lHg2yO16aQ3QAZ3FHJPWrrr
hWB6e/SynU6Xz//kWAMIdpA/AUO9NQG3PxN8deJ/pja7+NBgu61FcRv0ecMDrT/DmbYA2XWp/sJY
7GOIwTRHxYbk9xKQttFWryZXdLdZexk72aEj0F03AKspCZNyAlImtEyPUL8tBvJKMNNyLi1Kiuas
ofyzAVaXNXrniwzdV2AO6FuHMNLW9X/yNXvfdgPywuLSZwZ91W7cKhLZVzK74J/GSsGsvVQsabq7
Bhxqjvulu+9SnqwmY+1XA48kc8ow3ATzimWXRgkt+6BnWk4/q5qaxtwPTJtBQ52zj5bBsnMNr0AD
5XtRBcicTrLbJWohsfiVkpU8LWXnFIZo3MshmO/JCZ8V1sWQ/GzgHYK2KA3z/wjgY7E8cBj+D8Q1
/Cg344GbY68jWQM6Xg1/XfLx1gsB61tOPLWcORMA3DjM6AQshiC0O1yrnvX9Hzmxiy3gyKVCLN0l
z++NBEZd42pwKO9AvcUsGx0pQQZfK3X5fjwBHANy47PWYzud4nETb3yh2FKdEl75lEAfhKcNH+PD
VpTQwJlSeDxSYfxL/Y/cpIPUyKbAnmXRFwV1Bx2Uka7jTyCaNoTIEFYnf2S+jJg18K5JhgbGabyb
bOcvXySNsA9dSwoCodN8gP9GRwb5xWMGj9rWQ7M00LBiADfI46CsxvyVZZJQjpZT0U7JgFuPC6ms
jGdYVHq+zJ/ftNSKadRl90g+XJZBdARUfMAkcwzzIBTa3lcIZP/yjdSwZBYj0eQBh7Zm2yv7LsID
Jrt2kFxjrlFG9MgcFP0t74QH+TwZsjM8kMOiq7x/zANfGyRnudVWzVTpe6HaJvDNiHvIxssbLeOK
r9HiIXDnBLs0d2WffWFWx+u0h9HOyYekZRX3r3lCuVOAA+uWo2WPxtXrDv4REpHlUozmFz3qyS0k
KRJC6TvMrPXncT+oP+B8vEr7HQtqyclY0SjcTJPqwcXtfsy7SccYLlZORmofXQyi45CFR2Gmfs9h
PLMgMAb6UaxidajDFI0IXGbb0p9ORtTR4ZF/gOmQyGSao7l68UqSyrAVDEUn77dCSNeOrHJ/hDBM
Bq2lYf1+EV8RiwoSQIg8QB6ERboiwzr3yZLV/OCn0yMTW4ZH6zQ/5Mrn66AA16KP9hvmtIu4XTl7
D401xuNqPoxwzQalJrL6Z/lRFXgJS22IXxuxRHaZ6F9uYSrDPFW9DjOpiJRbtC9E6TliVxxxNpQx
FLgTilQNwBwAwdnsaim2U5KJAfqv46xJTEnfLcD4tiK4W2IAkJfFUADW4wlNi1t0MlFxp59GGBrX
M9kP2K01Iq7cLy++yZQI9a090MMLp6Al/7GGtumQCkcfg230Gx81Sopvn6H886vU7FxozjRst4G4
P22TpeCymGs93a2rulCvMpNtsfDU4/DXxXPL46JGC/uzA9L8Oa5GsDhQJf0EgD6ssJN3aC393gIo
KiCAna+pL5kg9gMMSFomzAdSb0x+vI3Ba8hXEfkdujoKkgABpImKW8yE9+ellUHJzaZ/tnk1JXx3
WY0HBMBPyWEf0P17J74gBrWmjaZMmHcNEwWW+QLuDhdqyc44l1n8wiKCt9Fajl9O/ywjW4pH3oY6
P6VpXt+YNySVpYTij+Mbtr5hGVVeRCKHpzckh1NX4oYwtXGAMSYO38C+YKC4P37Ge1ZWAHbwsYc2
aJoHdwiEudQQxCLUA5d5hPOnRk3Puv5N4TJomCft01F7a8fmMEDJ0GVyL8noscx4KGUNiq0r7PkU
EiMf1nAOnUU1A5v9QxRxqhov/6qJjz6wJIQyvOYivmRgRT6FVzDItvWhFzWKMODa2xeszwSZZsk2
0t52hTwU58j64viYIg+CWSsvzuuM3bwZW/lm74FYTibV+sHypBBRKyEq11hmbB4jPQcStzV5ODNA
3GEXrmG7NgthTuJqNcbR41W2pYRDxJsZojcQgpKgss/NPMbADmdnmqiUC6EcpREE8o0jsIQyZIk6
1V5UsjDKTMFB0EmzOJ2QQ/S/JiHYfUzK1f0YcBQxJ8Uj0IoymTOHkUD/VU+/2nvJNjm9rP3iCIcQ
VIe4oj7cCvg5yPZq1vba/KCmhyR9Pou9/OUHO00jAYdusNBfjhLuszcXgu7JolIDCgAh7GMU0FGT
Lp2PbTPj85M5tEgFys8c7SPb4ZbtcYXdi3TCBf0yAGMt6Nr9Brg07oGyE7XIjBMIYePj0lnhoA4X
cHyY65s9/1mJWJZPGW1mlKjft8N49hy2n81evFezPegM1AUSx0FUWFc2QwoAih0pcSgsGpkD/8Mx
7hN2Hz+yt7RqRs5Z1Ulg1Bo/LyFeeNW1LZklVOaIKcoW3DhTMRm1nCNRZrBGbrp5kLRrFYtazF8L
+1qW70Qp8WZ7gQJbBVidB8qRdauMhKYOPfDfldAGrYG+K/aj3kmLCWTRnYX+KGD5XUJaudIQmojN
4/LXRRTagM4x0DUhRBMZoFq+8GxQy8GlSy0WNeTVfUdEOqPd4ZNYEgCsQRTn8vg9Ufmm1pLyFSUC
ptu+MlTBlgcRsq4diC/iz0QToqwYYsY5URVYneVI912+1MYwwCuBNRdduC3Yprx9xKwuJQz+5meN
2f7tOFRNJj6/5lbdy/zTmsI2PQGuVLIoasjSz2L6QlK7H0A2fZR56i4RCBjxfo+pROqvcDqoS7lP
tfppmtF+JoJJTEKW+RHWNjX85h+f6CTlygksAfLY0k/ydTpkqeFyzX4NbxekrcodtDs0S9A+eQuX
srXtgnZVEvGHkNU03Wy7eWkYwNe+2SgckQhMAv8yFylLHIFKAK1LGd0FhQg9uw8/RKjmlLuNpz+7
IfImfXyqhOjXBzCL1qJco1TL5S/v/6O0CYvHNyz+b5xRoQH4/3LAZhMrzEfg4ren5PJ6DEfqIixX
XTrcr0y+p9A6jQ3Rbntaoq7gIzbT2tTDxib69xc0JD/CtJeG6kYQsQsWOaTE1yeYR/jAluFvUqOJ
IBAPIkY3H+6c3LImvqjW96b0kSsVemXtiJ2YVUNh18yCY2hwT1eiRlxb9Xjr/eonY6dg93JXZjNV
vCzPGY1adXKNZrczUpVyyJtaoN3sjl56AD3YeE39sUnTgCjAc4mOqR2GZuORPCrDjojc87qk8Qyu
FcMHL94C/7unmO4MJCsXbTNpwQO3L/H5rQWqKvVPg1cUuLv3Eo2m6guO8JSV9fNIZhyiR2qtS6tU
H762R1nIG/sz+sZMdWbwM61hr7JOS/sYjNiDakKtt6RmulRmPa5Ih8JTu7beFfMcLOtF4cDTzF1N
vFtiQ3hgxLn8w7bZCSt0QASB/fqMtp/CSFsgoBPgza8fggopi5P67ICY/m8JZmgyjXCCTe4K1HXs
Dv1BJ/lMNJgteV4DHcthovD+HSsKQAcGE7mTKIiH9Vo0pJIpZR+Bd5ZjbAPIv2ts1bEc9zR1u3j2
zT9ClqNfmIT6SJh5xqLF0LMQb8A4DkqHmDKqhzXZWkD4qXC6cmMN5zwTpjN6EAlyrbameD7H3sd9
J13t7zdJlagYt4LNZFmo1wEerB4WqaUWLxjDww35ACU1eUlsnWr9lCvcBacKZA4zdQ6gkOvqbDKi
wMBf8lCRdW/itreqDt7Qhv/lJecenO9Wxz8zxzYd19PKb/Gr5WHo4fCvi98rxCLh01S+br85tg3P
YqzH/Ms2Y910obrLx+edxPPsf19hjV8ysNloUMsgUyIaIqsujSBnA377diAfuJiNsl5P8WQnxdzj
7ep2m7exIzVZtrhxszGuZROc+gss7iEOjYPvbaGquTYj9X4NQ0ZbOkJC+mLE0Imqn3m1yPPYEiC/
bYgaFYjUjHmV8K0mcJVUmkJUAK4OH/4hW4hxS23dvYZETxBb6dwCvlSQIW5Gl/h2EzY+DFOXNa/7
poEg0Ig0svr4NKZORdsv8SU0ly6JU+iBLUEyUYOwAQOkuh08yTsz5vhUyl/6pnXSYouIMoEfS0zQ
3VQV4QvSgG2/F1HTAUow9+EDq6+hDJAPjzoFrAOqDS44ciMIpo4IzScGcctB7385ISbw3WHnq0Ek
GZGCU67ezK0lo7kNc/lWKcXvjnfNhTm2nGYtZ1ximNnCg6ToUSRH6uhswGH5qI8EuiWL1DVgVE8+
W2Z4WfgYJhU8zzsPSBf2WBlEVRuG9X9GWXnnlNoLpmg3ERkF1hKN+3R3EHUS9zXYj2QF0wCPY8/i
YiEzFTqCiXPRxpHaOwEyIEdIr/CzUoZSZDTZZ+xpea9QykruHmuYupfFxhd7EwmrMepjrADSx/Sa
lz05dLn0QPrDL8lk/iMV8AIl1h+I0VNTAx1IdWWAedP8h4SzQJI02h54r6bnghyllL86/lavRPHB
Kwb9sqa+7Z80uKG56HDhtihd/likrzv/72L7CP+Zk4tXZDJKtOhu2gR1h2OPeVX83NZ8+vo6ki7h
MIRGGNudIgsgIGWN6eKHcn/NmhZRwdKI/Yb0OMqmAUO95KbLuXrQaIOtG+0lhHHs7WZoWmDr2PM0
28XVZ7aWKpGI65BMnSobsQs24gbhuE0Zd3Aa0JscRLEhyShu8ba2pKBFJXgvsVbrx/IOEbxD8plJ
k0wSvT0M6tG3fhDNrW8wIP7YBowYlXSBWs5Y7ZjjHuBjImZGl9Uv/zUPQHrNBvE8UhiUWZNDntxd
8AylYVsTjSu4689ajUW1rxcegjOa9WDYc1+Yv3qccmKVnMFBEzzyWSfGg31N6VQlh+kSErhBSPG8
7076M1i6CnqRhr7fGTZ6SBOKRR3fSXym5TqPPNsLVWDH4RzcQ3ZYfsvRTxOA9Nl25rzarMsrTaAv
0EyAFcU6fB6bnDUMI/FPBhQPe57WcghHL5odETiwaeiBnos9MX+HVXvbAL/OuxrlF+H9D330V0rM
ktfMpH/3dRWPtX5xR1yaDHh56PQ0EySukoSKJHKgfETw1/zUg4UKiLV/ZET8WYK4mT4yolsahC1M
zKW4pYH/5EID74C56g914IUg7JTbbbCTLjqaPJxmlCrXMGZtszGc0mBtNw5HRxA1JX1z3D7zQt0E
k1fZCTnzNKLywldXGkOvdBLmswlWtlwz8at303B/rYHQc4AEnWUaeHi4eikmXGdA2YuhFHiOdqr6
16PHGSTPTw1pkHNWPsHJKJt35OBHCu1ECdXwEh2ptwKCIeqfi2uMDOqIxqqOOaAivSUxPWR7C6sx
ZDexvSO5ElVu/U8X0sJPT70IHPpjU0LBBj386ijhoW5ZeFwY1edcIAqV1OFhHN7x7Q/Ld7b0ZFa5
Md7OcU94z2noDT+WY0qnmsRoxFtQ155TNY+B4mQi0Qq9NoiaQ0lwVV6NqW7BUd85UPIvnV6/WfTs
a29IHa3MoCRBB0c6qy3TUu4polr3PZIQdn+boM+GIjJ34DKkQMVoUHOCa/IA4ZSHMKQYEZ0w6e3H
dMwu4dLUoVclsyNB8ObW+IV1hFSY/CME7S/WWuSA3sWM1I7xu4EH7IQBw1r+yoaavz/hcW/mKPHz
vn0uFELZD4GpTEkjayzc0NsYxQoW5yWaUo9CvmeMuVnIOFlezP4EoAyAXinVjj34bitoX63ueVuJ
xpS46Uu4CxtNVfl8D8srSc2if/OptmkACl8EHQizP7waOz8GvIIOyZyWfdFsyD3o455RhlaY0DYl
4vCReNMYcWnsevHKpZkmQduWTy5wNYmZGCoUQwxg/uacirb4NydPgNs2IXJjxzaYFAwbDKKaiw4k
Y+Ipfg0szGHXAhBHx3itS5lXN8pWRGAaHj/wYQyJ3XbPGd0taQgXBGb1vzo7frZwDl3vUOj7eRN6
WmRBFhyK2awOzZvorlq+x/NyUtdZiXbQl0Nb1pZYiAVEuhFH0qaoEr66b1jecocxZGRnC9TEdpb4
0wJ6DzRf3MNTZg8jo4EOwZ89SuuxYdqG0i3nnvbo7cFJNwliPwgou4YLP665/GPm8/2xgH20f+6d
9KWpD8C8Zpr0cO31SGkQRKyIm19o/dqCC3/TbTCcJCa8x7PSl4841qJHtmi7G9WGH6EXMcUN4OaB
rZTAo1N6jWig5TqPnOVAIYuBrFQPx0Mb/3xZOW+iYKkfAj4/sDo8qbl29ENOLqEmNWLXr0SZT65u
7H5O6SjyoxHw1dbs/deUOd0yAsbDqnGcH1CMtRk+WpQTiK9QDlM8Gr+XWUc6DamnufWZrirYFum7
Sfjq2TDVlryjDgx7tIKQe8euJr6kOykAhxQGN1czdkual8wdcAS9VRWswHGQ2LciihRKkx6JNYeX
DJ4lxMPSq9GuupH1l8QXOjurPJPYUN5vad0CTTCXHxVbc5Dv3iWn5c1kjpSffiV1MhDSE4MMroa/
SVfH/vVhx5ebFyER9LtwhPgf5WHbUspEIN6Wg6Ildcp1IaVhx+VSbmyDdCJdcS8qZssSsS8S2lSs
FvZmBgMCo49i9bv5p+nFOe3PTI5JfVNx29YwzZh+U03UDmqhn8U9PaPEeE5qMyaA674r3xK+/smr
cdQXO0zw/HVabhiw7cu1DZZhcg0JihcN1xnTrYFnN3Yq+1mKPsx5MjuvJX6LU9NAY1WYo/PoQkqf
o87iOF1L0UWgrEeYnR7wK4uBfWdQW4oUPmo6DsUvc+4X/8mChK//czcdjMsa4p76uwfDfrW8ZJo9
TfV4zkVIxKKce1WnH4RyMYhmCx5j+vyj1HJ5DqFL4yDW60aMR778cs6wTKiw0evtuh4YC47RziRN
ZAN/+Zw0eNSTvVmTHm3yNe0la9N1nNtqt6eYSPsfZaGDXc4D76rmXtH2JMQtjB6QCZXXRBiNeg79
4djqqulHYzcx+C/0rxKgIvrxhpE8ECj9YXvg/av1I8f7afN4AgVXaXzzx0R7vBoYgWXuUpyO9xMT
1QtGgaYSHQ3DrFy4pVV2Bf4wEz4SUbSmtyjr+e7EBoapRbh9FjuAEc3WvS8sipxWqUxu2yRx3mK2
YWihGVlOybnP9fyngMvGHYUOzkxnP0xpJ8cI86EQlpPNjldD93eQ+zWRrnw7RYf1smsDbMuC/8P/
VBHRNkvl0PqUC8t5YraaUkb6Y0xq6rnuOtTW7/inZxNWOBXF6XAQ1DIAMHZY/I3QIiUG/1bQ45oA
YGxcg7G0llT6c1EGI8UouiNGIbXHMp1rzf3GIUwiiISTQRr9BI4j50SvP98AyZ96zbWCkEuJdTjW
XHbAlmBqkHxfxzx0M7hNRXvm/RHwFVoclJ9DRMVYdXeyv1G+SdoWQx/fOw6fAkwUH3cX8E9kTTdb
0Pzmtw8uhH4mIG3NdeHQr+CY0wXtMx2QcSgF3SE8H+sz7hT5icEdrObSxL5wqsWx+MEngbmsH7sT
t3MHDgem2L1XoJYmsd+mlIsF4z6bzqH52+OpNt1rpC4cGoCYrWVTzCZDwW//86aJcUrUMCdar7nW
+ROnLsHR+WboolNJfDl18/AC9uXIzXWRMhdh/UtZxPOBOj3fwhh3eLjVHVILSYjja9er0xDA9hfr
uQv+ruI86h3pGrr203bKLWqNLXkQUpVlOloyp6X0oPi4lBzTkLdOreBMDgo7smXlOJDjAX2ryCGY
xojZbyWHWAmKhIKOcAC5AKhq2sI6lJKhJ8GgHikhx8k2Udny9FxHy1zbliCsUtHgE2q4HzjNFIUU
LNk5OhgCA56psJH/pPAUqeGnDcbvc174cIyFyCH+KvzC8UHE+dW3UYZmRP2CgK2QFdeEfK3Xx9Nk
cUkXFHqD3EXrFrcjWgBi30roP8B2LjNJfAz+9Ey7RmNc/e1yqzXaWougythuLOpnTfWIFczlQapV
fuXrpe0+AZpnd3hoADvuAr1mkXWD370+haHufjkBLWE6wEC6TBzlPJHzpZu6rOsPMRRbWEJqwhp/
Nb67sAG6IEckQWaMK1vUdW5Jk2NN2VX+9PVuf7+X4WUbBFSaKzbWWxo/Dy6UaRT9LV8/L5ZwOaJe
eUXL+IgiX2y9v2ZcLqFetnr2EiQu+WI9IRhGIJm5yXGD9Mof+bs8hQltdj+FC07yy9g/YDaEiHkB
ejVjWEb3Rk6lYSB/h9YnJyiJDwBfLaG3ejAnBu1iMcwTRoWoDP8187Gulo2PVxOMZptbSvIIl+Gl
ssAqhLl273SI/ugQHKenN5msSPccQcVRm+fWHjZ240n9Hn5XXxorPkB0YJsUA5V3huSElhJlfb8g
EJwo9VJIsRZK9SHio1SP0hGHQGiWnws8lc4pqopzmSgu1x2ciqAW4lLwpXRLr+Qf88CUEqELx9tr
7frh2KdYBxdAQXlpQlqOh1EXo4RPg6AC7fRahb5cEpq+aCjveOu4mJTZIkQBIcBen1KuP+grspVk
pfL+N2mam6SDH4Z4YLjoxmBhctuTLkhzWZLQEP3Bovy16poP1/LX9CbEo3thbCVPyWmlw1mET5UK
ehzot5IbeQFvYzRygL5eIZnRORhqODyZ/o5FIxtKwuDkkN1xETShNRKwhSbiocUOo929m589hoii
1cydW5wC7VLereAvVyXNHU683FgP/cN6fAgiWF/VNk8ZUHHx1gW6Nd6/kVBXLxf/zplGzxJo47+x
rkZ5BhH5OvxXwbDexbJoLzlsaVH2d+gNsQI8alUvvi59K2dwVxYwgPOr1q/IB90WWmetr1QlxK5Y
06nC9+4JNlcX6ukbaYZiAQiQXeZdJmZSw1AsnH7mmwsJO1H4TPJfP+rOXajB+XUQ33o/OrXCRtTv
R74OQzjxMAlu8QLhNc76HtWpuqnnvEiUfjHAd139uUvdS88vmp0VP2mlslhlSgUuPCa3X/ffE0e8
vsZ0bHtDyJ1FzQYSYhNVQMQJzPvAnETtdGOt+osoRreJuR3q4gNvigtEzQRXdzBzEMxXWrmkFKy5
Sm4wshe73teMZoUB5iK6SSIW6eTnVqJRIAmHd9SeSY7GpwtCXXGRa6rN/5l4jABa6WWe2AaaEqHR
n0AXQ/pN3eTW1tSRcLs7yH7fKu3JYgs2hksspmji8gpch9dbJXCMjmAch57feKlAWrI7a1zud8P2
0JVlHjgfHJXe0wV1rlZ0HWvEpPFrY3OK4yGOF8H9ORxlVAseGh1XlRPs4+xm0m4VwLrTmPn6AXTn
gLu2Ieh+dsZevlF2RDZS9s485JLrE0uoGTVsP+DRkHSAQ4sVLb/wCaZbrzjZUQUIWt3vB+0O45Rl
Tdr5gktuvYuO/+bTqxxXEP4xFF/7UL2EpGIi5LDbvcCh+dTC0NkTf5rytsKkQ5BBeYkx1ayn2F/c
NOu1nIkWxvRwCWWPXTIwklIFuI9DE0CgBPfxq/ylFpvhONj6e9JMpkxdRdJCTK8KbMneZjSoGgg2
LpAgVCD1Yssu2We8zCxZ4K5Eo72FmaF/1Uk8ke8pHoApBhM7abX8L/J4K6r/xZJzUin1nK0Xierg
1JNMI03Kty2yLgIjz53Z4qfvI5mf1KWz0c9VtIOUQ1tuE5q/X0BqcaJRc1xCDoWr2RJpcAeSosW9
exTkjvGC1NORiLxRUyfugdykzp8n/Q4HNhMEXD4FuIk3hGtYzpteE5/AqVDIwXJUxk5MHrKu/cFp
7KD0Xg2x0iVRQN5F7U4oKjJPRd0w0iJy2eO9YJ278t0g+iYZhn9VDAPZu1ZT/3T8G47lgCeQ1MkD
xCAfi4ss6xtQx6/PRkagAj9AVoApjPkOOZ69vDnseIPgGv6ay3jzYEr1eQisyiHJgmzBpSRScOpV
neWMz/n0mqIceOMt6LSOngOtYBL3tTvEtSWH13w8EXGjQq+8nXHku6dxANbPWsmfYB6o2dl+iZyU
pCKvgjEcp7RRFZg4JK+ZsU8OWm8EVUsYLlyTqQlqV/ZHaMaXXw+zkAXZ4tepRCl7Mi7oARL+tPNX
PdvAlvI95hUs3VEem2CoHKwStY3d6EJe7+/bvbWQXILs4mmViwJOQ6kfseeMQMJMIO3DfxS14l3h
GdLVdmksPGz2lZ5YuFmWJ/1dDoYHwMyGFBkcbPCW9ULwUy0SZzfaEAKlLvc40tEr/yMm7pq+Ikm9
7irHWhdxkcmFH7g9Itrosp3o/dj59q7p/76vu4d69aDCrUlx3ssCqpjnQxgmS6mCzt0HAr8wFQSZ
WaBh/VwNbZhtIEeuIQ1EuQwujQHCHqlg2DXuR+sGXPt3Cqz4c39laXNypqrkl0ZuWEGeWqeGsGYQ
UCNX288HYy/1TFg6SU/E5PykcBPv0U3WKVhWrJoKikdjgjBRJ2NPkOHs/W9A3ufW1k4qA55hQ6aG
RPRlse68fbOHScdRFBhCwXkPW6zJeV+wVfsJcuFdo381YCjc0t+rw5dat3l4zJQWtpfXnaPIGuqs
PkBruL6rZt5wIY+26EVGsZwv4RqAOB4eRqwLwbwRAkmtXf/4bzBAtA+xuUeDNFrSqoaxq2x1fRBv
m5hDKFBO5tLH0ScrGNEcBIZHjgh5tN7MDLh+HGwY21qoXhAvdM0Iy86+019O3Zm51pCCKfGxgil+
um6tLyZmqIIBi4CW7L6uLnvapFltinQP+mtI786ouUXPoxFuFQCUVQng1Bf9M82yUISbuwpPLPNI
D3Ki+t06dugpGETqnkGxEGQEtFRJ8VKwwHl2Q/Lp2l++tDujdqCraqqrBtNFUn/8S4nyrNqHC9bU
1EcBhQJC0KPCzIiqOsyT9ldW1CxcaRwaYP4m9Wlt50PB/0CBYc2dmTX8MZNOxBokSRje4SGl6DYt
jefI0gplPTB25RYKTjTAyK1kAf/foBbqMMWRgAU4+19Sg5NYYxmAsA3gG+b8i+QHwBbiR4bYHs/e
/vdpqXr11cD0krKsEkqUhTbq3K2pM7F3r5gP0ovzdysbDvfxBKhBxvKfuASVyyoV9zq9txcRrlAg
/DizMz7Eg18XnNuvZWTw5qxU9SNHC3R5BZEvNi2a54OUilircDj1QuRnjcRgLhs403gkeTcdEn/Q
4izTvJQDIJpFFiZPo+nQ1g9Pb/ApOPmL1xo/Ckoor0KWqcCbKN5nIiOhqjrrhiJCpNA9JwxXkmI4
mJrJD9F+P+AeBGqd0dWln47sHj2hPeGNNHg30JPlQJcPnYKARppYBRhyrQ1753HvsDb+3bXs2V9v
Ilb/ECUwLalWTFr4I5FHuUZGBdpzE1k55XWE6DtMNd8NzOn+6p10C3gPOoK4bgRsZrFMRs8r6pJR
udUiPcpTenCU1vZuQvkB3tgTTlpxteKhsB8ObAMs+ih7ltn7VbHVACQghI6SiGhBvyBSpJ6iKBL8
zgaP8wo6jB/1dA/8am1XTZ24vZSuvkEHKZ96ErUlAq38rdohuG4s/7PthCVIinEJDSbN8v47z+oR
O7QDBrImVSX2TN30qhRHojb8aQYvJWMVYxVfNaQdqQKQaPswF00dZ/SophKMACSKd+0DHc0PsRbd
7rBkB2JY44dcD6dkbRj0YDo0sPIDjYCYP7Sj0TCd0RT4eMKARAkjZx3HmaX9Y4neXpU4qMa/A5iv
h2PqRtDVXdmCxOxqMvKL8YCVpp9Nk5ZhPNgbnWz53AukwM/1CJVwH+vmV3/QTdPRohJWKYGoeKH1
3FMwmsPJ3GBWZ8XThV6B718R9S81mRDgPSHRvxPx5oh8QwYIbZAODtHocBsLYXpW3+jnFlQsn0qQ
L6TsiBWxHzSDjZE6rwqV1E7+2oWHoQSzxoIhBzGBXerfpZAeXhV3UohPtW/K8Ts0jfE5VPab1u3Q
MkdEVMrdYl3bxSjY+8z5qEcB8zhNqafFiS3HelaeHl+pSfJvBg03u38qpLf29C5mrKKLI/VnOvb6
Ma47+qsaJ2L1D2GrPYgr77p219+e3sj1jC7bC/RZVJHFYXDq3Ggh/T4/iwR1dQgav376JK2V7HMJ
EaXnHJYSVoDS6jECtHgbw0vUxrgFpH6VuF96gKMoIkJycfHjYVfnjtE/8Xlh80UWkDidS0fTJDkA
n1k4rbnOX3mvmWq6uWgcjWEOqiGeNTonOPmYMKt9PDAqYgoL8OXi/DaT3BkpISQsiXz+YYs7lB64
R/EcOaek032gksIm34BQbwPiQ0mMuEBnn/+w1C4kOF4DsZqqa9Y838v7Z6Sqt6aPtAxwnwN0n4CT
vGYQyFTvttswJ9bXNQd5KVUoIEwTgEGL6sMaMucDVuANFsrT2FlwkEjX80E1samLxh+hj9wIKo6y
54Boq+ACEK8uJiRTfZoeH5Of+K1Yd9sC+bfV8/8jth7tQ+Cwl3LaZfSq/72WBGTC1cvW63+CiJKJ
jroB8BW8lAXTMwYqFPacI3ujN7RsrUzk62hazsG6H7/lejcPYPruzFbQI1swZmx3Ans78tRuSLi4
IEuZs4Hb7ZUSrY0SEcuTWL7/eSKCs9eEu87HJj6VI7JIpKToZGd6x9IcMrKrHzDDzhzvUNSwSMWL
jX+LcR3tcZqhY0rTJWBTNLvHodLz+AijU5GswHcBqjTfIni0ttdG26YfeBmVDtJnX/oQeXXQnUFY
Dwp/0myx8zEffdM66f8Y5SsySqT5QPOpE3sK3Zcj2CLarvYN/rB7cu8uI+Mu5T8wKwlVinJLXP1s
ksvlwWTtqI+XVOmROrC9/+cRXAPlM0YnXD16Ha3d3zIHcH39iLyN4V066UIQ9gQtVtk2k2Xby/oC
58UCpt88Hr4JPNS6tIxiqhoAyuhIvx9OghCDTdXMuerTupBbyuPhWDvcKicpO11xrpJ8yrQ3wROe
rJgDRI7UYZP/NeMCI8H7007NQC/HGGaGBlyuBg7rrOK8UmcDb62zXzwvUxqXDvYdb4vC/ajcjHpX
cB4U43bxvFPtEJ2Ggy2VvsO8nkBZBag3wjqsBskpIYTDARhZPWa6jhMAMa8RbLZOhMJHvyD3IGyv
7hmXWy6HPK/TOjI3WOhtJuv9WCRUtr7ZfY+/6fsPfY+xpezSpe/BfpZ7vbGA4/0ZFZQ+wjp/ERRX
y8jGAqfzGSPxrD4iswE8R5MrRdVTutyhY1D+1R/vFyG30r4A5pL78lPHz9AgJE5HQdXHCbSANDVu
Vs6h2Q5g+6dkVQL4o25co1KPjvCJCKwPyliyH0f1CWaFPTu6TowS9vZgAMgOtvIxninZLpQ2hbbM
1busRWJAn3oAinI/1TY5Kg3cg0iOAUxrcQxfwbtOKorY0wW6q+mB2oe7hRcDBKUZaNqEwNi7MnaJ
u0YK6ht1PnypuS23iYEwx6wOv0bYttR8v67ehNEVcK2fuZDGQ/VajQN/pCHQYlq2O/NFMpvnwedm
c7m8Dcuahp+wUwQV3CWvgNZXZ5v/PNbWskcnYtEGt3cfu3Nk5jhrE7ubQHPbMaX4/4C68c+X13I7
SmsM44iRgnMJC5yUtI1uFUYML2yjyRjSEH9uB00JkR4rrq29nRzdt/OQMb43zjCwMq7ke1LYkgJZ
JKcqDWYiMn/dIltWt4bV5Xc9/cRJXPr6qXyGJQgeNLvrJfolX7g/3YpTIxqRY0/tOPAxGsUQfRtt
AUxLoyqyD56KAqP/1B7m7msyd8mxHx6D3+PE+JgbGPltAN8S8opbx1GJoWvK1j0i3+zZSq2kfnje
X6GaBE9eteC8P7qxaDm5wxELZrcgLnuRl4DUqP7Db/Hxc607VdE/iLVtaVLdexM0DBCcABauLKbU
p27Gv0gfQ100a1cDh/Q4suh/xkLXbnqU4OVozJgHPzkItFzuUwfBqMOed4k7hmIraSBBuqNE+FrP
Ru4J1rZWVeuoeVthq4nKijSFRdKkCfKepgW44vFHPT594vhD8jX9gd5vVpyB/mTgll3v32mNsZ3a
T41WNjjlQbj36uayWPEHiCcDVrA4Ub3CnDhfqkoxp4DkuXXjBpztIpI67ew2A2y7Vm+ycDTk9D2X
JRky81WsERsbF2hxpvGtJtSrGRXHnewnukVOjsm7cgQ6VM8irF7Hc78HKrTHx2SRp5VezbA89pmA
u7aPgHnAblIdLsE9pnUoRis8zzDmjRleL+bFW52xBAChNgq0ZQd+Sg9CDuahBZry1kHYI68LAwPL
IZQKEo3OUza7uJ7FWSsw3MI/Bx1jX3iGN91xqEGLvWjhkPzgmPu83gY6FPyK+f2Rb7uXpfRGwFvz
ZmKrQNLiC/O1NlTwmAZ5DRmmOzQCNDegbxaTbRza8x8bkX8cIOmZvY9FEMpsfAeA+vdme7mmIEgF
McxbKDecRMxs6r7Lctzp5LCuJRNUGTBtHQ17Ykx6l1KlenZP7zKwBlwNe/lBKM1kDySXPNiKWF0R
j48nm2G+/ASMvvYbpTx7FXi9uCn5i+GDq/2rIyNRXJjDSdVdOpKbsZ1T8ndKsNh7cftxzKEqDKqb
EEwELI9A0y9R2HNufBrRGPAQR+2QxStX1hu4bk9fnTO4PK1v7pTGbzWOKVqygKfK2qnzE1zohMsi
i5igCHffS3/jpsxjsW76xMAY1JYyPtdifTYvnJOiPuoPIwZdKfHdkXrtMDuEAhBZUSDuqD1mCjr4
wLPlZTwD+i6PhS3GnL3WRdBn+xYTnEqftWEDZtsFwgWPtgvzrx/S1PN53oW8PcNb305prjmne0Uz
+l2tQPwg9QNIpinHgY1Q2Ap9hCjdWBCJGtacZUblfdwcv41sLEh3eQ0NE0UsLcnfl0Yk23Z+L+6d
b4YADJpLcGuOmyX7ayjHWOWSR3hFL0KyReIx0j4Hdgor+artagfBYpRg1fxiWYFV1eDBBTOD7D8U
Rf+D9o75QO/0Iy2mq7xDOblxT/AXFvK3bVE1U5MS0qv38ij7w7Fp6FARq6urk0/xCM070znv2DzE
FFqheEToj05hTXFdNJ9KG+zqym4xyt1/iAPFnoGVJHz14WcUWP4eAFaT6is7cn43xZUlzcPBYBkj
7OX1Me9IxqfIi8gizx4iNnULeYKvPoQxB/+CdoL789Wro6JPgkgswU4bodvxuiSUTzpgcJgzdyza
1HoL89x6/XkW2p9NfYm0x6eonQvp898J0HcH0ARIp/knCWqcVU7fAMI3IwYEaILRirmprLPqRJBw
kfZyPz/wmgibDTV9QwiX7s504g5BZAM20DH2Kw7ddi2fV84FuCSq2NNWsKBPBocwmXUfjLUj6sSR
51wF4TIJzKEx+fnbi5ZkKUaD6R9D5muO5kjnyUjWwinab5GfDi67BN3zDDFAbis21gy/ufrTBK+w
Sqr1n5hTqzLHEvNz2u/CKVk4UuolbUji4CWlKP5MZ6xiw5iWgt/fIDxNxlveml/7+Foi5eCG1GKn
ZUxMaMIF9GQF/lGiiS+s70q+Cq535s6H1Mi2YPy9JpTFEbvjt2ztBUCTcp5lQ1xvMROqaClDi3jJ
FOjxjBdy83iePF9ZeKW2W3LlSbCXkkQbZ+3pNJxxoA1ibP87DYvq5nI9Tnx4lxebnzpmQbWotk/l
GslFVOvxUsP1Q3+Eyi+n85soKkShxUpvWj5UAyTwsT2hj926ooDdt1+9WnqEfQBHbzmsgGLopFIl
4yyCY7m7wrBNxY8NwI7Kt9WAynb9pNPTG36U8N/vgWLfNdJQI0SVF8U7nyL0MJvfSVO/Mz5PAfUk
gmQav3pF5Uia/p717mjXs6yLh4vQRXsItUXxE80hybUtnDVryGkuIXnA1/PvEWl2yI98urb4c1gC
ifX8SIDwGTKGj1HnXUBwDLJ7DlaMeHxjzpjJzMXq04Z+g7m1JO/h6YYUNcaGwkEneLMrKErKnAYE
K+KvS9sBx4u9NNE4t6Q4XuLL8l2VV2xeKDsLJ4Y2HIW5iyhEcKK9t+3iqMBlSqdTrKozi4sGh3zl
1bovjq9+fuY9OS0cO1/MFdyryguQoOsnMLeLs/ALVWQIrwBKzxBSnfnMjamjJpSRcwukKvR4hKFx
huhshOhRs7OBeV5qmpXDJzMflOQihO0ipWTaryMvrXqwMGBiveIljJIh+J2vun1txM2IWm0aIHxC
zoWJKT5qGHjtg9pV5musU7xSfFjUdv8SReozrhO6iR9VbVYMsRIeGkFCbVrZzrTyYfh0arPxCME+
O/rq1WPIkDkqmeHWdhY30KVnhPM5C22i/c5X6PZSVnoWEt9n+ub/0x+3dnKLvC1RYQknn6bXdh14
X+BTYFjH9WTsnMyqhsT3ZILBYDUdIqafGuYgVOqIc+qmSXX1htbc3DfIHsdrnvPgozJofzIqTToO
399yH80tz614PCj9Avyf62f+ib+0ytOmvWeqil3xN+1s2B4KF0o9TFciVPTVOvw0W1uN/eCQ4iEq
kJHex08u7Gd+ArUuG+30t6wB4wIO2d4/RRv9z+pH1ZIGBgsjUHFCE5dqpWaKaylmLdGyUTUGI9Qz
h3r0RyNtCMU0ZWiaxI/hayDmSU5wyKiwzzdy+OX9Xf/SwJcafNU9P/Xxi+Ui084Ze2ygzwEM6Nx6
QoufpNyviBJz1ASxHAZmIYH31DMukkLubX/jTtKyPQdVzL+GLf5XjuSp5w0EieiGb4A0E0lWsxvJ
x7t+0yFWU3adZ03c30QQP/YZZQEP5MgV02hAowGBFvdigs3Lt9O0lj6sdTTc3W98M9Cv1iv0XTgJ
wH3hsWvP+zPhqOk6nsFc0n0/tPKKVFZDH9OUa1O9Q6CGjUKTmlR/We9GPyJjzi0PTJnTKtxvA5uH
MykNT6qY2toGSzUt+ZlpB9P1alOGvwkb6DSSpvcjK6yUTkiJBHxq7adYvj7ipXA3sueUXWVnodjH
4e3rJk4QOF+ij3dF8W/TJNpyy38zTRjRZE2OHUNM/ySZ2Hn0wMzwGaFk3XF5PCJ2RUvxSOHIerEY
1ledByqVqTKYrw9D1GK+o+dW1IKaCEYYZg8yl1oadhY/DrhCn6dg/Y229L9SDYJIEpKtryLzvhSn
Ph2FIHe4OVd84narYUezRDnKXGntzDnnfJqboZX9SZi8Ng6NYev/8aGaGgRcTIZCQN2SxxfUUEwL
cabiGggn3R9i6b538NnBlGMwX4eTRdxgoFPNXsw1SABCNRLBaepX+QPdffFyz6KIqiyX/Zkl+EmL
tIXyP+Fk4K8iKEELVNY7BOztJEemiKzkdiQkUMwNuGPISoQICt+gpfJjmHusNimv3rXVKHrPLkYf
7qJ6BrSJlSqd9FAPmDrwV1JXPCqnQwYwxK+z2kyMfwELLeFbVX0SuGGdAcEHWEeTWo/vPkHeVpuW
PzE9C8ek40Dcf/nnM+C1JgRQ8QIDIDbsdW/eyH3cUfJvHEF3I411TPD+bbJnUDtzhap0KcW6IkS/
ZQcwNlgKHH/AlMYOCkTe3bO7rnuWO17atKtlpXjcgJRC0I97Y12evEXVX7HzBBHBW3Y1MKawNL8R
xoL0cZe2RLvlucDHL/YbswjvHKs5AlBA3KitX9QS198/lzp0AVBaOB4BhD7kD1pzAKglgI8PvSGd
244l6/k6RM/gyS3C/zc1aLbSbgoCtmercriN4iMnV8w3o0FW71xj8UlVWyTj2MfbI0FAyHuoqtyx
tZyCy0aBxBapkyxWuDO3whkqi1mR9TnmFDQF56wz/IQUUkwtih5tkwLX7SVPDXLNTe4oVTU8UR12
XFsesdmybL4QIMm+NGG0anwvI9cmT6FT/oCya2CackFx9OS/nKy0c5RxFSeSimUVtCbErsZukFdB
EHh4iiN0gjhb1izIM1jWEueodoNYq3b9G7D+xmhKS0hA1NYhIcTzU4D7LY9djGZtQarjjOjk7ZXO
L/X4FwmLnQJprVsz8bBmAiowByDLQTKFfonsstPZblPOd4JAxhl3wkb5kFrz+IsaHjnWIEcOI8rZ
twQl3iaNRwqCh4LIFuZ5vDvaetVYx1WIdkTnf8SqGS+PRvBIH6cyHnVJuOShBwuPe2s3X/bau9AY
0PpI1XhoARk/KFlk2Ludp4sIgfiy5bE7GuMaeUCgXuLTlBoKX2xh7Rn6QtGwWV+lkH/dV5fc03Pe
mqJna5ZdPt3z+8tT3fP7a//oCH2viM0QWXykusa3UjpmgLB4tywlFS2nniwdYC0VDKTO+aXor7i2
fH89XtGK6AwIZo0hhLh01gThJm7ZsCJrRy7L+Ujo5PRvfd72DYl3x0pfKrWCyRqPOCxzKRH9Rje7
8D3DM/iEnxL2JZIyiMaTfCYCkahTA5xfxqFYCzXtli731VrpszE2FeyzTGe3n9PDirdlG4c6DXyH
7fsYLJ8S1K0MwEvZVuuZ20+mg73R5ZbDictkwPxrYtBTrsTr2R7yHGQWCas0n5FA4T5zlBcUA6/v
Aa1ru76Vc9GZ2Jqv5/xdTabs3cH/+GCeIAC4Sbo57Cn4cq/9ew0YI6x0fYijx3BHo5dBSs5WkKhi
TCPbvHjyuwPRkX0YHwgeBcsmuKQHUU2wv1folc+wGXxwBeLfYSOLgWCChOdCuLzUPeGKAmUDb8nv
1ExtqLKi5I6tDGCDYYDqJ44+fTQ8cYHbuQpRueltH8dyhlQUAsFkf/C09yN2lK7cSiLkoV9oUDWS
vDSvnr//yJLyCxtSZNuFbx3sDA3q9B1uSsEFVJofZ5lc3d4g6HDUpTsjJgLgpq3haKru6704qG7O
d1VeejRiFY9mQXtPABZ7m2IYXdfHHH9CeP3TWwwAL140+YTDCiYTvLn3YedyUFtDOFgDwUJa5k12
zfFUWRK7IDOEUc2z9wEoYbcBVcQdfHqB0ikSrB0J88LtwkOFZJlhILVIrvY3sM7dOKpA4TBAKpBP
Dwds0dNMqkuP4EMUog3GKEdsFkoqAC6zW6etbd8T6kPbZa9UhbLnZqwXal25hV8Ul+NawFF1JZA/
1YQs9TqYarQO7PAOsO09mLXP66CVcPmzq4SKtQdjbezhJSdDpvPvNZacwtS/Dw0fr4Q8Y6FQnVIv
ZVsFdcN2qsewaHMTD2rUWmcScPdTxSADolYEFQK7aVTi9nENzCu4RE9jiZ2aq6vqepNc55WIjumF
+adq1uq18dGjl9Wc4Os0KppyNuUBvWJw9+NZsoL0TTgzwtLcw6sLeK6EvTY0DYQFyhus39uEp0UW
txOmwzjuyu7CvEQh9GeGQe2lMQek2HIjusTF8i76j8OsclUElw5p74x6XZ6i0e4LSanMnqej7XGL
1nLZ9ak71oGMxYbe8fXKINNlM9zx3257cZAzfl2icfUdrFs0xoM/ptwUJcYmH4HF39+dWiiKyQmQ
IAj/j581TV+2f7H1xiaMBrXGnLsEKxsE8PziPX52q8SShLcmwYe7YaxNb44ckjokjknK8kkaOStP
9A3UJDJFOPKT+ghkrPyNGhT/cmlaQuFXi/LQlDERB7lE+nmG3kETdfvjJAfMeUmfZc+bgKaGFlN7
4Bt32lf3T8AHgpwcwqq48ZeUK1Y6czoqwd8RmFbcuOLX8/4BbF/05m9pd5o2xLlbjAE62GO8P1Wm
egh/6xQRvVeYqIMImlbmCL6TqSunHampfr4s2Jfid9IrtvX/Mqih/XQOgf96IN4AjpPA7Mfqwc+x
2j+EXJGqgS87oxF/MdDqGGRiy4hgGiTyEiEQTmxWrv18+ZCX9KMX9Uexz9lJJv+9zPMOat0mq0Th
NP25c/m9Se3GH3JrEXP5iqTjLiyRWxvHLk8f3T1FxY9barTc+yDYu0rmtpJRnLxL7yZELRE8vaeT
1+iHpuXZRDm0Mo3w/K+3JXmRA57mtv1Ck64AczbnyC5N8757EyluYRYfukq0hldxcRDbSUtW/5in
bJ2STZydjnHTNfvJAaswBPpFDtLxuUkNKN2xbgwczVaxRHy36PZ4wMj9ive85Exgz21o8fjWFmR4
qx3afOzhMrT7lxCFc2OPXKmN1DlhcXDQuZFAx9rWUPBqhliyjl938BjcHwhPJdbp+naM1eKOz0AS
ElOZhp3JPb3t+5JQfSbH2ESW0sNNX01iptuJblZ5DeGVQQpuDrFLK+Us3DMOFW7H0sq1JRgO+lrb
twf1XCgLzgMTviRAVk60laf8QgNgmb4/stCp7cERpqm5VaW4aRswDCpbqmk8a/Ix+CsLF8z7zY3w
WYKqpYDWFk5CX5lYBXe/3L4I1KbS/aDGefTA9GPHhEIKEnRFqh74hSaZh2pMvtSrppdev8w9N5jP
0P8sletpCZd5ZIM4KFDQCMTbprBP12ahyYEVwSaHImnewmIltsGQpQMJEwWdvviuqyNQOCtexGkt
bq0ZtC1TraKrKYB4BH0Ljg0PXtn69s9DNKA3xg/xybNe+IvdVIVWFfiV1dE9i1a6Qtktm7rbsvsf
/cFiDaiv2h210IatEHYmrBWtjLBWpZfnvFSL+wvUppEjjr931Pk3uT8SaMphj0waKxFrYt+NLoFN
e5798UpDtOX2N1jWU2D7ebPaiogysaiCm8XfZy13XILkVsJUlc+X6/rXFmq7kyLYEkEycmnTzFL+
OnwnpAwSKSvuwsi1vWfJopWpjRjfIQkZWWy1JmmiTE9yY0fzJR+6h21+rDg8/oYYjGju9HkVekdu
5cAzjTNagOU2zFL2qghf4mUsng+rnTe9t6Si/EdI1aIR2gSTRnZ5vIouz6qGyABEY5d8kooA0xfb
gGE/Wwavo3YkXq9RYZv/tET/Wz7Z2jv9yCymW9CXRPUkuK69J0sh8Hiuf47L8/IQbNtp4dU1S/IF
TzwkIAe0XeQDPxbF48t7BilZy6o4PGcc0PIqJM//eQdzzfdWTz/LBFDJKo7yicujdCo7EDQs+Fw6
9PwlwtXzjUEdRclzhoPx+ni5NZF9Ep1/mqq+g9PgGGb6Xmt6h7fNupSBHP27VWAklHWdmkfE/xZp
Y88nCOn8jhPrJscrK6czXZSudPWWQ4xKKQvsKAeV95+CLjegzB3shgyCQ4cKjEUDmasZYkwxXpul
evKE0C1vPvLYvoEKOFJs/5dQctZXPwerhm8xgLq6pDJlJAS99aRH5L1mWAh2ysnZRHFfSCM30qxt
TOt6y2SMpdOVwa+D0UbP90NRtW7qHTpJISVIZSfIp56esKaahnVgr94zJemxRx2sfZ68KYGX/ByQ
XHtr1CDQHNkwPiNxy8KGgieS+j0MgwaOc1gmj7yKYZZG7TzN9bM0GS47LTSMFdRwM9ZZBXOBvqkh
21iiTXyr4GDodU36eDp7jtm4YO9fyUtQzd9GUNJnjJDHwxTiFrKan1Pv6fr6XHeE1xmaRLEQjnKY
9mZVlUqsBLTyeF7sE3wFhcdtrKZ1knSfgWNIIfq+ederLEnZBTjl+ONCKrS5Dltft2uYnxbr6c9e
dqYG1CHLJtbrjqiXe73QrgUXMXHbdi7ArlTH88gU5B6gjiBJ8oKtSbUiVb/NbpYeNmXqIfHrvQfK
Z2uwig8uNcBxP/d71feoQ95P7konhS9O7pYQTPVQChhbgwy3oLPqMgmf3hjC3mO64XG+a9NVeKsy
T+DtDMpU/wSo5x/KWv4VPqU2Jr30VeVvI6gvp2ehnFzcIz1mvtHEUr11kDOr/kciEXmrLn+dXjqo
shImekWd+1/EJGDr72ZLfeAAVY8OE1hioU/JjB6jX/laJQd2S+0Su5ElMt1yrp2XNQOtJg5iJ7GQ
PqQUzWPW2Td1Wqn5qrotTv9paItcHomjUFFT6nfVNd1fEyJt5ETIDPXRYxdcdIm/RE2DrkeDgt6c
Lzntqd482XyVr9ooMkFshRBCsPgFHAAzr42xDCAi0UTHozeBXGFaMDThN/961w4pGHn1bg1/ap8L
vdPJALPhNDvGo+BzeQyl8lrL6Z61aYdC5zzT5CABsMCZ+5yzoGPXaAIlXFuMht0onCFyWNxEKJXC
0oq5XPOtLvUUoBsz1ZWM3/EcygPRtp1cL8rpQDQYm4XP1o2nYHDmfDoz3eXzSnfJavYP+MSrWYJF
oxs0OSGWb4DXjkiMcz5YHl3WS0wfWjD2mc2sP3k9XPwbx4hljEHMXlxdBee+Kj5VsiTuJlwCr3jJ
qhhjMyi+yH17emC1lxaUCZgffXOuJINv3xad6eKQisHfDd4zzO7rs0kQ8hiN/m/zaRi2ArnI9X3l
T+tWLxA/emsNB+Z58oGAEh+wtxXRbsmah6nn3wvajsxXCMAkm6UaFev5bpx0JTJhgF6x6L0nQ/DP
tBMU2QINmdD2R5lXyFz9l3eFv0Y9+muSn0ssBQVr8JVPwKvkLQXHaQrFeme63jsxEy9A0MhZ7xyQ
gU6nq2cLVMqD0Kss2XrtOjwjycCf3x1f0gozwqiofTACt4reGlXOSF9uhKJx9Jow233zfQEQcwRn
u77WSjOSxz6heKxRUwMp0nZV6HaX2ZTHM47vQkVgrIcD1ernQb7H1nzGrjak6zKcYtYrajPKK1PR
1dz4sfKEAW4IpHah24J3ERArE2c/6AL2KG4I93DVXVk3P+gmV41yHd0q6ID+5P51Qx1vHjtveKyS
nsyABmHfYxGfyEuHt05NBZhNT90VSsiXTEsoAV50CcnscZHVE6XZGGBEY3M0gOp135Vn0c9bXLPk
goHjw8iH+Cg32v+J4yBloJi92tnqiXEtgFPtOirXyZEiHcql9jXXZe51j7NdM/Ud0mvFtIp4OqZA
TdwvQWcV4j0jNh53K2czEUHgJoHNAEtFEg14lRiPk0BY/X0vw+FbU4ymj26OS8KIH4FKo4ai+Eov
+Cfw+m0hPOfyP6WBDpC+ZyzU+Fk+4j+j6o2+O+dB0urY2RUP0P8gICvzGOTpng7swj4rnOGCos8r
mNyVHOwAzzCDmWlr40pqc6muTTOHV+76CsQpB+WRba35TPV8UJgg2iqo2Rh61MnViNb9buQNHGgi
7Awgz6OMopF+iprnmgaPWqkMelXlJvpsoZsOO/rPo8+DcS6h/EaIUUYLxNhRrIaa56NB3jIduQ0n
Ti/78VOj12zN27N6sVxh15bup4xJUS0K4r3ULW60JX/vVReRLqRKJd7Yi4DVTknnVHTgXNT/HVgQ
5zkNg/75UGti6kuQ3VAgSl6zrvK7l9HzIJAqxuasOdT7JrBIsQ+ltUjdg+XRp3Hb0yaeUlE8YMFa
kVzfqV9pj8esIpm6KNuvEn1rL2M0dFTj5uTf0lPb6GrMR4zQEMQINZ4rvldX0RtjWWXses1isPHL
2h4EyCi8uqbwuPzgtFMDu3OdcRtu9ZYh3U2YYCzAPR+3iadB9hQzQmATIF85HPcgYoP+jdAv57un
/6jA8lvLOk2aYbStjGB4mbsmHvrIaFzryFShbNqcLZJuN1e6dKCNthJBcJlLs1Yu+7M/V8vmsH8d
SZRluZfhuQT6t3HuxgFziJP2X5M0V5q79ufTYRSY9l16x0bZd1fPkyUJkEtSZVJjzbRp2keAbmKT
UlKsWXT8d68vaZYsTKRdTAPokBYc9zJ8dQU78METdpA/kbcR75zdJ26D5hmsioqCtGRnfJKKhvIq
Ht59IWM0zJZmcnO8U9uSvBZBK0PHxnmA0U8LxvyF2mwsTRqvGWGjTvDbZbML5ud5XtrEb+/l5zmk
VH0Yb8rTH1JbP8imixAYDo8UN2Gg5fLS0gRN6Hry1/GzN+dijCl4fXbgaDTGHJY5kVXYJ3IjZXkJ
lFokKUeyn5hlih8mYgDzt+z2APBinb67G0inpFgVvweNNcuZ3BsP7N4/Kk0qetw/fIXUQZppOXC4
OYp81w/OZArLsnHCNjYci5uvloBK+ne1WvghvnHBWxnubfyJH4GdANw7GxBvVig08lfMzme7Ci1t
/0qm0939g9qJ0TY2BbGK/aSpvN5LJWlxk0Jzr4DfIgT0Z3JRIWT8vERzn1qDcjW/OqnjX4TKCDna
KcWOsIRkFQPjYU7d7dDBs97X+Cm7Hk5GDvwrmL6tfz1cl6ylkA56hMmBjxLkuULV6lVwomN1LpAV
/h4G15kmr5DoRsX/J/wEfEAvNMpcdugM01HzlfL9f1aObn2mwAacz3CC1i4ORqGCiUVOtiv6Lmjf
ngTKAtm3wUzLp6YYdC3BxX45L2mqgqsnhqFtaJUT5NQPIijgcXl5BQJTE6YCV8Yqp3csm4WstY6B
bZJzJpHu2rQ07RJsbf+PptIqK7LgHUUsSVmmFjEzVdZdISdQjTMWDc5ZjUD78zhE868jEm5ioQTD
ge67BM41Em+/rewtMtresPb4h8eMfXi3UVSdcYlYVmDi6jAxHerIen/7qBNRKuHFQ0JK46TvlxLr
h0CCTLTFuNK2iq7JxzqiFZ/Hxi/c/5o561dd0lf2MSYDWRSOAq9LVAFgjqwh8aSUMye8xY7VYNJk
cT1YqaIutV93D3rhBoA7cw2EpRb5ueK6ggcTB84YW9xjj/pVWU3B33AJkRBzX5wSNy8UfLMC3chT
noG8pUms1I99TwFPAdJ1gsec+heb2zyJkHmu0Nwt/Se0MCIzLep3YOaqhcifpQMb2NChDmp7ykNb
0GaqxnmbiAhq2ka1pVyf2J+1oC/pH9H4Q3f8MFSbeAR594OuXI6q+2q/TkWFVhjo1j7LcGa3AsDv
yku1NcTDLpngcxOl3FItOhG6Dkj61ase02TEzy+16EPmTJzneU1mGqEVtmAdEmGlvD9a3Ma5+cOT
f6Ua702Hw4JozqnczLr/oT0oCWBLhocAFOdoKW1nSvW5T15t19PRVx8xVlf3w61c5Am3VlCzVB7H
m3wHRSykxu1Xrwwe15fWqVR8w1yocBMcaBHSqadcl3ehh1XTWlRJNkJc6HTggZNEdtqNxZH+idGA
4Qer5xsWrQJTPoG6YfOlHUBkGhieFXMMT7m5nNt9Q5eqVZRFU5SNMzmXemrmlLyuxPm5SrOt8lWD
DMq7z0nTFOSlZQdrQQx2w7uzkQLJCdEDanjEbVkGxCMj7k+3w/DBmYjGFlyoQlHs9uiAlxxL5q4S
QC00WjTEPftk9f3uHN8YXIGZXy4ODLbEJfRDUoeMF2dTxEg0E/GJn4LvATssZIT3DBCADo4MIUuv
mY7OaVpOxezEQeYSa9SdT/Z4BfgDasrGiFvnsUshCwv6u7f3ylM2cKgc0yjVV9lYRAJWHZkbjY1J
rZR63vKeki6Vvunu1to3vMqOXlmy2ReBFYwjrt0wpUXYTw1AOo/64YWXnR3V+EOwAopKcJYmsaAD
JSoWT/gSgTO7jK0ePbpfOTEOmwSf7+KEf0+cTgPbvrsgyRRdh3qXXMxfEr5P+mgB7XbGzcXm6Y2H
/R3kZJyxGcGXCQGW7D9j++VEDUMvQHY9q7Wvze7FQa4TqUdgpL43Y7q7niTjesNKGHvlGy3lb5GU
CaoKlv2xCxUdatS6ITRk81haCF4QIw8TaXmA5/MpyhvaS294TgF+JmkOos8Zw5DT/I8Cg/sbPq0b
QILZIll2KhFBtju73xL875OCltJxK+JSKX08NkyYhL2pC7qL1ZnHS9ATGUsAS63CXdmX2dkQ1wFP
6dX6+NfY51WzmD5S+soKKKeBz/tV6MCtdYs1ICO2jz3W32adtBNEsEj931SKnkYK5Y8R8s+G7Eaz
N+3uClZsJ9YB+qZkZdnLAUree7LIji2WpCQxZAff6y3B2ZQx5dxiv5VEttg/TGr+GCXA9JGLsP54
qxeZ2IU1oee9cjJxZDC1pYZbsauvYuUmiItvu5U1ZnYvl43G6z4rBWA7WXLbyiV1h/PSL3hu8n2U
FbHT/acer61oym52FWfLPXOoBTNvhcNuWj6RA7RdK8liaCga2+dvVGvfdZkJN3A5yX4ESw09XUEW
bcmhj652lWB/LQNBV24c4edcMLAFKgv0uW2CtAL9SI5dg1WWH89pa/+wofDRhpzS9HeQ/dq+XJuN
AmC2y4o525p9m7PbfdAWLxY4HLDYVNnnCky/H0phH9xZ13+uIyiGvA4AQHwCUyFdGTSy40nrVWNl
JqRjAkx7mszlE/PkvSMUdzoR7AnsYnVgs3ceQncckYelB9qmt7dlxob1NR6sEcv4QvtlfgklUCSd
adfMauDErJT4y/+BrWRIfyBk1rjT4PiX0UFlYBRvY4+n3PWjSBZ5xbqZiA2TYXTVuCyMNb78WQA+
1i6FC7429Wqnw2tITAj4Ju7ctqWIgykzwgnDEYHnmm1njnTM0rzP0Jthy0N94kyTtF2wxy16S6Dr
TVPXhsfjswA7Lk93Bn4Yo2hp6HQhlaRN6ckq80Cjoeq5eNs2gjmA6rpRk5KypxZBvmIUxu8qbk3Y
oKqoSfC/xlKSEfZPDcyST7AhSmKuIZGnfzO0Eb7HZZ+pOfHtnmRkYNIfNhqzW9x8NW7Tnc4No+PE
bV+w7iPnNA5uy7W2yFmyLB71QwzAGIOG6BUIhSmIWD1H5PSjCPcma+Whexxw4oWeEKs0YpaPNeNV
iUm7peNVw1gsgRlcgOF/YtpcOolMdnKxihH6UTkVhl1dtg6WE+jd3bhhpCJDSZCJhF7XcpQOstZa
prLd3KnJTMcVIvNzCg3Sfjaev0BTstmFpUJ/ue+JrKp95Gzizgxw9DuP7EJgU+L7J1bTBOOii1Jd
cjmRuwEmW+z8MR7viwaZxTedThSylqsGdspKpnCU5/el4cYi1W/mNaV0UQ0V+sbAn35u6hqJOhga
KI+Pq638ki6XzyKrjb3ZIAs8Z7cKufCF7UeQQVZvEat7Le0mEC9YyvlyKMBYbALAMyZAeBMQLBo3
DqQ9hmX4tCcIucBsD5ex294Ia1TKNHE9B3i2cpsthi5Wxu/7dPQWuTIa4fiI8cD+saGqlLj8V7o7
PQ7EtHF4kJqm+ndx8MLIRktzYYe6T267yQjTT0+aUEP3CnKq12CReWzqEPx7r6+IfTBryfZ8h6FV
WaHhzmmKNK9aj36TEzE0AXJ5MP/7+8NGHvvvts7oaiBSwZ50Sw0LMhS9G7r4X1HelkXWlZdzB8vc
v0UETR3fH+QMmA72rO8pvwlVZEy7bxL6z1FwIoUV+K1ALENxVqcCsklYhxNaFDDvxga8KHzrBVO8
X++kRsDjgpTNRClb5H9o74gd5VMgfkq0QN/vDMxGDLneBcmXE/cEUm6N7GRGjOIVPt2F5YRWUsN5
1jk8TFvzjqugHQZ9LxKVv99WRT/5ama9MW2hwjYLa/utjiZ96JzikBNJWq4eBSTLFI1tkM1AkYus
+NQHOOB7aGv08NNMGluECSMviN9byFE9bKcvlq83cMRDIMRgXSTlGJPl6YryvHyEtwVU4tMXUSiP
VD9pvQA/uLDsmOMDVg6vvmiIGsvF5yb4qeWKBHuVEi0J8BOA7LcreuCqfvmp9Mtt9Dyw1M/ntR9S
0Q0q21Mt+EiDzrCNA5l7yrVspd5qIvmhTUN29UYs+8epKogu3JMOKxqpC+gUBSHcxPzEKDoHwWK8
9qZO4y6Dd61tDOdwlDOFKYSfRyKk2C6IuAjqO4nKUrr4XWv3A3RBTEffuqH8PlX8ZQW6t1tYV07Y
8iFoLHeJP/45/HAHn43YXBNqGFExoRosmXNCOFPs8N730yDNy52pJ45Xi0lcSqyGFTDyVHttGP5u
VW93ZjT6n7q98ObEZTXSW+eesdM9l/EIR8cPDs74foMNVHZ1Fb7xdiuV25bEIY8+g9uBbo3SeF35
mX9+wpz6DIfL8NTQ75K8hsw6QtzFuQhWcgD9gL7zlcvkuNcQetpH3p1cnpeExwu9iYpXBJBTdweR
P+ozPB70AJ96RM1V461/+uV5hP152kQV8wbj4/iS6eW/TLmImgvNL6B7XFXEDaTpKRiLYt3PXGmw
6scFUIGN/0wgXcGNk21yt456NP7wYPI5XsTiji3ndsw0LmNTUONlqeD0oeDiVp+1MG8ukJxgrd6u
0O94MfkIPT+j2gIeq8y4wu+87GBPEAP2qUjLG8nHR7RdGGp5Edz6TKtexAO4fCzv5Mxu0w0wq2HF
3b6tIeryFjezMb+LAEyDIfr+NDFVeyOnAlPWE1SBT1gY9FqLxI34ctgjuZfMGjMTUvVQNz8ddNEM
tcJm/6E7+hUcTkxnQ28M6l3EoFzTI4MzOJTQqbza/kZdz/yo+zG2zoiK32GXrmDtF5j4C2n4hj4S
rBdoX38tIKKEs797PdZWAAkDbNIUcrG6z78cztB9rDptFSZ3UoL9NrvYTVd9FeZhoj/6XRNaH0ml
PBk/1+u7D3FsVTeSbX3v2rrme/5tA68AyTJ/1v47Gg6Qb4aHD7ClaI4iXVn0VeELCWEEWs6G958h
lnArkRvotrF4/D40C1Lbl3EdR2wwmBKD9N2GQ2KQ8B0hJpPzF4TxUbTQT7agaYm8aJkKR5Y97aAu
NdtNjgfyAeLCq2O28xXoRL3IFpaJK6d5+5/KGmbkJHn4brC0PGlvbm745QrVTVKeaIlHmySYI/wS
AqP0GiH2sql7mpEICvCldSWDZDdGVzAMnq7u6mQ3PSwRGWaLbUv9cCEcMgyHvSmbRhD3xtVRece+
0SjSt+U+HXVHQPa3lOAA6xXstclmdM0TpRBd6syvsUdmDt82G1hkUVo+baZ1xQPVwzYN7jSP8ac+
iI8PP56ERQOYsHkbokOt+Vl+W8gshl7uMj8J0TftQ3KMO1+/ehgnGpPl8Rez7u+UXSV5AJ+wsE1D
9tojMon6vGbMK0ra5ZEHGWpV880K8fs+udBaHPKrrIGqKcihFAAecR4hGd5UG5beJdQL3Ob6g6Gt
7SN3f0bxN8loRIu6UwKXq+yKQAgZ9DoB14dl4BnhjMpTRGbnYXU/zuttD70B+CCU9Vanw1KzNiUA
dN9MCTNf+Z/RcCVDGDe9NL0u6FfluV6a2r/OZF/USR1Cun88T5w28dudX+8Gc8c4sc0WD6NnHO/h
0Vh9jQNJQ6a179rK9aErcUkBx6ob7MramT22Od/jvw2By/EC7XL3yWw4cDMVN99YSivXt7HkrcYf
gqcQ6iBBXOn0AEPW7JSi5vPWSbbo/LAhyJH0lQrfHTsecOR1ABXS6Wq5zHlHw4PJYAKnUqoXAhX2
8jI58B+4LC0jAXj6D/3vyPDKmHutDi1pndWwzAejj0XdDiaRHbOR6VjqpypbKk7dO8JciK8uCLl6
lrFmYerSmCBJTlHo8teKChNhWYEqfVT+Un0g4v+vIrfzoXPqBUGv1ShQVwP71kuVlbqDhd2RTCbN
Su0QmO9UqHTuAQYe/7H895ZU1lKLOquD4Y1En5m3w37sbg3ha0AAeA7iWRrdwRbKBJG/4m+ryBxl
2n5MgL0vL5T+XrG54hP9BjUlcM1/0eh7CtPamW5sxPa2hJANfo0MVvhJ9rLszwNHmNsH6gLUpIm8
/SboLk5JbRvIB4icvEUBrPH1XQt410vDqZzWP69tU21O0g774GaCKpZmBurvG0dCCf3yAvCFSWu3
m65TK+5fdWfWow7Mvmj5b4PyliZnHY3EJw5YcvBLCuELDTyqEObk70NT1LOMcl33dJIf93HQG62E
T21Cbv/VMjFdEagRrNMuvsIWX3PpuLc3JaC/xO8FW75CLN84+vGJzhS1HfN1pqzZG88OOj/3uKOt
XKEgxneRt1o7NSIJw/37Z9Cc5N404MW/lGqB2WJdDHSq8VA5S4pXMy9pM5/Wr9X/6BIBUQU5jg2b
flee1I5isqXywo7vpEg9r94lySuTW4ZZP/BQpLIPhZTw2T+W5kQsOsKp7/lIToYUydwzkucrh7qf
a74qkQKEiZEGJ9UgMh3Xgh1ieN0i42SifoUEj2k2ocVSUsJazQOMk/GQZs8RS+yuMxM3fPdLsMir
TvdpJz3W8MbPuijEtWofPKBTFoXPp4erEbROdTd8yWt9+Ql4Q8f71EBVrUxAi2ONtZjcgf26UmXf
DE5SroxaZ6bLCDsDrX5KHbnE3IsGXXx5vH+jrZmAd1mHhUurqluMH1rPLYNLL1WKI5upYsdtsK8I
gOJSmNuNQAcZz2NPGY9DTOjxHkllc/TMidthuPVvBpI5e89Dm5liz/ZFuZzpih0mOqj9yUERbNBx
lQkVSJ6Em5lwKvBASfdoxZZtwHgsjjgSD1IxMtKGTRzEHk19q9S4bHr0s7sgFoekgXCrHYztiqmo
tkMp7f0i/eJd1bOh0sPRnjQ5qWhZFCPfFegKVyuLjwejk1wP1A3swATI1xw7lzqwULXDkQ+2r7Qf
Em2tgiXqhxjGehVm9yQyWPO6H46PunRIvazWPy39pqgrFQtvYwO02t/EP+tXVaMwqdBvxPctd7xN
D2RPdXFxUCy7DxdE4jV0g5Ht226c2gqnd9W1FFDTKv4tLSyVI6c0kWkXw1Rm733r99q/+OBUDMiL
1GG1LL2ThVy8v8TFs+LFmRJbej4P0rqR3RjnKesRhpbyQyyVYa1pjj5FBa+bopkRN5MAIt5yHz4K
0pia60o7oinIi8l3AV59fu4BWf8zt6uqEy6Fz32hSj1fhcJ9Cxcr9KAhyzJOYvq/3AIxSJtJTUT1
4uOQzZvCnX5MWmY6nRcMIAtYSM6HpdOX/72GdQ8iU5DlXSoUfISgfcD4Aeiu55Sm4EhWptSeKXXF
PuB0dKFi9fHgQZu8N6Yq9yKeJoUKIENjGzUyVEYlZm9GK9lNqqUenT1Ma5pblC+be+dYEp5AGhLB
UTtWqcaNWHqCFrD8Cf9WgcQuZv8ccy71BS65oAtlYvxC7ZR5j3EqAC7B6dfpj8tHXoIyR0hlClS2
n3oinYHLuOzL/Q7REaUpOerSLydH2SJXXC161/BFmwjaZvrqqVmBL3Ru5lGb7Fs+ZRt2chu9aqBn
Q4cPzoHe7TqJTcL2RdRcDyRuBl8YE/v4JcXqr7TXuouPUFaAI8N/stwdIoxeY7/66qBYsIpWEXjV
t/5fJlonyYY0Do8+Ifava9K3z+DO7uViIURe2sZwO4wFWKaVnDgeyV0XfMzmGcJm+7UxM3eSfG+j
dE1A2LBWf9VaQSEWXg7n/1RB1O43PW0Po7M84ok0mXqqM5r/RtdMfnGWwEPo3vWPZLwIhL3Lsn+I
IpjMDAuuyzzLYeIBdqOWIA/oz76g019kEtMSwW44ZyN8FbsDS9F8UsPjcbb2e1G1fFZ9TbxauRNK
W2DLHxVKVOivNx2GutU//vZgfxKKSujO0EnaJI+v2GUY/actISP4l8ultscGJ87FgvN8DFWKljxM
pwRKO+FK5n4papW/BAK9drUJqMjyvwX32JYewK3QQBAdQnY/jp273LN+EnFKb1O754aS0MB8xPYp
nT4A6fIcn0bmv5NDq7clbxzhzS9JwEkDx/Cwyvp0cLdV77HjjVOVAIvECX8zyQE+8xwYWrzN2qw9
VJ0FWXQyJdbdjA1Vse4nITI5B2ZlIDMprHYX43YX3IX2410cKwzbTVY+ee2ArzUZ/jIRw8r6460Y
HELdU5vpgqU152wLJ61CUi1etHAS1lfuPraRnq4TpXICCHEb85mIqnGDJMZpy0xQnM8kagDg0KcL
GUOjOdIePRLHR+jw/zqKs5giMKpV7Vs36yyP+ixXfiO1ZQjQ4yv8IFj4nBN/+MapeyUxfKpOdi6F
MJ1HspoLEb90JhRMvIfpZ1fB13t69FCXHIOqQBQlFKjEE+j2cCmJ8jLubC9E8HmIfoUhHxuPQM78
0WAN8xZh0AbJU+pxb21+PgpIvOfJNT58d/Qf1nty61FHj+KOI183Tr057KEKO+hhZnmmbxLOmFcB
Hp878tUQrJ6/QSv6RQHDI+WG6hRfeooOp6s089iGLSJ6F7FYgjSWU+3hcmj0kqp/FfiMWI9HuC7h
bDeYSKs8FhIT/3JI39XdmtwrQcoyK974z1xV3cllUzHM8tAt+K9TBL9wQrTtAO8DG+jYEVQSn62B
0sxnPUVfVL9GcSVT1T/d5jbJh3XbotY5H4OZCVras6S9ba9zLb34BLtcIzaDP+OlgYBdbG4aK3Hl
s4EYxuM3hfJPDjRiXtHxp1gtqtnHYvUjN1NIsclcuPtEobwvtYTWvPLhFhYb1RhQNEHR6f9qlVAK
sO22q6vHf1BLshKdkRvX1ePUfALJ+Y+5AcV5PKpxDt/+HBYZLOh5mWL8hMB+7OJbAqVFGsv5TpmH
YjM/dPlcsJOtOLDO0Ma+2xjox4TB80SHm1BHvXcjyi3LpvXWWwmejg8x1Lwt1hzNGvEsiuFD68RZ
9a8lWcOz3ldodGs/KGtLLpP8Stvq7q+CbpOiiSXOXtbd4N5SrjOvVT/F96MMPOfMXyB0tN48X91I
JuCy7PL1zfsKTvOT9OYE0PW9N3igGtunNtO1hyQ9uVEm3GAmldFvNZhSNLT0LIItApP7igBgKc3W
sZQc0EHp1fA4oNAziRHAW7SjwW3EzlseW1gghg5AiT6FDfI7fI7EXBBN+knYr5x8FBhjrNurOZoZ
vBn+TVv0oJJ7IN/0hfqAzOJBbnkEGWjAKpxfFsiAl0442oSgBTfil61NKeI54ihep962bnTKS6+I
HO65Bj+wOTGw4oCOxeMyekTh06GGdWKrT4KCI7XzNJAhBXfRNHfMaZ3PUzDhSauIgxOjlT0meIz6
us4H03gAeSLJ1QL4cyGY3PUl50QrdwnKsCuKEPa+k8hAyhXZV+WB2M+1iq7Bx6Mi6jmrb2Mwgjha
u1BPnuM4sl0fa7MgZSK3idKkQjaYkK7G4EVInnFI9mSfD1rWKM+FZ007dz0q7+kPLQ9jtKUPvJbW
8aJ9BXgCP5k9ozFh3scP+FyJuQBcYPWtlBfZ/gPbFQHx8OS/58/x63aInrWizQgp6RSPKgEigf7h
BBmIJxhIDgCR1mpnHplhU/tybYj5ppNL60PpDaNEo593KflnMXeThmDQNq7k+mWzl3AWMj+MqoXs
rbOK+usOSBKaiAz+TJV1ujYuNpuGl6NnqU4c8aT85lXrgSHbVkZHQe5LQ5lDrqDD9srFcxFe4af7
b+7yPFB9Cu+8d4L+pS6HTTyFpXAm/+qCA5nOu2nYcXyAleirB0Dv6+Zyrxa65dz8b1MsufxY/6kn
X3QNcJKtN6HFdPqu8IYZRjqD0i74v3L/FUoRu8L1F1ZYxGIJemmlbcJEdWLEtXp67/nPBHMMPZX/
nYmixuRrIeaC9byupQwDcZdgYBEaBur0Z9R+Esbb/L/fluCOzWEGIJ5mkq4DNoQ66etZC/9KjCfA
pxw/kW39TJ9doiXEdVxyPyCAG2iFzSUmaUqdGUJtSfK4HoMAHWQHIE8JbCG1e7kSar7K3i8i0H7G
8Ucu9kaoYdMofxiqcJyN5D1bT+X0jhDW0WhBuUln6bQjfgYTnr8EBvuGpEKp+qlvYuWypTi8CdbR
vAAkGhma74E57/uLFtX6jLLAdzmo0QbhFcn7Xefo3kT8LpnNkdQ9tm+ehs2AaFCPUKUgvpizIuQZ
c6kgjpBf6+gK2UdU6Ys3245j0Apzp8SCkBbEvy+4sgDl/PlDThQHBXKOqsxxu9k7Gx5q7UdiA5Yg
J3r8HJdEd3CPZckEFIhnxCFKOkQImv/3UQ0Mn6DjtHrHMs2PdMU34j6E8wdn/roZdI5PASMDS6Sc
zE77aJsvT01hserkyVZwvCEGelVBJ3iDV86kg/N5zRsp24NHHZRumn2SD6YWXAcRZIY7r7Ga9nnL
V5VMr7KRfJQ7NVU9t65qQwO9TihG4Eot1+xtwZ+VmKK3F4ZN8GiLN+S0pFS0SGKdGBI8nQlwy6NB
qtxQ7nj1CoI3rC1UPnXPU+el8KxHGfMCJihOwMKA/d2Sq0qwu2ws3A6nWmuk/kayQh0fyoRyjQrE
By9o6zsLbVZJC8bJFFbDTdOqx9NBCa8EajQ0131SNhdd4fkJL4QIf/O1hsWRHqVNJn+jRToID+uD
vOfrH0mc9X/Qmi/zcGUuniT4++eWUxfayiR08O0kmsi3ITkGonk+DxK1YLFtGpWPakNaDXjulXM3
ET3RnYiCd2EJ1CkuI8t0Pg4xTl+zqmCDGm8WC/V9yR5HA9iM/jYjnbfNOwdDPmvYYHY2KuJsSMYv
e4DLemux9c47ljvguiQWrffx6ENgapw5zjstX0n/D8xxXM3IMgw1vW9uVY9UWJrbTZlVCjckCnCc
CJSBrpRW3TEaTRLC0eBqDCHJ9dMMpRB/se81V9A5c/FMXlYhsyFQzF//1GLCIk3QNpEn4uxeOpsN
gnw29OTJfwufm12I2jUYMSzEEEL+J0ZgDrYGtn/9HM5PkW8wUFQ94CyG9aKBrZl818mWi3JhJgi1
DMwo8zJ4i0/IMxSLZdqUXILigE8vqDV/y4p64UEjfBMjXnAkKu6VoJ0UWJFWiNSWVsTb3TAzqy/E
Yao5rauU5i7Nwtgd1Poyph1b/s+c4OEvZs7F7xO4vvcgMTAXERBB2d8P8jHT6/kfwh3zfMQZu7GK
2QE3ifVBanHyqdVdS+tpyToBoE28SJ+pG7h2+WyuCUidusflJIIaScBrpkmkaDBkXbSRUUrANeML
tQddzZCfqQZjlBhLoKVpaXIr1Il3Hn2LoWP5Msa0mjRWnd/I4jLxqD8LsIQPyF1P2qM1+i3iX9rG
/OJT/lV2ROFvuLd2oTDDNZ2qYGo7Pi5VoYi+TcyWrIdWBZqNsGpdehG5TgXmx94AVS4tos0LCbjj
1WxeT9SRM725AQRiW0Ahd93GGv6xnjAIx6nC34n5/lmu+Mz7zdC5aed2wE7VozL+v3tIU7PgCd9X
IfiGDIzFyuE8PuVIORhPXEwWwY+pFrOfifUrHODi7jGWwRYzNQ/kSKehe7JxZOxzh1WE7HLJdJiW
2GsLhL/l7UP7v3o/ujBKujnjwqdWAl9u47zATHf7og9mGVdIwQmVmZnLb2byQ6zrvgeUyjjCLDIJ
jXwFZxjt3EIBX7d413rggu5mQb4ePwnY1V/Z24rMA0JMudberpAC95wNac+ZmS5VZzZNGu6EISk8
gcMMUp7l7Rqi1rTGwJ0X5ACPUqrIEQFkWuaYnp0LdBnfqB5yIAV4WO0dg2lzz465nwNXoZZDw41Q
DRs0kMtvviM4JASVx8zkO3f20W6DWW8EdiEmRmsXGvb7Y6LLs2t8fytgoQhfEwu27OLveX/CMVyi
Yz4xPwNBltLI+qv7VcwpmoxhctTq0GOxgq0ASeb3NOQPbLwNpfjrDcT60VtdfZr+2ehYdyMhETmf
wa6gN3frW/iPM7rLbxK/82HM0A2cSB2M72MeK2hW40RgcdoCvZHSHCZLqtSyYTT5L3Yk6GnE8VFV
Mf3tYGDqkiFujE5UH7vtKSvCBSO5OP/+c6EyVFUOxjS0x1V//HzpeG+3+YkXHblEvyVx32zvbtD/
UwMBQk36Ar/o/6GDGMUDp3aCmi9eiunYDyKDx447MAxoVDkdjA/lbEUGENfTUwqtHdvEbpOKkRSi
qxuWw3+NyRAFZH9rLYEKaQhUbZC5HbcjRSmGBv9dt4zOHKqO9MoZetVFYwnXGHxt0uyiLFPBdZAw
MoiBWvBVjMmKItecv3rZQi+80nVM9XAQRHXlKmCIDp3zJZ7g3V2w0/nZO/+gMLMDuQNku/q2rcBQ
6N4lrYp9078qFgfrsMBABt0bmrHpgH1Ox2AzRzpVKVABPXEgRVJ7RcrKtJsmklcpcqyGcyKdJxp4
Ju0XbXq+S9GlnXNz9ehSBRjSDW+QkKRXS51Jz7Rm5dc9uOISWlGZPg8QOi32qKFUBoPxsPIf1p0r
0ZxWS6e9G5XmXz7wDQtxys7UlHrr68LiCZewdoaExQfDHjkV37kYkD+RSOkt6i48Qhza1ZRk9HgA
B8KGIK5pZeYupys/7aMwJX9dBDo9wIzKlBOARSrQWYlBW9vMHzU1ZWsyLa+P+JD+YvCl7VWZ3Wv5
vFJEkTonCL21uRPZLJ04Tq/hnvKTzaS5g2/UcgCfCBpj2R3gocDUau3hRN7B0duADbymf5YVdQB8
RVKtMysrvDM81kcIInkZ+IU/8OwLNBGbB9L1avi/pnc2Eesmy8tOinGZt8FYGe1g4HDlhcyXfrFW
jF/56AX4yKVJ6FazwV5jv+7btaN3xufctz3KnepybDVrhDlLlwlonCEuP3g/Uc9qKhaF4iVP2eL4
Pbro43YTzX7ycdXFyikejL+9sWNaXatAjgVHdYQ7sJ4y85YZ38cHLienu4fnvXby+KUM+LWlB8Ww
7FUlOmrKa330qmo5KkpbCmXqwBiKgzWIzMSPhc7Bwd3I4mEOwIexFYFWGQu3/LsrpBDwXnCFLDVE
XAialq41OSChJA3pfEN3ieZI96W7/9Mj26Ss4cCi8pv4ewUVPsTMxZZ/r1g5Ue/U/izzvTFNlGsm
al8xcMWqoEQVvznoKfz8a6Vzki7qhsR5+iZDGoBdtSlFh+CV+gr4WBISpACGZjMC+6OIXClVdIEL
qlKD/6BsiBZWa1UiGkrWSUW7QuLo8b6XO+26CBWmRkeUDNONMimvjo0ExTqFnb/qkodtiWv2V8OX
xNm3ZSB22obSFJWGnybwlUHhEZCelBjWkSLeeBBbv96WOsqORplRNRGa/RPPcoLyL3IPxXxlS99K
NjdyijY2EUGzXZh+7f9gjoN7TPEbz9ZgSVBFZUd3RDSq552zPxiDBs57SHAz/jsC/8rbKGewzJfq
nzc/YAMedxbrCNcGX5mRY5jqAZ11izpQnyIlR5WGOxvIVBPUQdTCy5DmID7N4r2lTjqg0UbWzY3k
6/9oOW/qGl68NFsLlMHuE7uPFHYLD17ux8StdHRkAciUu3lQgs6Feykfs0+exbv0mUQORajVLtAE
Sjh9lf0YSUtNgwXyRFMZWyVBf3u7ehZnNuNFff02izsAFvIQ4ihGQ0k0xQhZDJnLZgctN18c1puT
Al+R5zAMsEQ0v/yK5zDLEnCdFmrjA8VbMY2tEbW2REIU3RY3xwLkcdhtzbuG03s1osLGjp5EO0IW
MjnrJ8xJJ9P2wJJZ2tYvw3PPaiQ3MYSocAIpCDYTKdHOA+FhCpogRUt5s2dASlB6ekrTxojKEWmy
NuQzyVRyD1eRSo8UOKZ6CTMPOB64qUN+z0bUeZlJH/Aw+f+D5cm0oiiDWmo2++3ri6h75eXmN3R/
h7QG3h+fI2zs2N64ViZtvcLYDK30V8EAYxFJTXfQwLqA90rj9llBSCmTEgXi9m947jkOE9d8U5tu
kHD4fCsxc69Zs5tptiH5eAUAAs2HL7h8My+uFWJ7vYV2wW+1aBBHvfszAL2XjEo1CLMd83Enbtqm
uNsUgGs9nISD/zU7/D20d40AYDM0yC7z0905sgKTfI84OZyAfLI/A71yvB+pRX+UchSVCLbwg0h+
F14X/jAoXmfS9fjW3CRov4LUfN94gp3O1eNMwWJAxiR93DxQHW34Wg8Ue3QALxjf9FY9oNPGX0Vt
COhSligmzf12KX+43HcnelUKem8XGjdWVRlPGIDjXd0aDHTE6BqzbZSsx8rpwzvGe9YY1M1Enidw
lGfxmT2L2wIZaOSYdzwN4Gk2NG3qIEJrzQ2QAfEStpQPqw5prdzT7QpmQ/MkKRD1HjWVGA2EuJXk
T1Brkr8Go+18lAY2B3K36oTWq1uDrCSlhJGRbWqtonNRIaDuDGYuhXdCezRpxVqPI5NhLf4Y67bB
4liWQ5TQFAZugEKtXNNuMn3QDPl1qpRcJURbzzOjlVeHCIHxA8Rj23IN/G6lu1hglzSCe1tlAYk5
7aVRTXUNGFedtbP48tXIRxogbSiYgsYZ9RtSrfFNga9bL9cR0QT1xCZvDbaoz2NVB3ToQY1kwuHO
w4+qYH/J4dzU6hXnYueCHM0rXhEp+zFV4FjqhrOQxTxCUKfl8vOvZY/MkksNxg/zutY3kEneLYu9
Jw0Xu0rZ/p5Ei8ZTkkjNcYs+3f7auvp+sPkebfFAzd5rPMgEaKgEEAc1iN6J2LS3A1Xst24nmBaU
o0LOBkxSaEzDaj9gVo2rcz9GrMqM8Dauy0jq5PjmHqZiYO5781e7MVJ64cqMwWBWpCr4I7/XyIN8
lS0FfIeQJW87YaRMGKd+8IoIqamkgNxvtnU8UJaF6gaxQT5KC+DKNyVa4VkrSIc/HkVIBDPgxcAi
dTA05hqLbPVur3fc+9fYp1B+Owo8UJC/HjLfZApxIOlcQdYXJIp7d4Y2WvWAp6/5zGdGugb8aKmN
3WR2O9YhyHhNJTCL86eL87CkxyS2aWWlW04r55v+ZdiTLwBb/D8vBVJy0jSwiSgYwdvvY70b9xZ3
IQQZGodmfhNlPdZcHtZtrnq3rDMa+TtKDvkFmrTHmZA07+E+VwcanHQputFDvilRaMB4BSV66Ly3
DAxCYOwSRVyAQM+sLjPW0EnOuY9wjtaOsep0zyGX0EaPslcw3GFdE4hAbu7appcnb2pcG8C7DJzP
0ypO5V6FUiFvAgwmwt5yQpwF7UBxnUScbzuQXk3pY4kbvbWOgtJjwxdF4JqMg7ECSn8cVuHu820E
TeJF6et7rw7VYiwq/RkwcfEl73sASoMS4yfB4ycIsaAlIF303GEBtdSYyIak2JyaGvNhyGFhuE24
GG8/xGn4sdqWrS7rGWjRZuOYDYwol7mrPdIAKM2DJ3pRxQWfJDn+9e0jyUczD7nA3FRIonIL5h0L
pcdtoYeCOwOvl8l2THUfK2tz6GUdupUZx6UWV49j74o/V3B/IVe6g5Q1L0CdD5yOCLqJR68e7xbP
D/94ZVfTh2IiAZSzcwAxSUDh61W8VYBjgWWIEP+uoSGlnlKBPIugsbX1xAY8vdgBVzRzvVpy/6Q4
saEGbi9TzyC8jet4/2n6klutPxeDfyDbtyo243Rf3Gx/dIdeFKts8DVh8eH+XG2VDwL+TwYVx/Db
7tNoMBhSqOdcP3joRq8NFhCJf3m3X//M1gbxwAJ0bxWjvKC6PHGgTRCeOSkgqgGPyvWE5AyYtLy9
p7UKLgHAqtIAdDN2VuA0ySp5JMDvvtIpKPUbUyeKUdsd/Uu49WV7RAnjrGSzElzoF0yhcBdqI0xJ
z74V1WsaoXkdv0/xphDk1f/jqk9FuVgOrqJrSIjH0RXno9znySdCW9i9sSRUfuF20/1tx7pRuFQ+
PJbzesXRSFPthEWGruS+JartkxaeDfbpL/sEatHeMeVNQeykWulLIc+FQ9dmPuaZaYdrnWqrlDx/
I7JlDjXCcnRU9sznPWlVqcYAmG8NQwNA5a7SieOarwgCTtOoWtIKo3+4petBgW6lSMfxnQ/Y89uH
HKVZggotmHCKNmrEZT85f5RPeG2OB2CU9JStN2J9ugvTKPimtQG3aO4KrV5TCZlKu7SRIi2b5tgM
EvEBuHrlnGXlqnecGPupYf28+eKLlbkm9bOx11nvGuDnDnoCzPz9E2ePvEwsprq+f860rcGHtmK6
f9ebWYUuKhoV+POvq+ao4CBDc/v7Jdv6ESjFiOahefXmNFaZdweTefWp/Rfn36AuUiAYX2HoHYWf
ouj19DfstmIWMIk/ZQMOdFXkhZ71ItG3aqmeWrNkbifvTalWfhVV5RWTh5hbb8vZm3w57zpHv4SE
wKnkeKsif5VqZqM1Xrj+JA1dqCoTQh4xSEzMvC9OkxSo5wQnexGIRdTXXLEvsf6Y5yyHEKN6QBFh
ayzV/a95pXhzM+GRH8JxCWqFsz0mbj6kP4TNgaUZDAI4Dx708nHbnVVrbTeMD2C4FaziqI3YgDpM
K82Jg/a8+re2JWWG8QjQFqWdwxhBocCaL5vxgAcIfnGA5mMikELf/QUtZgseuecPrHT8VtfXjzD0
jRda0ykncBrthJ6xGBfTKgU3s73LEXiFLm3dLdoISB+UFE1GNd2x3l/b0GMxwjABjFQUFbXBtlWX
Rno2F9mSYSK/tcBRNhQ7gTEV+XoYmup68Awfdod9tm1gUNnlfiWeZkyOoBYBSCxx0CNcql5xNEMR
cfa0Q3SProuoSnvkSfiLnUsaw34/rFxvgbo0EYxy5EWG5ygvrx6yiYDY7p/m4hJ+42ZSfof0an0K
vye3H+SuOySSwf3pc7CI+6NuAHxcBsX1n19zteZCe4T1F/E4yu1Ik8NCg1qOYbNcbrFPS/clRdnr
ullSIkJt+dCI701FbhxqhWNvBiEIMlRSWWzR/Bu5C14wLAVJ1C6y7gxd0g9QhI4dhO7O9WNHV2vP
1wSv6EdCDsVjQsoKIxSsC2r6I91mvwS9f2zmiMALfLlTjEA/8zuFwZvSwaBTRugV8yV0fjudBnhL
rDPMmxciaLSIOQEDtnzQWCOI3nOj575UOx4iOEPB9SL5PwqrWzsFk67Fj4c4wAxiZpodOUHhFIXR
WLPmZ4Nfr7M7bVhLzF2vD+VSwvNhgtY87zxnMJs6UWs2I7OKFLF36PcMGB/VAIBz+FfrWJB33QRX
l1y7sSUSlu5ehYty8hjfRRPkcYU+gi+0cC3OfloxJHYQa5TDVsQn/39Qe/RI7F/Hxn/jzUMywJ3x
qEY9CGoA0y2kHqa1xTK0hIMHpuJ1fnCNT31DT4OrTvdtCuQ+TFnVkBUf/9FZmafkU+pf/GeULhm5
KcFK2djI4kYnF6/QgU1SK2dKGpx5Y83MnGa1Lo0I7Di/YlMnNnoi2MBjaWxDrR2ZjE36dHqqE1cn
qMgUdeAp7fIgKHAxMKNRdjh4he6H3qLU7OJqtgDswl6ZLDFRa73eoagVQiPXHClI7OJvW5XxxuYh
XKciR29DBQjjiI0sK8JlKwRCHbg0+SaaJtr/t01FZTSncdT/8eLJyj5VkIEYXJ9eG+X3IkXIZ0Vv
sN/co5FaMkPoysEVm3EdmdafjcghzPLRiglvjUX2hE9ucCLsoQUKq2s8dPxxKvyGWDGuQ6+EYr1g
KWQTzO8Ll7sO0iee7Pl6GfmnuD2lHRsSKn0LBfeW2DBB+5d0+Uc5XlfQcvXiOJoKZkc43yRdHqG2
jvA0pGoY6NFyYxA2TBNvNh4Tgc8FtwNOT3pkW+tTrVhFWLYZF2BMqH4zh0PETqLTomxBam1g0cmW
x+piMHs/kMZUF62w5XkM53BMct5ZfPMIw6hkljKEbb5JZDThTBWYIO6D/cy/s+rOoWSNXxLMZBMk
arglDRhS+VKP1fbAqOj5awTtUOaqkTUVLn/FatWy0x07Fe16ZeZkaZwb43h5+daQsMNR8CxAs/kz
9fW0zrCu89ITlRMvRlGcj32fzLZq/nOoXwMgfFBaox2eJV5ngzkM62v6DNTQlPwXd0ohBo2tkV7J
caMZAnsS7rvwQuLeUXPv36cpBO774sDKDHMjD81pSQNV7MZ4JWae8NgtIlNiSh0OHxGnxFEGUjUf
4d8ia1xXvOPzUw9+hfBFWNZbehIiivkUOcYk0SAzXht/GaexQDQeBe3nwWWRIQjpMjQb3QaW+uMr
MjJ0A+aslg7sf39VleRFKPpmKh5QmFGMssFXBVM4EXCS38hqsFV8vH+bOjXVWsEm/wIZ82/Z6jaK
2D4wSD4Tvyy+Svj7tW+jhAFPTZvVC0/s5oARYEc/5sjC5MtPSKF6vBNYLqjs09gLCAX1nowIkJWy
PvDr3/6UwZAVGUnDQ1RpQQa6D5OFs4TonDij9NpRL/M04paJs0wguCJs5n5+xCCG56b438raV8KN
cLHrUz5OKSF4SplX5k78nB1pvqsACHhcSEBCajF3wv7h72Z2cE2IaJU4ihQC4X5Knkgncdt4GONV
ky8jrdqktZ57FNhdBxu28FKXsoZaXh4BfAtvCBB3e2DJOcDKc3VN4umarOCW6hTNx4WVzETT0wT2
rsJfqVmdrudRxxIaEoz4WlmzxSXnm5jYMqzOSsqJ2misHV2S0nwfZ/Nma55e739g9VeFqMmsGZ6F
zeZ3pBMJUhlgQJ3+IooSUpBu2N3xQm6w18MOevstXuNQ+uKO3Gy6whtlsQD90GtYi9Lrb+h5F7vF
XMwOM1uA9JHnzkjqy8dwUpWgKNSipqOwtXsr8kHDxtBBJuLZaOZq8QRLNGN1v3uCD4qWXhKx5szi
sCqhk3VcHR6Ny/QLjj3m7p/NKS50xHWCuToJVBTHK0nJPGdan5WM832ef0NH8UZHWDg9UWSS7dlv
Ny8EW100nXoEa4GWYNZEgCtod97VWI436R75HGHrLiTAtAj09vdYwbe99bCwTEU8MJLora/YtFjP
01DhNM69jnxt1x4LgFl0kWfsfuv3Dtra0mzHRKgqAmWSwtJGp/GXVXxE+OcWFId+0j5KH3duMsR9
Re+ID7A2PF/UJ4MbqptKLMv2TSH38Q1USStdw8D1LnKvvLoBX1gk4tfwtVoNyY4BGG27nEmGQdSl
fLwg1ADPxrCf73DIqsWnmShVNnNs3szei8cymbszoinHeVCgHhSBtEuQLO7QsTzaYeHbMVQSrnak
GU1lPQSx/yVfLz8myLYlSywvCNlqgbgyMvFdCCghny7KW74gyUqQtnpM+FOZiLYSE2VJO16bkNM8
78VQcQPChUHaiMBiPHcIWt6CfD/s2+n/6p1W4lcNxH07WiUnbIi4tF3C6Nn2st/5oisGCNuXjORC
M9ip6si8al3EXOV41HlPDLnVlK2hkt6zvJEkLHDOu88P3CzqsYwWcdTytsGQ2AQ3ySyL9jmXiH2V
kXKtebTshh3btZ+pJhQqonQZK06iYVyaUTnmiAPGgOAVW0nYkq4Cd2l6TkKw52qHL8ezW8OgPSog
rEU3t+9NboUk/fktVDS17QBU7tnXqMYbX19ap/jzdZ5eRW9qCQwLDLC37IYbhYlZw9asQdE+MMPz
rMAJu+oUBgx692aptJiSErzZ/2zi340Ey21S8pi149AxacYEn4iCmp7sTAIzUi/em7tu0/YcBYyo
vXdkGYc8Pv9GVBFoOQcVvmGL72q+OsqLkZTzL8iVzbvbDe07wGFXwSbbuz8QkzkKTVK9LlLdDHzB
YBwqvbbW6mKfPWu+aC4ONLhBYCDdsDHTRMbRP6nF8JQ0ZjOJTMvOrcHOYcFjWg24UgnIO2bf2981
/eSg2BReVqxcd6tSgleyLqjOF7fv4YIZB0m7r/DSSf8/wYirvQXvyyLYypApDqVma7eS94KeSWZ/
P4NnrcT8nqg586Qd88aCqAzpGIv9VXZMUex8OTGvTh7agMPx3WVkR2EDU3HSRWe1K1ObmatftRer
uS1nrS1QfwCcE0oNEwn8+fSB1K2LoJXRonncT52vEw/8LlhahaneeudJ34z92maaTaqRyPY8RMA0
Q71nRHHhQNrqfoZlpGbEKYhe+5zaOBRIkWMhA7xHNhZrMr8MDhj+TKMgEmwIK23UycDgKLBihWtp
CXfg3OCEjVRxcVEW21ZCeLn+dtAeYVBca3G/0E8sUczNnLhMefGcICWP/uhtpy5Z6qn/n5QbdG0x
y+PrPPKa+NxhFFih0CPhnoXjhWRzRsP7lkwTuny1OqU+EjqlVKbP6ktsXYOOZRa7lYWXeYoeh8gl
YHgqa8scvc+DNi0dr2J8P1h5Kc6Vj6Ql6T1gnJUA/Md54b9mCC1Rg8gczDenvzw9lr8QlPDOURFI
akA1M3RAeamCFKnyb1m2pgFe5jXE6GVo37paIZQXaDll74LV3BW6vfShWnrOIq43a2RO3ARPBUDg
niSn+fzcrifeeKoy+SdqrxZrt9Nf7DoH4rFgWy1kzfqCoJHWnlaoc/x8c4kyXfmzT7Vi1iAiTiCb
B5u1Djz305c1cMgdaC9aiSbsFMewpqfQhp0NJPje0gHoC/PAEOAvFs1XOzJAW3N4F4WSQ9uU+Vm8
lLIGEvZAhXxJuQboMOxxCr020I2X8xyG7DI4++vFJosvikkh7L0ELxYBfFumDIRvhi6dW20Qe5VC
dYfGpRACBxvCjx015ZWML8BEQIZhAoDIpgDKnNQcsrkrryTITz4o7lU74DQRwYTSLKJC0sP9WDti
yYEpoVSVt3tAWVYaH0FaOXyLWfvActAXo9sIKv+IXedpqThqxftZC6sd1HsMXpUmpVJdyuU6hr/p
peW8RESWvEwifYfAonDhyoS8IqeBSlSeM5ZPa/kJzxYpH6J2vOgCWwFZsmpB4QqDFrMvbLO09l4q
UUzC2FCfLg4C4Xwz5PyofLJY/AGA5e/vN8HeKKj3sGGD+UycIUCHj9iKotpHYbqHI/XvaB2is5JD
bK+no8d3oUZB8GrycAwhIXCysKKoimZWv5JPNsKGSbJ8JdLiG603E1P2ZCW67DDQ7g0sVSsHghYz
JTtwsnVrOPDks9iQFv7hcv6EN7PkRIHnLs2odY80KMYhvtFLXrMZgdMc6YBjpDYhF0hP9e/Llver
40/VLVfkFFGpMSsfTPkKFa0CYb5v6RJnIz3YHOXSpyI6zc49E+iFzxhzpVdF1GoOxwqn1j2Wk7Eh
VxHMDNe5ni1ZesyphnPfs4nm1pI0/ZYd1yFBeqQZd1Lh4ELGF+GuqsHiFrVpBoiivkJtuHKREez4
1wgras2f7+vplsYKepgXp9r8MnWyyS+a+miAqGxVmgJmMLJzo3sVOGdo6y1l5MTg8qnckINVeJZh
xEowoBtsTfVg3oXoaH+49z6j/t7hNGl/jwvsveYPOcG4hgJ7Aax9/8Hzyz1ydL+e/DLVlRoFVtze
6uQEoWM9/oNln/3zMjjDuj530cFJ8sksM0/eG2h1nhGWbDt7ZiyB/VqEw0XCkowBuTgZrn+qynfZ
+nIhq0C/lp5FxPCDCpi2AKZTnL/JGE83J/GrWRzMPOhrFQtoY6A8Fu4qavkJjYO++AAT8CX91reE
oic/DU6igaDExZMjJnPni3KgBqtSWu1HwlD4JLPpoMSXZGIZDNQkoWpdtdCdGe/XkvA/uehjYVgO
WAI39zH6iJ38zMd6otEzoltn3nc6rH8XfXvK7xkpVYW8vsv8lNzGB6+ln1bDnb4zEEEYHao1UwzQ
ALbxzAK0a7xO38enFHOIw7oeA+oIiThtZVY8E/vom3mWCgv4CTz7zxkalUa1Bepe/BJ/3HEEa9tX
wAnoaUwYArpUQDqy35foHyssrtXw/PsaGRXQJhG8SOFJhgsG72zWC7UaAVwxQ0uQqocn2tQBDuaE
MJFwIOFQaiK8HQRZs4Zk43ea+uLFHOPrpyyCJleiC7udf2Z6JTU7Kim1ljcRiaYPP+3dPjoM5Y+E
jhB7aUlQDNfuXyL90sr1hIal9DhigNCN5O9Hix4O081iyAVKC7A3Y6LOgmW7xGna96lkV8c9qZad
jtG7AQJ8J4HW2xtGWwJJVtD2F8rPBi0PHUDPGdEmyJe5eZLs3QO5L1sZsLXOiKPD73LoONazLr6d
kdhPEmBjtWankL9ZLxwU2cJFN9aDaQZ34FVMDJzVGBtuJpGOOeGxYgvgGpZMclD+/Ky/BUrhopu+
5URef5ZEnU8scY8s0z2vk/X/O+y/CFt+zP3R99TptDUAsJGydoEH6RbPAgIyZgsH6FmQdr/7EadM
c2ZHeScXhi75549rhYnh1cMCfo2N0FQQc3VL7JwrMExxcnO6bSZv/rQjP3jimGlGcClH8tX7uRYE
bAiuGQ+V6L4J5b+tsk1of8IqTX/GjUP28rRfVL5BRY5CkEQIzNfeXi4SBFQ2q2WwHH2xbLMh8qYt
ClQ6dGaR0NuuirniYSuItu9XxicgMb93ZUVbh/I/V+7H5VUzW73hNE4Zd0P7Z601Evikm6tzmtsf
spb1I+c/0mGHdHg4aUIav9Xxc5KRd0pZubq3rJbokWNrEWE8dLBsTHcDzJ7cvzseWYMbE/7BUwK8
Ku+646LTCi864dI+7KOB/qNoYKKBjwkQIae7QCb5OiP8kxP1xizAi2MI0NEehiMUfUcqL28J+2Fr
1WwYepYie+Cluj/xxDPdtba5KQ2JpOUtvR4/wNSEakIPZ/sFaReJ6cx+BgjkWGMVrFt62o9f0pRa
H5BNsdIkHKbEhEHCrsNXjfBaF1YbonVXhXO4dS6KTv9i93mNtwaYIjwtl5GtJJX27lj+iWFS9nxI
ZZDDut6OrRycVJjbFmM/c9oSQmdnJKkNr6R1B88hsL9f07hlREo8sfsx/va6tBWm62+H3hqcTnx/
0V0WKdrn7EBOw4ghe9S8pdE6CanuYEIypcSRr8lxomikgY3nnC8jd2WkBwU2fhSsUSK3T0MNGbuI
i321SXP5rcCFj9P7Wfz2keZKJmf9hKWxeUZVDbhNEd/G6hJig2RSFoeV/bRPw3EGE1UzMxsUZD4n
+0Ohg80eORZihi2oA0iHJm9XF/U5dBloMaBmkOAckWwueFp0hCcE6+v2lESULTy61/NjTs/8D+jI
rjW0kTqF4XUbEeCFJDOvx5wgBq1PfOZf4H6T7jX+RDwP9KS2vtAisP/11z5ISgz0TRu4cIekA4Z1
o/V7reBk0IjIFFfxgcSXeIFluJM6eILFusg+63z9rh3MBu7LH3EmcKsEgRY/nNIrmWYgNMrZ/Lvk
QpuOSe6DN2qSkqTrXXSbhx/QtssqTjRJCKcrWrJ43ciUcwIA4tTas7Mgb4Njt/pPg6LJwaSx8PJQ
9eie1Y98vlC4qaS4AHAVRzjeG/eKEN7OnuAZ2H9BX9Qv4iYWpzpMun5blyvjRl+1E+h77Ua9eae1
9BIWPCJTrNC0I/WnOBvPtFp/Mp0i6MPGf4gh8dtoSd8dBeFT6cCXLeOv2dMdZBm5F0ZGYQiIe2lC
e4Pz6IeI7i/cWKPG4fpAr1dth7pQyQSRrbATQpPvQMODZVwYkwW+apW4ZxFjrZOV0Psq005Tu64m
yKP9rXA47Hq8S9O6ZTIjbM26/PncT5LdouV0cYF4YnHS8AVs5YcPAyURXs9iRgHiZDAbehNeztak
apq/IwmCGtgBz4NbsP9Dl4FCCwXJ5nn72N0pYBDk1Jz74DoqBi07J/IyCtYuqfT5alOCxbjDolEE
pIIilghP8MQeNzQmZVDcxyy0R/yHvQFK0zEUiNrDUtySHqrjVQsbBw7s1ZJUMU0WzcXSwwaTkTbf
dEvHaInmYCKfXRKCd80Jmmo9tp0PKU0dpgvy9zTDo2RHREKF1pmZLENxIMmXCmHbBiSTlrbHkPfu
1aQI2nel9jEeU06fZCmopGmVPc8zLh5dJFDvalH1VUJbGUhj7vL7K20eagsfHERHi82TrmU+zog6
g13J55ATljzuPXf+d+IEao8EHfRSo3rFn5o/8nIu9iNgdFe37JmAkugjgGcBclXdX70Em7Ljg2MT
g/M+2ZGKx5OXfLeZlWmGwiTa7QYOCd6CIP+QrlwD+tqSHpTMC+E9IzNMw383Fw/76MdjWy1G2JWd
G0vUAIOLCvA/KjjF76iA6LjvE5qLkD01sjbs3HcEO1DwsDagUKp4zDuKMYPqJgq9t9Ja9UOrKva5
91JkQY5y60yYEO6NK0rCX+gHa8GG1YLJ3wZA11a/4iZ6RgeyABy7vvXWJ0MLJC8zqfykonzWk0lx
k1BmvtJjs5973YR1gXBqfjpI4/GiCT+8kVW/7FXzSRwJCe0g7piy58ugE3A8c7c8Nga3IHu/o/Ik
iuIsBAF0Knq85EU0SmAwboVAWiG6s6Ukwg/bBrCZPAY2NcfV5hUWpT/G6WPXCnwzWszVNw7lYhXr
UWCGgJqrovteR9qlFdHHHcczaqsvzF0HTfRvUC7ACV/sYg24gmKHEdNpDbWJZv7tIJB7Xf28mQ/L
27+5ourc4yygPVJ0lc9+aRLe+zF8yaTTEvp9a0WNOaIfqbMJQripL8VYai0K6eKKiGFWlMt5WuCF
0JYOP/R+bLIZYUxcgwKauya8pFXTiEuSxpT3A5W8V89VsaPa1MCWaLcFJCUrpzHWFMqJgi4lnlBA
QVtsoLsfgMeVgBJXPby/stAiDlCEtEq+AeWua5AtwwpRoChZxb/+8fUhkq78xccbTvJUbH+M+95J
zcR7PpCc5BjnzNTR4fZbwsFzeZOfNwy3p7zeFhrLX0uznCmRWQJ5Me4/AU9+7gi0OOOS5p5ce0GU
9bVnSqEDk1gORs4fCMMB00kUhakr0JZfqN14JSs2XrszFsuSaCjCbkcfHSFo5RYJFK2TG3kd6REl
EFde6q9tacSIgcEEzGjYBwRSRu1j9NLVgNtj5YhOyyMblsqQmzigrH73/+8KQ5zyOC8p+Uolpiv4
J2sJP2wz6dfuLXj/zAI9quxO98yBGO5E198z9ibhgZU70DHMhKe17teiAm3bOrx2KCfK5QiY5D19
v4OFYaGA33ZTeMBmrh02KF1ZUxAaKh4GvBqGtgaXpxzwKoz+gYxURhEXIXv9+/OY13PUwds2+/S7
G4dAoz+PbOcgbjvLFJDelzuUgB329jk2l5Z1PMIk1UkZK079mn6Pe4OwAsuoNeW3kBe2plq4y0Dv
aTpnv0ME01/6BIu2fljrzxdQIXnVbc0nTu1rkDrj76DSgANR3019NZcHEyyFhEPZ7a0t4Ts3o//s
OUZGCnLmvy1xGK4i1UgbiQGIWdxZGJdqB04xtKjSXly19OomFWxHT8fMAjr6WW9d2kDGPmNGEpRK
upz7XCXbCQd3qZ8zzYXKr+oAkK8B5hz1+6mEeSa/Be2LwmT9smR6N73SPNjBwc7XKb5qH9ujquHz
mE12uhaokWdHbPkrhZsjMfIWKetHQL6V7725Adk44lcSOhmJTVNH7kepjCWU4m33UIAOx3iDj+3w
phY49LxCAIKi1DvEERYcvdzvt/X233DuCOCP/aN3rUasqIZ2gVCyLpM1A6IQEgHLSDcdjJ7rhIzw
YdxTS9mo1gSgXLS9Xr+B2Bwk0Gjl8ulL4YLAmGWNckG+1SGYlVffWZCElaGz3EuI+zj9pgMO6HSh
eaM0jW6bh1QQeGYUHoSknK8Kla8wuN2/0otkn+rdNN2Z5qKofKppdrk5ldgp09snptdoR0z7LLOk
1kASVZp29N2E1oFUtmfswZH3xxi+synqz+IgZnrljESgaB2EMD8ARTlXoEoEQZ1ydeiQkj1sPJTM
PtXN+jieNwYMeFjz/mc1Z+5EAieR7tWKN6gasUEFX/5OslilyvUq9R1kZqqWLPVPPsLGNjXJyGHw
XlquLjvVWpLVWJRcrU3fNYAmxFD8h0mdTq2mCZo/4h8rS0gX77PaA+wkTs1dfblkVecwEh5FX93h
dmN9sMpqM4MxrHcz7wdI3e0/764AzP0rDwsSD2ldhEbRhiUu/5NCHLgcO1fwLX9ndUAxWz/dm1NH
cbfmHLiHw7cJd2+lPBFakMU+FmbnT1eR52YeugC0/CCKT+X5L4CIvttmlL4f07rdFq/iCAUBUL4f
zQ79v44ISqvbaBWUQ/IOC10y28IosLDCFB9ygHz2WV9XkgSUJOhAxjIS5m58MaS3FMEapsHZ7NLI
QtmpbAypc8/vfz1nFuSjBMOlggEmVh1Lxer/TdNGbSXLmDDpTQn0khAk4RHfEdoHOHe/gsc89+hB
m8d/b+F9djHiHv6DfqZVMT1MkAFdXM9m/m3oStdx0Hr3xkaROGcYUNhADo+cjh0G4XNeCs43Q2fi
5tiL/HFeuCfUDtZRmS6J4HTalFEGXWPM2dVkmKbQoeS9bIWHad5LcqugwX11pYE7/+wMMHu+Nj9I
mHsFy1PY/pSsT24XeQXENRgBVMl/zQ3LA66NsSKKSIPw93hVWt2B7ugSfk1U6Hm4duISSOHajb7T
Au97P0hwCzT4cAkeckxy6UWrDTZeDIDNIzOCDmhZSRlONgR54wt8NUkUiLEE4mm/Qc28jQbwzNq6
bLkvogQ99d0jayIEbRuJH1K48PyxuNHNLMU+51KJkkHbFd+o2ORAwyW4pzm/dAQcVy/He8qhqSkU
KCHqAa7V0dShaMtoqn++85CovhorQJKsBtIlPS2BTWu9cReFQQlie+kMHuGL4qrASU10Of9yJ26w
Bx7fIpNrabBcAvaZOQQ/xxBvV6RCV01liqyInAM1y11I/9pNiZxUzjOz7xWnxeZU10jinjB615O3
JGqP+MsezbPUuMAguh+tsi0oEjnbWxcIPZ8sIs1lhrW570qCtJP2S+z3oHwh18T34Op8ewT8Aa/b
mq0Dr19lFTKELQ3Qyl74BVhKuoijo/YlVs76jeXwBLP4hH8zr77abuxA/0MfuLubJxmDqRXWsKfg
7BDf63Y/9R5lrJB39r2917bHTvi3+Lye7xy7wk87kE07SvlP0/JagLlO+o/n00vUWY0GEReoeOwn
p+xqSHun3AnXcMgIWYaz15d2X8BQbeTYkmMYPMG55mz0s1sK9vZtdo23FTCYsILcgPY/g6MURiTz
S8JtJ3kf6cp4xJEKupfdMVDhdkY5B7RSZwCVAx8p0QNQ+MHn9JEAjKuFCTJTrrdju/G0mFFSMy3/
e+9domzxj0cJwY8j0OTeZTQ4nakTAxn/GBKwiSflQcwMDueox9w/YopWumbtNNRgvmMt/IBTC0LM
670rW5bGDQaLivxwiNUm5ytKp3sebrK5YmYU99DwrJHPrlVJO+umIzSBCV+8vwaH7ypam4yb0F4K
7MWAPkZC2MaJ4gKrpH99stUslwC9NjvrFcLvVYWFmC+RPk/bzqtt9gvYBLFzt5GUfvDgCJPN3P6i
J7wKR+xdiZNYka70Cydr0HL4sfoTHHi3C29ShBuAxf6aF/MRYf7Myn7N3d7+2DANsHlzCe/cNPXE
0ZMemSxAfL99CBub34Ep2qthsAy4ZTYlhMaA520o4iJa5SGc7cmQvloqu7hj6vVVgP3P3oKN3l1L
QkZIPgsCdPmQ910N7HDHKYfrDSnc2nHbpCX5d5SdlLRO/q/TljOhNVj/yVB8uBXXeJzPqtB0NyNG
Y3Lx+HEp4Y3xNQ6bQGzsTNmOVnwTqAr++qb/PSyPEOjVNN304/yklC4BgJQk82IgMq1DDRHhlWB2
3WvArTX//wgEh+1MKtdpyiHlL8pSfHUNG1PKcut1AI0N9q9Tc50XvwUr1lIhlKgslFU2KFzyNuAn
dznPsuUV/HW5myXv+OyUjulXjKghaLaIytLpbudqCPzf74Hqy+435YkNgOGV6fajJCq/Qj4Bq6N+
GpNdcegiX6/UQihucoh0hxrGdbGh7jmWeO2VIoaI262KjMed2+kbL7SBwaRUikGI2LMlc3CSQ8B2
abNQvsk+QtzqUeMCmXJ3yMDJ8rjN/adz3IixfjJ9i3e2Wq+tIl+JP/2R8WzTgOrKo11SuGWGfzce
YQHt0wYgu2btj4nnJ5lwyO3gtCPzf40LbNYr2WdCMipS0r7GAXwRDbDX07/hKqL+aJ7piiNfnFgJ
xI2nX0FQtGU+ykaEYyZKWAMr8YhyLy8WRS9YGl49mUn7W7vPpmyi4oRHO9o/OomTzFuLT0KKJgaw
sv8i6PcVNXft0/6s70kMusGjlfZIwJAPfFBjqQS6kzWttR9iV3QCtFmXpThzng3H4F/9FK7l3i2G
/2oicidfiJrVpkQmhxi4X82zsYcwfv2/RIFvXtluZPX8ouqYepJ4S0hO1b+Dw9evYc8YFRtS3ywI
Xg5dFwq0m1C1Kb5WgGva3dz74Gx4ImQ+D+94EDqc2pQbVRSxX27PPObcJEDc0mJ/lmpHwsAjZgvp
nblA0kB10VK/iA0JRUh0Y2sNkAb11oNm0S74POTG26PEXANQHFeAMs6RuF8jQFG1Km8T4mbVDeqv
l4KxUqzQn3+TRPpRzAjFgUb42bURhi5bLpPbMRqmPiKqsaV/AAoaxra5cQDqZpOxI5j8iKlL04Ud
CsMuXtpWGbWnmmy23vHGOYd8f7OqTsQAG1nHXSrakqH/FV9Z8RVRLHEL/SQcGRiBTtxqjcWw3FxQ
MhsIwcPWPVDJkVGiJIsQHRN4WZyTNxMJiHhgQtuVUiUp3GVbY9GMDUX7D1/qfy9AhxU96l6BwtUF
8k0dDWT/+e4qwdl9cbCD4vZVBi4XyO5MXjk3B0SDnAKE4ahSzWxCkP0Bm8puYJdwkikScyJOmhT5
0wWrWydxf+TvN+H46oD0GP3Ab+OILYOP8D2OIQLnEEkmYp+SCziY+rdKzwOWHoqK9mlbkFNnsIn6
MHjMXBQ1Nl0XDjxZlipioglqAk7nfcqNdFKGajyCNmV5AEnd5/+MuX0HhUS+Rr6AsN103K8P4/BD
nP2yvgRdKUVWy1YPX4zDXFTycBO7IukwfciXxW+hVIVvHHzEeLjUtUX51Vo6dnjroalGcBAuVlvA
IzmWSsRKPlt3/dqJvcylT0xh3I97CL/z9CYdh5QCPC7AKzn7x//0xGBeuIGWs8OdrteIJOGBu8GE
GyxHNzy6MQXLMLLgrZU4Le5tnYfFFXiFPks3BnFH2Zk6dAzp16efvMg8m4Ll8/BegNf917gAsPh9
1aWY3SSoff2aBdz2oyri6kNejPdBTz35yRj+ZiUuBZi1pcbY7OeIaeEUQ/ALPKREg2eYg8S28K9j
er0mN42PPk0FhYUJq21PUnh9BQHpvdaIe7fmMpOkBKga16Z+on1U+jkKkdlFSXHGK6DIqmQeJtaL
lNL4mfOuWYYYB6oe4pbRDr+TP1vrJQqD8mg/B6qbaBJCXoSYeR8D28zuhapNHy1ocTgJUj/0HZoa
4N8rOoy5HgtQIIePCEeM7UO85R+eS+iY1IfJPvdUdD9MWIj6JS5Kao5XWmw9cRw1EUUf6zBjdEeg
q5gkwAGGz9vRKgSDwCMr//q1Spnvia6V05euQeFne2jgNurlu+v4Vvj6udilPumjEV9yLJMzroHo
FuF5mKANrzT5TZ4V0CqVbi6lMwF5KrE4C9DTvG7MwTP3n5MVh4FSFpzdbtRfcl4CrIOJjA4CtO/m
f4bG9n0ba3/HCftvurf2sly89GVGx+UF1MyuxGLa2nYH//unFsc2zfFZ5UZ2P+cDvIhZeXxWDtPB
JlToA7avad0OFrbASM/NEvd9xZbsUI97W4KjZ02+AVfVNVUKiqy69ZOEY7W0cOvDcY1fNp/NYJWK
QGaFyzFVDB2sUM7aTfVZ/ZHGKA599JK4vS/7PUwSClZ9K1k+A8OixW8k1MB/9sclqY0TG45I2l6n
SlrVPRDB7wZ2cnuS3YvzgrbLtkkmPDX8hAUB7RnMCHFXv5Gh+1/T//XBBRNadCkZa6Os9dO4W4Sp
mUXQAAE6HlkSYvlQvZ0HsEVOpDoANvlhl9FS2rZ9cBspSucnvGq8aGYksbqD1YL4b2MKd7SMVoSH
Pt4PS/k9ImYyI0n6hp8zgcoIksPK7d48gKdisc6oglZ1vMoIHdSUhpZqS+SXE2fmDYagOvRYfrKG
cLdIybp+TDQzrnu/ePnNYUMs3zIk6EfLyBzdcBdu0taKLyhRjy2b7UW0LUtdU40waJWF9X6nJTas
jnLbi2TiFgWcDm3mDRhu0qYPcZyLCvcvvrz/O7+UX4JuWa7tz93H0dGuznbR7nSudb6pwkdsO9Ut
KdlYUus03Djbl3DVaqJ4UXhwj85kVE/3+DzIp2CSeJU/nQIXLUFX1zAp76Kvcjh7MNJbe30iU+6G
Z9zB+E2ygzqtrqfyr34UlUOLklZQ8K5VgX8Gp15Q5EJsY8j7S86AX7H8mad5RXQmYUoknsdtv+PW
BMrYBEphbEQhomYk0Y30T/13++arHNAwma77n2T1BJVcUjL2sK6C2nSzdKECVjZI5IZlrjMXvlLv
6kPJT5uGJvd8Jmr/eViBI9se4+RK6sw/RWD+eelF4YBClgo1I1Y4Nt1Uxb44/v3MTvJVZ2GV+DXY
U6uzU4zGhWop/rhBtpFCULnMeqW0d+xZeFOS1pxzUDzEJU33e8yiWkl1uqztixKvX9NEpUbwMUqy
qjF1+UXdg9cyfaLWGsZi1ZOppQAWqwZYj65SsUJfCP0bC2xKz4iz7gJtYA+Ky48p1ZkT+L4OYn15
d51OnKhtncHLW01q9oMxXKI3bkT9JIJZ8uiwqR+n9J3CszLKU5LsBYPbrEE4Z57YzaQdFT/TpNHb
wLaeE7ugG2752ZVZD1Uzc4Ocqen1EHgLgQOpsVCTKOIJ/38dVr5rPqcMrp4PP1juBlQA5pcgQAjA
bB2mX8iN8y4qon1aNZFcGPXpe0HE9jul86O2M8xUddb7QXHLwCpgtCYNXqtd5LgB3k0iz4cjBAQ5
jdzRIBbds7aEU+GM8NmoJmDwH6/PwxWpHZ6Oj4NXqa9xMiWzfvuMX1syIKO7tjgxe4ros61b7TDz
sRz6t6xkZT36ZR5sMZMswBQP8PhUspI+9XAvhCXUSupQB4+Mdziku4zb2D0kJrjtWno/sT3NLoj3
W+baVlBHBBxBzMuke6v5qWeqlhceeUppqKLLg91i8CdG5dzphDMlhS7O5k1TEnR+v6KMJ1SAFIDB
b2BYk9YA34ERWEvFBQJLRkyIbDvoeSM8zat+4SUZ+TSiTEM0FGMXyjjs+Ibss1646YlusTo37dFT
7TVYNsMgYsuxim7JdJFPTDwlyLpiK0EjObiEWwnH9mX4n4Y7UQRueMUK9Pz0jqWgFl2xxWDNCKTR
7qZWV1ngFIAuSsLhE2B4QeI3IOpyMNuJh+adAGVMCpw6r+T1PBuhaBMh49kA9irLM5+A8CyezxwE
Q2daMyBARWIcNoJ+vIUdXLDct0hMexkIjIa9cOGpRQ2lLzCrBGdvPDGGaHmBapUc/80104ryEFBZ
Fxp1NQS56I9DwH8boWS4j1ghpJq/sR7kOcCYu84RbwKr/plFmLAD6sPqEoIsMx5nJVtBVybFBQMp
UROFXGiYqfmoTo4WZDa/txOrAy4b7dOfMumOuqzBjt6NYo845BlVblhm42gjA5LR0MqAZ+vGCcC8
HMoUzCLHhuUcGlK6Nwdv8dTf+KAej9Y4GN+C0JjVm/5IMDHt8TdLs2wXxCotaZDwa8TsZaXksVMD
CQC3+itgOH/WmEGZCePhdbMkC2+xpmVz0eht/rUWeh9zVP2bFOF2ICTXXxRNrcpos9PJ9mR4o29T
PfpXli4mzE4HXWbfctD7tTRsG5RdicG5RYrNIk2gAC/4rSLeBj/t1TCSHyVEhP9wajR9Dgcfthdx
SkMmR7a7poXv8fDP2pAZs7nmiOP97l/ZM5sqRLqoXsxB49u0+nGbREyJ7/XIYYDZgIXlRobsPRIc
XqM8a6oLtcl5RJ2oMl+d/WuCygv69+9w1OJcgWlMYbwzUeoajaOL8S/98obYvBeq3kQdniNiYnGP
kdj+hC6ciynwKKu0amG4RaL5APOmd8EU4MY8QgTTVy3YjRZc4loYMmXzlRx8bInc0HxuSYmrjfMN
Q8baHttcrqQdgxLNfC24Rki2KPHX4ANsGIekeJn81I4zj0eJ2E1631WKiEL+WNOtwobQLi+zz6jj
XEOc0mEwgY0zRw/IDTPmQPp2R93kNKhchDKvAAnBYbRAz6RGHek/XCFmjgSj5+44/VPN4CAt++ON
ju9KTX7fafPBeuOB2xWutNOmHmZaqh0hqjWt84sGoqsbau5EAS/OSwiKhrvU1XX/GunHhM1yR4Cc
88cU74IJO/0OfuOrebLu7onYvam+n1Ms9dKeegwl4INh4uOEdvhfUJLYTbY3CvgCpV8AUuw325vz
5lZTyyLfnAF0eRu4P20vjgAE76e+Z4on95Mr3nezw9nuDYjGk/aG1fPJOVZOnQNCFdByWBFiYhWw
rLxIYA/KJ8jex+A28Zb2dlRLImWZrnt/HydKQZoSE3vUaVimtUOMUbFViKGqzSMO0WpqQfVbB2DD
6rSr5rs8tTqYY0W87Ly+y7ZwWDGYoh4Kkpjt5zFK0STfq+DV03fDQL9mdfsFawIdbx0l59VLAl1a
Wt2y/rzdEVocAuBUi3M22rkOo4eHmNk9eQzxW4dUM3qdyjveS3Emicxe/teQp6FhilO9P1fIVg1D
xiHs0RRmp2oMDaCy9nQ7KtY1y3lozJjR+WRmg3nTkXaBmVqeEY+0q02z3nXmTZrWK9FwPKQ61P6+
fL9oFut3yLAER7MzVnC4qBc1OfhcnqTkCoWSl7sIGxZdkwsOl5aRYm1NxYflKp3PbwHUsj6H133k
z6x3MpPbSjqrtZ/twXXkYuABdljSrErPGn2CdmxDuBt9VwaIXxziFaQZ5YHEH0YYNqU5M9G0A1JI
z8MVJiN9jUzGf8rwYhmTP/g0T5cs1nD58jdCXiCfq2iO8aG/qp3G4OVKzT1pQAOOOiGGT8j+e/qJ
qYSGfmVN1lRPTlVfh4p5aHMDDzKAj7TK1MxBBe33e4MDoHMK9oBx53zLg3uBgL1wvqOC+3OoUfy/
OyW3EfcDNP+IdfM9JiEoJURodWzPsqVDVGL2JGrQKCci8WfyyoK5fAAp4JjBLFiOX7yDDM3XSSxN
NY3Ofq3UHmBa81wDwTcGWh8lSxSGKvo1fpkqfyFZRxPP+UvxYyrfHmp0FI/GZGxAiNzzte+U9975
Ctn8AiSV8CO+uniQOQEOxnEgRILEtUt3Wc58R4SQJ30RnJ5EHvamxsE4TLqeXelA65OhLEIsqfHX
8YQf6iIr98anC4+h5o9G5H+e20eLRnTBoAjDofAQ9MS2VoElXo+OxIuSZ7gO5L9F8uoCaSD4oyL6
D4+SK0VOk5KJT29g4L/03frsIaAoxFS6DIFvcrqEUc61tfWhra2THw1AmRn2KGVdhsWAMSxqUQD5
Rrsvw8L9aH5dY8JHmlIkUfcUh6/UP9TqmOJy3nWxqS8XkeWRw4q0YvQdTQNCCVOiIldWvOAJw8cJ
DG0JotOh0EQ+OyxE4syLTmCee9Vjcfv/wtT5qI4xRsu1rPjur+U2BN4Qh/b8CtRtSFuHAUSod2WY
0E6ZM/HV/M0XtIckxNLhQVf1hnCbsNLU/RJst0gHgNTNRYDD6bs1ERDfAMU6s8Zd5LBwJ5flzq5S
TPl/SPphWD+D5YZmXDicGdoF6bIQjXwkRp/ibKbnaNnenIW2QQlNyLJCroBq/WvzW2/epgdRelvz
e+3bR0a8QJnmr9Lr2vleMMYOJZnXiSmlyuL0a1myxjSUP6J2XAJFAZuZBFHKH6sUFUFtLy880+X2
Obd6hmfsx1M4tk5lb9XpsGRetugzVQ4+4vNGeqGz6GsUrotPOhIKLdNPj9Jtz/WJ8jGTG1RuyHrR
OTBnzz/A/iLEXH7Lqr8Z+mPVtO085eY9oU8qUHIOMqIp+e7T3MI6U8YEtsdoOR5KanEycwXqekRX
Ynr0NxWfK4oWfwMp3pRtHwh+jJdk8xd4TPDMr6OzaTTJ/Nk/awgzAfNii8WnbSVKt0fYWdq5yyFb
+3YqWE4SM4aawxl1yRROleGNEwPD8g6aztYErNoDLwUlBkYd7ZbA+0bN4dQs1Q3af2nRTxgICif0
yjH5LNwU6lG92Q+Dj7hZJRl1AHY00U4psKRqNOd0jGwYU/WWaw4a9AOXeEZyns+/VtL8WKnFQArP
VuRWydJ+hPr7t0lArrxQgSugIHNPb+rrrHnAMb34Lv6pvCGsIwKGN4KGbCchMylQdLZKQu3K/OFh
CJeBB4U/2O7ZnSeMr9TTsl1s7C+I9G9v8H85Cg8oS7fTfZqJzx6TnQXSWX3IKqHTEPj4A/8yc59s
9itplaYJtbPlLIrkpl04xCbB7zTlE+P+t3DVAk/VppXOum90iA/MkNBAKNBcgT/SjOo5b88hf2rl
FV9ZQu/VttSE1OUv4R/NnfuaIKyV/D2bQV1jjIN+OJ/ulA6zb50uMbkjkHSvUuWV7CJ+Wz4saqqD
EZoFvOdFREF6Zf/OQg+tWcmDz2nU1tANLm/xaZhwGhsox5zoI4iVj2zOiQSyUkEwNUgMOhC5FWXO
JyzBSSCEaHk7iChxDHxIeNqKH7sZGGJwu3p9sAieYOlnRbgLqLYCcXbE81FXCDhdQmW6KJpFuYWv
mePhxWU+gqWpOurAxomgEcL/AMusWV/BsvHNH9Jg9RZiPB+1SDiEhDOGgrb6FcOO247UkmkV4Mih
9Fx6699MU5l9I0x95eZjmAa6skxRcxhcdJxtZ1rMdc6dDk9g1BQ9QkwkyVUraKEhX+hHrye32Lmp
Mq/RPiakzqp064Exn/NSGaWgQoeoQlV2lvCYoTcgxOo1XRbv5ElQxy1zPqPY/WsKYA8tFyTzzHnV
VieleG7iABbiOkHIEj8oMmbRONptbHlLVrKSi2WX5NYiV8IkX9eW8HeV0WStkvY5OAB0Nv++5FNE
qKCgsA590nrmWHeMqWN3kMxmAMW5/TjCUFGhDkHT8SFS6TZSE8dQ8WIpb3P62YL69m5bNvWZbbeK
oeCvu+35VqKb2QAxWP++rSh3n2rBm2OoaVAmW78q85UJjwojTi7GVcJBLbMKRqhyoUEtErhpGWsx
aG1HGYS7uNXcDdA5cSC9lOEZL+2SIIR4FJ3utu0mTixTvOw9vWNGUfJKR53wOxpyVk+C3diyJOl2
D/+FENfwdVnyA25HAU38JeTxaSML+AzDamr5gnW1sjg1PqzL8/C8kb5Y0TaaCaffWydQpEiy5ieG
9MZs9tMzf4QoG28AV21uz0XqPUQNl97h7ar8x9wQMPrH2tVJaTn7FFqsLunjSX1/9F6IbRxneuBN
SJRkpgvruk/A38950G4W1lZ8SEQgrMOPxaIbEAkYZ5/dRnjCJWRAuxZHOJcE46V8QkNAYCVXbwI3
mEwVJJw75K7DEolrF0GH4l9sf1Rgr23bk9TyLDlmWDj8HOeumKZzJYwpjNKrnyn1m2to/0KX13Vy
WSBxq9P/24hAiBaRDYgk9dtodVrSr/+ViKeQaxWHza7GSI6+kSdEp3FP95Lb857sSSA5fJGiRGUY
ioLNxrJ4vHPNg0NLKk9WtzM4dHGxGKnaIuH0Y3GfZe5jcy+ONzxFdhOEt6t13BgDhrDKgaPNEK0o
+ONMflXTiIIZB+hrkjxaKeqTtoTNYu5lhpfo7A+tcT1HPT8m7+6g3dJKpovXOvwQSIZ1ErTMOpho
Q6t8900bW+bK6Qzo88oRMgIFNpUewn+4jK0aV6Gu3Y3MQEFpdj8ZLx7nP12yvGHLMw/IBM31HvNa
A+Dtc+Fo1zFiRNgTvCTOft+doE7b3aGNEGLMjaIH4tGLrOboKDPoIgbc/Ry5wN+EH8BjzSe7YW4p
XaWhVLydD9BoqYXXUMiCpiHoEZL2DKrLEwjXl3OWkngVEAVPBpnfBOhbuyEoU0k56m+dEUB++mx5
tGOdT8vsM7HxT14xjljntnNua9NZ/ODdJf1rbewL7E4kRSeXlVcDQZDYpVRg2kQ+4WbGufJFTQxh
zBciNv2/F+LPMrsmU7W72sga2R0ptVSsj0bx05kdOJFccglax76GImm78t5y/vUfXX0IrEXIH8K+
CVdQISNx7Wy7AIO3BNpW51x47LbBAnRbGj5Lp0bibrOGI5gXtC1/QPBg8pl0wzXOgA+k9tBThLn8
ITdc1PUkHvy+NEYBEvdOJOb8BLEPx0LxR7Jjw2CnW4um8bHRzV4rFKGXR2aIMiyrL1jeq+4jeOL0
jJX+OHQ1YUryNsG+M7mnZPrdT9HmDCoioeQ7pb8JFQXL2wvU93iP01FLPoKhqv07UCdu9B/XtAae
B+Brg/U59+fgDVTCEZBSWGzyRT6iby7S6yGf7BI5WczaTnJDD5xHRq6NnAoPfdrAwLPfDYhygxvq
hr6o8nwi03hANu67P+ewAdw9O4rD5HAvg6dKY1KBGC7tMrlZ9/4/6XqT2kSlNAMhPydB/wkyb9IB
7mRTACzAx2dEm0OBFZd/dK9wmVNLac8nAArJqmXhKT+ftgyWv4lnDp3AH5AVYCid9aIsJm65aFTy
5CfQ0OPL6pa+xe3rSqrYMj27UDRk0FfupApvtzAvtHcA1LQePW8f80/ZSSpso+jujAKkuePvzItQ
6y+J4AubVI25tCa7iCcR4d9Gn8p1cRQG213s42h/cQmFdraJYzMATHxJl4s9Xdo82Ml5Vl/dp+8k
7OYbpAJVflsEPbPOEtw34WWRCnVtWjb7dmd9mRq0l4J13xurG6xDiC/026e7FS1T4qgNDJntzWOT
TNj0PzAQcLcL2wBoPJLDRLBNhIu63FO1n5mEztx0jHG9AHJDn2lFmcPJDklVDQMLbz9iKc+dP8h0
aBUw8lQ8rPFhl2dO3AysKfSey16/Yy/pOrqAig7Q46/h1PmGz3Dn3xdW+aHr0YQNUkbOjyMV0a/G
hK2sgfBLtdDum8e9RPYZ+u+nmRg36jIyh0uyhJYa83SXx6U5/2zFW5iIgMyN6ZLqh9lZ3UYgtv0c
NEYn8NWPBZrjk3mvE+U/r7oU2IwzQfflRSBnRYgXRmP2KxZd+A56LwYKmyqEwL0pP6Bat/Ll0wc9
xh7OetAIV7t20rMI2LFyfUHyOU9cxhAuyjTF/lvVgpHKbg8JPR4oNUjskmrDuHyTNGdswYWqKuY2
PNtFTTYP4eG2zGTLcjXtYKW8nvx6zfJYxr/JmIqFpRAF976k5OPqF1YBcVHdUFEWH7wOhwWsaKqp
OmOgmxULjS643mPf8DU1fwR/0UgUsvZgaRDf/9w6h8jv8fygkFHR7ZURm00QP6X0ay35na4Zug2k
A30WTgnAl+dQnjzzd55Z7zB0RSpNVv5ysh41pl0j2X32WEWNRxbZdyJTLSa+1jKjc9qf1YV6I5i1
eKJ/q/bKKe8vghQEtpjQJrgtI8eFkn8g1VgJHAjHbbRueXcjbW+hBOrpdlFBicsWAk93nXrMKRyi
dZKJxyovDouby1HJkYwEDoK+L+mV2G21dthjihkzJreIIpLQIrxOk3xYAvP8qead2LEtvmDRmq7V
5szWRBTpOmyeQHrD8NGci3wT/cq+CWJtOKekgAgkN8gq/cgXWxvQ1nR0wHqbjGEWj4HOXe20MZZn
cwCfzMHvPAa3KbFDAa8fuU7Q80uiKPvNOuufv/I0+g4oViWWPx1/c/rVvyhFbhI99UHhLVNWdfL5
JiDO5mvCq8ICL7UMyDBj0uWtE2v3k3CBPhEPws1cuOTxIRPUazR3ZsZhJ9oBAae2DJBKujwc5ulB
pve8GSQzAT85V9UXn9Q5/pVFsG8EcAAEOivnQwYF1jL2wGI4pifVubOcKl91ZKXvK5eI1auIBE0m
Bc4oaosx+VzyEmfJ6IWHOkouhMwCxHE0XSZexITgMXGSOUE/7UIPyuRH6LqHGkGEL9j7A4bWGzcm
tLB9nJoCIx5NaqX9S8y6OyonaRVSOxvQpsVwLMYs1o/MGSWIaJ13Frut+0mCfVrmrzX+mVfZIkkJ
xMnv6BpE999yG8DN91HJw9AY5U4kO09PUJfF3ipL+p1Erk0cs6iEFULakDSf78m0URtN4lcxpqlE
Iu61ho4Fj61h4oQrsQ9+C9GArXwNPRwXMpklj14N2iPl0KRlg/AAFebqBlO/pxA44J01bA9bPN2V
EZ5p0iKf0ZmCOiRB/xYLbXx3unfKACtlNKHOJRrmhFy4OcmDU1wFMdpoF5BmCItLC+yz4xpsWjGc
ids8HSdtT+uNb+AcyQUGknmVha7RGDSqHqIpAtvO1VNBT7KBKjJB35i6en/1O3Ze4vmXQ29uzbAB
8ywn5fe4j+tkH/op3hfCN402om6Ks+hq9dXI/nPDLBSB5Gyo+Veu8blhqQtgMgFaP/+CbdmTR+vO
x9ik/qHNEdhcZrmYhbkeOhAut3S5LPmmUK2ToLtHMyM0xqbwkOWl5MjzI4c8oDLXj01hQokq5hU0
xqfRHPNd0z+bEnGkFkt3jgp+LUyDjrraI7C83agfqgOZiPlBMun3x+zuljAKgZ4d38kppd5QJD9C
RpmBOZTfJudmdTwQbCYFY7xhLK6Ou+MAegsUGz2/cv83Hk/31n2DoGTRAi7u3WtgOf0sqJzo5oTB
V0X8M9Hw5LaXOAhReH4sC6Gr0hBlacy26iCcwRgY8eQuaIFrVfX31uW52Xne1/ogWZENlIJtRL0P
hsSgEO2qNZKPX4zkWC6FTpaJBzcsyJnKiDal6TxFePXj1TE/Vh8ygcsl9eBjMXljwzxS0flH2TKz
3VOYVKjAlRBBprZbLK74fK/sWOJIXy07ESre4TpN2HjzkQj0661YHjUROVRNB3Y8kzSiDUJaH799
Dc4CrImxkuEQ0lNfBqF6iSjeNGrTmm6Th/GbAC/NSVIfqvqUEKBcd7QS2qL1Kf55EJDLBuF7JSEE
WSTszO8+Gna7/fxtnYpCiRx0khr/ybNbu21kxmaAHxziK0YpMkjEBGCRUU1e8zKRNVnObrQ0FfQu
3zbEaIG1e0pWJHUKzAkdUKIXn+uJNflcXN5h3cH1Jhw15HE8hnZQsvhbPq2l5salocoiDXVydTCf
WwGxbjF3sgthavIPdLHxGcn1vNO2qKd7HY5YkCrnIkf07dGF0mXQH/5JmI0j4G4jdoTOwqp2xAhj
+wre0MA5Io1+omly4SWG8hNDSqCetYfp6VRRdNkBTnVBYZxUaOMGn8QJwcL46FyQuC7oeC6L3b8y
CG9m5+lQzVZUD5GnbtYgjhg53fZDNzVRxqfA2OkC1oUMTcO+Eemq9m6tddmb3o0ITg6XzOudEGSB
ahd0m7L5HVr7exbvXsCXvjDeDd48AvOReK7KE8hNPTTg++L79rbhObsMuxCsfW9qQLwEy8uMXCLL
SPfzdFlBb9CjgGWnKHdGwzJzTxI7YrWgVar5yPhpPgB+Y6EV8gFXVsA5YxzRsc++5MqFVln2SYHt
CO66ttTNQo0m92cxBgVZF7vE6r4frrbIjRCN+X0Z+4y+mzjz6JdTGEtq5P1LHi+PjGIE5X9vGR1I
5/mNFvAQI3h0GsP4Dl1Cs1+ujVK6a/6zzKatuozL7KWoqEVFAATtS+6Nnuz+GmtkIK51ENZs3+O2
xdsyxU1HkiRG06rHlvriZTYqyOT35jjxTxv6ka08wWT7pGOgZ50ra1a3V5RmriixbJ+hjHYiWxXC
z8EgkrQSibEPNxaBfeXlN0XN39SwJBGfGJ8E94Ch5wQDfyHoBEoUCOzv+cDSMWNGuAsm4IflljcT
8/drr5L4qNEld/cROtFqu11ioliVEnnbS/yye4Dk74CsNcn7Yu/9HNrKeoiLUZ70y8DYo9DlM81D
X0eHWFxLRXXmZ907KXUQfFwG7SOJ070BmGtWGe5pDVYNlMpr/mzY9lvAm/dG0ADjyubD4jDd+nr+
FZpTIr7ZMwcpyoIgPhfzssUIYCZ6dGayEH/ll5U0I+8UH3IoVTQnCymTt0fFQlbpxtVKHO4o2HV4
JEtDe5QW4U0CCyZLmh9UwGCPhu8LZXtYafLF4XopfLszP3UYEuMhayAkNNZw/t0xSzcAu0qPitFj
nMfCEgO/xIfv+Y9fbCIDQ/mucbDB1FUF9n9HZVeMk5N1xnWfdLQp46Ef1DCjSmDuPXDo0bC466iJ
DCYLelkiJlcG0913ZnpS5DfN4BRRTTterKf0bPrijyCXcQLPHj/it/LqqYkAXdXJg+5EH0vBgYK6
9aeDh/uu4qR8600Qj+9/dXfxbxkJqATQP0HV0cq54dkarIja8G6TtokoPeXGFQHNYtnM11khzUb6
VZjxoudk/y/I7cpQnncF2clNgBynuHeF9/9r879IuFlPcDNhG4CibInQDT2xCByxnQej5gvt5LMs
nxeVcklgCXJKQsmZVsueBX7Z5YSuuVCji6IG8pXoovDBZVZhPNdOpy80lnLnfaAJ/SjEXXZZj/ov
4f0paNsxSSe3vb6l/LqqJbXWGtqso5RYmpCcNDysBxzgYd3H1GHVEEC13nPnsxLq34UYuaJwYxky
j22IQbCBRCU+8xqZLK7ChKXcdIrVdwiY7QEE3LZK/RGGWbqGOHCRrgmDTp0BLVganMW7gGqWWlhd
bGn7FfufyG46rUj9S0+0rRMK140iEtzsJ63IOQbPR8/98lQms6CVXZwtXH9VEFuTLvKyxAn8bWxI
I1vKmxdhWTEwQHjQW0VqnwlTSXMGxvGqKvtTqd72CDvEvTWQu0caSQ9A6Jdsmcv9KEuECBtto0/A
mvyGxtx1HZB7Ei140GzKP4D14CshgUCiyo3BuoB0eIs7Jq6B7RC+YuRSaszHNYgoJ8BSx2+qubRz
9bQetVs+UQd1+60XD3MBRKfUS013gwPgEmul8hRNjQhLvVPxaCQ7IioV2C6cdrIO0dwQDIaIYQDn
vLdpipxwIBZiCwBRCPr4VHHOqvbj431QqXVH9UbwxQj1qo9ttHqzfXGK8jlLQrDsLBKAVPV3gUKh
5DJNw+4glu6AQCim/g3j9/dmfBqf4CPklyXb4bDF8RyqC1PCj+uzHb9Jp0pqXXoDaRi0SS6CRQyM
M1aZphEvO3WfSWhGvKYNs/c0POkJosEYv7xSsqFGPPz3itUZikIftS+JqpuMETy9U/pqW7IiAVMA
sdAcm2YeqEEAZyBKBIwzKrIAtOuZWicog899y7TKj8jDBX8lmDjv081/La/sCOn078uAO6KaJhGu
AtbWmm9029RjMU2NS952Rs2AOic09ngGklnVVxtoZRholOcplbR5pX9XocYsdPHJ99LfAbBEB3UA
QXAy1FZ2I2LBnhu3lgyZUVob1OVjyP7A5ppFbVpIigWauprSDIkdUr/+tDE04w02GmJNcV3pkL9n
EDxu2AcOAp2I4K8d2rfeoUsaBl3evXeGSmHSknEC7hRc7L2ql47OFV+oVr+MPZmyqMvvmbRc6Qe8
3s/Vg0/zX1lXdGWU8bcIxWtNxOEmmQec92FDnKEFhzq0HojKro9pV9DMsy2OpY66iYWdW0yaLNct
ZUzFwpZKeSySCpud6TLZ/yUYZRvV3rJQNUW590dvktu9ANxCTwl+ZLc64UOuxwm1ciYD5HzB7/Me
0QSKoSstkQ/Mo0BZiQPmZQh9qD52nrkBUT8eSc3aV9bAoIkSHZOoR7aU6a/2R54PKgQ48C/naf0Y
vtDjZdDJyQBnhD7I/pQDKC56rTGt0dwkedmsT3xzezDM7wO0wPt9J9YIuzkPQWHG001eRpypBCdp
XNaQWZ94TAdCOGQWsWVaETAlqdf6EP/rZTInYjqmYlYsde9aCfUd05I9JzN7pTbsXEFLmQ5UT2n7
oR7rJBmvzkohMd2nf3xSjPrkL0mrdry4hW39F7EzVntxcKX/J2nfzsgs4TLRkJmBXqo6XxEt1oqz
xTCskim5tZj+vVv6mN7jbtLMuvU2/LX5egoLXXuh+LkrRj9puLNhcJeNR2d/o8886ksFbrXgzBNl
8OnotsnDysfqhSIUebBWRtqjDOfgg8bIFkRqIbRI8kIxKpxWX97avrsNzv0vSgemaF88uReZUiba
VzPdLYUj7K+G9z23NKUrlkPf/b9iQ9nO1GTSQtrDZZaB3XnUuzRRbcliGLSUiFZlmwX81u0fU//y
xR0ucfIjiOtm82XR2Lsv40/0xpIie1cswLUDAxJiItbGsSKi/13WpIWP1vQppFZOucoPSPG4Edm7
KvSlii6yTDg0aS2w1r3CLl6OggaCnDI9KpKDG/FcZEeCl0yHhZhyC4viSFLpLzlZvPTq4NSSHp5J
5FsrAzhKNS2cWxx4auWxN1e7kjapq6TtCwqoEJ3qAl9x+UoVR7/zavEmgAnQ+ZPa3zXsgSUKTP3l
VgoYxPSnEpuWjESqp89/Tz7rtwZGl1vzPoTtA4yx9l9TzQXQJii8xmMw53ktHSSTQ78NDkxltAl6
7X0qtpFRJ4AJYaR8ltn1e6SAAAvxLaFz3a0DZrFFoyRUKQ0TFNGFdmilPSg52S3bYhj/3Gr2hTWV
WjJdvu1eANjemUr2/KY9pym38EHmWXNWPdj8UYTptTR44yBuGw+QhkZHdlYh0MAZh4Y0uhKJB6Vm
5ux1YHH/YUzTGXooDM6VoFaJvOBuA41aX1iRAh77mLpt4mrcgoAg8iYMbvlwO9k2qO1lTcg3JkAF
RP66DEPXtcMx/cP8SKcWBhsbePJ16VAKQG18sZ0pp/kN62L7N9Fg8yb9KCVj4/WXaKqxrDQSjQZh
WE+JNl2eujBfNmWCnt3/ETWkGR89Hak2Lv66tOyuTrZGnCyV52jvk7cBCKLIrcdz+VZJtpnkiqsp
QNgK8WEdXXgpZ0qfe81btDiXEjthO8LtqshB3AXhfS7/fhO1QT50rGUoMXeB6+9nWFSiu+VQ3avs
Leq4rq1FrWddzxkIYEehuaAe/3w8OfB8TThIUe1p6bEq3pK1Hi216OvlWLJC/JJo6rnCPU0lVQX0
57SBzMDVZ3WqngsTfWT7vMeiqaWbVU7li2bvb7+EvFuIdnA5HAzpAdi5GReECetVouomdK2+JqHJ
NTRao5/+L5hCWMP4Ofh6PqbDaSmWKSa29GXQqSCuihlXV2lxuZDNRRrRcQTa6O0/JtF/mpgg7vXc
GnesrhYoXFiLW6jmgFSVOX68leB9DZbY2QcSINVhYVTH/DXTyU+ouGZ7+GBrkZ6XAPIJzjNzIIbf
I4anqMAz1FXSG6pfW5D9ctiaKewcMZ0xZ83xZiKhU4ohVoGKwS/BBZraIFhHv6ZEwKpw3zteWEi6
XfGsOfi0efKHIshyhbz9Yps+uziWHvv3gJ+3HSrTvRlZxpi7O0Nn4pWuD+Hjp2BiYbAXcVi6OLzR
tRqdRC9Wvzg3cod8ex4zJefsueSYzDNc6hmpp39onEBK7Q4JltQKhHz+R3sUmuLa0Szn35TgOU8x
n06AooRwawfVySZKZ2CdhKcZfEt43rTt1WSC1v6ICKUF5H7QZ0+PPc6mRVwxGWUlGGhAxNUCUxv0
dtWiXIYQLGyNHGELAlk5GN5nLYyjbOmepZilVxYmp2OAQsmJf5LMUleReLZooQEgMLahqPOaUfwc
DToOpx8Sis6zTE/1nGtY1EBRZVDKWmgliYrlP6IpZobwxGDVU+DnTL3kdSMwwbJykXdJX08x75bl
X2nIIvduZ1iMvvRsGocrWvoRtzevoLhMLQyHVcfR7/b47WTjx6KTHGVTx0kZo+ASj0qqdzM8OG/e
IH9Hb17Kn6yJxnjqojRcZADel017hsS4av6yGKsVAXPIZ+YOoWD0AS3ZSdMgkky1EiFxwh0xMKzm
dapHMzk5mrG5TmLj8nXxqOfIrcleWNSf1APvmOjJhCFHfqmurENIlvT4B4NfFaDnRz4GF5H3h7PH
9w909+MPAft5z7cLLWS28Nyt++zhgZ3OguW6hgBAc5fYoQj3PyekCMet1cJbOHh+zeQu7VTJ0oX7
Ye0eIcgBiYvgn0VQqpaIcUPNwjbOtYZWBNFKcT/nMWCbc2mF9pL1Va3Hr+pjpMeN10osVkyBpkQW
GjLpHYnIWgd8uiOjLlcjmuvxe+6PCoBBPQ3I0ZVeXE9WK0FKo0ApoCwDK3RD8KhrCjMoEnLdKUOM
eyyJHRb9P8kmtC5fJQZM7W9/AbIoppQnxlqqG43kBEBAOP+wIPzPb3lRvZQcUf8NhAOMC7J1PhWk
R1DWYVPMETWoqYaZjS7rKhz/ti7dYi+LPg4BNtN8VW8rXT5FQfKPSjmvI/kDqwASfjN9XYeXlOww
ZguH8XEA3zrlqai0Zvzw8xupFtQK5qfzqDoSAFSFZHr5em8tlvamQW1LeOzDzxsWdB9TlOSGIg19
VJODqCQSe9qQZEXxF8VguoBnVuvztdbs9tgR1NwPrHagKviTGbFg8KAR3BzuPVa2NM52RiLPdqOi
TlHGo5Wx0sXt+gtB/z0IsgpMTdhSao8RNtMLkikZxhxCcdB0YIVkLQpiTSy26xOY8FAl43gzMFV5
zgIbeyN/64O4iZgKa06SofL6ALOCZ/3yRv1mIbML52TQ/LtT+ChuL8io1+0TgoW0uGIEsPgqUChl
aiantjlTh8LE1/l8EdL0Jf1zOJ+AL4RD58WOW66SL8/Pjqae4YJR6N4RDiAuriW8m6geg4Qqx9uy
Ys/9DLUC6mLX0C8uTNLMQbfo14buWqsTmPNeKcCnwBQGL+EElDZ+11Kacb1T6T4OgY9PDbdMdDhV
Ide0qLhTNliIi8nC/wu4Bj5IEa6ES6X42IYGH7/vCtLd1bmSfqyVVJu4uHB7DY3XK9xqNLd6IceU
DuQ0uPz9LfvhfFzYPOjh+m9/xKKQfy6cBBtvJjqOamqzxmwbfsSN4G4DOqIyWB3Gn+1Glh07RDP9
yHV9e+VgKBOF4oPerm17A6uC2QZto8qnUc7Mc1jmBa2juWS19iywFnMH9Gt+iNHxRG0P10CE+GsI
wFV+mPOu/c8hXjZYHty3d85aqhkRRLH9RxsWouwvY5/1F+zFYRh4rxf3x/o/otRg6vxw4eWdE/Et
8RP9jiR5D5QGR1l+LLuaowJDvqgl9XjaJFdziRyYMdBJNDqBRI53P6USfDtNCMZkUmnS1ckyiT5M
Wzv1Y+nt8PU3Rz19zff588eVoeCKN8U5u/xOTcPYwsMVLH0E8FVxV9pmBjhkE1tvAVQyREr69iQY
dwyvUxTe0kWOKBAHA1cD02akgqiQkx8W0mZII4Glgo2ftL/h5ARs9oHMvyauOJ2V3ZcbB7WibNx4
CVHdd1WKA5aqO+XwSncrwX25vNBPOAIGIUscMR3r9ocmABJRrg46B7kdcN6ewXTcjrKhzfqjBtuc
+p4F7o5N/2OcvXuAn/LX1k57ou6+A+UVz7pZ/bp2Ty3rSG5QqtfIlK0/a4mWectzrjkz0zNtf5lD
35mb/nJvb6wn80gW9+KCduQ5XM0Hepeet92EK1MMzoBhXU85xL+FC45K3BuyUCmO3U1crVI8KL7x
3VIm7SjuwIDalMLsWFBGJASiIk78C27ncl/LnuZ3TQiR+OgI7YhJXn9m4beKTqeZb0u/eQq7d9xd
QzA5fB2vn+ybBFKNIH7tYritAxS4IAYnxLjvFjwih+OYvWYfe8iTsGN6GouKJcHWHs+EKDDm3gYk
r1P87L3QRM/D5L0cF/Xaq44tYGXoOQ+mWX/1jILgNUzfq5CS8jDSWde1kXsu2BaFi7tUEUiXyNnx
I55FbIVgQTXoGLGM/70b5t257vZx0Z8FLgW4CTHzZ97jRE5hmo0uqvMdlzqyyzM9HHAhaNzKdv9i
E6xuxwRGcD54i8zfJYSRv0Aakknr31jwIUTNhsHaOSO8SY/WrZ6I14Ag+t0beonNDx3U4rNL+Ey7
eh29P083bu6uQ9Nhq/Ow2Est9T5fWuFmtVDoaA5IpTMlwvvbEr6RuKbcp/PMCzD35hXOTJlVQvZK
+A2Mp0pR2+EupSgBOJEuHAGz8sdEc8sGzwYvBf1YKyY0j7gZT2Qs/PaL0p0Lpd2hfB/feSwMMrwl
in0BmfvP2TRRK4onGug5yEGUbPppRSNq/0mw9xcXg6Ej3HagPlEejUxd/ybqSuEr1NfPshgIz6B+
qQJ6PGnQXJqTEYzE8ZruSO6pFsqvW7B94Y4vXkBxzidjeUANMV+oe9Liabxko/i3vX7y7km9hksD
4pQyjc2MBGU6L+Z3ItON0T0Y+HMbs4nC4DwPbd2rCflNrk5p+vJ8aL71d+coVBRp320ohxkFOXKe
vYKFoish0jQwdd4EZueBO4JPYj2/gjHhE4VN8nYLBNvO/+ZKfQpZcyQnc+ZU0RiT24hNOoBP1JeW
umHPCjk/io6Q06oAlxJVLN1ViSXzP9AoFx+lzvGL8NvGKlj6+3HRzw1mKm7OFRhroMv2jsuU7VPs
dUUhzpn4vTbiGglrmyDo2w5um5XKANBOjE6nWIzt+U8z4hbmjNpi/BH3g9FtFkWfrSbTEtIw7lUM
m8aCWUme6ciXERslGRLFW/NEvvz7joMDhKSJWNS0mLbnCrr3e1jzSAGww18qG+bxTiSKlKBxNdhQ
dDDd6PEVDFdtYRcL3PsaDs+sz5XaY4OZS5mwsPXFChGO8KzNfzjMAHXG9z9r23PHh3LRxxEXIoK1
LAwFo0icf+4NZutcVHUy/dRIXEGIjJ2tJlhzOrBQ3S0oDodIjDjO8UqIv6WLj54fB/zWIX5I7RpM
LAJZOwSlBZPyyt/R/ncR3JBAX4PjjUatRShN81o+yo6w0nuoT8sKB+AvhP3vui4hjBO7x1i743rx
aos4xARjWYlDhiQeTCB1mA9lgW/VZFl1D5fhlAo+QIcniLmKoF1QO/QEMa8EaG324mgAHsnP2KkN
BrJheA7oBioD/Wg95L5p8hdTdvMG2KWxvSz/GUjMDDb4Qh5Waa9RX9M5G4McFXasY93gMZcKcOxP
QL23hwnLLTyVzd6dUMPjPBMWwBPZ9QZkyNTBW5GkdUdfN9qFukSSbjoCW647iOHedA21p5JHWpTN
boHfm1fnG3hPdHe9EnB32o6/S46U3L/tAAyLwODIwL5kUYmRGwJqLulYQxw6fOw+n559KWIYftwM
zMdaf+7GANx0F1q5+2MysFDO+BD32zd1A2Qkg4ph+MA0VJu54/B0oPb6bbnCV3csfWL/XuVQwK5W
AHmnq/R1MsvdHrGrYSL+C32BGNozZfiNEGOSqWo9MjN7VoJ+lPadsXvGcYX5C/YzyMHFDf9bB4Jh
cDKpqaqrwU9wfd0Oy5t3R4vGVIqR4aAdy1gAER0Dx073/3k4rUk2biUSoj8/iQfpNaqCEduciYEa
WlyriHVtUTNs4HRnhIp82+TxYRhverr3vHQqqeT4NX7rfrTq6hKf4hmPQes01GVp7dyUV9jS7XBm
QReI4C9gGb3byrpBNiW1UeQyjsICNMJWj9UwqYdCTEUO0OXFrJjBEX75Rp0JLg/OS+c+lLo3Thlb
9UyM+oR6gf+RS7eLfudvcuqjRol9QJgFYrY/dvRbemb7Su5HFRfWyQWXa8ZAkxc7ryeRyEl2di5R
PujQd8kRVejKHJB5X6UAsN6Glff3qQiEkbYopVVmCVvxWEd4bsdhx3iemCofhDOGp1h9HzZz+VXN
jYoJtauZmC37k2ivse8GdYhtFX+cnmF4Vr9fK9K5+7AAByM9OoZufvG1YaU4SRPruMERXdqV4FP5
PgVn2X2DChiCiyqdf4ont3+PrDLuNsMvCGJTnnvAvsYQ1AtOol3IGvxVFShscwvMb+HVSd4UUHON
LU+X7Xluo3dHeaN2AV0IWRtpPV68/UX4GXf/eX6VRaexqiP3z0A6moSRlUCjTjpGMpHzcnTSxeKb
ScuRr6cvcTEcfZBIWZmXLgimAjJtTYaz1kwvzpV5vAltaw4lC96sj8rBHGr7jYYXBDZD4/DcUVCq
9I3O6uwg03YW5iW/aQkiClWM22bIvZFh3pPeRooOJiTnR0z3+VVVi/JNrfo5E8Hqs79r+vyczn0S
6r7r0dfu5nDsjgmktfbELdp7ya2YCcK/FvaJtu7sKQzRtejgv94qZklONdO3OuefZ1rb8n2HaKn/
Wt44PWapXD1DQBW3kZFAsedpuZU490ynVXSpRtRrRiPLjGOIaVKoP7uCALD+PQXYr8y32K2RDpGI
BfY4FqfC85/yPfe0v0G1anROwueQfO0MA1oOLspDBwcZ3HMyPx/Em4BCdHNWdEuAeG4H0qqqR/Vq
h1XElTpzkS/usfSLe6FK1dmY4rMhnOnfN04bJwoYM8bgJJwK9PDovXMuzStQdthrqJaujK0n3JTo
Tup0pZeiHI/SWuXXlAxQ5Dx5S0LD71w8HWecbpwU6X1WhJpmXCV2qx7StZqmtuilm0ME5L1aEHx0
dJTGHZKsQWmm+zYBNziM6/GamOFrSGN6vwbKrq1sYr+iIF6JUAnFgr5YI2aQjFuOEOVeIX7rSLSU
u51y44T2CCJ473Tn9dVYj3P4VQlJvA5XAgW0aPe5T37TbMjEwpow5N+vLQistrNvvkmYXWfu9G7X
ijizJ9/URCxkMUTNINaM/1ZCjppgJox9+R+BCDraiYvNUHGGsP0O2OcdHg+bcg8lgu0cEshH9+5p
iFxA0ME/WAIHBzOoBRGzrpPAiR2qDi27WUX2iNGxH3zie5/6LuZOP/hNbvyef3J4fCc8R+YDnQIY
wul3QLbA+CkdV89rGLpBYqF9tNQKMoijvzgygPrnYRL4vxfkcEe5xEXAOnP9KGNVn+JOYguAz8Lv
hBbq4Mfxh5Iki22RnUa7GsdPqorcPYV6qWCUxvOtY/HRIBR2gv1EoBm+HZN0LBFI1/dnF9KL6zVm
v4FC7FAHktrDohYN467Ex+KWKlh8GsznDt+jDN0bS5CEb0RhTjyLc3oII7sr50y6UP/Styoxb9vo
HETzWYS73yAzTF+OIa9Tt5Q7UwWz/C2V8zxQLvzZwoHL9rPHmciz0P95v/NsBKU7nAT6ptddYoxg
J0WWcNW2LJxYWZyk0BldBwwhCXRFip14qz8wdBK9p3rhHgCLHPN5rcDe+Ui5fwgY53Gej+c53HAV
5h2AWWi/JjVDg1TpghyVWEmkRzViMgSkdnzVQwS8VlugsVA2Mbjnfw/JFKSkHbE8gVPHWXlnV1eW
oAODVY+DWS0pyrNLlwSz4H5/lzcYNUWc0iMXLsIqC0zrV0iPSavGrVshx3d3eAdAcwkdermvsLSa
PqUFISNBfNYEgGHdgrZqTbHlDFCzYGkN3Askxb6b1fRf/ALLsUkOVLXGbVigWpI1+glQAF1TwdgN
7k7F7uJ0oJYcw0t0aKn1nfMdDLRuBboqPXIIv/6DdT0ojQvYoRu3MScBe2hxPvnEq5c6u9d2Q6YL
ZS4DYgm8LXWOVKh9g71+6chFUNAkKEcnHBILkQAXwZEnH+TNbxJGxntILU10e5sr8Q9M/k1VfPac
lNP+pYOCY2N1+U2qOhbK4AUaHCRHTw6Pl0YqhJJM59gexyZlNmSC9xaL7PBoed/rGGY9Fvww12zs
P3kRVF2CqIkTBoDzyNyNwM5XcQuJBA5/rXotjddyUMqLUUpk1gYVBdp8ShiD85p1amb1kobJA2N6
EDnIc/A3e5UAM+ESF2Xbl06UXstRH9DUYUnBaEdFfzhGmOZhBZA6j7X6HEYVJ7KSBGtmuoS+5zHJ
vl3EGKdUXcWdU9n2FVl469wV63Mdkc97J0pj/U3ktUO5GsVhCDLWjqliBAXOXxcWzYvSTgexQSGM
jtHPsMY8ParNunENVmNceIIhmFdJkhB/4lmFvcqaJjlvDzFfoFGXWisx1eLYMXJQcseRiAKSNFug
WkONa/g5uDk8kfbydQ54dxg+0i664LxefZCa0/bgxT2u/tKvXIZtuueKXFbZbFH4gc0Z4Ts/KTTL
rqix1hdhpao6hY7tmSj78iCShT92nbXpcpLFkqIWXarJrHQ4Ppt3AzXaIPhaydFAEk31Drz0zdea
/Q63JTBCZx5n8xk9UH+9uGsKHb1gXMheGZeYr07KgtjWhzbAYz9ZBPT9ribTlNbbchqVjvpKH/rp
zZtjkkFb5ojkfjW3++9lLQ81Z1VzpcXEqbkozK4L6ydfq8fE2+MnLWmsDFXHNM3sU1HdKez7y5uX
CwoXX9OJs/8GUe5Ey0YgG+qTNcmj8YYbOJHz66I+dJMExSLzR2SAjhUuTxoLlqj0eD1Jfwk+azVH
8Ic4pJ7ngpSC9FDhjkm0g2i5u67QxNQdmfTXlSU+UT56YOINIgrGfrv1Y5qW4LtWtAYMYb4R/kUt
X1BDT9FnAlPY7ucunt7vvjlhlldqZ5gU95+hERKDq24TFEHPwhoZ8s14lhJU2oqcW1fl/CG1D/7D
j/yec+36fHKV3fI7uThUk5fVXZDJRpiLkji8lNfcdjTgtSjxsao7RZoDbgzBUHJnopw0i4Ig4RTI
Wuo79PdbPyC74Fq7khg46WwFTwwNlhW2SRGxroLoGLsgs7i1YCT6oP4e5WuUywnD0Xei0M4jEbJU
Tea6xI2jOk4dA6LfBaVpYb7aM/r//ptkGHeCK+E1Tuo9uZNLgwJNUwCNqTim0TdS8IxYwYRez2NH
QToL7ytWIdO0So9cm1W7uT7auCNRH+xg1Bin0Lzd5IPdmqqlekgm8TDv50bSz4y0f8IJVFsmWvwJ
4ER7nancV9phtgx2Kpl8y6PyPBJjqJ5/hi/LHpbC9FHcFyV8p1lQv9It9GT6cHogTfk+waDV1itc
7YUhM32yAqLmGJAVRaz5d88xEeC3KE+OYcDVK6c8l759ftZuj4IRy7+gn9pvhuoqNgxCgMjNNf7V
iFBD1u6b/U0mrGmZv4NlOO9vCSGFrlKI0yeX92mPV67+KfvQKu9Hy1/EQhvPPs99c+4L7VBV24d1
zFFP8cZzeNtT/DceNG7lJtCRkSXwnA4TnFs+HXgtmywDbwymeFRaceebd3jv/urbp5F2xsfFbDdt
LVpoU+LlyUWEetl59W0dkFWM4bzy0TQ3g1ZMPuLjtZrYoNRy/qFV0QH+JJK7UW+lQ2RsDOCHbJPO
Od5SGh7zEnICqumiqCmj7qrRculoSV6eHP6UQI9v3bRSEZnZ33gb2DUFMQVKCcEMbSzfY/eJUCuP
H6kNjLXze/k33NXDJrsP0UGLUGP10sKQKxDACPl9CVSLUuozR56huEEoZ8dgRJL8vTLjD5e6uaed
oXqsi3UFDojf98gblmH3bZvxgPEZNhAFxNHnB/h8kuapvmz20u7P/oN2ABAmXSNCgo2zKECoItfr
+z7Qmx+B+ykaIqs0yCHaSxa4PChds3AMf+hd33XK7R2qDRjenuAMPBVnH0GSYbYrG7eeUoUlWOLl
aySjn9GqJX7T/+Y/ouSX9a1DKBtyhSfDRmjfn9GKd9qXhTu3EkZfAkn5XKeA9N3sq0OdJG8wJJfW
h/dANWbmHOYWLLJ2Vw77vpC+771l1s3hd6ctRujeIUlAB9iU0U6Qf13SAU5WfP17NmIlpZqAorPY
LrvqrtFKhg/jDdCMeJrMOiceJMdBX3uQ/m++mj08w7LDVqa8jRRN6eB1h4QhfpI/jzPO/jAw5cdn
YDECoL94QzOEIBM1hd9Nc0xE8iiV9wUnocypklpxtWrhRhvvD2AEFaMQW434sDgWy3DbzwFGMfbd
lqRG8SZZ7WgxFHXScsG2QIiJfi21pBPiGIQTHOgUaUUORV2l2kIoqeLELnf9KJHhYNA0UrRS25Rq
kHQ2ZEkW5NYfsQ5VH18PzNWxhbH5dVpjpL1jmoe7OUnBN97m8wB2MFrmqUGdgZEB9lf0Nt1MgtPS
k4lbgALkWFtWbWTvDN9AYG7Y/BnFrxIA9aiNkXX036A3816qB41UIGGvgNQm+wREMsu0fCXXpbXh
TFsSqjKTfcVzi/5AFzaB9EwRRe+l4m5ozJqV6Uonme2NcTQAO72FuSxK3z+nLW7LEN2+4ZQw9wmC
AtWRcRMMM+A4R5rtW3j7lpAQszl48Y+DDme1+tFScWtZjG5/SAFra8oSKGWDwwXTy1J8p6ytRUeT
YAAIPSz5j1FzEBi0PTA/+4uxvrHear2v7krlFpA+H+ujGXy5NETGSAMCAbtmT5z6x5hL+N62/j5u
n81d+w8kNuP2e4DGTcRkV7vf9K8a4aP5c8soE19FiRN9jM/c0G/74twYEpOsi3L3wyqgfR8dXdCo
QSHIjN/e3/BClMXZ9m7ZYe3DJh+j+LL9UK7P7SADIYo4NoaKVMhuPLGcRdJ7pDRpfEtWy5QpSqsj
dI968PxHEiYNfRGuoK6Zb6Z7PkuEU0CsbpcfPj7We7Q75Cbn4p54zVSH35FuDi6E6C5qGqR6Q1k2
7s/5nMa3Dfe4Yj+Cys6q1/L7Ew4bSrWqyMTGaoFQ44akCd925HsWOXiS5J5GIBLILk5JoS3EFpbv
LgluAOfDpjCZFtw/KA+OWXchZGxVUmXXLmof7JdL5ZqLqP1kbnIkr1nC3pe4w9Ic2DJMumZFArte
AGXfGKk3EEJS4HBqk2mHYK6ATkkKAr0kzrCGDrTbSnPMQDlUXiDpEtQUXAcuO1g2tfkVSIDEo+Cq
rDFJjYbC7h7R5RmnsR30BzRDGN0WO0wPnSWah+STUTQ5Kfa+kVLqhjf3lFPdn5tVYmtKM6X3edaZ
OvjWqBUKa2Lls+SzK/0MvbRLK1yApNORnZy7PaKQeGbnUOTs+PG5NPsYlptsNhLL5apmdd8eQGC8
8UhMPN3nsutZtprISlDip7rrAXuCPN8ekSdlHgvKx/oHxKuYd01FMJjltrTE+2KH5KNY0dy9Ue+c
2DRiUVacWrL0c/egcsP9M1+4DXI/Ckom9z71BB+/RKyyg/y8ZkI63wKZZr9XBzJxXQUwWTYZYbuY
N32PYjpaMDpUt/d1cVlCz7PXQR10wzfaGPqkj+4Byka3rv9wJlm9Ru6yXwWRNxVe+gj91DjnxkpX
oQ6lbeNxnxE/psEvJ10CJX4dXnSvIytfF5SszUPIXRdewAd2BAsKfUbdg+C2zWMW/lgrarXjRqP+
XsANLj0uDutjCDe9K+Y90mAc4CwjnwnihLWnSilr8bi6xyKt2wxVhruJj1qflnZjAUFRxihuJO42
iAaBchTRe80HjGeixfE51NGZCgBVzxIzr8wI9SFflmzoGC8hUZ+Blk+3/ze1ugxniLhyEoKsu6Pg
gEWSpMuuDyT4VJO/VHdqw5DDEqfTxb1KGtVlQtys8Ku8M0nqxAGuZT4zWE1elGwmSJz0COMI8Iuz
u+bAL2wjagB0uJf8HWWtk8KKwMjXme4lbAvPk9fbV9sscJxhiIa9Pp7FSLlj+1cNIdwHUYKGCJky
0cCoaWaiJWxr52zuetl34tVCKqjahyRL3ygDAQ0qdBx22O7BRnSS/EsZiWellsIC4Z21PzBJ7aWB
MO77oNQfclhlzSc/jKG7J5q+uRxhLsdOlUC7H2i8py+THIGd112yFhFkAEWzAxuoSNgFhc5kXdcX
q0CaMmPWoThQtS0L0LuxGHsTOPHpe9dw93ikzgzRe2cSQXarIRdPi/ibeSsirY8YvcMDOPI15xOh
gwv991dUnY8kZ8H5RSh++feFzubl6f+hcq5ew2SdVI+4gaSc0mmBC5/iXN8ojQFqwdSl8I8M1sez
oOi9Au9kcTCwxZq3rodNyM7mMxFMP/gvmAKV2tE6yKKBT4S0AMb7LZPLRZsETjO5easjv1KJqHnc
hvqj4I3jzJQ33C2lw9NjKYlpJENVtRlMxSkw1btKhyVvUW6ffBc6KHkJtLgzbCtgOSBqIuyk9h9R
KKkXr0nWyGHHFNEM8knDTtuYaEImYeumnA73i7Y+0cMgZGT7mL0Iz65oi3ehNFPe/wO3Ezb8Cg/j
b0BOPUzn5PfKK+eYHFRgNjg6BJXUk7ccjo/1+ZYuyicscTPZZxDpoVcM1NZ4dEafa51yJqXgQU9C
HMnjyuAQ4gdQ0+sFPZTImTQ/ta1RERU/bZpCoUM4QLU/xgbTZ/nfgfwb0GcIv5JyUuglyyxoPxEu
t3NdqB05Uu5lexCx1YVHapaLaYZxfehOV+aktRVQ4eZeWmgoMCoaZiU/bELMyv7rh/VAC7F2Ji/p
UHna261q3+XfWuNz0E3PNPfBv8xOhbvXqlaEYwaP02m+o5faXE69I0pe7GQjSZxX7UMyuge21M9A
ZU0olKDbJnZcm3+T2MeKytkCYcF4yeccnEm2cipb4InS8mdA5DSsPIRsYrLhItxU1wSYs2yyjl5J
aZWorNLljHyzm2L8fxv0LBI/jPt7KzoXla8GIKLiZeeweW56i3RthWhDyXT7pa3sVz5P+s24+Jb8
6lgrarToWGes2H5tw3cA+zUTpHwgUK4DDjcrKr35umO7a7QEmh3dLQtzJJNOYSu/WPWWLxksyMFX
zKh7K7bcSaJpK6sysM7gU7rw8YLeFUNXK6qmVk8bgdeCjq3OXrI9UtsCiIzuRIldnPAwLRk8nSCr
TNN5W6DF5ihto91cFYBu76AkCC3AbkpRc+GIzFc3zEthUknJYxRVQzAml8k5PTaeIt6d5QabnKHW
Vo63XPgMcCuJ7J0cUeal35EnQwc0iB4oozD1VDRFOurn1A20Yv+CDWj/OmMRya7rgv4HQ+YFN6b4
VIfpQZVdUlphP160kKIYGvznCRkWzII5WuDCnGxz2R6mwKx6UaCNrC+ceNpWk+6oBAckIK4w3jlr
yPQnLKrKj4PybAeHhRhEwHu9DkuJpE2c4q8sSAHUxdz4BTKlG6pZPlJ4gwX44E1H8ljr/vcNSGNR
XPpZEqrL9YMVifonu5e272XzHrklM9tGGU8f5TvdHkdIISKAFRz1t49BYsJJDpUFFgdXpwfQXLWc
lyNfr7D+xLJdzbz4z3+npclTLmUB0XaWt4HHIVqOTl+6kXrx5gAzI2LogSkFC+N+WJ7MHexwGSbM
kQEl3sXuoT4+aUbqternPD1Lz+ZpZHFCFmP9RrBZYmr2YIj2lmhMUR38nsaD+50Iuwom3CQXziLu
UwqNw2ggsyYOxjFNMRK1SMaTfdGJeYzuRn/Gmt/DFx6e3jkJc3oqfA/UZ/IxxfliwlTVTt8O8Zgz
IdUlRKU9VY7GeJDXQhkHcohOrmKgt6Qtz7TDnZdBLNwA+Fq5A/+T/rL2OPIRxylrzpgbvcw+W+1x
wpnbkZi7VLalBsvJjQpC/4e5oA0h+k5N32IgViOLA3zYs4/+qKYMjdViIIxg/rOWSS2kR6UdJgr3
LOtwOQf6+TS8T7YsSU12Pyt6Sjy7y0vPJyiAekMmu3F7rbiNaYvPknZk3kZslcjgAcLTk3RfLwfk
mi9hlzQRqi6C9VvT/YT3WzmvYWCvDppH44PGgGMgrSgkFJN/QvsxfpVTSwKjDSWpE7aw8wwEikC5
NojAR2BJzJlBgR8KR8tyexodsLiCknAN7tds7ANvsuD/uz5JROFMmjbUrA0E+0GQgrG/7erTAl/V
3jDtweMw6rAxuTuqucbP8abEUXKMYT+BXFQXmyxqHKbKgIXezmjk574gwjlJJnW7SHYURvEpz3lb
5TT/ZzsmpUiv5URdwEMVnugflb2ZoxHiEAUrBKx9paYl7v0yKeB1s+2DrhWoqK47mBmhkqpJYkA7
51Fj7aRtLj5AcnTY+y7bF4/1eB19N6w4s6cT3KmCPtXwWvzMYlrN+HOJGCxZNW+CqTckX98Gr7Au
wk9Ll2xhMfZo2DqstTSqVm2YdJv8K/lNANkvaU6DPkz+rMGjRZAg9FYuOQQ76PEUWBlXL6yWvY7R
7WUBB6TWL4TCgehsg9zn+B6FlRfuCYP+B0VAy42f+mKpr8mgrI46ZA2ygzlSKDp+yXqrdh3ByQWi
0K4hPYG1yyHfbBBko6DXh+v+YKwnPhOw8UC/WeidO7XDZg+aiwjXS3qmxK0mATpM142AvBcrKueN
CvPGpvvqApAVZpJI6Y4/UGS3tnlhcqd4IG4P5C+Sdt90Egescg5r9Si0J1MooQMdo/JRIhBqmaCX
hL9PpbjlwNQtrNkWZn3m844GeBRfEvCDaZ78RhnfhrUO+Gsldj5+dPztCrH8vO1j5Tb8YubocGLB
o9sExnpHK3V0faCZCXvYgWSORt8W6BeWeWy+gbKzTweuhsUPk22O5u3pQiE4BWrvaai2/9OpOyxO
ZUliGZVk7OpDGB/hQpJspnPhc2Ues1FBn1Ues36SyVINmT5eJXvzUlmDc0nucPwe+mljqO3IPBFY
Wcg88azSXRNPYH15CGFY6Vak5xWDOzNOaa/k0NG7/g+HBzHmzA6SgANqxqcB+FEf+SWSX05ncUZg
qMo+vhAW28NkAqwG9iCy5WX2jz/q+MzVhNn6qeG3pzURrMfewClruxr1OLG2e+PVvdSBLakEH8BN
5crurw1ggXnPee6JgnExl38Tw50Eny48xYX5I33hLpw4CKOkcChvEzDqHwdxAm6VXyh2zZNTPbZd
Mg8lguIr/0PJ2h3LPCc3r5vfstOuJ3LLWfcZyKWjOs8RHuVY4LlLaYyg1MD9JSdLHmYbWso5O8vk
AyOFUh50GDqNvhDE7cizoj8cYU8sPlY6YH0horPK01599ZM4YAymQOlzeWEUIvxA7Zy4lfRePu8v
Tg1CfwfWX21jttEzmqdKVZPDwf41vMT40nyNYbO24QSz3A7+PYDNcUnujczY78II3UgN+nny1pIP
mh/XRPPBl6y8taMZ5LgX2k9wq7buQeD+T9ZOvfhl0oNx4VrkDL0jBjaUrlzS2gljKzN5EoklyerW
CSAFNhDMQB9p0ZiA9nawTX4u6uXtF7d6Ztt9nv35TBRJ1miRs6Tz3NN9MjTLQp5+14DA0SqMSqze
ETIovzYRaStBcPlvILOx0uufgQIED2U8+kYMrpjhmmMXAtfN0UQpT344BU+WT18CygCy1V9J5FCy
Bcihxwh8F8BHsbgXr3RUT3u1UU/QYR4VhKje4vwJ0645blx8tZhYomBGg7cjeLJ0qmPxuDld5Fud
/92trNrBsJdnws+S3460hYthnAjLu4WV7Fhg9riY3tjzCTo4k2IrAr5+HrOuA1P7Z4gIN468/mte
iENuWS3uuiEecewI3iYYHT19l9+v+ppWaiK8qUzxz1lMHdEKGlCooUO4xW2SwX+Zh2R1NJY7XlZG
Y4Ua8qhQMP1fVmzEFyApVKFYX0wPY2Rzkgy4+5Dd/8wkrqZ/dU/0q/VfHx81rvfPcUVdijEFL6Tb
t9XA15gixqyN3+d/fQZ1RZ5pNbu0YaVKOFTmyA5P1zDMmQ4YQK40ywneV17KzdCRefctTRcPSEgT
e05BkoIjRgUheihofi6ojSa7kA+QApyFcqfzU7ZQdptA3CFE6QNzEXPuZRsXAwdk66uEPV/XYqwY
mivS0CfKeXrmBN6QMz4+iov9uMUkCB8Xy0eUfCp72lQ78SeXW8zC8Fc8KziC7SzW7PknRM4IPsvI
nwawl3kbOcdSG1N0e2T696p3LSdI74dSHJWMkyTkIXNikm3EgC8pETWk221LS6bInTFRv+wiobwo
qOG1x0chefO6c0XoLZuu06MTyHFVAfyHik88ewID4tpidREhlS+kxW6F0Q1JH9L2CAvXr6v3GkmB
MNpi0bJemWDqVXfPF8Qp12OWmYfJilo68S5bnFosiv/ehMmWLuSJ4syFyUUh41BFi3j3AX8KwuDZ
vs8Z4iBVmQceRsOwIxja+lUwkhlAR4mh6VuIrc4ydLCv4zkFa3jE9Fcph2Pj4lcFyRcUwlFC1EW0
lnT4K4/KTtajExazEw3z0U20eirOXGyWQ6nA7eghf29KA3i8DeAeZGV241v//wAyKsG1PA0nC6qf
Fy8q7ZJHIRdCVcCQTtGh/5hcXf8jNmXEIJxzWvgc4qDzkWk+EzzC0aJmPFfkwy42lgVQS0/4OS50
t+aCITsNs4bun8wI8xgUlaKfxqaSvERbzNUwMc/st+XnFcKyFUuEFEfJMcNXMJGluVTTHY9pIGEm
z2twM46LoeFmdca0eDGzOQsCA1yuZl5Pn+hlt6HnP2EhzEPw7yY7qaMTkOWvtDvtvT/7Tm17xCJB
spgyuhaI6aBfhZk2sWOmr5ISSbafCtiK9Wg07jfQTgbETNcYvm5G93TR62KFvu0uUU6Wnxt4gWcS
QsWSLgtrc/Jyb4e3NRePibz4pU6egXAzJbt11WKfZ2WgWzXMBckXswT3/mqqzTRvf+iewVDchaIN
mCUbTCs8Kk1w1tNQBrndf3fBKiKctoUZHmuDP9T/EJjQmzzTKGmqtrzk7QjKZ12oZf/PcKvjeyQV
3ZEjYV8SB5KwbTuXEvKABLl5XThV5cZoqPSj7HHwJYR1fIpn0SCEz3pw3K81EmOvx7cMoOCPfasA
wT4PC/MZf+jYNpS3Vjc/pMMqJYdyJeKz3wyvlAzRyzrR9//1AB8rYZpomrZFUAvZyRO+UXT8J/qI
/cc8NftYWzf5E2r2ELm5IEiqJeX0Dcdm87p47A8MKQ86DcxWZMovCGDjx83T7ES6sAmPr4twp/sL
1PBb1UIdxSYkGV9AlFVR4A50jRfvOXQw0i/n4b8q/6TgTRnAkoziKZgvn57iK9DVNrkGg5X2QxMJ
QdBEr0q1fgN1jVYS/IwVgdv/BOoGiSWkJvHegE7bcCPN17JzFc3r3XNGrhkdyFHMRWdcOP69jDQ1
l8lI7yzXuN85vTXAhzQswJnQWFHn0P39hK4a2vYyTjiiz/j4ouGUXIjH9DtYzAMYxOI3vGKDDaI3
C6B4GCwZicUHL0kZGssYw3xzm16P/mWRMTS1hH0bWHInqc548Z7AqpSrnUrN4PGEc34365eQ79ng
aC1ksHWTOdK5jstAIQ5xjggxwqIhqVYMKv0Wh81A2WtX26/gJYBku3IRviiB/fNZ3iCqQpVblzA9
BTeB4TjFSfCqbwwbgFl63vVSEw2JKy1rQMwbfHGOeRoxOuW+hebeuPfyoJRHJ+KFz4YXCWhEv+Zo
sonTue4XxUE77vqjmW3KF1JsVaJRl0S8nqwiGQwScD8sjm0J1J9UDUqqvHNdTImWvhp63xmoerFa
mM/IyyNFuHjWhSoQ3+QlShqpeDNhkXksTJ3EkKXErYCS9SnxIRWZH4AkyJWMSFPxP1c86T9EO6Rh
hxlrffbptLgO/w7iBUjw9TLIW+Mt60fKhUw4BM8qRvXrKvgcfc7fFZH0xho8CXvEXzEsQCiAlSen
a4qs/W1x65B0S5AuHZ7gUWZzDJ730H9WlNDcoQFtHTt/6wQZhPF9hQuy9KpMYRG0ocziagJ1npSc
JRMPeiNS2+nJraQDw/BgbqlvninpldGyK8B7wcjK5Nx2CPs4RVteO8IhViHUPHhdy/2kB3v05Y3d
qQ2FiLFAWif577O3jZKYhbFUP4+uK6a5AwayQ27bKVjFGCqfKD46rRSKDw6pTB43yZkZdA7zo5E4
sZNf0pG+nbUXIOPXpmIAJGG1eaNoCEv44bKAEtV9omZsFfxmnYqfBwyJsZKFmIiRalltdp2KOVsR
zQt8qxuKIw6KOBx5P4fKC2g04vDEzn/OLN7qxEJsq5okMDpZE70057l6LVJ1f91BN/0P2J+9VAk1
evDVtx5j6nNPo0V34eg6IL0KBdgoSlJQgO8D6nUZejSViwvsW8nU82e0lNKjsqeD+w20fUJSHR75
VpA5hjDa+kR20ZXW21eF38jBNvgEcsD6RWpQkosO/pdw8IBoMqJcgjG3M3PZtdhHFIdRu0xi7Hod
6mS2KhHAeQm/XaXIAnJ8Pd7XJp/8R0UgBKmdxdyd5OrGgkP4PFHEhgXfO5P8245U1aOqCUoNF1K+
SgnpJQyE10NDPM6mvFE3h5O5/FyLVrsyjJqA0XPpOmwBV8W/iJf4rhY9hHs/2lpNdinKyxSE/ca/
1dMQZWQeHOembHPDihbBnv+nqMBlsTHZAK8+VgeVCwPJeo9SR1uNL+J/e7ams/Thc7jCW/P5SScX
O0kjqrptF1bMhByWit2yrr+NG19Ktqx5OZhgRgWIzhOuGiPZwHAV8drZ+7hCSTD8+2dLzZJdF3SZ
U2lU2DbbWquj+Fu+3C1yeiXPP20KXzas55Oh68J3/NWcV27TKGAjPJ/jvF9q9qERzYoCox2mPN30
JYqi6+Ps9iJgUrlKPDaHFBEJ7PKA4wwlcYPJv3KPphpznJ8D8KQDHhJfYFkiyv1ShLKifVoEzilF
+EV0RYqxvcqKHukpr08ytPu/dPUp53pla9mUuStWXmlBhj49LnUOFBG68Nxto3jEQFWJiJfcE5Fv
B4kIN2qkg7L3LCDG9nk2q01Wjm6TtWPS7KZQiGU1yrqfrIOx+yiQBJ5wC59FxA7CfMXe6KsgTVBj
1EzNWg4sxc4JnFnzEf1Lc78Fw04sFMVSJv12ICqSatGZqjgvJ97sRPTX73v2qUaXsWe6xJEw8Cuf
0AbTN0btxxAYkdf2lEAVnlEtSC5AT4PzVNNvG5a7qut3jkjeJlBdcZPISrgnh89gpcYrJzzbTuHa
viNZwb+2wLYgDLaRWq0kAP44qU0dfgnOVXVeclt5gwcguNeWO25XZIF8StVmwaw7sOWWfyToBtqS
25z0jJY8r4Gozs1s3Li4W6+Hg+GPyNT1piIhOqXLDLhxnfjNPgqsMfDw4hnpB7J/ZrvjbSFW37w/
PPgbkSPoQmNzzYEy5/1QCBO9Peqf8AZG6aeaDoAGpSW6VxhtXWgeRul4hKNuDNG9Ysycq3SzU7pS
O1fUMIK4boqXnjF+9lnxnDnISf0bYdsdkf6/1wmBF/7ViLch4jdHTaxN3K+mPo+/xMpRbLCRNTmV
Sv+n081aWcPRXN8uPtjOh/upjNJE7w+KoQBTvGzPbteRGAM4dLIGkxN3YC0jK5b7zL7E1X37etV2
rIm1AfAFYrqqUspVmbtl970ej7lL14quqqnbCwaCjqRga1OIonUQwo2Yd2NI53DX3aYMyX/ZwbUC
6s+bcqTrw+8hYSauFQR44QFo/etXr6N/Ua7oGX3uG0AUJHK0yJ3dZEvPfIy2sIdUN03DxmFFil20
mcY0jodpymn5axOswVsVI/+0z9aIEC3/OIKB76nI5QmQKGn8cuovL+sovBKx3UjlyrupXFKPtXwr
iTwajTbV1QQ2iyiBX4dZD7CKNsrFo+L85avN05E7IxQK0ej1W9JjMfdc1UZ5d4011qtnlA5sFcgH
IOOL+MJPzCCoCzl9kmL0rXLmViAmENy8V1EaQPScC7a6tFRPSSAMp398izjmxr1W8jhrEOHS6956
Ngh5GsgT+l0OnqA+fDGxYTtayCOwPkLKnfar9TIgdbSecYavBmCPUUOADucEvoCg4A5t9qj54i7e
o+fSuZMkWrSTOYjxK7jxVddr/TbkCopGsStAok3aEK3MJLzv7U0kYmYPCACGC4H2nSkQAxhOTEQb
yx2d9hNumNoDAI7lK8cjOB9+32BlFLElwPT9Fhxjw79e5W2XotDJa7mqSmFefqEaD6XJGkv/5oh3
UWGZW0fAVgD6CcfgxxMXGtbcqyRKYUCGaOSxVP+Tpb1huuKVk/4+H2K6drqNIqwEf/sy9/2OiINy
Lk4tc9UyjeH4xGuFIJh83YcAaq5s/Ff0/wI6ICrtZWqXJxTF9tfD9NuPE+cfcXvStMpDZD2S+x1S
9jkfcLngEtd86wUvGuwIK/R9pxS06aj6y6+VHBBcMIRUitZI6q5dD3yp5Hw2/zelB1zmOf0IcmUO
5FPgkuVbz7zfvZ1VHs1tQeUYO4Gkw09bWM4odQVI3XSafrATxg6Ur+ceg/GX4m3eA0ITyZeSpZtX
ssIaIt3of96udxh/0AQgJnOFEB2Tn8iaavZN2peX3LK+cPv8bx/+uT1DRipW8wLdwb+dXKAgcqE3
xXLtz99HXLwiBR6rqipLMO0be35djlPZdQPMxLwlJhiZj0ULnMHXkQ6iywtJIF7SA0JlL8MhiHkc
jHWPlf2uTpgUDGsVDaWnu4GN1D7mrghgSYYyZZVm5EMFV02GpB4VLkKRIYJOwQR7vfRO1qJ+exnv
3HsYeD8sb6fdOlnlH/oI/XFUOHHbRvJWh+3RscZyKviRB0CBVD1S2EGlFjs6wQhpORb7LJCgsSMd
98v3R+Tbona/YH7K/uatyx+UKD1OHrvV+XxiDXs8ydI5Fap9OGmccREc+QqvkHa+cFpauVsqBu8w
y8pwpXWM+rvv2DY4V3EgcmFZe4tmSvpz4hLy5NtZzhilTEL4J3w32464kQos573fTS7aWPw1O4D0
XEH18ItpKwQBeTcpsU2em0wbZNAwPvfv/GdLRQ4lgTfHGrwFvsjA1YI80jyu2JR+MG+ARvXYoBsZ
e53JaC4DHLL6CRrI3csSdVpa8BtUuCK+2PNPwZ9cE5epnRYwBO2ffMF+rl+uv4OUFnj4qr1I1p8y
FcGB94XdB+w7d7HzK4WmbLUMUp6lUpokr07Mj1Nz2+kF5HdKCLmzg7XMXOrPfssafHOxWCffuveH
GDLTaq/zxFefvyUC4EZ5Uxhrp2yg9pJw0U8dhOeElY4hNJkjZwf7+AArT+ddnqvSIMDhuNpXe1/c
z88O7CPjjZzu5gs6u25xHmfKoy8WSErsXqt+zNYJ4D6w3Q1aHLirDkhewCEHIq2Vr51umoySrqL9
NxsRFmLcVKJuXi8kK5hLeFCh9zEYU7rw3nKDyV+vJFl4nPvx06Hb0U/g1bIV24+kayCEq0L65LDe
z3R4hI1MUtT0YJLbVjYbbQmkTXJ26/iQ+4Q0rnISts4Ub+rG78/KUUAdxlZQMHWJ/tgB3OCm1aH6
3vfM94hU/PEY6W4+5P/ZdqRbnJU1DD6YK2N3nrGJuB/aHw5ut9T8xb3lifSoh3K2jxceJipaPpY7
fXurAOcxJZKFIVWOLvFRkPRv9o0jVAQZjkBv+29hPEyq0QpmQjIGzNrHnmHb357TCBkDPuXePYIW
uYE9MnIaa4VGmhtHwCd5pttPTOO9m1DCcnRgsA+2KPVFQe1weFufaCaxfzbIs+g5NeNYosFwOBa2
HJovSMlvvZQ7hYmtCfM87Kvlpy/g3XLsFjO5bZ2qkTVxH/t9Zo5tsM1rQH7CS5Cql64jJQ9H0WsS
F6ChU2VWSaTNs/Q01XRm8IICDeX9efW1bMYa14PcxrNRu2LWE8RtoJUl/xUrOvLu09LMEme56u72
DxKjWNgHH7j/U4D2rqUh0Bm9YnCEkyN03zuurfm32cj1JeJX48IA9mlHDkt+/4LJnMW8fn6UoKnv
ecfGV8+nYVl2Hb4Aquf4X2vKxYW1WpZDUuJYOYnD5dQxThSw4nMNubnYAzX5Mhgmn5aU9e3WsesH
sn9k/TftD6m1raif9UpYH+PlvOhmBJN+6TL/8wST4k2RD9HUjY9LhLFKOKONewOhwnAin8j2RTis
xQPXNJDWoQhukmO5XzAk70faB4ZVQlQY3HoHtVaCpdnyRUSVWnraHJ4xMBuzUFqwnpfjdUxQNQHw
d9BmEpSd0p7HSUlOR86hVVsWeOKWX3v6wwrWgkLXdW2HKOR+batNho/FZVZeknfrFPN5GOQ02Eok
W4FZ3bpGCwseVv1XbTkQ5jkUfcrHssJEoFhh7qPDsqk30X41E7jsVsjjGqy6E7QA2OjE3tfLmSL/
rb0/miA47JQ3EOYDBgYDqiFhPJ8kccWjNe1IBJeyHCpe4+gJI7hu538OZaTyDMusN+86fEVAyllJ
r5AMhAE3i9jdDxIy+0R/vt9xPjTY5DC/rbKpVPyHCweYmpGflosYwCStg25BKeHoo/899mE8/QNo
XuwNSOtVPkT/G5r6TCvvtir0jT43QeYEbo1dbtl0TfkZhkEqe+Fg6jACGdY3gYxZW/KmGexWcbIp
3mw3C0HpmNvyY8LF5OIY/lc9Oy7c/lqhp1qMmQjYB4BGyDLDwUPdduZSM4DOhY240PA3CLBamS41
3GEUK6PxGUdO4X7a9yITxFxvoETtPqrCrhknOovt5+pzmox6PH48+VY9ucyA5pl6XbQCk9GhK/13
9+zUE+MKexglRu9Uf/sNUW5/vISfwNNqRHoKeiU2x5C7GWHsccEeQewH7Hev3G36qeC2hXpOTnR/
iCLcAnydD67V9J1mrnNvKAVdO0+6FxstvPKedHJKNJd37G4VWWBvGyN02b57W1HZctuBLrXZf961
DakrL5JJDTrH+fNvq8DVet0TrTIQrOSM8f4oZ0lHY9Xai6N+Fbfw+n0IjEdJ/0uFGYrnaBDgFbcl
4dIVwP7WrKN1HbobMlFDDRlzFMmuubj/SKTZ3Ut4MOpG+2JD+lOKSVTIy+NkUB0p1fk6BEjHW6sK
FuIVqhuPn+pZp9k++Uue0KWR6vE6T6OnAwAE6dKGNTyeIWQjqWlt+TPy8KVqFCM3NOG4Qe5mio4w
HG+o0UguMcq/hZozLWuP82yGvxIAsQeFAbgKZ/U2oMwudaQTUrrk6hVNN+9FOW01NL9NLf3rjtNm
19p/DaEPHq3Wtf3G7oPaUY+BetH962REHbtBfMf+DegsVdKIb3nU7psMMyEarJtp0Y59rBixouyu
/ltBTQ/kwqll4LA7PEaLV4l7G73s0JKnwBcck814RiNhzt9MgXnyK/C4c5xZtlLgZ50IygebinT6
bzQrGA33OaU7UWffWKCnPNyW8oCiHdZgPQ/IV9S2bv/RIZOVirCbq7I7gH3WkTw95zSJbjNpPhBn
bM6d87/A+7ML4bdLOJbDmWO9czEa4CQntQQ0LVRwPGGN3uwL/43O7ZMna79KbLiAN8yJ5LFpbo3Y
aff1xio1oMaaDtTQroFIw8u6sT2KUDa6LrVwylCLH42uhxh1TOa0Ae7pDKNjYH081uV7DqOvuFEc
or9hPxlTYW/UxJggd2D5Em4IkQ/BmjeH+wwQ90R1P30iL1RbQpQbzOt0sj1tQoKtWz2l80AOMzxY
Mflm1nFGcPS9leJhb0c33CnyUKorUkU79NxMc+DAe4XyIGcKslH35Ef6S42NmT8OPjtYnLyfvIBs
k6yB66YJmoK7nsj0LEbTDHiHCcRgnb4UXyWyDSjuj1HHrSDsioc1YLezVi7axCBmLvfvDH3yES6m
CxDnwquZiDkju2IyAZ9wOiWThMB16ueMFSrvPMYPZG3eCqlBuqQ/P6U8ZbTaVIkDmpl/ljF1NI62
fwDj/LJ0Fq79ru9s9i3qnu5Zf/9kjkoFGuZvEsy0NSzIuEvsYAsu8Uj0qcQnxdj/0kW4WyCu4IxH
1/h1tf9J8vDcxB1QecuHlqIVOT+Cipw6QJA92YBpA5MM40be3xLIy6Vmkd3QAA4C2Uf+nLaeOUMO
9KhHRa8w8738dYe6kVxtPF25Y7x5gfcOhlxcsoIfXhpiOLzZ8DXVavWrPDTWWSYvCxWdtwfLBv1u
bgs0fF4Zsm1uieQY55TO/z//hezR8ePB46lp57I8+e1zmE+y+Yq35iYBXZ2CbncNHmcj3G+qM02F
ri/SadPUpB74QE6K216ori11ccl9omegrXLLXftdYQVYwAsnUq1GOuWkVAsxGDPgrFNzSvc1g9nv
Tq4rSg+yPwUQ10HjkdNbhAFc0MKy2GKAtAliJqAavnEInMC0UEKqP0kvJy2VkF729bICN0sI5uH9
xzpQEPo4kfbIDMQBvA4IE8fW5sr0aU1dMX0LHlZWYEOaNCPYfZczIO1+CknBjXfd7PR56KUQIn9K
4Titt+5F5JGAnJ/zPEA5uP+XRp1H6D7YjQ==
`protect end_protected


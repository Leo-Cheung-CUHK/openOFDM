

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Yec+F++z3wIQxkNq+HkCzhx9yvE/toYl9P8STGqXkGpEzsQlr62Udpo95rMKQeiLwSrHQp1fEznF
Q1QG7UM5qw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FLoX7yR6u3qZTIpzLbZZChDcZA05TI1JvCxNNDnPFVjAl+AjxcgzyU8p1UBSFMTEGUi5CeD9qD8M
gfJteYopZbD7/jA+X2ARuzQn7sCP7KCyCrlgs5JGjCpHoZfpoF7tdfPcIP20QQu9cC6fDvFxBc4U
i9l9zf1peW3zZGdD2Nw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FhDIp6nEK0DXkxfcJ8PSgwm/Jqm+lRY1eoIdTiu9o8ypesjgXAQ/cWZmEYl7kflFV9Zs2VajDHsi
xlsTJQJdTsKPBhJkfDlpsxtmAzoZX0uXNRtqJuCggKYNnLiwCBYdOJ1rVt2KszpTMigRwW2jisxg
lp6x2GHweoE+3JNMnMtv7cWRXA0q4LHWGqx8obWucGcfhktk+6tnTZEJ+E9k/GNBzE7F7Fzq5IV3
FH79RBFA26ZfjIYlRlBCZdHyIHAZNOUVVpMbdymIVYPW14bICgYnidAe+wwLixMWPhQfgeHdQ4kV
WCsEDryzR2P0ml/L3YYiIJN5ju+XrKREKO+8zw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DS+a9LtI6fMXCE/r+MSJh38df71DFCzFHmmc8S68kc4YfuQ8eacSS3WyQAV4j3fn+YnMdb/XsXF4
ITlDtDgEsyBfPKO3XASW2Sh+sYU1QAcjLmU9+6HmNDrjnhjdQ5okw/t63HMZDbt0eAwk6pA75Wj/
78GqSF7EGJfIsyMUASeAf7yKijcYOOVN47kviQORymwgSYNGIra77FoBBxekP97UyuC0E/AsO5Qe
ZlEa1+z4VJhej9lX6cg27Omq2ax5E2lluM3h4yHuaNZkGcVUc37t/Oikq9149n0+zpNmaZq375lr
1nHMCva0KGtUI+Mj5q4lhaEAhLVWejT2YuWM/w==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dAfCGzEoG5ww/VN/CcJgGcq02nC6L0VDo5sgtDHNJ6Z7aBdUBx3ALQRgPu9ajAbO5xYFqBboe0pL
FyVVJ6dLNcuVmaFDz2hlqiTSyUlz8JEg+eKLE6VcFZvURC5aUH74nuLpLVkDQlqE3OoYk3W/ry40
H01SRdWvVrwFAtsJpUriI6uEm1lVHiglFNZZasJvhw28IZDxpy0QrT78o7pcF7uiy8R7jbl36QOe
lhsEUDHUGXH1M9mB2NvUNxEwvhWzi7PIivDWdwMwQQROyTS3PvhdBawYM1actxHaFFqZpj5rFylA
57qsfqOe59DuRKVoB6Ws1yO8AErTQ8gnrUCOcQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
b+MNc79bqGCWayp07urW65EVoAtBn0W/y5D/Iw10hHoNLvwNI9DlEOK3rXmS5CkeqMczuHtbc5kR
TjocbD9VFf+2zr8PZwlcxTjhbE9isnRVt7CD/g8VMx5WetuuDz3byQkasl0nomjeISV/+Ek0TZ2G
BcoeTSJRJWl8/+q/MMg=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ml5VaElc3u5o9OQAeaoKZOzSgxAT/UigiaRFr/0/+HBzYBLpzRT3NOQ11TyVYec8ZZ1DEXPADZON
gafcUsq+HhfPPJfA58Rwm4+r4olpszW7jtewYPPFKExevpgPxWLkKhWIOmvDUuywpIy0CR7JWy8d
/U0EEmOApXNSFB5QpgllEQIAADHuOzUX0w7d5CzglPX+5J8D0m2S3FK3gxcO8QCkSQvPW59HGP9F
TENSl3ykpC+OrdkS8jMiNhyqWL2R5qIsjsKN9ANHW5u5vysFm5V1gREL0fHk49uLmxW+2VJ2qii4
53uzbJtr/cu8haxZPZkc8nDZkkEEbVyQ96xZ6g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 175280)
`protect data_block
v+ZmhiOiMolzbJlbJ1Kl61CzkobMqUx912Y7oDmtAHBJznpP9MonTkAqTY1+PGlf+GrfumjSw3RB
TX/9vbfOISgc1OmWfwuZXOHNUW1tQMUlOkLGkvmYIbSMJgJ0vj36lJa9zfxcqlV7Ve6g6hZUjopZ
0leObVMhJF9DNjsLRiEQdkvjbN2uN6sMvfZIS0V+YHluykwYLEOiBLTRT5gt6dK6pRwn8Nyz2QNc
Z7f90sDF69DcpWsqeX4ziklTEVVPz1n7UlFOLSQYx54RR3oV3/vmkWU6ZOetDG0LdbbZzE9rth8d
g/e3L0Eb+m+pqjzMxcuutDN+Gy/el/8Nkgvht8Mbdun4i6785sC/fQYlXbVRuPlQCOVKWH2XDtZO
biIVyv0/GFXnAtpwQ4r8yQDnewj9g1haxbxdt7XBdt1HnTdcJq6hI6uu/9TulyCJeu+Bwi9xJ45J
jv+G50oe8sRZOMuYOVHRxAwtTCCnpz19+HoVBdr6xpL2GLKRR0P5NWV/+hm+5gvOhl8bKPfoOvUu
BcZrITUM3M2D3+M6ie3OqmWffyy1TA78Fsd5frYW5v1A6ivMNNViIy19H5cvewfO/aS1YDxlaHBR
b8C2gXEljwSubvpOJebKZfxFMXlmwHaCStW3no+IshBeJibMRZwMhD0EuZjbQU+Nc1eD5/XSPZqj
ZN0cm8R7ebAAuPWRqN6sWT4c5+VhWRgtfOPMGSt2fq5UAe4Y9JujErxLTKK7RJvV7bsStC7HNvko
iWhN7H+jUnhx/urtEMQWF7tOyME3/oJoaUL1Pu28B8Ey3HXx6rKdfQEDA3ll2iNAuDfLrgvgviBv
cRLs7f7OWx74aeyksL9wp9w95FnZ0mH6zKERmFEeNG7L0V2dlVE7ek3ysknNgbjMVXw3dRiwYGao
3HfOvPvB5I817CgvG7IXyta/oUnoYWU5oMHbriZ3aXwnKr5HRV4q40YcASW2/kQT3QQaCFczQRur
rDNUVhNqEfr/ZjU9A5LEV+HaOnkxhKPtk6IPK0zXZUjUbTnrm9h42jVb7E3HdMs2wxJSnMsqlT9G
vhZNXJV9MNJyWDMggyJjYqlEd5gZ3/VpOfNHf1DPUnTAB29xZAvQnxLZmdPYuIuYMHNPklss3n2R
YTruJnjBsP16vJ11XGJKdTJ5yuCn+YEFeNdQApyJngWr6ah30xvuTgAZnKk1eQ0Bsgt94BKX+z/2
VYlcAhhjNddPdSbufwBq5n/tfHSrn+Wk0Dmas1enhRHz8a2ENvT991MrHgfAlo/7yHW8KwKSxTWL
0aj8GceQT8u45SNJZ0SFzA17cpEsOeOC1sQWY2V7y6nVcdDKSL+nZ1A6yDVSP0yGQfKCzoyx2q9B
NGWYPVjQLeY04wPbwohDc/MVJWSIjELVbW6fnHxzIFAu9AGNCsIrTIw1CAO1C4zG/i3sPPS+XTVP
MKsHtJyudHlrrsTgAN0R8dCai7padL291FmGlCl0r+zEG1rUHIsgGltcXN0nYy3Pz8r4LmaBMsp5
ncBh2UgvqXA8DSA6l2LvGLtQ2pcLzUFaAfw3EIFl0V0b98N1nA/rmEPV+w8KckNWIE+/PJbAMYLY
0wi00bMqfQB008XsqaIeh+vec/mAn5OG5wPD9iSLn6iErJ1whG85qTBRMpQjuUEXC2gyzSunHLXy
QnsOn9SG57OA+Vf825wP3OP/uC3MrUMnZ49GtC38SllOxafk80IfWqEX2sIHadvZVZ4QSHHMIFe7
40s/UUNmc1jqCById1X0p51//2g58vkd6jyX6PfTPIM3tjKlfGGPjO6YVdlgwzEZGPQov5KQiEag
6aznz6l1cHS3WoOjSDIMKneRhK7QR8WoZ5QAZeNLy8CqUOqUs6Nv3I1wrJUONxWw6seaPqaQuWJI
v3zwh90JW/QdO65i0mVbyZQjca/Fbsexr8yQK51pRh06RiyAMBtg/AygOVZnvI4z09WZSVrvoKHp
3zKiUy7WtSa1vC8qYVh8z4dEoC3W4+I3NScIJG0JsfLoBeVZDD3MnkPFl0V1LoKJlXoU52yztn/i
hWKDkrAEmLA7xs7pwi/O4zOCFLk58O4oBQCE9rD0UqhDsJzgfi86nYrL3jUQvDDNzQjFvVM3pqM4
f0yUSHV8nn79bi67CnXF/SU6AArLaRhjJfw7AetBHfVDTsGeXD1/S9bCGm/KKbgUKeYMSLGssKWB
vTa+Ru6/yKLogCpGlJQlG7M2/fuInQwFqtF75tc0OXB2dwH+4P+evqBs04U5uhF7hIDZ7EzFCnPz
HkSUXzFUtwM3oREYCrNAZlbZaEPqU4BRXt4j3D3qxLA264Fj2E5ZPMNsB+HBfK/YeBQHpknHMN5C
3b2PIpdjtlIvumFxQ82a3pxVn1Rpm1+ceuTUn0NbhJAvMyHgpdb1LgZzmwPRbzfYwZWudAQr1ZVe
8ArlPPTqSQGtJgD1hKMOfnDm5XiXx1DmX/4y5ReCjJhzJNrDB5jlrGyFsRjozKeVzOrWFmT/sIHD
QkC4uoRIqoqqanayHC7GPOdkRfIDdR8CL5vkYMvxrqoKuLhHLMMqhG8RV94W0GViSlgYt2jqygui
sVMIMJP28LKN7iYN2+xSvKXIfqf44Ma9OJTs1Zwl2HoQGutbxcxNTx94SZM3GCwrHBrSt1YOkM0R
9uWTVxLS9DWBMbSID75tQWzpqUfYsxcmjbFGD/QzMejv2b9iBPlk8arasJIyLRqCPp2gVBdU+kmT
LKEQQgD926gpmD80tN5g8Q5ZEQFS0wSIeAnomZ3+C8FJSmi2mLbS/VChi/GB3KMGh3ULhKp/cVah
1QChRYEjl+BDylQLErW38hixPI9ESdSvAWWCwWw/p9uKSCC6TJJmS6za8yXy8xb82uOUnv2xW2sy
Df0ipGM4lYlP5uPg8NzxRjZWmHI3ryf161tHxTvnJ1EVkc57uJkmI6zpvGWm8ptqbW8t5gQAehJv
kGpMxusMCVVVg5axvl426NpauvZ9RH87DOc5TPlYC57o76PKCvyMVlo+cvr6W9Bln1QdXqa7zDQP
pqYWCaxy+WkqJGz8JT7lptfSLzj6w1zaVLcoEnjSzwpNeAzWFB/cSyTQeXnM3jUFVugR+n42rJjH
DOxKpL9cm4mfZyj7lW9K9pIbo31io+fkxS4+WzMj8E5nvKBnTT0Hwq4/Q+n/7gtpVYm9lt0WKYMy
3mbDAp6gHDj6dmsvWcn51Dl7jHmV34sYHpkomaojTT/kZfnpxShLtNLMJf9OpFKMHbZiNJw7J/sr
jgmAok1s9AW3e555d+A3QsAf7YL8htrTj0UEFpxpNuGPCmfGBqyDA2fb9EITSVFUMFd62iaZ5OZ3
g3f569UzNBBS077Wp9/ckv0+etKai4p37fYNj1gwAYwWNRmqrGfgUb2NQkCwx09VvFl9D6k0T3TG
/P8VNr0B27jPD1L60K5+m4m66yDKx90AlochUKyHR66nqQ1xUWXSnEYcl5iOGk1RYWT7jZFTVg4p
2Fqt2TJImlIsvg64ZyCfeNV9sKT9bCVzn14tfvjWsr+1R5aRPQlDEjX8tIEv+MJfL4tMSdbiJ3JK
39F7tfBAPtljc9VQQKrcI/SAU3/05fXUsm/r4UjTR6bjdqGthYcS1VEGY+KGyleg8oI8zASycaS2
J8Dd+PwoO8p4mz5N7qjaMyZUPvEiOymgfIoxoxv5mVerVjpUyaavp2Q6TK6YjGBGHWrWP0g2qZLl
NxGKY2ImYAcuTDMrK/J2xMcDBMJ8/IM71b6T0eoTLSuiTO393b9+ky/uUoe045y6/UCWzuoPpIPq
GfhvpDgHuBCdpNEzkS3ZvYPbE1GAHzbHraLikO2ud3h841XOopG7ci6ecRCYijS6YzMlnfxTFa/g
L/MizQb6gsSzOne9gDNVCuHLmRkr3PrDGVXwOQNMfGcwYqeAsfk3Hz8fb6zW1GqrxX39qIWeyfD7
SIDksPGtFjmc78OEYAKk6QmVfX6Wuo6lVJ0Guv2QWCHZS0Mx+iDarNWwZm33jmwSCy9i4gQ9ZmOM
qN0+y+44SVqOwAfUyKNQA/eyTYgP8FEfHx1BkdENycrBKoo3Nn0PL60hYDPLZr/1VDbagEwS1EzP
Aia4GSmXMg+1JmaEZFYVG1xpChURrCWBTSDtV2wmUe4tv0svQTeIwt7OW5Bue38UBT+dvkUvPsa2
Kse3HiXI1DNI9Eac/2btHGqADrGvoZ6DRaczBt7Cn8medHfK/kwhCy6f6t7RJ4ZvF7M7TdQSRYfY
82Z6OFs3NrDpvdZNMwUyl10Jksh5w2AqNs67a3kanMClfRragU7aZ+aJPMwJNTCFkjm26UI30KTn
IL9HHlHT4swet2553mtseY+pkagOTLfeif29t6ChjOFfW8J9vHBcjACwDxAWeHyMkRz0FpXcE9jY
M7/VCQyG61o+XyA+NTjThUmWdQ5MhpW3R6UFVxVcl6itQr79ZiJhJs6+HjE1tZqpzYdQoVFfAl0I
VavqibU1LQP+HFpNlOby82l8X5vIsUae1yOkG2s6L7DYXMWhzzm4IebA/n9CSQ0jkhwddybeslxy
7RhgldjFcBTuhx7BCLxityGmqlilnmx5rDwvYeOfDAZ7xKzC7WsWYKA+tE6+6KqYZUb8+F91kCrK
DN37P2rlZ+3C8TqW0W7Nmk0KFIpoUWxa/Mas1vbSXLp8YWCWQlV2+/Kxb9AjLPELkIX15lhsjMxG
jn9V7qfVjJADYM3Safc7yDnx0q7Rzu1/oDE8c6hI3vhScaGJ9eBx+10Lf4Blhj1t8ZzBi/AEogT7
KRhkPF5z/XLtuoaXa02H9kg8bKxFU4pkK6gtGNNk4wZ/eSU4EfLyYiPsMT8N3ofRu9uJJTunUhKW
y8z4NsoDDQJ1F+3T/RJwHD7uqYQ1zG+57YCL0qNleqGGdmAcVUx/TM4TePl40sH3TctO0nrEQgJa
SMH6uB2G6Z6bvzXkjBaSTNZf3ztZpR33tKZy4/GZc8/isgnXS3k3Qo9gHT+0S6OeK2ixv5OeqMzF
BHiLA4RTfpGyW4HdIVsmJh/NlqazsHF5+r0cfQ2oRk0b3h52C8P8l+Mlh/X5Mi5S2pdz1P32m8xd
s6Vna7DHThVvCt3LTihYceVqHg29HQ/YG/icfSgONQpyNVnAn9yTiMfjBsnPvaPMvgq1XJ5j8Oy6
7zXSQTEVOtqd1Cp7BVtA7435PIv7YVB9WjB1awQCKiKPDmCguEkgHtQzvcMLokcwm18BTbOIdzCb
jvoQ2h7sq+qUmmnBstXrNY+joCwlALO6avXTkhEKA+ro3zmstliZlsVjsiIFl/WiDMfBy1tBp9gZ
rK160/FYaCIksUSBIld6KE0g3XnhVcpAlqNLREXDbwjEq3oNa0v2vQQi8q4pBLF3TVPn9FXZ0Qz7
xPX7kz5nqznlOiH2LTrf6oBbQYEW9DjLOXrsEwDYHsao70kZcAsrAM6J9T6T6ELPlCeRAu3ynE01
bG7X1GUiJcGBnbM9CcjujwshnD+gtsQm522txZ6lJcR7gbYfY9QhDgY5pkuVU1EVFfxuKF16cEtG
X9fCqS633D2UcO4XLV+/5M8fpYOmQioNC2vkJh4WtY5qRkEuC8oPy/avROAqnmJl/Uvu3UzR6SwI
aG2v+ZXvjnIPOAO/nLHgiakYEphvRFEV1XOZA6FFhTos7Bu7uUnZ8kYgz3Nr0p+X+EG6avpozuy7
l+jr7cu13ulKQ3FqJiDlo8KAUvFnUMLszTCzXC3d2SWGAiatQSk1SvmDhe9PYLjTdWjj95LRBREf
Ip+ppZlQ2CkvJPPjKPOy9Jnot44OX8V5xzGDspGtyNyvD7IBFHUoyLAPF2ZdAf1xiuce1qoiexWE
mWHcKNQU2dpnCDtMsqG6gjkXQ/sncP+f6U8cA+tNWKMviOpmw2ELDUvYMTkuo3cyguVXgbVRL6Jw
XHxfLRkL1AkfXWkUajne3Wbe/7ZlWgayYidktwSdvnaK37Rj4n5S8YD1ey9GmY53rd8Je7lgOw0X
EMPF4WhwsRJ1/SLp0tbeQ+k/3592SknJ6PmQlmDdfILy+njb0MFTzzM5IZIaFKeBb3sieE9wo/uX
BEKbbSFh4QHeRCwsmJvgLjYEJ59qHh9UhBGWjQNFVmgzk8+5HxC9KlVoffVJUtKnJp65ESnyvwpK
OBKem+O9UvwTHBEModg1QluVQ4bn5c7iNqy3uXjDmBriJ/VAyIXreSujMvOAPmv6ZEk1NBjapUj3
uB6K/acfc97ELqwdyvKhXe+yUbg6CI11ma6zchgwQbd91TtolyI4Zoz7eShkLLc8hDjyNe8Ry1Ko
NpVxLNHyYgQEo56yVVfTeYospd55Z1BUuWLR/sKqwdw6KWtcbVoMZJh60ut2eMIo2jq2/dAbA/Mv
kKlWTWFqa2fNGb56YOU7HwUHAbXAYAZvptjlNCcd5BsrgPNq2fNCJnLy31oA0VceUpoqceqHqcKO
Jov5Dr7fjsyululRe+zecAizGIpGj43MlSwEvvucteaISXqIvRBQTPtwHrNNrAjK2PAtf0tLaW69
6D1NRR5N5dSCvsMaBXz4ymnXTNIIazLmjRLZe8bHdWwHdx3dpW8WdKHxNkEcUym2K5jHmg1tG526
q0fZE9kxXOrPcLSQP1qim8QUQMBtnW9YWGM1d5R6fePeVihb1hc2OjabBvxnEisENSuOIAPeyLQa
SRO0yFlsNrmiNHWhuQBznjTgWQ63dmNUe5KucsOVrzMTQ9xIJrlGE03clkXTiifcqf4ANYqUPDuu
9GVaCwlBFt6lfwWRtaU+1eTrqQNfBJNr9j/Zc+2kjGUMf5mWPQ5HNT6iXuTnbK1mzv9g9Z7wsrbY
tMlwDPeTTeuHt8KSrNToBitkvlUHXj0EEJB92qNYe6vG3GFmbsl608FYvaHQv8avBhGz8maLBV7b
bifXlv2DPHJnce/LfLrYxDDLipSt0fKnkMyQsI+qBf0Csni6JvsH3lRLD9UH82+BjOErmrmBqYQ1
IHT0XTMny6CItMI23bf+0YDcaSQLfjcqgWb8DesYRGAjXoOzVgmt1qETwAcUWeg0+Dl/G/kvWZBR
gw2sZ2O7+GKYb/v1vvoBouCXhWCeG4Ek8lFO1zpmo3RI9lOrvGT3rWB4ZortDXrmSsRy9DAJt2gS
2PZiz29GcF7/4xfn/AUJVgQdybXX6fdP/Yu0HSrP1VP8JQ2WnFI1hQOZDkBytduV2SMIH2sGNeIQ
hupu6B4cKrouy+q7s/DzbwD4Td++T/l2VQ89A1IbDqpIyjoJsbdJcZtXsZXGN0Ci3pn1n/Bi/AcV
xXyIEgFxM2yT5UgtqbUSpu8NYR9fNHvgViWoNItDpNd/xYH9hijA8iGyNIIKmIS1AbORdUHzUjuj
2SqZLA5dflJrtBQtxzZ18XVxknowuj5pEbKgOtpXIoYXc4YxOGeHQoHAc4KuLvxygSsQzs7JaLWZ
BCZ1S2OxFHDLu04fE1s6ZrRkI1O+TH/Gj2mZTHaUnYPlSDu5vQiHgcIx7GT2oyvAXmp9O+AutPSX
Tw5leeWsAPDMgniu3FWhkUiCV1yybZ1pQCtr5Wzc2kbQJewuPrmNM6SymWS62wOOrGOTjTPU7FPt
bLRpICxXX6PA7UtdqJimjxireLhWDdCsFJ8yj22IyJnAKvAFYUE52ucRq1mdjXO0KbkdomXkd93K
BEbzc2MqJCRBs/gxGBjrKylILEE3uIeh/+zdzWYFZeQHT6Ph4+e5GXbtBWHqwU7hDrv3oN7vIFNt
rt+lBxDer8PhjlFcV2dQOLj/n8CZ3Q7wlq87yRSm2HN04UmzlP4SS411BCQsjmn4wCNhICHkpfNg
pbguI8MdQkbpcPcc/4DD+u7EA79C0+XcLDoF0XYqg1z6HQrb5H2AorkIqvBN6aRnA8Ltmf4vf2Y2
aTQJ/f9fke9Am00kbQl2B3CKDYvpWg/0hKQZ3UeC3bNIGI+mL9NZEtNyBDWY1e6yzX3JSRudomxh
kL/XQyZRi4Hv9AD7Acr66asMG6rgkJaw7Auiq7/7Ju8v6dNcDGagYoLd4i8khdEKutyBLHnCw302
g/0mda4SBHOQXK2+Xv8GruY4NLE/ANhhyEVoWFpFjGgXFazlKpPgReYSIYa6b5/Go/LX7qc7F2vp
gvzrVowsOnYSFqBdK0Hc8rPLGuQHGGUPZ+Ylwvt1WvwXGkSC6zkCbvMRk+LsWIEAoQbPVDENP0F9
gY3fACLt9qc2H8yWjphYu3gZ5tlGsDWFwa3o+RXfZe7xmseeDIzpmksBu8tLYLEGiAXyP9LdKA5W
Ox+tBdBuoRxaSO1BrXrR7gUka8WZm5+EWoLPXKLWHfm/BKXaR/5Oy9/ABC5qZFXfUBvVmvtdtv0S
iO+KZ7Q2BcbmyQZ2ANHJp5O+2NWnE0Y7bTlAAblbp57G6PGA5Ax/94uCLZphQfqgRYtJdUE/PBkt
b9EGWZng2siKLF4MfWQllZ2ZE3GjHjOgzGLg1GJPqCXdQ14PET+wJw2WPzByObiNJgdudjmqMKxu
1W2cmKDIArMTbcps+ypjGBgByf09lzPmxZJgCsbsbAa9HVWuAbAea1k7EsAr8zcBiDzoHAIsl7fP
WXRu+UIXzK1GYKMrMpLlLu15MOA2DJ6qwrn7AZ3euKHhxJOA8S91kuBBTG4/P/q5NBPmqlBU11p2
DYoYKO+gGLGOImQjcNwp+90sC/FR1TGUj5tsdmMB5/G+zh4VTMkdqj6IwxhkRgx0+euPBwZDsPmB
dFcrN8mSruQ1KL15SBX1oh37hrIaNYS11+ZHMuMqqXqDriLZPDgnI5Ti72QxuFCW9xXdaJ4dwpi/
3OdYdcb58RHGro7BecfwoYgb7jclwyg4OGknmL6Nsit46687jDOOHiIffQFC4GveDPVTQGvSUIUr
QpqXZAy3MsovHJCKEzzzcvRQWAz7ruauOZSjAfq77U+yTWMInmvdQ5B+YcU5SxhJRjFffjXBnzdL
pG/KUGefri+7pYLtwKe14zanlM6h3f7FjC9fxu8BVMs6XYuit3yGagR4Gnvm1Kc5BdMhPdlY11K0
LR5FfLFWz6JGwed872ZaCE2z0Nn4aQVjCzNVPDpTIRKxV93N5Amt3ZuBOnvU4eXncQOng/AQxX1+
S1JtXuBfH3BRQhIiX5hqMXNb4PX2BiNElZCZZ/y57VYoq6XgbfmTnUgzSyJ4zUJCBzN/jkBJrNkO
zIA6aLoj1uoHDrEFGEpS61B5I/MhA+J9E1tRhRMtwWyv0XeCK1kmFnLK1OQDwqaKBputYaCWgt6t
/af6IgrBUYzTTjqrTfcm7noMhPxG6pT31yweQk4UOB4rXN95kdijFIiYbX8d3k4o90sFh3exyDcM
dRAIO2CT1V2Lz1FqPGjmsTmmM8YxIvH0IeVWvaRKFDZPCzffDDLFhmpAmC6MIOH6jZYMNoX5u9J7
t9g3sOg/nLAI+3Eu5pyQx4Sw9o8kkt2m+73t9n3CH6/CG//20Zv3c4tpZDkK6V5/UhmOIW5+bP6D
sMaY3xxj4DPSPsc0YhYNSZMgMdpOnoMCTWIPKpZiuhxqDrGpWd6hgVWoh/NTya6KQAOxUhxZ/JdV
v1PKbYv6Bk/k9FvrGBEGlVP6811gXWU8RD2BGC47SOSA0hG1UQGks5LIbB6gcZ9IMU21wqreP04/
wBUnOEWWuONMZmyORKmzFT8QBP2L0+b0LvoN2kY2etK2kZf3UtPrteB0QAQN33Tu4manyrOrYnoB
QR951uU08yAROZjp/oNLteaoXhG9oLnhrIJyNlUwA0wBbrPmjti77z+qY6Wedy9yT7QzTw7vzD3t
/fohPO8LQfNvn1yZ/9OC1mfOOmtpZNDOGUX9iUBBZeQNWtXp6dSLJbyK3kLqsDsvk9vOm93kS9bj
ZL2aNB1zl/hbEnRW7WfuCX7POiFh/qJokqYwQ9YkYz+LwjYLxPuCr52mSFAYvk7/6iJ3TLvHL1w9
XlM9zAK2G3tFOiVvoj5PUBT8aJ/mpUFmXYVod2bYJMkTb6UkRhN2x7FL+9cTzvxU3dbm/7mxrC6W
JSGIFui++9ydZNe0VP3AdL2zebhRJzn2dofMSp0XGj2ODc4+i+/IYWdhYbYsY4BWz/qBgUXgJz/x
iz6UBPfROP+6E7EpE3mqfS8GBHbY6AqrjoXxEeKv7vK8aSQnBcH+y1nNpqkUQDBnGTEKp2Lv0X9+
UXpmIJGk2kIViUDB/WSeTp2sWiQTnkWKec8UCEQvR3iCGES9ShU2ftS+/w5Bn0iZu9Gm88g4eqV9
Q9pbs+NFEDNDvuq9RgV1wxhKqUWh2ValCZ5EX50pK6MaK5S7lUtA/MFeVCHeqWOrhiRlmkWD1KaU
vjPenKMfUbcqWLrhiu5wJ+jP0Noyh4EK508nwUASPpUQXNaHysgitDmPDsvbzD+BWgw3oOlEHHYJ
jELLxzu9HogQ+kvTzJ8UzPBHthO9Z2bsPxkZXuIMHavHJeuLYwdsIzXF6hh28iYs1W2N6kg+JhMc
qF6Wy86010ZesI9MKyiGCOSy6DrDFFeaGwLmsc6hhZp5KhrWynlRUEWWo0rp6JfcmO7UeyzXH8xM
xPSgqbCNH22IvEEfwNGbwx0f8AALj1oyTaB7C6BTVSjfehfCIaF3Z8jML2uTG0bU/S/yLjzHqrEf
QqfkUHHUrKE54sUbeaYUXziaSkC88enAhjff9MEL81g53joT2sMg9wSA4AkTeHtrgg6c1uC5O6ac
mpOwaXdy1DjXbVySIvSB83IepvkLlTnp3FxnFTALF9g8oS/ay9l0TP+W3d56yIz1FFkkS3IYoDmJ
dqInK/ZgITcAEnLHG7ynpLu47lGIXmaJPbXuYNLRC/iAh9EHK9tlCdXC1ZHjhJXiUtTmt6AoO9hh
u4XeS68yLEn2nZf7DwkHsOUJK+sS8ye9M43+IRek5u4qhbxUhGN9/+OCTt8QmNb0V+L6wIXrsw1M
Y/LPn25Um2TsmgoYOu7mdO1e1tI171tR88kP0aRgDmwuMxowOlVyFt9VyWOTaCBD8n5K9MrdOBXn
OM+ki+tqROXiTsF9b82xxs9B1fJKu88xSDYYQB9oYugASlz5fg/2zhtPKkfjEGlSy+hwi82M7FK+
eaSzsCQ7liSh6Pktd+UbJoGcc0zrF1LAUm4RhP1Gxmw0MAvArFIABLPoXrjc5RSqCe8ykhytEEVG
mfh0glLqrKV2DAUQvA8iipTyRHUBv0T4Rrdx2iXgXb7fB//sObZpOBrhbxnFP/MMOAbwymmzGFLU
TemjJKmkgHzD1Q8kj7phTzLHBUAp5+zaIBF4aY50OrLFiWKU9FBzJ9AFuOFaCTd3WWe79CA6fa2y
Tqg6/eSa8y4nxUMvtAdqVMHttk00tSgTiWeFcmDBDgTbydPq2O5abToS3koKeagL0KqLJjVBYvO2
GRvJNgrlQs5MDZLBMFaf9K3w4JL4lEMdy5yZg/DvRSYE604IL5HSS9QkEND7ePAcYz7C85whmnaT
7mpFVOk0qd8qSUWRnz6uQUFA9j+xXRK9UOaOMePOpeB8d8b7uAaPAnnyRotwyI7wY/ipBpC7mC1z
twuTEN4PpQ8uQh8Lvd0yaLX0snzbMoEU/XzOWftryALeVjIUAqiTpWnznM+KxIHj9eaXTp5EM6Ir
TiJ8BrHXaMI1+/3c6IHasBE81gw3YiirFzp6F2s2tKZQUXmGgzqxtUwNO+KeL5OMEXDWu20kRwNs
aBd5JlIWy4Fzae3mV5z3h6E6Gu8zbE2PyopItPqtfmWGyXgPJZQ3IxPlq0J0nA4T1Yz/QZyid/jy
GcVlkKrxGCf9EB9BKrurz7BtO0MMtNvhL3KQdhVgmsqr571cF9tPVdrRNJbZjMJ8u8nais1txGkT
maZjxqakR5TQFzDfzrtbBt7bYoMyLkZ2FqJYUL4Tj0qDLINPFLF60/oFRVyKRJTkDpu2abOszy/O
O5Qa7yPNpxqSyl0btgYlL3dLAW8yB/05F4y+RYs2wyRGkMAPyV/ZOEOHLnY9kQjTxMm2g3AsV1ob
Tfpw+SHQpw4qcc/P0YPiRKsEQZ3RxdmLuIP3EXglJxb77rIoDrDnp6I5YtwVt6SMJI+ks3nEpemk
Bei7CaV/mBq6NabW1GGmOsWRpWqPXkJvT7iOd+WxBEcK9k790XCbIHJABYLOoDxhKH/3uu416980
vme3Y1RBq8DlqPE/FjlUVtgxsn5oySEf6ubc0D5XL4RXO+Q4GevQimCOPtunpm+vGU+hwRbChuNV
+tIaat8uD8UwsfEuE/IlfSkNoUE8+HUz8ZfahgLLf859p21gSRFHQAxq1Q+1f3csqBXc517SnnwE
HCI/3ymT4+FJR4WZBrqKstye/V8TEJ2IM2oOBznMfgy1gLVXcm9EJGqf7s7iKR75wJwIrD9kOk3l
OsIId+YwFTZ4Cb64GxJ483SUdt89kaYBXJkbfKbCIKYcqTMrx3JK2bhD8xfTzCoktsgWmNIiG9ix
KGfKQKyuZL7nwJVbZZ4bju+FELUhfCETXQSpqZB296TbHCe8sUJKMvN3hHutKjIwZT8wVsN1C1Ib
gyMyDcQ8cPwQu3cC97f70O4wa4mM3EkIcm4PTFLty61jieTWNyNobTYXmBJ0Ty4zbcKCHsMEpyfu
+SA4s1r0Tq3yy4pTxTGKW80viLOC0ViZpNlYvHMxX5Hu45GMe5fmwig7IjPwze2DOU1xkTwHuL+2
6YfvPdyjxgz2j8GVQ6o31MHcWC7xsUP562QgOZEXvAtNYBqODbcPjtm44pwxs8FnVlQyAQZ9Cuqu
AP6V8fDZReDJH/SQuzobZSXl9NoBQ2NjynRNrYg3ORTw2T/KzgqG8hc6UeIauz+3nlnafjHrjjdi
EZYiRzm2qrjl3MPXm/UgBjHEqMqqTskS2wLMxVoEgvDUhFRRsr4UQ7fI0piumcvvfpLSdymOGfim
bPHmgbhGlI5KpmuoK4lzUNB2KmykCPXNS5FohgpVXEo442V7ZYYb2fX/mUp4WS/bnUug9G82rOfL
i4FXGO/2ClFh66tM1fKPyLrRG1CG7ts1VhEXF/wT8ikFrYPy8aw9owLazZFOgig24ycl0Sxhuzda
leBfjeqdKurHuZx28jVWUip7bUWBziawPkJdDxgk793QQPHWymDSD66kLWtuxh2j9rtAUIccvlV9
Ny9K3vPeooDQPYhNuVZkdE4w7TqsjeoFuxwfwwUITZRQELEXaE0Mujv+Cybf+AtUjWXKElHhyUjL
3NWYbW+2eDIAfaVwHkD/HvwTxRBMKUxHitA0+qE2OHYyE9vWMMilWtmdj6P/HBRIE2obpwWMTv0Y
uxl0rEOnSggR66hCyMX914xPK6czY/j8Fni+3T5m4uGgjZGc5S2RL8wmigInHgo/nc+UoWGi047y
ZwxGPUP0yj/T1La3iy37QwmPirXLZ5BKWUufcUKo88z50ZCUqzU4hpRn6cNCd9VINNHaptUK0l7u
wbtwdnH/8sd18eYruJa8BQFm8FeSRRdiPLwtAhZhfR+G/UuGlGq/giHtGHR4J/WhB43qrJmU9QXo
noVFgBdEnR559Pgk+LlE/m4YYUs01h3oT5P0e4OqSPQo4tTeMyWe36TZg/DDkMKYZxvVjVDUgeAp
VcyhPYaiQfxHPEbJ5ZYp+PlBQpo+BkAg5+DKXj22H9FZa580kZMRxjyg3bc9mMMT/4MiIlUAWCSp
aVdgZWZFTapENKFbyE1lSWWJsAAjBfSaaWj4eqKo0xAHG2PKC5g8W444+Dyfsi0VdUnen+ICBkFd
vufx8cfc6HTp1Ne/GDrKPUiKaM7Z0cRxk8sszlQ8Vee8V38kiJIhLzcVxAyDK4F+8mN2epgSH1Bw
fHEnPPPiHq7xh0rIAn+PbMAtHwkeUzHjJG6faoSUCZ3wczAh8vUx6dr5/bm7iKW/opW72UfOnW1L
MMpYVns3dSHcE7+ebRSVQsBaR9L45WkG/2Koqtz0E8F5JsLm+dwU6nDK0ZNU4G9OoD/f21mKqIjY
DoNTxh8G4xQ6YQjph02ziMLBHjPgvKtQIzaE2cvU/e9TlzwONPZ/YG2nUHx/xDv09sxyUtChz9ZS
B6uyh1TWe8T6pFhCd3QeHwA17f4gRwi83PrASmmpdxP2sD+jEL7ia7ma8pBoL/9Nltl/fWkwvXUE
Ny+opId5AN5fywnujEHPvQXN6F8n6JQ1NPG4cYZApAsiEzAWhuUirbV1oeCZ33UIjpWC/oNK7NC/
WAMwFfujgEBUS+Wo5sWzmV0wvmNSNTow7GLtMYxYTzGHLS63Srw7bR1hGg8LNnMZCWoeXB3DY+I+
FzqNNJlt7VYvsip7fi/D9wKmIUGcg9eA0HX+QMuQwoCLCg4yqo4qVZjyBh2vYJjcl1Mn602yr5jo
8BdYbOX3hPnlkWoNk9KhdbCD1AAMM0yjkSkQOaEmDuwP++kMW+OkFnMEP+YrmYprPFiZE+YwXAOz
EYrSE8Zil2DFkRHH2uRJYTHfg7loeeGofaDAgKqqDWy0lp12haaqEaC+Lja9BBRWgwGnEkO4+Hag
kTk5HBEAzWezmM3Yr8UGqhCiqhGZCnQEyRscsppMUGgPVyG+1Q32/dPv/zVpohyvLL6GUyFW1/zC
nkrmJK3gQGDM/6Oemz7y95xUUFD8dkmfo9zdi0hF+joRDJrPzRv0pqATHL4iTZ35Pred6h0UKUQw
Xca+keSRgdNz6ExoVOajMhXFV/QRS/ccz79BhwfH+JpowEy977OI3BJN9chlKBHsClGLQnugOIye
jZz+SM6Dv+1TdhJtYHhK9FwzdFZfDo2GWrzMVItNU5mZxl1PtXM5+HeoyhNHi6ZcFqpp/qav8Rxn
npEh7vFxxi3d+vwVNHyyA4/w9k+6Gwc8VbjLo7sxgpUWXJuaUwCmWXY3+tJPrcTtPbx7jf7x72q3
7anEpNO9BragCAaGAc2wbRKhiw1fiZxi2izDv2tBNR56/W31orwcU5EXxZidc5yYbxE24PCed7F8
Hb8Z3FallbRAXEi33UF+FrTGpaXYkBNFqhFwm+YZdKNWYKDoCDSbCq2l4gEVdF1yp2eqgK3bE+xc
RBm28re6ljpCbvJ4cd8nZyZrvTVwfyyWmyTcDv+p3hkM+iOyYy2O6q/zdszBcHq3+6yAcx5Jm74W
At9Dl45OeOCSodnQ6IT8MHbXn1JNEBivpIgwzKNX46CJjJkonF8wuVnWpqSe0v3ATBlPyMzfj/Fr
P1o1U8Ih2IcwOeHN0/aJOEpLwPvkn0kD3kd0cWS5UxwN9y3lUxg1VH73wYSH/MU4oJvPx7dAuPop
YOMHxKzzbl9B0vQZ42H/SrsfM8tQFc6HfP5WvBVwNl9wQcDXWijEbzSyjpqElOcR9X0S213+DSVc
h5Z8Oy8czX630lYyY8S1LVDCmd9XikQgfM/KutN1Si3ZvoO/xiVrheLpQ1JJnNFoma7p2eJarUIP
eijVuNZj/IlPjqRiS3NHKlC17DqGiO2qHS40EpEJhMpBYqL9WC17LVn5WVOS3zbCOxLaPcAQiu5r
RMkm3rzN1PiJHzgg4dlqfpkzCMWNbCvuqv08ZIdX4p7JHvJNPl/9XgC7yQ0SJrvWLNmpI59VMsOM
eNuzrqPL403+vPIbA7g5s4RbcJwY+wRGIoNNLc5YuUYAaIQ0r4euNo+Y7arZHSRrbm2UHr14kAJw
segRI7WH2KMt1KRSnKqMmT0yFmsZhu0etP/NzksUgPDQAAFNVJaONlfgRNEFtXfk6IcxY+ar7ZNX
pHvLapiaTCqrhRAS+BCVxejqvkXHvuC7htSeDVeZzqE/TwvhzILhXJuMUGhr+GdgGlSMAzFXW32i
iRYU9L4wEG9FinIg1plmDyUGArGCYQ5o3Fedk761/q9J5QdhhBsB7WwbufLf279VgJiejkUGxOxm
a1RDn0pV7IilF1ivAsPO0Gq6xIkgJMN+C0hLCmpMKLkc4UfuN9S/9eoqhYPdR99gP2Ki2Jggnm+B
uyGQ2Iq6Tr+jieJYSony2MHB1f2MVifWLeDjQrEjyuPtdsEkQ+t94GH9Hp4Tz4rgf8fSwoVn/i2b
Trymv5W3CNN85GLPmsB41SZdpqBiUWji93Ss92PXj0FE1Xh+qu7Heg/Dx6Wgt555kZ+qqLtqTyJM
9JDkk5iK7jlHyXQbklDRgL/dVYt4YqzvjXqqQ8bmbaWP4a2el79DMyJRd+u0CFuznyP8r+wiTc/v
Y+M/QgpGAnu3zVhuPv7JFLhdtY0nOIX+c8jlXdikZ+yE9i3VUb2q5qZbP5ywyT2e5MQFds69RQu3
UzWT1sGa7/2PjPehGCdwdoi4PhqSbOiTqikBvSmPNkKbF3eUpDuIxtLBb9g6soygXaIHqPCINdhG
G/PpzzzBb+CRrJM7Q11J2NXsvGboRCOg5Kk5Kgjx3DzRio0YvEzAU93qO7Sg9zetkevQxf83VdRK
7GYP27CS407eshMLFwg11SS6fG+PUPhZxpD/oWnd3yDX3cVsXlz6q0f+xv+iHmSJ09XpH+usszz1
4w8JpCnybyCrIscSOcq8XLPRNB9+Qm2nuzjW29WNSOWOdfGgyfilTpmzdnfobOJ4+AxCoQpy+IXr
ypg621Xa2Udwii1kBH/TCKPFdWWrgcC5zHnd8q3DPLxrMJiJMJnjSCq+K2AgJoQTTXDoZQL6jKzo
KOX+RvD9bn6drfHYuTJlCFDP7/rbAceicKlXwYBowm0pIpHVhukxGvmX6hYafHEb5wrgR1zoYFsy
Xm1zTvOUbNAMOJVU9cqp8B94mXuKwS8EMI10HhgxnWdTv8qWkDD1acsIPodTmLgCsjL9jKMJqU6B
s4xNmG4GVAtdxVYTEoJaQx/tPi/N66Hp/sN/46zTgNiqq65Saut1WmC+ya1N5bV8Zuy+syTo5qc4
r1Je/qD6+nQer+cLs7LQabgzmTQfvF+j70T/H7X2HXQRtNVgxtIEUVykEWbPZZD+RQj64mRNV7fz
9dDU2SaNqD8QROXoKV8u2bHalcMCMPPO2pY/9Hgs0FURTiHD1al2Ifp/yp6dZaEGzThgJ3wt3Acd
T/NCw2uhwMInhtDWBZE10OREy3arKBLxKvHH8GD63yBGTFwTTuQuCzclAGATFe8aai0yOisrzVAk
fBA+KPLqIPih+pIb3dN27RkrbHDtY+Vsz4IKV6O4a8fj2zcIc2qSZL8m/Ae2KKUnvywiauSzlWIL
SWSa+Xt+dZzC8FnuxZXQHNAjxy43fua3C+Qd9qaGqUKdciB33MPnr59WgJ3lrFiVv1+XvcvZehXV
J0dBisj9m955VaRfixz3KD6PRBURpJOjf7N4pYyiTaIIVq7t2XxyypE6EfPMFMJr/Ms60x2U6cwd
GkNZUAZo2Zw5csf6Cadq8FLPpVHAJGVuOFB6NyBsCB23Qui2gd3oibYtC0nPJTXOVgMq5Rj7hDuM
xn8x+Xt4uk3JK1J23rTsvgHPjyzlXD9ZO09omUone/rtnM+pgXsta3ea0DWMhGXmw5iKuGl31srT
nqBk+wTns4kq5SkNR9hQ7HM57myQdNJrIXpaxMsQMFz/lJyABrsJCEBkwvPTTzywQRleNtJAqZvB
j7j+ehx8VSg9gHf9bJP1T8okBTE7hhGQjg1fkOVW8mMIg3x14AwKQYJ9hP7YpYgTJqXboq+0ZI4b
Oq0a4KdMAr1+p9M82Uv8hjjpxyss47yeCC7DIckyKGe3LL5ktX+Diyj+WP8iRAMux0794tqkquGd
gFnou7PCHuqZI6t4L4h+cKKIDok0+qEncLFQYwKbJTnKTRJ5aAXeupqpsPkQwxQybtLOEZsC25lv
PqT9WNDCyIk1TayFOPMi7d22KcTUdSGRgCfIFzQIYKt/QLe137A0cKg7cfKYsKQnfnxk0rg8tHr7
AytgBXnVgGJ0YNHzXPrVqC575v115mEI12I4hnHEJmWViCllK/DfjY73EPr26/ObxMq19Nlh3Vng
PbCF6UEcN8PbHGnpjV+XJTBTZsOF6y93gE+y/QBKUcFQ+DQUFZTYEiur7dYc4R850hu5X6zs7AU7
ntDcJvSXcL82ARGQS4L4N3eOvjJUHifXA9Q27R/02wnsPYRW+MVUlOONyXhHIoL7qrSwJ7kGf4/M
DRf5K3fFWBssbPjxr5dMJkSc4Cl91YVNvu2cDGMJPi/H33fyPgIkRQRqQNoStPE1RwU8lI6C/7BJ
kjNDYh94GdZ2E1uo8tGzZcci2ZNbc9Hbatr8w9L7Y9acX4MYwkaOe7uWnG5y3QcWXilC+FTk1P3s
/xJLQLAEcPhXS/l2L1uh5gpDnIPRZTA8BjKvfT7Ufy6MJV5PHR8LV4l+Ab0UxNDziai9qO+jyRdK
ufhEcokxiSTaAX/GZ2+fNtHBBsVJbZoLQSU0uIrYIjSjuWT4PEnp8t67XYts0eQi7plWKkZlpPuk
FGunNiYnKdOyXtF904Qs1pCLXykzsmZQ5l58432XTeiwNiGdmWwrM3YijTg6/wjtbFyfnJFmZo2n
GYuL6++H4gtQiogOWUrKmHgPeUd2I7X4fwfrwAhY0JDavwwRPNxQK9CLQcX/IV4OcdDuLsvUUILk
HF+RhZgadMEbaQRzXfbWgv1TORCPlcRb/M3tFrxTDV/b35CQOrkuMx5WpDLdK7g6Pfj7wAr8gHuy
VXIl6UgViKzi11hKbB/bRhTmEWMnjA/gQkvvPv17zIFB+do0vJD0xO1gTHNXO533h4dKcigaj8pL
TOkdC2Mt63PeasYef8LX/3kYeb/yxUuN09IfOcxlvEnS3fiHDwFSVFV3kClbEBrQ55+E+Ut+CTrA
QASvTsbXp7QvMFhOvCzoYECJvPbB3Cl9B0rO/HdaF3LjL2Yi5G7uFHDXIlz2M9BBGdBk6TAdZ9Ui
pI3iw5pRmZFjWmP4zbSBb7ep+7CWK2NL1AN2Y2hMrhjTN5seoAI+0IQgYJus13Oky0loHSAVX+Dg
YJDmEO2bZOmkE4sq3lDlWpDXXH+G20hWrw/CjtqmFNBSTB1RLfpVBheOeMulkcYNJcC7l0m9QtXp
RS1t3kDQ+Lc2RiZCB5MhLDjZza7ZZ7bn4fJNIaSK0R3SVEAONjr9Pn23z7qBMoGBDxDxSTZg8cp3
3YZYLnlssZNCTwF96gJK6AMcHhf0zwYgUrXkFrOM4egrmjYkpfh+C6imt+8n9fhrs/+OErX2BZ+H
C6vMrMxOfYWa1XA04JDyMR7OyX1/LwIRKGawoz7Z9MW2HHfQJJDNH/oeVykXV2bLoxj0czJbGrVU
/0ahov5V+9wyFOCm6RwoF0OAulBQ3bwPJQ34NNVn+N46HwHUpBwjEqr0XCjc4BOwQRh0tbaYurs1
7rcHkAOetfLxbQI5WpyDc/5kiGzlRjBFTQqPWJLsau1/xVsLRcZkUUGpRjpKJGHr/zR2IbPYOeUH
IOk9uKqFFb8Uu51kS1c8sf82AMDdGz09dYDMXzPbYqCMkyYzbNCg8eVj5JnrpZf4quvNIUQSX9v+
swZA/6kvwVJojfJYiSV9474SGKi2d86zWorXtvoEvHfd1snur1K4aGNvwlwbF+UOSX/b+NhlDSw/
Zc7E2gjMJkfvOPAiSBnriHkEhW1Wajvz6c2Gp2XDNCrTmB52ImqLtvFe9M+y9BZqfdbFvdG6gbhD
UfZu2yzEl5aLoPjobMLNO88nKMhM18JNrUk3fZik0dNa2ttCp54uFTiLWrt9wGu0lHMX60eQnyS6
Uia/V6/dyd4ezQ2jnbwxwyqqZCJlpNmdVHqaShcmMJA4rh+6QExjHqVaewdjeY6qWl9bjFZvYPNk
TIQ9sIc5d2yd3vLcJcZk3taeN7T+dzvV9KOqHbIYY3ASZGKm1nhRPX02XoFUbzoXk8PewWxu1b+Y
DMiiGB3Rn/yvu16Y9nhh5SWpMRgvIPOv39v3JW+aB23e+yH01DhQ0g5zgRwtK1/GuKo+MryU8gvy
u5pP+OvptYCSQ1HttEwnUY9bZgWBgIXdaN4bPItGTIfWEVnbhFLypyJulOVzJRSTQybwRIV7wr7z
BwZ/0SoPo3JqDQBqj/fnUFL3pOqoI2ri4273FCxj11XjoGo/cseAe5pEUgqguF3CPInXZqdjVpqu
GGCXeOVj7J7EBxecUagd3Ub4DlE1Ncbrko8pIGNB5GB8r8r49FW4YmKTIgLziYKrv4weAbPukWtl
GQ5Yi3fKDDmB6ATMOweZVNMttyMLsrnJZO5lT43hH71hQeQZYnpZ+Mlt0ufmJMV52GX6fKE51c/U
S9KGtmK2bjqL6FF0CXI2xjZkLWTSUisFUJm57QMUObB2F9aixlMoYECvwWizwD4GNKVt754gPj72
wFC3jiTUbe0u52x7b9upNs6s2yo/X8bRA5uFhFXMMDtD83BxZHo5gpV/628Rwn6qAUHyd3MbFVUD
woih3TjbpxAlz3wUps9B4L5sQOjRQUT8vqfelElHNrueK6/JEIEDDmSMw65ZGZUOQDrexVAtm3Cx
BYz15HWHYWEZQSsABqjom2ivqVDKku5OohEjqrr7L9vveSJZ9n7D6wocmne71MHIwTypIk+aDrbX
uQPmwXf7LXGgvC1vSmOeTZfgbvVoUXne01L4izawbF+A4LfEIA1/cPoVfP8MCySCif1fIKy64yOe
/3VtrFc211x8E27j9SJ2dyqb+HniHeCspUyrwr2+r7alt2ab/v8j/D7bI2JMnhzcXLx1VUH+NMTP
JEWPFQpTrMJjKB1kgZ4Vsvr1kv1G8W/qDXl0IzSetnxIuQUC0ar8pWFrGzi8tDDFssN2CWEsrGBn
AUlzTH58ek4lbjVRRGa7YvtQsWM3CmNaOsRLaEb8QesWGmDlnst5bCfQGc+1C5rWJCXTINwHIMcq
92ypnIo+786vbUS7y0O4lQX2R6N1LU++fwbfeSVMXBGAHwsdyX1J7hwt+s0HFmCQM3bNrS+ysnoA
6JEjKBqhQiUh1nzhMDvwwOvwLsYwn9nQBYNWZPjBJLR3fF8LolGrr3W9kg3WdEWJWIwPCdtjG/Qu
iWKxHfBP7TdfeuORT5B6zUXCo9YADkhr841i02m/6cyYqDuFrTx7cNLovtvGbgFkb4dT4kCZOpGt
uoD6qNk5JRpXCo5DtofgnNDrWJJCBhSSPj1/0o/2Ewv7eALp384IMsVsX+3aM39jF/8zAanMopGx
o5hr7xBxNejWBfSQesTuMq1N8cbk4owXgn+vl9RNdf9oouv6diUQdNpzAZfwQwN8YneAi9r05+RK
kFfI9DrNCLejKqlxxFZGx91n1Ew33hdH08CaUUGU8R20Ye4oJ01jg88ik9xBkq70u2abg8C2+DYS
pQrX4so1lw8K0NuEJeCcfQOtDmU/r1NkjQx8yqFpAX+NUuQAfe0yN572r4I8kYhA9jUKZ5KIutxz
pnfInfwy/s7GtGEz67K//BHRhbZAlFxm0Pi3c974TSaKZT8lhTxFXvEyQ8dBQwnYBqT7qjMyVxP6
XF1Bq0hULLX/8BUgLVZJt2kbtATUQcl1tUazQOD6h3MWYxswzAUpOZ0gFoU0W8JFhOU+uvgDVsVp
LKKspADK8v080gr09xAqs8VV1MFJoVqmtCb5WuNOCpSRY3dIX/RTy+s3X6JvnfOI0ucbO0iGZ5GJ
8bWZkVriuv0dVahW1dvkIMSgIU2lWuLvvH5xS3vcYXFOWB4gBV9oFCJ8OpD+g/uMK/l8sgkT1pTl
D9N8FAS3Cc1gCnGe7fpwDotNXl1RfiA1C+rm+VBRvC4lSFMdrlvaMsKjAKWnav0UlWD9a5/BWW4p
OGo2avdBf2KopfxzzIkdNnfMrlCpQnzgHrBHuF7xIEg++KuFLRNjpFwr2RbjEq6Z2yn1qNPgQ+z8
FmazyhnnPZkxW+1xaWm8HWHTe4YQ9pnnHbPlM3wQ+nk8J1x2UT32XCq3FiW9bc3XS2p2Fq7UAYYG
7CgBcopRCWberHfVPQWlc0aH+moKHcVdppWnqZjziHUM1oentYECqffnVk1V3DfVZxwRk7gLyKGB
nI6BkQsnDGE4TF+QHUosA9mR5hUpmFw9D53zj9oaQpHSFKFeC99cZHvWeoONBUCqSZ2gLiunj925
5UAoBUpvsDkht89qex+s/cuEkD+8VhjiaBiNSJ2lFVo673NbwSJk+5b9MEudapX7mFuGLQm0XlZg
YobVBPrEFFeGFMsiYtZHa9hxKYZT/io8sm37o0uadCKdJL6ZzxpWc3AcDVb6llPEzG6yopZ1w720
HKjUEMxhsP5lC84tEr7ODiE3sfXWTyePawf9UQTTYvIvY5/xWb412B3DXGNe+MQZbESlPUJbNj9k
jWAFvJOHmUl3TmcdfrVhnPF5H/h3sPvH+i4OM7UX5mntQrSD0UpUHFYkoxGH89OvGJqZyPpKNvcj
Pn1dAAvMoa3BFq8qYg/w9yRil5KhiC73O69URXfXpIwowbj0cQdCWM09xNnpO+6a54pdUsJ5Yn+z
1gBBLDylWx27ikNlLS0yid+1EDMb0ymlD6jtPGjdVLNw6sp2IU5K2m/t2TwvS7CyO129dJx5QWNk
LYoN0/Tb6vDZ3LeAlhLhOWBnKgBulBi8GGBUIM4qWlaDSxxS5/dE/Mptxi4KTTw6JBsuVSEfUrai
ub4fa2cPkotc+l0vPn7wjPburPGda4RF/CUsVOUpqULlb0yU+/rPTwr/vkvlnymitW6iT8IDrXHo
U36MfFDx+cDA8r8tEIjuRIfCsF1cEnEq3b0KbzCxVlXuNE2vEsvLAfwyC0/GH16Y8YR5qCtDcKji
2Dk1WhaJTz5e2Jn7iP7SYf0A751IYY7GZdcbVkUX1LFwqM8jKKzG/A+xIBxrJw5yiH1se3Fdz3az
gySfu+KSToo9C+lRHYkNKSZ1xzPt1KdWc6LB/FbjAusbREPQfKzYubPlb4nNlUW6fCb8v2X9yeP7
0Q8c/71Theh4VDxZWHkKkzrWRR+QTBWjfRCzmV4/MDixtMy+x/JJP89MnX3pi0riH3S94R5ehYOT
Om9aO9ftknSMw99Adu1/b9AxoBND2TKW0arNWZCiI9efWWTyJZrXdq+dvCgRfOj3THI7+A41vd95
3UZRpNsOZx3kbKEjVtcaZB0UZdZpq2vUZG2E8Q+S5VBni1j9ZRD4ddQF0VIpXFl4p+p7gJrvpRDv
27MiAPRwI8S5qtAF72ROWuheMb0OTO2fdHRveOWiTicnsJguaaBfCgafw0wWAfMcDxcbZHQZVxa9
Och6sfRL4djPzwITZxbUAFZCsIGYGfCwxeprr/6vGCIRx/wQmM2arOIVRguhbTzecStOIsgbzvb8
oTJUJnRmk4D37Or4mMeUaXprZEwwSLS4kvf6hVpC+exN9yk1DbSLd9tm/QrU1aLw9oOrTZc37PLv
WQpHsMR7ub1Xro6HEFzXlYqXgpIYHE6cJnyBm4lKzl5MbCPwrhnrI6eLupk55sTgo0bZp2kkyunA
dkS904gjkKnwtpwGljA5pS9LTM4o0ScJW3HbLp/0QYfMBlGQmog528R96aLozrWOWlONsJCg4HYH
gs+YVzgXP8D5/5hnZ9N/ZE3PkF1N5OQW+UdhMFJSMw6+QJwU5PWkzDWaaG4HEuQCR0Fh6nP1IUiZ
MiWpNclvdpIO5SiLZLyLHSeM7li9jke2JpcXlQM7C+9otBWPtSLICcucr5G8Zs8FGg4/Z6pIAtbN
dHBYZOKBl4od/071s8jre+uqevPva55ygxuMryQTiOpswvI4BGHhv0bBSMCeD/U+WG4lzwcKEnyE
nccHhoAY9VPYd35OQO8CE5xllXyYiy8LtHexIXG/F1Iv/d3TqDKCXUqBXozJZ9Sh/8U8ORLKgUfj
GL3Q+Y9ehvIMKKGZXK9vg5bTHQU3Vj8ako10Jf54qnj2ysKybFvp41nty9YD6Ql/kIu5CFTXsLG9
kdmx9VNcx81KT7XIs10CmgmaTPJsBP07RawdCGi/b96P0ex8SStzmiFx0xqtujXOEQigB8nvyrrP
Gah7UonsB9tbb1lG6VrmnzWnTyUkZ6pEKrvcrmsduNqoldMe3iPFoQIqqt9AdNLH3stV/ZiW5KYM
uoN4nSmg6TexIo3IPzii7xyr4h0j1zuI3Tc1lisp9hfIXISDISrGNfIsLByx+q1agCcPqqqsdJmo
7RHw5njtTnYfDoR9Tfk8A+qqNYMSTvfYzomC/z/gOmO0jD1bYt2E1DnKSkWn4mrT1drqRoRRgUGA
knZDGoZRlRJwy7YeQm6YLb682msbIIeDPFxnIJk6ObwUBXIoND2wFeSBruDsTouF8uu+pdCGMeNe
+fnFQF6/AF3Gm0+WFMg5O1rxp6Ld6YHlxsYXZCS2mr78REIfq0zPzsmkjOqln8DJAQEr38lPR8lJ
HKouEI2AsmtbOEJXytMte2gMdNlQ1mbaOXXVsVk1AUuKFudXvzaQ2+kS35HrvYOcZb3vNIRQi/Dd
496D1pcNAa/k4nt0ioiMn1qAdwXVJA5etojdKZNIgYW8mSYj55ijtUauFD17DP5U89g+MR6lbikq
7FclUbA7crogAODaxfdQKjvn418sf8xUQg0QnhyeMQvsJ68Uoe0GRe9b1YXUmqBmC5PzmeipM26a
sz1p5VSx12UwFTGq9cmdNm26iOq7dCMdEjcHcXrbYFEFdtFe8D77rJTLd5n0ec1UztvDhE6Mwo+9
iuDwU5QCsJlS8YnzaJCxXxAFUdO2Gdt/BovehpDAHijfYNu2+CWLNNlgCtLSW/dKzmldYz/Tddt+
J7nSeHKz4SnciTV3nNL7pANkQYJ+/ropdNg3LKRHfNvp50nfaLCVOcFvXZTstTtqIwPBVXJ3JpCG
0dLIOpybapKSUr+0nf75F1koOFEc14PfxmT9Gb0tPm36l7DtPZa5AILYRAXiNoiZsYW76BANc7I7
UexfKO2/EA5v8C+UJzqDOt999bjdDfm6ke9vn5dI7Tkj5NrsmBW6HKLegAkNLl9r1KKN+uRqIpFv
VHTxyCKXUN82D1qEIDLRPD3eR9G/Q+7Gx9tTxU31goKsIiZb6kQQzxWQxdXck3qQ7JfyvFYHdv9j
Y6e5Rs4gFwSsDkz6kFnuW6cQQ+R1t6/uzO4w0IccOjWx5c9yOq0FcIbBhLx2zAsc3RaD2YaKwnnq
AxlSEGKGL1AoRr61SCR1EBdLtTUcA5UF4wrd0vig1IZButN1jUTyuJOy0G1hrIaICny+d4SHjdzS
AIfhZpKEuZdmz2xxyCu8FfbXmf1g5tQ6vgRKsjlcsowIpJ7A7VTzIBZOOwvLL+4JlQJxD4lrlrdJ
Whi+OYF9u+uMs2olzcghC4GgZURUZFQZEAd56JaAUOC97Pk/fop/8g3GqzOfVnM5myFP6v6ZbJOM
b6z8lzWrdcQNLS+Gd855nvutHnl1wAot3De6WIteVAMTwV55L++w8lypA9tM+hVVwkvHVHsBoYBU
E9B3HWFXGTfX4bVNm1P45S6ID4uZ1SJXQa93wgfBMIN2uyYQmRlr+e8ydcgXTw6g4axb50Us2lpp
FW/TJQhRRtZ89825hv1+T9HRcHK8X6G4oWsYKbZpCXNNTdVYw1Bw7Mpv5kOJsnQY2tr+srmX7IV+
vBPoeD6BksljmvXq+DTb8NrA1Yxb6OZUjRRxQliqgh3d96Xnyggg3HrD9wC8loV0dBySnO579zRK
h7x1cKxUGSkc9LDv9r5lhL06n4xdGzDnTzePaXpLUmrrsHYo3fd004joupMlmsDa7cAnfwu5PTPR
ROhvKD3ms+0Li+UwGpm4+OscXSyWncixgmAd8lnL8hSMUJ6rUSyrg8QHYQJAJWz9Gn7cOMRGJKeY
VusqouxLud/SJHyyq6krLElsFQNH37rZLr9gytoJhUJzPHZLdV4XNt9R31UOW1q2uHnwoe/YQvDV
W/UFtmIh2oCg/N3GH18uEVowk/qsQE2OPdAfhjCu+A/wVWfHkMb3KAHTuZeb34UvX3Ca4AaaiZgH
qwz4ts+wCeLMfm1pai71ApunStcwNi0gulfzWBK7jzqYGZ57IaAKLzCQdqY+9DASAoH1S1SwJU09
VAgetUxsCOwMKxLDUzFR4BVSNcMq2oyhUqe8QGofQN4OGEDIUX62iRYERh6DyehrzbVTEA7Zp5pW
WjX78VioXOsjgh3/RXOr4SuHb10jLh4+Uaa5YVWsqIcVB3YAV8P8jb/Gt+nk83u/zFwVIGBB1yD2
sjDoGxvbeQjMq+hnCwG4a/mqSCnSOPiOIJiRmQuQb6cRV0EIKi7NEeh5aYkAl0WzL4nKZ6eIliHd
jKU7rR0N2UqlE8pVAWkU+mlYRdLhlreRsWEDcfn7Bim50V/y4u7Ftbu9NjLtsub1o3UBzlC1qQIO
K4L79z2gX64bCIxqJ3h+tRLVNqsJNNYCe4w0ChxRnDD9haNWHE9F6R4zGj0FqSJbg7jeS1X5TkW4
xP1ZJmNev4kN8qyOYfpPdq9UBA0VVuG1JCb2IbNlsHKaO4zZ6i7ebs5QjVPdLLGbNM7hFKBRVCFa
V6Oq56pNzcUjEf4l65aPOIS/l3EhmtlqoNaAPxLlZWpywCcTCTmqiLMDOlPExCqj+rGtoaQ/2TAg
laQp5oMlKvkvVUu9dHmupOExjQDr+W3WARpHVp01DI8cW80KrUTW5wxAlucoikUGVQoF5Wr1a1TC
ej6gY8ieMOFlvBELGNY3qgXqWvAvI0t/RNKDqLRNhiT6bGkLbx7A9wueH5pKSkthqhssFggfSESx
y1IrpH3PbHgYTAnhd36uS2MwM1zTmgncomAQtH8PsVowB2QZqergtxCZzkaIoYZndpESOdfF6jkH
ac6guCccQnRjwkhpfOWLSNCgMGHx2tx70TlkpGWTqSzPivIUyiVjnurh/+0UxAjV8E1KCV3T2ZaY
P8j7NcceGQdXCkH/sZXPgyfXqKhI43oOZwj5TX68hjQ+scvEOYeKzrgF+i6z+XMYshV2UOksgh6O
7ZWI1q4ZOl2b+/kn9VxQCgc9xJ+AFWtnbT2iydbFlCfIe+Dk6L1g/l+FiCX8vS5xx0eXVLrAsFZb
TjE+ayOBM1NQ97MVCDx5EgDZzjupybtGjTwDB3k/R8daEwb/+9lVuMusSeGGGWxfwo5DLTAu36V6
ljd5XoLqvcSYdwPvOOfHAN91zd2ZuFRcNXd7bp9KDlFPBqHwlBCVZGnKhLO5BKHyFAAN/5UqA8oH
P/cpu2toCHAfOmTcd1PBRcO89KCXjPYfL6NIXeTGMsCAF2rPXUncLqxwcMuseM9y2C4N8DSeqoAH
3O98QOqrVC95cizty2g/P715g/pmAAaypXx0Mh0zs4gS5RZHorYpxJaHvPnj8jXGrJ7N9+fGcfPe
WuKvLhyfHCfgZZuOkSpNhk3ba52yCpVklZataLq1o9tcXDTsi35k9SbUm7KMc7QzFBIfLTVZ7Sqe
2nQYiRYeKLRc97gq3C05eAboEksUijICshCd8TjihOygiHi0HWtTVA0yl+tdjNHR4xBuEnLQNd+y
rdm7LUaYnNAOQvmIR/9KL+S8ZomVrqD8AbkDip0rooWeXRGMkk4eHawnhVBq2InSUXJgX3/7q3w4
bYGzkwNlkxwFhFPUCLa0wRaJgzbiMU5RDx0/4zeZeSDl4lFbvRXtjkFwKMsmXotGPwx+/GfhWo9f
Xt/5RxEMxozMidr7ytchox3L4XXUYEt4XIaSsDQEufjT5Y9uD9Fm532EgyHGw94vC2BViRc+lGwJ
PYNTBiSuEVcN2ZL8uVtkwYc7s0+q9uVD/O9YvdfuTLKblkOsbqnSO3+s3uaykpD778kGAOGvVQtb
a1RxhZyB+Lu7IjDsjXyKIebPgPZZ4KvzzTr2xjm4YmvLSuTQJdUnUcB3WS+1JeOILAkZiWbKiOwN
Tt6KPqlh+TLnpx5FthtAd8pNQ3cAz+dW+ybqON2jVXQLnij461PnZql0jfJc9swx3FatyhIin9Xa
gvw0K0FRSgHpfHdgPSe9KZY0BGDkMDG8qcKFvzpT48it/J39q7Vj6o90QnVWLYXzBLVb/b0JRDj/
BbV1bVtIbl4rEgrvQsjOFbmxUra4TYRyAeWh8clx+0QF6zhdK5frPm8VT8oEqS1w9GogQQkP+gfT
XXke16MGKVFMtzI7Ej3PXD0Hu48hIxIvaikkHCQNkE8okoZ1gfIy8Al5mRrAD/sk4YgBlFpZK6GR
SzbvIfgOSxxpMrzb/dBqdP1yds9kdtV0K9HjCAefB/HoJKpnyF/i1rDPEBV339gpnU7r5zg57NuV
FsL9lExLXlHWOZO1MxTCH681cdJXhTEbLVRJp4cLlJfFkv0LiDxO1u/IbT1v9Q2FgPMAn+2KJvZJ
voWOSomEQLifaG/RHWNN6x38MImYxuhKnUHWSMZosZ8LlT5KavsWDOPLoUx6xnpEa6uxGqy+I5VD
aQSjFY7y4CgG7pr+b43oNmGYdTqMDrjI785m+Loa2/R3m+HsWdzY2Aonsl0L8KXubAfYTzrK8Jhu
j45kGt/wrM2PrhC4frTDHKYwSiVRuT0B3j1Fx97kOP1QbMU7vEf8QQODC2YI9Y2kXQxwbs0p1lzD
g/JMSO4Ht3bZZr0Yjx/wWe2BHO1xVCmvtnoIWWwEMaSSya4xWPMldMaEC9s8LIEgvkZEg7R8DzD6
Ct9cV/nSPoCrUsAurSkuNH5dbswNeR2IOGGqBNvpXmcmtMY2ILf25dbFPjErpsU9jadbvCGAnHPt
Ye+63OIIV+3dUQ596zM2lNCfnOAOBRsWR9AWWJVIsznPmLAUgfAY44nEWgKv7+pgsoEqNEM6RUBE
ONQ7C+uoUs9X1XrsHZgWI/Y9Zv5rPpWOIsCb5AQeY3wkgXvq2Qj3t4lr6qzLaxmyJQAUXbPxGUSW
F38SLxBjWsDf/5gkpT8lpqt+RvC925bi5QtxqenrNhSS+cbVzCmGaQQBxd/MQPWRDZVH//69GfgP
AmW78BD3Fc1stJWtj5pzl4TnbQJUHhBv0JNGIiAQl4htdQ4khc7qN1WSqKX9D/KntW0ViCFWddXX
Sl0rFkjxSKtwMxsMhgGlnE54VVXmYN9Op667inEB5w/0/iyenJFWs1lXCufc+f4AjnaS7A+Sb1j5
O9MDVqQAjkXFaIzmANKQy9Wysk1DO4iVFYcmxSz2hLsO733bPeT9rWaIdwfwZA0+s2HkrWQnly/G
H0IdbL3NEq0P/6zKeNp+k/NXTl2NaaLvy7jZiXnI6Pt2gR5277Dsbk9ebcqhL0FnpFtifUV2dCjg
qykGrRDeZAr15hdrgh27iMHoGkmRtk974YG24jbEpSVfglT3aJ81qDOvlikR/HdA10uWNeoS0QqY
Cn54o/NqYIHFwaMGdWM2yuVD+4ZUabxYDqhAOwdciD9QZ6qDl01c3ksoHyPw1/DQak5enGewRJGn
ShJylzOcY7ioMRLg4Udw6sUq89J22CMhZZsqEHldY6v/kkFnknK/+xzsgo0S+Np5mcLDwa9Lribb
G7GCfWqWNOz10USmGeZvEk8jA/GdgmiIjtN+R4ePzJQT4nqM+v/66KmhS41F9s0BagxLqJXZsjvV
V2OvB1DgWfCCkQW2UDM9a9GoeKFWUw79hct66BWH6542oGJzd11Nq1uchjKvMmYQd7+8xqqKBpuq
6LZSkeQLZA0RYlVcfRRzhPvDBCr1auPfbUE+AgFz9MeShR0fjf+bOSy5eW9cEaVmDZfFHCf5qkFU
41rltdhI5h64bChYwYNhmn65bc1G0bjs8rXjX2u0yxpEaJsK7r0esONQ3HQwn3ztvGwyhTNegWkY
zYd4E8Aus/PzK4pKJpQlEgIesCV3cnZWu1vWuHJE2ylam6vytQt0PHo7rRlbfi0Q8Q0dsN5HOE3X
WPuEByLdQuIqmRNPfguHgNWxzioB+Tnrwi5h/RNUqEePJNRmS+lPRv1vIid3UjBW0DCAuFl33yva
ZQQTES2Nus1/kl4d+CEZwsp8BxcyKxpuM9hl+3gJrpEbxkPqPYyFW7T6DsKlq/WoSYE7AacsT0W2
c4J6PLnbFQpYkhE34UXXl7kkvoJz2xS8LJavwGQ76hnxZ6ISG237aGbchitG2Z2hGTHkHsFyP4Yp
FBbu02MuOn745VwzAmpE4Y9JnmWE9tGttKcBQm1gJjjqAThn0q/cc74zMK+wGGzfNnKNYdmy+Rzy
tXeg5cQIPVCJ/r5Le0MspQ71Xcm1djMSirdhJWYqTetoTm/SzJouYWPc7b72GsAEs/0pCiNraX9W
v4EQZR1e1Aq4XpH6T2gj6BdQUh7h85HvbEmM4+XDfNQY5G4HOQwj2Ha4bJDQ13w1FndRCpc/zJaW
Rq/asndktcv02sLiDWfRbi5vQU3+hw/l8jOfPetkQnisD+Rdg2Q1ozZMoxwAzDHBv/xbCTQlUXFZ
01/7fFHkUsUw1RboKbhKIeW4PsOubAv/o1pe1F4JLqxzJ6lWBcchpNAMgxfGK11FP1w/7S7RXOCy
YGE8xv4sRDeeX4aWAGgxKb5JeO8y6k6CwRRg/FGh+lq8d+I6zbPD6X1+LOg/zxYPLqTSMOFNnkM7
3tdFofDJmp8Pg4Tfvq8iFAk9MuFsTqyeo1HTLT7iQhAcEKk9fJbyYzEK6ISq+4xuvPyHsXvIvf4G
VV0V7/D9ZmBBsjEmz6d8EKp4cPi70e62DcHSdWncNnZ9PTsRbdglQ1AI9A50tGAUhxbQ7hiNSOPG
Wmqg2/coyGO+Op87dmjJUfeGJTSRnnzcTp5Yrw8owCjIBLvVJO1+MCmAmcqRspnncGxe1KvRxSl7
nJwjioBS2vW1k4N1Wx3itLGENnyQNeMfzpg5HUVaFyFPV2koqKg2kPqDzZ19wHWT3HXF9wWp8QIn
3NeLCGahAngJE0IZDCwVOX9L2MRA7xbTOWsYESt/C2yMaeYmXRMOWZN82vYrULzXU6N1Mt6JNlOs
wCCDUbi4GqDl2+5k3Xvz5c7EfCx+cX87fHiov4K5zO6Mj26KUoNXyDiLQP+UbGJZXOvkBUBj75S4
oPdclqv5gSFHcgPscCObmKFlqr2X6Ktxe2suGb/fj8XmDKv2O8x3evSn+4XSZqcc7PLkyPSDq8NG
fmvjGRdC7hUdbUl9YB6iHgz5kgkY5BRGi8CaUNMFDupqnkqQ3/dxa71HlEGtJ0JjcA5OjogCH594
u6liP/84D+YA+2gfxO84Q23pPPoLLdj2NFpBJ8S4q5+FaltZdntAt8Yx7rZVUOBwbNqk6WD9rfjy
0GLwo7nyBLHLhaXpdTJTcm8iTdInlnioyPlAEIndZSaE7Y07sBcj3bBxG5tfWQVzFZoRNAo6S3oU
NPnEjqtJBNqI0QPXQmxUTFHwqKaRcrg9u9KdZgpsOB3T40a+yBV2UjCtMfPCyn8ZIbI75jJo58g0
KxJfh+Ya79qXmnNKt2TtJ86a66gAHgtPQnORJxFomDmdGqKysMW7VSiSVqShgcsAtk01nX6T10/E
V7zQR2FbYDIcD85D9TEf7s9LXMgBKee2FvcjnfO/cHLeXf9PfP03tR/cUp2JdmoSoDy7CiMrxVwm
jUEf9WeXe/oznB97QEPDVMTkqjDOdn7iWKdp6oGGnZlHkOgMFzeljq40U/NH5JLlRuh2v81BCVLP
410knpvGAyG46Mea1nMMLIByvD0wHIJnLasVDecmYp2W/qVwuSY421UasEl3BVS56C8WwEv7QjhI
CaCaEvvzS0SLesJDL7oCzxd7ZYiJxilCGabHpfS6nsieE9UBjgnrDNdc0YgrIYzyNJbssOCTt02f
lYEHKFdMTVp51JyRBszrxIuqYKP52GFBSyuwZnFaL/mJjZGW6/oksPVGGT2M9FoF4Q43UQW4SzhG
3FPhCbWap0xbTMGSB8Bwd3xYOIdExx/Lk4a0ed+l81Xavn/7Cgwi27ZrTnFMsaIFbppAkkFQEXGM
fAVckTVz2NHfZF+NpjeaAksdAHQxyfGgkH5Bs8HYEB4x2M0FbqQDJaqH+UEn11/iokbglfGhzK32
+QYF7/9CLeycsBTCgKE3BrM1fGZfgx7NmfxmXzYo13Yo05y1yw4OogVrQErRKMzZGf0jovyWwEap
yo/UK6Ar8GLVzDrYIjQUDhVBcLfXURuTgYNe9slySzqqTSmozw0D9Kv7vORUqXEHmz6FIQuzIuiL
Y2aZd8n2sb3I/T89bmnBfMUVXHa6Umg9Juz8wp1TQMTUxPpYLAGk2M6KJq8H1QfPesDte+r9HH0X
t5IXFwWF9Pzz7prKpF1gvXXr6hbHclbMjbxWu7dhcx4P+LKxO15Dlk5pq6k8z0WKVXeDa/0MWEvq
+u57rylQKxrZWzjFOruoURyUmt7jP+DL4TCvytTVfrGvSjG2wWP37JWsj5TM3Pa7pqF055+QhbZS
/Up7ogjx/OtQ6soDfenst4Hg9sSryi1ojEskGYoMfaOF75vNhLlt+xuMfKtbvPC9wq0M1mZfYhTq
O6W7iXWCbbTC7T1GkOfxtwf4byWNKu9eE85PyKbwcYRWgif1HCDV0jeugOD/5mbMh8lOdkrQTCh5
jRDPhMddlE/uNPuiDv+oyMhLY6u6TCylSHy9HgDrxFxYM5gk4EubQK5uY3BVejlxHaUKgSVmh8n/
BsNMkorwYzKJGypnYAZo7vWuUv7pdSsCN151rV9ESB4qJvWs+XCiY0KgMi2lxM6uz5RBmzBP1tUY
X/wdPTgP0PK2Bi8Hj0eze8f+Sa/dL08DLYl8ica6uKl9L4ZqDlEJiIxr8vr1l4zzRUrPVQAZLPJ1
IGI5na2SNfxDqbGkNJTCDCmdUcfsrWLpfFwF5UjgkiesBgsA0+BrP6b1tF04C5I3n51KcfgtK66g
SC6uqs80wWyfKrtdRATu9tZe4I/0usVt+3gUT6/pdyf6uYY7WV8yJQ/qgBifeJ6OLBV8e3lzTboK
OuyyVFUjR8SW+PDjKPqCs1qXdga2Mb68bYOQ/EMhR60ncSMr0UnOmRguUP3/v1rsCNgQoahXYYkc
RjMrfUfmNJsnoH3+zm2EaaPANu6Gng/WDRA/dFX2zcSc1KnUwzBC7/bI4AL0YjMNqF6XCUz5wNLW
eVVco8mn7hKZD8wTRSz6wB/2X8maSt1qM6UEc+5BQp7BJt8yZQLKbOTh3O+cloFGAOaQ3da7uXsz
+c/MuqhEs1aq7NwEJgHZlm6yx5X3RLD2QcS73K6BKy8SSQwXfBkl2NXftVSBfbC6zT8BNHDk1szX
Iv7alg589rldbv7QjSLeFpo1oi15RVM73slpVGX++rpohPuiEKEpECm2dONDJVoVKdsTxOPAKJm4
yz/F2SAzv1wrH/kmDmxfRLGt45U38WpmiYlrgtlauUKx9ajD6puQYGFv/QSpduJfCevbbWL87JYm
NQo02wXcBvjXFS3XVwwc/tXqEnj6SJogiTztio2zreKp9BXlDjTdaNTaVJqgI3yAwcZQmkqVZYp+
b2EvqqRYlYjamesgo62AYxNiwPbkwNMgehbeYilcqCsf75EcDRj9QrD1/RvGZ3iQ04px6pNi9qVE
sLmdhuq7wUx8bFJgqrSc0dLOuvEIxWyqIZuRuUIa4+RRgXyHTD23mX5cjyFVjgucIJX1SVUspWyR
bCIImZGuEY12zPZ0z91VJsNjW4tSUbWuxE3McJBgu45f+bBYp8ZzRNUl8EgoA9rVLC1QmuCqQxCq
EY1Jjj9T7e3z7t+1YzskOaRwGRNMwta+ycz982PhxIliQV6kSOZ4ic+ci/7JyWZ4/ai1CUd/NjSt
2yiAlegtnvoSKnqqy3iua+OX/stN+kGE58kr/GWNhLTHWXVRNQhBUqhiubI2Wc3hfHLAnHt1xsUD
fkaezZ8u3xtz0HKBuI85EzPZKK5eP56ARnzDbJ3L0cjHllzMW/K2GR5wQjOmKdkF8fRQ/cxQnJyt
g/MZxIuemjsx+cWPJPeiZDcgCTaSx5u1uz+LFrPow4euVP7NZUfnUIrIOuzsq+gSNbiwfkITjM/q
mVgnqObP9IxFO5UI+7HXZbk2hcBDweXz1TTA4P97nR4q2TNaXTDpI7N4YXFSZw98n5b9lxcO4VIH
qZlpW6NDQuAa0Ia/V6hliKKOQ+ByJD7LVaeWfPM/9ina7ibPReIa6lokWREaNFap4Ju8tKbeVVuO
BcAqa3ZGRFDr9wjYYcgwjMqXxmr4b6n7P+eVDlIRWCMlPGOFC3/IgWCpzqZmfZHRVWUmB0uMYD7i
NilnOTYC2netwYtYnSiURPXE79EYH2Wp+auRAjFnUhW+AAPNrIbjVf3e+6fKVB6i0a70MiYom0g8
/DEB0IZt0fgeocNj/yDZc4LFnz/XvBKOOpANJ4oc9KvoOWR5Yk2k1Ueh3IwGwlURAQQAScJeDvr2
ahu5tNrKdAxgS8vmB/jhg4DC1KX07CP7Fpt/KQhWZ7t1FPZG41OKq5Ne43KjnA+nZVvqVkVWKYL2
878axU0QUaiqKPWufVzOir2R5gH8r+jIn7BKIvtFwMwIEMcb6ljcxMsa8i5wfDavAMi/fm806aZI
t1bN+xlOq87f0iKo+HSz9PF5tKusSGyuX6k1TOJLBz2DZpJ0IY8d23xmuxF+pfvZLZMQLohgPMTx
1kXt/6kqRG+0l3wsd7tBdpyTScOp9QVR6Q40Z8TA7JDohpkVznWMOLCwSy3NWJn/S06WS/X6svbP
u8AjotGLIcEY/pY4AwXiQDIXW7ao1QHeqdHFMkFUhKNGP+IlSG0+mUsLR8k7ewHB7NVycKyVU2At
oC1zSCMeCsO6GTejGm//p9H5HVSFAQvb8Je9pb68RxGEGFYiIHw5ox5eA/yqZsOoB7ruwB3NIAyr
wyFbogpg2xXWyiykwNXzQwe4gKCes2uC6tDhNRMvtiyzA5dRKf9nBD3DAxT7yau35B+Cn7hu4NHv
lbPduBUMLLfx1A8YZzCByYMv0E7gxB5FGmymCLj2Mf/zhQj0UQ3jHnlG65I5AFKWXWgxAlY9qCAk
8fp4g4s3uXEd7jxSaq5PvJxA0sx5ELRmGPRhVS5/0ymaguH5ldEoDIdJbSPaNVjeunxBMbjLHLI+
lLTu3TIpVxIGNZ2Und0F37NFx/H0VFDZrgy8+8yLeUJO0Wq+kzCF2gQPFGHL0ln+ZRn1JphkqgIO
MEMs4UFzNee0WEOA44xXw+16Zm+QNv+FvI/5cDZalopDWLx/TOx/uiXlHcIB1WU4MM7RTuP1G21c
k5fdoScAND1eq0aLoXqalGGLseUTDC5CFdnXAunuBrHkkJDN3DYG8mDEABJM/p6+7mkj1DiO1nZ/
RkEOyKg/Mrm+CBCZddsMZAYL7g6LJEzyZTqG5+7odi3pHge/g6Rbnysm2jcZYQbrrUhGzf8RWrrZ
Ls0OZ7s3hSzLVXTSTuBPwd58fToLdEqBfD/XGGTg3hjQTNn/HlYyW3arjJnIH7Ba6rjHdBdmSHtp
LHppdYUqPa7CEUrC9A/jeR9pJBWoi+L1/hIEtVT9JYwadSZcaF6+riZJPt6gWD9+kPi76DoNWhF7
IuM5NzS73IDuMZp1DDjVPSI/qNFagQ311QotIZZ8J48SS1Ow8A2oaEkzX872BK/3q//62H4uFQKG
eoaE2dgfXSOJCePIj5tEl3Ju0MuuCNSAOxbBpP6TvnIYG9zNfiO/ZVxOLxBLMI3qhl9ATG4fSRkh
jJ3t6jBQXJUOCzZtHmscpmSRIcpaSQgP33zdU10mIvSljhn7NbNPhwvuLwEROm0cdt4QjGwWUlGv
KjvPIbdG2Nd6yKAPCTCDZvnotT3ogKlh4qAFuJJ92wcjIyX6PwSebWI8C3nq0WN+RbaaX1ezTN44
HvGY6zCQUT0Ghz0IFW0AyxS+9dcu9KCpCbkieDWiP0KxSL005vWzZ4tLgIxP9e7WMEKd2ZAy+unw
+SGXgyqzTVM6FotIuvJSk2YhR7Bu9SXca0zLWWHpX76fbU9sTnBjaboyKSsAngZCBJ/OGKhcnINZ
gO0tMJifLG+9uogiH72t+zifrdq1DXDL5B2j7BKCJZdxTBY65NZ0tm+SAwkbbtoWCAeZPx3kyigT
DkuZ33bv0BBiHpVHonXh1IElTswjTJ9q2f/R9DgPdpD/+6DfSvniFhMBNNOzfRklYlgC0kmFGFPn
9/xhvRDFAingF4NCIwDQoocsK/daxuugHIL6Qz7XlxU+buU8vn5Pa1dj2xKAE/zP6V5ZapwH4uAb
Mj4aKZZXru89qeSdAzA+xqHIF0LxQlK2CTzURj6v3DqtODM66zCS+/gTWaWMba/TrqHREdtXF4ZE
QrE9JZ+Wl+UNRAJTfDLqL7gb9zNfeZ1fk9y5NkoXFOEPSDrT8n8udvKo4PoYUkNDp4EvaiXtZpEe
rBGOSfKGxaSLAaAOuVuTo2ssUpHggrsPMSsjr65z7x2flOnpSx2tTY/RYOsKjEx8c6hzUGhw7xqw
iJaIqJbBduuzh3Xqa9tkbvlxTYxA9+syiAkxYo/HmCZoCEW6rzoDqm/rt9wjmR7JRQSlbCfUd1PE
Mqv1Y2jO7kHo2UJ8Z8oaqkAQrUtqnhswLyeBiSJDmunSgafo1IyQyaSHOYP/JUd2Bp86kJ6jDlWS
+9F09QIk2VrV3RV3RDw3j5sA6DbptQ3Cp7vLG4v87DTjApqTNaMAElGF6nE6tSMJWQkKY/hosTy8
TGXlos42pHRr+PTupM4yVNEplMUz2kiYcIcS7Bi8MTR4k/vsG4ukjP5VgfwP2QAGvgDVwQN60P7v
ZyUFuoD7tH/No6CH9lCzzdhZdm8v2hjxCRCZcKklVDfmfTFyDA3hcdeHFY8LhvuREczrHKrmTS0O
Oj2X1wsAbMaRg8i+YUY3iQurRFf/EDnPbFcIO7PJGTDo6Nz8wBOj7FwuUoybBUD3jFfntVzEqBNE
okElLuK6Qcc1DzEb4MgBbFvkSc4L+SoIjd4buFasevZ8OrOGA63KhIWusTTQpfsbaKJIzX817Unt
Z3to3Jdb3jfIiMfruDhw5DHEgeyD5UK4ZTf+LWLOjRtzXdtShaEKx6pTAAi4qTeap4h04nzkz8Bu
l0QCjPyMSK47k4T2Z+qEFjGnsnkQAAr3a21LO6zeXvdr3KYkhZrIzQ56Ia8VD5Qm26sgICAH8GNN
3NFAiR7FiP+x9rcK7g8vgmQAeixAfekHEyVq2FPpiZhdXWEHNe0HassMvZER6DuPcA+Zhe3WoUTi
+u7YUEZpnzvzPgS6z3BhR4OP6VGEx9MXbyN+cS1sAFYrJ61zj0sc3gUUB0KRfPYSrkmG7SihIHxw
ckdk4HwdyC4dR1OxSNjd+wN/ukONeWsQyTMLYzkrt0Q5+3txz8hZ9MKrGFpbyFZKwQskREPKcNZS
UlfUgXLM4sQ/2D1R57ot5cHQq3UgnCebqR+xvvX7I4tXjOX17XruXQo7DB25udgyZ3pB3Hvyxcos
falXrgIO9vsRujSeW7M5dSixwHHP3wo0bfTauhZ5flldXmnzdp96HnOyrBr8Vgj48aWWN6vf/oAS
IeVUeDjOGXjjEAMuxVSrdG2awUFP4cBPcWCoeCNTgJ+0pLpwrormGH+B2Ohl6qxwtc5rQdAdSbKm
0HTjH6f2FXDx36yqJ5bHkKaf8jqnICWAkPKj44th0blpMqNGLn5DhE8p2EW5YJ+kT9hbroG3LCMX
+UUvDgePIdPy21rZtQjseOnUKHl1w2fYR4yCgoPqUzxoxEowfn8akJsTRLR02Cz5DT6R+VEkDICj
J9GRetGwN7L87Upg21WpxKXoRw1swZunSsrQGQBkRa/FGLwrMGMgZGejDd9p022VZxUEUxJ7D0uM
xhRagLa48HZPBYfL2VlQxRu99KVPUGVb2haxTUlLNVkaBej8TGlG3al4BU3vkcJra9vYJpMXx8aQ
jbBIp/DohIUUD0XbxYN3KbR1v2YJe92jeWDpGYQA+V3wL9S0MDnq3mv6R1Yhp+Gynq6zf+b9yC8D
EGBbc3Vz1C3KyjbeJjOYN82KXCKFpS1Nku+YRnivKOqAoyLtoUQjA6eDpg+BT/1idtNgdczet/FB
KzB8uC4fpzwljJ8/E212ZM/g51dr9bHcQyzKZHZEhiyAk2KMZd4yY/1vagw5Z8/eYnIdKAJh0lIc
f7/z00nbMKrbDy7JlxG0V9u6/ciy8SjYjyIq8evjFkFCm5fr8RnmOX7EfHf/+b4ny5jo41PEazpX
/neFlrpo4LKfODVPfJgqnHFM5TUxMvfs+F7sfovVeEq+lvY28XZGAWOSpMzWhCkGHPsgj7yzooEF
A70kPOQsBXXKsLXX/WfclcIvkLU5cKGDGkNilILN9maCwPtqUuzi0OdSrPO/y69dIwb4Zlrj2bf/
NcAmKhKgHE4X0WoeGpXNriF3rdu9IgNei/1AlJlnfSs3DELzpL8aQI5qYJiW15BYEnVrcVwdSyLg
djVz6DEp4l7qLRkjYwOP8azpTmrUkDKL0yJ6qE/pjivhxsc5U4ebjBMzluBbA7jgIuQhPronVoia
biikQ7w2SuYDP9ItWc+KDFWsgR0DJZ3lTgDr80UvGvz/4dTigV1u5sWuqhAQbZdP5ZW95KQJQXZb
FAeqEHYH5fEg8TI/PB4Wjjs1PzAMyWOatUbYxWfonSc6VX1n3uKfM65iosZJ65HfLdpJKeecYeDc
EvCL2NFvvVnKUBmqEc3NgoJ9IyRC+2s9tg5G4YHzBH8ihL1eO2MXfUqG9V+ZXj2xNOlKqBd+9DtB
FgjvLItZ2Gw+acgXm/TmUmCk2H8sriU0x3KEVq8FNu9IYFE1XJpYiAtiJCpjPWJm5h3BgyOvvrxr
n6u+oPio2uoN70lMvy62FuKu2yFipWfEzJoibSovcmRfwOc+VZUFxopHsq3rsC/0lb8LI2uEUoDa
OnlyaZBYvF6gRezTUyStbPxtbO7ZeeQl/PM04Bm2Q/2a8YFjezmOLLlCCsR06n+ouWl0V8TP/nXL
T+R8v2Ezp1Y5rYc4nwz2n1LudWHtFvVKNhVrWHETjV/Fx42+x6UCywMbrT7M5tkFgx13uUgOC09W
TRTaUHugr97MuK5KstvmN6lC6NaTd2IZcge2A25f9GeDg+nE+HvGd6m/DtZPlPWnnulCpCym7qcc
5X+MALdFE/48p3jzHUuU5imZ2RR2pckD/yJSH/91oUngNqPy+F/HIW/nfae93sp7GYSGCWRNCGRr
BsKjcuxdaUqbsmMd7y9sUfsznlHYAQCRuCdCAQos0516M/xly3BFZ4+DLdC/tsv3M3Dafwpof0Pw
l3DUMG8DvCzc7Ny4ksVItgdEYZBb4c6oMZB/fGZh/s9QLd+kkVapWrXjOM/4y/hqZTxuD3sfWLcm
T1TgRgDl0rf9I08O1xAVOz7zuje7PthpjGxs+rPox8Yf0nTQiA70aC8ONd1J1tEAH/uqD+eN7kfy
hKWh8UGkFUrLi8lqYnW2aH677fr222394NbSj0FsPMLqCHI31vzZwbapAM7mdxV5HCMGNwn2VseI
amz7dpmmS4tCBlasVXCbsUR+1zxmWt9ZeXku6XFtfJSayncl7QvTcVRbFdxAwDQLCWTXnytRyUWS
x5e5YXrinilVsa+sCZ19OmmfJd0cyp6RvNgJ4TnmteAZ9h1DkZMfm2fmseICH15m1JssNbSP0NMz
tDaZmJPBtQmn/AC5YAgjci+VZGyxigF4hRxBldaOpn2AEJeM50tJJyfSQs40PxzqKR8odytjYb8q
HMecGWAsTA/+k5hiHUrgMxejYudnSXPi9dtrpgg28Xfvs1pi8Bfr9UTpWHBNE0Q9OzMAT3zSvaiX
JdJuFVUA07Aiky6CNZJFTrfaSh/G9sqQslx3J/Z/iKnRISG6wHp3mlnOo1Skk2Y5fcNKvogDSOgs
9hArd8MAkcATrPvp9YaqYonuCj0Wb1jOYaDC9aRG1ohiap86vGv2WgFIzJxZziCIJtX/cn2AUnvZ
WPSVM9j1uokHnXOHBfo28WlHuSo1/0TkSYolf9lRj+O+l8Jk6Zl38V/9PpGNciL8RP3MsGblCeOh
N9wT/BSDpTGfwft/fIJ15jHnZBEILIm2VFpvK/UddJVAJt7te0g5UrDKuzLNybkhXBwKrvwresnp
76cw8ODt1HIpVWSHoZqZc33TX6EraaI4PIIPgSrD4AABhDssZdSAr3jI8jSPP41gUaoevX+QNYZ9
asiIwXhpCHzzHsPDNA120XuMzhm7kJKgMhczuaMHO61rV9MRo0xuAFtNH8bhiTWZRsIJe0huqtCY
CSYWsOXyyx4Jld8sEZ/oUNSHlDa36UWrF2v/+LcN9V8suM4qICHq0/DnyPteh2lO0XVx+3cOseXe
R5P7sJy2YETzdXBv4ORKMCzVNbmv+6urEBBHc/JaR9pnKClFCvBvGj6pHBD1RjNMigGJHCySfDXB
unSMa4WNJH5vJSTr1KqjYHoud41VARCOn//9wOfqFuAtZkwyAMI7+xP5eq018bKT+M3nm3vwIt/1
Op9uEGqdKdBBAardkwOKgn1oNdoHZP/Yo3OFjAQ/YxbsafZRnYQPTKBn0Ffqgwx3j8F+cA00UZgU
Ql7gsBkVlXPsUruidYaFygMaz6PQ1vZ0KKlGUlMH84rLu2yh8Kcb2eIlvg7G1WOK0yfUu77ju/zi
UAseuk9NgaoSYiUPu8VwW+a/E0js+NkO3cyywU5Q8l3CYCSc0BOIYZtpi1WQY25hjw0YmiEjpUMN
G62+ghIlxiYiT+Cbt3qxUgurMpd2NJjcAK8lgtTbMwFfqWFcsYb6WseD/RfO1L4dJVBEV4wyAfQ4
IpIMo+eYJkK1tZxXQebYT0aQh8Qv7mLWnV5b0jlc8PzUUJwRDRIVGfAes+nCU4LSxoOhXAU8Vjel
9FqVOQ4eQeY/WZXvIk8LH63WY8o7D1x9mSxOxpuOvxVnUE3BpdNzrDmfhM3ikY2IUp1cnq2nk386
JDEaq0kxfrH3oESFn1dl92aDsL8XElIG5uN5eNjZcCWKBQTDSAFpLOOFnnYho2+IqWXw8dBjnbGf
qoWLw3MxnotqaCKDLCjqReNbUk5nh6p+DnrU+0aLQhnspwEWqsL5wtgxxNf6tx3zJNbpCKSkeFKu
lAGnXLbZOJg1HEEeVRMZadDXx+GB1OgMEt3JOh7hKYsKC6aOF3c8nXHgctmfjusvfMisgtF0t1mR
dfhvzYy5Sm9ihhG1PpN8iNXWg/ZOyfO8VHa0YgQmPZhViP//NZtW0CYpIu946rVZzSYE+lX/uYxP
0UrJANlfGwFoNJ2Zak8Zz9Vun8TaBV43TsI6p6lJxTifLZVJAsApWlCifAj9eTHOWMFUkiHKZi28
I+ukHLqIrjhMe6tutIHhLJzG/0HkSvxfqedh+e5FFXc1Pg81bKX3wgWsxbwocTjBsNqcNLK1OkUz
KuW8BFiyJrEdTzm5DrKM1hxTWR54rzgWfDR4jZ0vT8Po26BqyUA3IlASB1GHbrKbxoAlopyUJMaX
t4zwuj9Ph0MFHqJaXN4KgwSh6iXXdotLyR5k62PtiTlsiMgu2kdpQh954ZXGXzA5Paj67vFGoRbz
yumORA9Xf1EnHKIjXiQK9yzlsPtB9+Z380r2KMhBAz1I0cRA+ymTbKvugEJP39Uhoqmm+/MP/9eg
OENo6CdVsamNdKdbUsKhjjlhigQ7zg/Wbnx+lwbut2rgukcp2ydbVkczAL5OTr0kZ15jB1mAwe/K
vWuaj5dFsi4V4/9HuUHGFutkNu5orUHn95XRAh+ki63zRF6p1GL58tTb6G9BxZtYzN0fy85UzGay
kGOlQ79Ni82+BR4WGah2R97JzpAmhh8mVKFxeqcYu6sFMhCWLxLPocIHyDrGVimw7oxACBB8B8PD
TXuMJNeiIoUKtJZ0DrCQJtE6B8+NRxgbOY6hNbNsu7FM297DFKASkAfGp3xD9nZgnWZMTi9peRIi
m4dqgzQNmWhfkze3guCvRDia4mCyB34q9wdt/uSCn31qvTofzOIZbbrEs1G6/FfsdMxgp0Gqv88y
OBFmrP3JlBXEoPDfuxwQnb63sAPvY8BoMehHAn+QMPGuK1koWUadeRVvlOhbxgCuy6OGDHJ0WF/K
T5zTQlvGlE0zXeIj7WjmvIx8j1T9x89gJO8xwpw92x4FEsnGVdBacvvAqNen4E6I8/O84kZFA9uu
QI1KszYDWVIwbRKCA/IkkqudHhXswEEM3tSDLMQJH4pFiGnJovcCD/Cnq30eps5Zsek77uWm2E2w
gwLHZR26HIeNa1qYKzccrEoOHxI6BGaenq5v6XIDwmakDZFkg9A6n9N7Wpnf3b8GLpUEnrjG86av
ksSF6xCsxbYzsmjsy+KjWv+hhlORcpzC/3UIdW8fv1Pr7a+GQPl1ia1Yp920wJu9ouMDZ6dt3zhD
GocZfrKURu82qUWzboF3Fj66rdCEwXEgvOkqCdYZRCnVewup/BOJNKu/JrQHuPnaIeXEA+p6zHmn
AmWYe3SiJcg/PKaZTR9x9M6h7fBG+2cMzf1kWg5+k40Rm1vRZcvReDCCbb8QwaX69jXPd8WMJ8Iw
6rHPz51ntQp1yaiNQEZGhWNo00vUamL4rHu1pJIB8F9uJOvRaBRIZOMa5riBUqlN9K1R1qph1iht
OPjfCEm1QW/oBkW1sGIAngv2Z2ZMVpxosPtlgBQSflwIndtLV8WnuZ9cNGq6T8j0bHEaooDWd9lh
fOOGgzHvJsoc50kfLLyMpqauOiEJ63gYO7ZABiS5+xSURcinOiImutnp6r8yEMd9tRw9btZHl6Md
PwwMXuqnhIlLRduVTMJsihpeXEoLDt3mM2i6BMlMi6hXkqWCBx2kTIQ62GHjdof/OY2om7snyIk4
r1ea2VLpr4cOFVADYwUNnAbuGcIhjsje0oU7d/t3CkVy6+0tKUHj8CMb5YIkq4VRx+hSle7IE64w
2yVimGK0GHc0SkLYt714MfMBpt3wSovQwRgZF3DrcrZ1ur7mLhOekr+uWrQmhXBByZGZ4aAFJxva
b7p0xFS5PBy87z1EnQjC97Ctw0l+yCiEK53Ky963Dhmbn8h9snJIiVAEvO4hIEVKu2OUWnGVulM0
akEgRdpgR2K085dn9/88StFk5YQGKCxW8jxEVdjpPpATwUSd2sr3o2OsSDnCoRxZc1GRiYJPX+2h
zQclsuAzYX0jGVbK3hYQwM51tUUBkasmqg9iLNpWhmgPJx/bXczV40ubV3yZQTF6EFs+A5VroiaG
fNfO7WcijEwZlyfY5jH7zk/1qOwL0ajWRMqBINw+00NEEAwE+bHOb5NpBWPiyodTxXR/b0UW9Pgl
AhfrnSlcBoRgU5CZRG8Oj9VhV7nfdrtvLloCFrHG2q143wKe/1Va9wV6XbJUlpPusnueYEJa38ZE
SIfmU0l+rjuD2F8KHzQbeRKKS8lwc1OfV/OJVV2C+SlsXPIsUQuXSb3xyPiNNAhkQXjbGDXQ+SGU
yeo1J5HaIT9x7vmApY5n1jXdue77rmflLDLQ9Q5khUE7KwU9Kzcj/cnXTaQR7cCsHefhPqzgvkeO
KsrhFa8wYdv5D0Anym9iEYChtyl7g6h8dy12aFJb6nvIB7+yjmEKd2SaFcQV8PpUY+6Zj34HUUES
UY+0hDpFe3EgC5/15cBS3VC7c0mByo/YVzFAmr7sZGpK8xdIfzTGDR8fbIGefQlXoOHicjiBtzk8
LEoLPTpNfF3A05Swx9Y3Tr3jfxAJFDdHUR4aOtRzgW7Qe7ch/ouaq/vs9rEOy17a0qHdCu7MF8Bm
xofZ1MkE2w0L31fubClmlhhrh8SkD1lGl1qpCQmvBOYHMXdVXXJ/cuk2DbwA2GNeUHbTcKl9Ps1d
tN/eDg/rDa6UNlY44JwkG7WzWM6Yr9YVda27m5iDKDLJaoFOq+/WTy8csf4EyCHqJIW+eN3re+vU
kKUxfU2E8ZdZpM3ytBUgVLK1Im43tXS4NKsNO/wxcFfGP6LM4R8TGhz4B66BpIqAA5hosoiRnEgL
OVp6hUattOG+rGP/TSsWNk8mh7nom+1F+Bpkb3mEi75EPcgaJ4IfN1r+Iw8brCdUKbNrgn1R38K6
PAlwD7BUqObdu0KowB/SYnaReIu38+UVWVIrtPH/pL2x/ECrJlAlT624To4dcDK/d8LXW3JtoJ+j
lM71bu72S7s4XQH0u0VBoaTNYs+wbi7FtoYf9oGiLyVlIUZ0oB3NS3gpJoiEKkgb0RHZQiAaUI4+
ZZHkyj+9miJiLiKwYmWbsGN+a1/bnVjykc1pVmJG50QcVhnraDt5Lf6+5vs2KeQzKEHF3+jh+27v
pu3x2NMZj1OMWvNPJ3WEM/m19MgCn941mjpdX0iRLdt4xd8++36vTgdWCwtkJOCldqj7QhYJ9S2m
aXlPogE8R6DKLj3PFHA6xR55Z4xWjPIgUzv6ky9wiRCl+V7r52pdoRL7h/WpQ1cJCuJwHpO3LsSN
P6EaAuo8R9B/8hV3/bqxkmHsWN849qNZUGnn3Xpb6uDo0jPHiep3Vcz19h3p8Bd5rpNsj59toiSe
IFIawj2gWoQAKqWRZEO7nyN9N2y35zgwNPlk8YsN9sg9mD9BAJlEnWnpsPM4BdCbo0rwuEUhLpCE
K2VCudmdlLmVdw7cEXjGlTWUeEEjQT8wZYGhnCdITZnKmlfQkUFK4if73v3Mw5WgPP1cGw+cZTF/
ZqvesaCZK3q77g7NLnAuDeWDweeeEpZlXnuHh13a7hi3MJLyvEGppdj7LBJqTTiGT+NhxNQvaVif
RwdHTJVAMV6MsgqaEh2YBKAwaJMzwaeazSlYD3CeNc5Cff8CFGdnyRGRsGRS+rlvuoFGZRNOeWCX
LdqZNbeo83+mXdJvOLJxDbIew7XDgKgO1NdHqhVUjcdSilvZD49FDdc/ApOOWmLklwaEO4IgX+Xj
qO3Ukj+hc808jZ0hd4Z7+DUD6sAGCC5cGKhDJThtpRrFYAfwyXHhjC4rp+hyRW2tuXF6pX0N1oWQ
TWbD10sPhYq9UCZLc9+aecWAQBq56nc5SA9tz0N9LR4kLN+O34cz9B6ebiupdy1O1ivzhOXd0mQ/
xLezgf0vMclGYUJCa7E8HvrOYCrrP7HuZs2MHSet7WbqOsuJ1d0unQ9MvR/ZFI1NI6d4UxGSRdgM
/Jo+hkAVNIEPVUwl9irssJvdXDiA4vC79uHnlxktGjkXBQONynI/ETT3dCMgdBfXG08L3E2nTtrC
bJku5pYnC8e17qZMD4SChRtk0WSMDhJeckGYvalFIQyTc9/SuKvADJ9p0h0y1M8EIzhQ1xJdiyYz
Qi12o19SFVN7NlB7RsLL9mpPhO8qZKIHfNVKAh3XKJNvZXM6RWg5cprZgbvWvVDHZtcRPCf1VNjW
redeN6AEmM6GCXm+RAi6UGOix79kIPHResxiMF4PnXe0gwuxgHZaujCQsInOHkwZNOR6SwTiZ0FS
MTDGsoy8k4ZB1cikqFWtbbTPBmIXy4B85unt8b1gNVniB5C0EsIg9/avGl5jJQfaiIJZAtz+2iWE
Vzjw8Gg9udN7N+CB5YXtaq6KeCwx8LPJr91j8+zquSJBg9HJIhBrgssVhg2P6uKbyuvPYPwR6Hfn
i8E+RysJ8bVpJqybL8bfhN4SvGBwvjqJRYoZVpUouVv6HedS/dNSu4qM8nV8pxRU4E48AaOgRTvZ
us6sRoMMcpxIDxkdfx2+UUOkMu/afUrcHyHxPinQx7gKx4n9x7ds+i9Q3t0NDQqgo+a+eB04RsPw
nfZWZdcwfPUX01Y1wdppFiZPRECSsfeoeG3N7nmFjcnOjZFILD9VJOrek/g18qCVsh2vxFoWXZWr
yRyYN1SD5BcDqvx7gjOJl7TEerfA/HwwKapGiQ4R3prX0xELMEyEFYVeW/fZJqbqB65b2jhLhJo7
NsLnftswZyvhKJcRaO8iNoJLX8HdJqxLu4owHT0EBvtlZjV61/T/chhYIqisj0BK5vqe4rySzCDG
+Za2pKZaCAkhZyoAhnDt6gKGAWxnTse+R+H099CNq7sUUQeyuu2F6VVD9CKQW1EDqR2UI2Yy6HTI
52uhaO07IuCFAEzg+Vw8fHynEPgu0yRft6BWmh8WfXVG0LkfViUekz61KgJrRdXF1EHShCiPoibm
NsKeO/0hGY5iBODmv9Lr3AtrL2F4wLBKFxkHTuR1B7qcKnJDI1l+22hDXzniT9XT0iUsBNOtxx1Z
APrInPloH161Pu9hKHXbKL7V0Hh3XAEurc/Vpahm/K8wiylUfsNjhnKE1jeg0w+FjbjONi1XkF9o
dYxgkUAarQDRG96e3pDbjQuFF3YzrLi0DCKo1idMATed+OGa9+zjQAsMKYAaLmx6e9/gKgIABRvG
Vp3MMOEY6rueozZSi4ZSTopFNs13yt3uMDHk9Kxn/5dvXojjX0bipvMZkMAd3LzmIeUupjdNPi/6
Hb+a9ARzxE6G+dhdlp7QOSjv9LzZUE5uOvYOvg4vAKGQ5GZOF8PguIsKQYKXTX6h9k5inRtN5azS
v/MItk+7M3jbig8A3SwC1dzjKdbv8UYtBqJFA7+6x7AZzagSfBb0mW+n+YDZMdd243Zd5gu9e6xT
zbmsGu2cL9M6Wqp5YBvDMNQTkigHfqBvzpjXFnOCISSbstxdaKVQW+8nOn2pXM1AA8dbMsDn3I+/
3YA+XQ6akQ86huHvXGBPe76/U03o8+4OMY1zbpzQme/d+PfJd6xED7In7mw3NpoNFrv8b/gnJ2qk
+Hw3/snw+Wn3y9SplfHvpUSyUMgyT7rFsv5xVTRVIp+hrmid3JooKzxw6SoNU86s4VPUhLDXmMve
eA7Dh3llhJTjFFgKUE96GP1ctHylw7R5S4hBqZ/Pq9VnjAbTI4jxVFvEKIgjcrm1Sur57IHQpX3s
FS3fyLqIZEz0mMvuARRVhOT//Uw/pTBlkfVvLTdky9NypbPIIAxiwNfjUmYc3BRs1gWEjdTuPKLC
nMqWLTdiHam+E6K/UBu/+hyNqG4zvo79FB+B6ynO1Y8gZVoZImcvweWlzeuusZzlxwB2Ra9MoODi
UZjOFyHzOZyiP479o/5VqY1+mgQTe/qajW7FRtL4irzx1eXbheyu6VZvFFm1soiHlQZGTv1raVrn
rlgF0bUgPV0Lr4h6udrjCJ3eAx+8/PzzTLIrNV9E8/d3UeFuM5j+I+IResDNlHx1jDGH3nTSQPSX
xl39CilH77w6xoBTncwenHBHGbE2QMbIIOwCcqK9FJ6b/DZf+OSTQI7axcoAj1SdMkh5x6RLGpzg
nndKz64Gt9yxvGkKuQwl89KmFo/RIuBC/vlRcNzQsgeCB7MsIGIMsYXk55O0hVhgJn2heOZjPgzE
ZsjjB8/v7wzKTf+8Evni8FoRxTk+anpN7iRhhQdpcver/VLNtOcbpSMZr8UmvE2+0E6bB89gPnaf
/V1OiDup2WHPTHZOZ+ww2Ztt/CetGhR8zNiRiy8b7Aq4VxUTV++d59p95Z5in0WMeqGCz33VoXbd
wag4qCVORuLhsV13KMBKELRqaozEUAAJwEd5ljxdPA7OGYkS19Ci4K3/6fXHKwXA3Bd9IbyubsXH
JXuGnHVldKTWqDJynAV93fvuc/erK22uacktL1ZrMR1rYcggEyacpdLdLS1cejCKGOhdTz92SdcC
RFhFV3bMzbsOa3hdszJdEnP5Pm7/C/m5AGX9iWQyF1DpCBGTGViZofNnsUBroJQNwXl/OPk051iK
hzbZuVL+1uFVmEZ91yzfSMSPaPeLoGpRNreZcrlLWfrECARy/FnTwrqtd7VJmWsXs4tf0j91T+rg
AnDDFz+C7mk8IBgfR+iNxTEc1hR76yWxbOwjI553kep+I4JM43jnyJspWXo3RAENTia7n86ZNB/G
wv8zx/ErD32/QAbAyydLCxgkCnlIVK3hvKofojbMhDl05LnQl5PbpusPuCgkIlItnCGVRQkULRLf
AiDRPcYbkHHAWEP2z9t7sLR2Ni25Jivu+0cLJ2BTqIq51gOzP+XI9tIiTvkI0WfBWTwH3pUmU2+3
4xRcgErWpZJtyHmgJ5hOPu8V2YdrxCvLd8s1N1h1zmElnJXT4poixu3Ir3X7o5f0ADBIdc2mhaWA
tFYMJoTQUbZr8pBGF1dJj37JtrzFJM3SBoKQCrarfuni7Xykdu7e7EQavBDEnX3d+4OO5nErXpff
A7aFopbnB3X5Krs1aHckMzpELy62Aks9afY690ahduXNWdeGxu/BGOZSvQ3QdL2mKQXFAWag0kHC
nFZL2XIeFQxqmI8rMcAzMrcBr+4iJxLYkS65QJjOeAW9L4c6vBbKTnDAiWw8h+p1niLI7zbOpgcz
8MIecIbaD+emq+YxTfSnX8s7325AdPk27LBlStkAEgKnpfTcKEZfa3Bn/Didwae1OfhuKr+9nGrH
+WO76cm5uaCO8U8D6pz3UErryeKOsrLT46rlRdsgvrWVEw8iGTsoJiyLQRLnjpV9pIyktz50CPPm
ecBrlrU8znA+dnD6dXyCXAGQhugADTejy/tMJcxm+Gv8qRBPclhLMexOFGOUwds1PXJXBzoZeqWl
GX+ZR3aNEriAy98iAaKGUqoFpBZp77a+4ZisF3n/DSpRsKIYpHY+QT9mEMo2o+ipMMYOa5TM8Wql
5Z5OGZR66Xyp1j/Soq99eMy3oPPBeHcKad2o0AHIotNxpmpuwgcdNJY3yIzegi6EgqQhOc9+cNPB
pwjwIqZRRHpRwnBAFRs70M0fUCA3UnLFF44V3XU4FvcCE/FgkodAP5hOrE1OTGNxHHdpO4czc10G
9P/MweHhnvIbGYLZEQ9NZCDkEEEQYOAb87kf6mhl+Wccskvwp/PIp9thO700U5HVRg5UVpRwJ1P1
/rLiC4hyTZ6PkzLnlOkSd/x+3a0yZsBfKyukt7OGFVZyXDZ0JOoq2qEDeqfbou2SslCm2hCqyWCt
p5itwlsixPIq33mOqg5wwb63NWwN9zpeqmWKF/gBeRi347WuBRNPC/stqtX2SVAmfRa9O1Ju2f5e
XfbGno1SMoGSuQGm6gz0Jfuvoyd+kdoCpd9SL0mlhAlbelyGNimXTy9Ilvc5mxMhJHMII/AvDWwi
UsLeC3fkM4G6Lmg550psnLsQxFBKbF5CYKzUGURLcrm5CPF7RdGHm55gCmb8bk4f98uLLlFjrySX
fZxlFHuB4leRPP3y12FeVKjlzk+yFz9KMUZVNQOs0ASF1El2wFQnPizkpoIgisIkvUm8TgBgpf0I
dN1iaOgYt9pS+PawYdR45M8vR4oAM40L0vGhXN7MoCUID5x6lXLmbXe13U8UjaW5ZCfxxSxSNIIW
5YkUKC6Vfju/7QhEkvaC2Svb3WGxF/8YCiCz0hoIMoLEEFqnod+KXl1dVitvYpimhsFrj8XYlOEm
zV5kEzAjfxqMawjsE0TnzDIeBdbxYhiJ3exLex4EuOVKmFRBA1jaZUHPC502oW6YZCPppchs6Iss
+xGsV1drfzlv+1VIY7dJq/NyUJZgKR3Mp7Ba0JcmqozfSdiYFQhY51ICa9mNzQ6EsLmkrPB9/cgk
4VbRyEllOQepEl+M9Z3HtA4HfOL8DRFljMv0EEILyTiOQu2bH9AQZOB6lRHuL9AtpC0Nz0pb9qZ9
fF8+A668XVozpNNiQvjH71M7b8bDQDgtRtZ79ucgu6tf4Qc/dbtzcnZdBX55BeV9qPxTn7kxhwht
SaWWGhr5Nwajoy++hvjsowl21cC5hTPeo8QWA8r76iFmmoYhe/eYXRaQGFnUy8I39I9lQhLHlfNk
ed1MRheVvbPPa2gj8enyl7FWN1iQaxyJK1WpBuU8LRBrG98dn555+GcN7rdjFBMGg2Bk9gTlEL/r
mgVRKUp9DG0+XYM7x3KsIDc1zydelHRBcSdx63mEutPep/ObnJ9wzk5g5rSaq5cYHod/rS9q8/0o
j1JkDoIG6HeakI370ce/I8Ps+/K6BSgENEj4jtjUR0EGrPXWXUyZDYcTUwNUQ6wimUbsgBpxDVfK
6hoMj/HTyrCYCDvis2S/sULp09rVbCrgfEfAN9XrsI8yQRo3guMphsgPZxoRCKUFyFbaYMCAp45z
LdUH1ymRA54iRvC7kFGJ2zg1DH1Xh8DJX99xBZ8l2u4XWl5GOXhNLCbM89ncMvi32J5PBFpkP11g
ywwbP6dKOeLRouKk0ZYfd6m3/cirWY1LzlQ1SGpZJ6UUdNXQrdPTKsiC5z3JgTAxzOSM33IMS0aI
hjU3dghLkxEbAacGVAIt2xrooL1mdUw/Lx72ovWt7BOy4bauZP5/Sr2EAAQvEnbuCE3qilJxqrl7
/ZBEyRgIRFYJquThBpb/5qp2AMcjsxWKXJyT2cjI13mfW98ksd2vhjxBLRLuKy0bQEg61gCPTBnC
rfii991NuRyKl5ju72QC6ZoHrwsqip+RfbCfGJFofKuBq6JrixOJA45qwfaRxjN4MJGcksSCAXAb
5mhd/3anmfrgMczavBYH0a+pUDAp5bB6L6mYwRWLx0fFgRANdy9Fe5kTJ1H9PLvk2hu5OWcQ6/KC
cDQkwPtlAwBUnyOcKFAbuXSoc/pqExeCsL3PNse0SOMoy0+BjCkuVR/C6q3+fk47gbnA+jkFN5Oj
RN/EXM/5bTSyyjIvz4MTpCTte0CN8NICLiRiYPVYcuI6IJ2Ow9zhJ/vFgblbRLyu+spdvwxBuX9I
qlqXPYZI87Or7V7xYgEEwP15pRfg4ORVv91uLCbIhd2oBBAp1SyhhNsRk2877ZgN9h5IRaQfgUll
0zcIhuU5DbU03KId7Tv5V5T9+cIWmserZ9xdL3ixa4Kd/aiIhNqO45qryntKP/3d9ze8BkZ+EkIH
0zvB6Hp0o0/Y7cFL1y8YApnR5Tm/lIpgKIUaKLSg2gNEpP9lIAXWTOx5Sqe5KIbmDuLpV8QMb00L
YguAh2eI9exZDa7NmskZsBSJu7/iocveLvWFN97Ex7+DgVZM/5BKaFJbJ8OckR7gaOqMVvVSDOLu
1sN/o2F+qyEE+pVHNsb6NbvyThW6XvIj9Vv8QE9FChfVyWBR3PovzD4NNekaBlSG8ZRFiQVu4OA4
Y/ps49gmPgDqUgftNqb5xdBbN51VZMl+FNYpwzNRGrzjr58TyFbUXrynvBczm0WCbuIMz6RqxJ+t
5C3dEk2ssoM6h2B3AFNZyg3IyQyDCTworPtCdvKPrpnUaM8+V/QAPIhvFuuL2uHlREJDFnxPo6bL
NIQZLxP7rl9Tl9MmpFTfVwfEgCiALx+akvP9GpisY+g9JhCdnEEVopMMS7W55J/+leWLbvqaPdmE
uemaL6wwgQz8PFefsTQ2bAwFZyGW5Nc5FsUTT4PONgqnxdnTqQOPfIEKjAaBLzfqzkwwvtUco/QN
n9o6Pm0L4Oh/RyDxzBjIarSkhM3OdBdNZQ9gKoHplcEBqt6R1TKjBowQaPXNrW54YANm7QIuanlP
scMHfHVAaRBMR5Z9aKBizJuI/DlnfJETVtqpkfnI/nq6FNLugpGym0CAksehK1tsvpVoyXvI+TjB
aJFZm7dbg51ElQdX17BKPugOXgcEHAEg+xbrbHTF91FPb7Tris+YLSceoHCLfKOQ1/Sotirc49SS
uPvcGRMJlI+/+406vvwYZMGz3KNRKuVqv0hyzZ3ybyIcjeijSa91AqzwmL6wcAqKWjD6yKboEdDW
5E1CIFZO8MP62l8FdG/QHwi0REyl+WRLZt2AQjNWrHvWkjqmkOkoCKizoSPWMo/FH1dPMNxmbt3N
9vCa1bESrRIh7WWR21mpip5ovzdomozgvwN2B8J3phZhUQhAz4dHmDyzcbIoE5EgZYixmH7PYwLk
Il3LGT69zXDXw9vI7L+lekcC6/uFSyUqhi/eRyuERwFrVqgpH0N0WDC+jhx/+akTWoIStYYP34+Z
mCnQXsAJuK5Pc0cqoEayNE7yY6o85GqxcakBGJ6sMf/1tYQNymZ1V+sqPV04KwvBRu4GHpAF2soB
oLK2WVrWlwBnEnZ12Nhqis2PjIWy+AQlEPAX8EhqLSJdg+afNp2LNzL/kZO57GSG+nRNYEcgJrvh
ir38wCr6MFl7HclVriIwBN8w1VI7BCKWJIciIsxilt0AulmiPl9K9oC9mW7Mghm6e/DDIvOVgV+b
wC2Z4bP3o7YAaf5dOVLdmdWOdYDh3wcTOtCYqHNde1WFV1qjS+H8/YlF+Kwp5P/CwfcIVy9tR1ty
j64L6Wk7AC1bL8GUT36k2Iv/BlzVivlVbgIbtpC0isx+rfJjvcCX1jTvw63aVAMTFIwRJiDanEUK
wlUsly7z1fgc/JgFHDOLiqSZWbPF4OrdE7gOYS71JSFLN2/2u8k55nN/UVelFl+gOhQ7YmlZixyR
F2VnsB9C9zjMEg5MmhbmDtN+LQi248VOxM9UchRgtkIdFW0RqHDPRixSY6P8YW7vQJkdpftf8MU3
Ymd2p8qvNSO2IklepfIjHXU5B43jPVWWnpflTYtE9pYLYwCrjLR7sjfk+O8vGVKHpi3DVSET2o2B
7mJt9asXfYX84u9dMVJ/yMblPQdVzKZ+kowhlp0JymDWkAtI80TTvrNGYfdZgcdyMpnAgUUKyRc5
beqS2sU6L7Ke6ccPe2ONK9+2GH8Tr/n7VXV5yR/pwP9nAkyfM3LylKkfDuXaqONaIUzY28028zpU
NdnGRXCRGM7E1yfqlxV1phgdGvpMy9G49VOCESPF5pGvUbIPVGm1dE5PUu7fVPXVUJqQwBCPunCZ
EbVeld+BOQq8UupXrYwAC24qZX1/WOCaFQDocCHp2G0BBfdt1xEplc6X50OvCrKQsPG6hUi2rl/u
ejkwnizEKzvJawS3HpWLgroDDe1M3aIf6yr7ix6Yk2YGKkG0AIMLozfMr1FK+xYlHhdw/WUoDooo
nPlSXiyHt6DENRMCJUP1BwM5Ri1mKd4TFzCOmECdEAK9IiaV7ZzanYGPsIYjUAzhfp3oCrFwsyG+
IPT00XwQWjj7feQwAg7utjizf7BCL6UN1TA3DcGWn8e2UEw49JF8wvDj4sTTIPXayXvsapbd/axm
iHyPg9DISYXBfTLsy5BQQ2lNb41pXrqOAhNkJrGe00t3Zyfiu4amjJMLukyJV06oDZxcLwxQy7UE
6pqwRc8L/zJ6Q/WSRudkybeTCcpDweDQY74C8TFnKacWDWuouEraA5U8VuCpx6nsVqNOmiK4JEHo
yytJarpmf+oDwsS2zSgs8+TVTcHtZ/CuD26P0Cv9O8o99C2+PHuKNfmcO54Ws0L6WZMcDbRwsnuG
p9q/IS+8C4XwzD+W508N9AZl1skAd63ClXEWL1oRLT5UDh3RFpkJZOF8cwWN3YO35gdgXQ+N03Kg
OlFh16YHUENOLy24ytOEJmGlErrCt6GVS3ppUlMjRiEST6/PN7bg146O94U8unX3xl3opZ84n4l8
f0eMjuRx96sGE45ZdnTxPWQ01cjBkl8Crz1ZCxy63HIlYxpbE49OHHvwDf3HMFVXLnND2Gyv2VWX
t79kQkSBhXaoggZZ7X5x7i+A+xcbUCDk0i6N7YFU3F8Me5RNf+HMlxjbWITFHQA8MAL76189OGHr
6B23j5qGhHxrtAcqhLIbZDr2FE0ITE1JKhH9t0X4Tx27IARiXOUCPqncuSwCRQP//DXrgLLk9sVk
u4nxsTAgE0tAC+ua6o5+K7DgF+oWyMBdkW3w9Zba5N+I5zA4IGxkw1gSktkTi1H1TyBM9JzfGmNY
+pYEe0D/HvrHkm6J5HgAji0XjS1WZL7K0QNcNA5aL2uMkTvYMG9U3n3W43X1qrjsQfoiQ8wWv+Ri
bQoIxe2FyW0WqXT71wXUwe9JNYFFnhEq81pj22KLI6JnresnpDfYn6ATESgj6NVnDnUXy7SWyZ0G
AebonY3Q/cQTWrl11iZ1KC9bpyTRkrD6KzgewJ2XFHGxEhu7URvM+UWLCXp9+jVGMQClCMNf/0y2
2bd9gonlhT58z4SMFnE0+k4QdPXfVM5lCe8+03P2c80QlodwSegYiZpBZrqrGNeSaILLpUTHnxtF
jODP5W4XCFWpbB9HbsCheOd0u7YXkgxk8gPSokG3xN42rEBtPmRv6L3vsnv2ZsWvQHceGORRWvdM
sh4HTQ9NwQjsmPxHq06ISVGbZtPPJ6VSv6yo3Yylb5bVql4TAESuZ2pdrAwICWsT9gfUPScfRffI
2l3J+62R0FIRBVNZJM8rZKiDIgpjKcTOFf/XXn+UVWkd7f77mZGENl/dh+LhgWXOsnp4TsSkdWEf
BeW2wparD241mP2AWBkCL8/zdQgyJQA9gCT5yb0DamHqfzRgN2rJwSQHym92wmiGDjiHCkbiI+lZ
UGrE3jGzbC3CunJ4fKuCp9enFGJjAEBUOYY8PVJ5deAyAOAzXlIGIDixQXwYoVrla8Dv+NE+ix6j
u2XZ8Ok6+RIkdCp/qFpa/74GVDdJv1In/+nLg8uKKFUgblHaZ9laP/pX1PA4vAj9o3XVUw4qjnlU
ftYzJGCUMhj+Bwt8opHlo3F6MCarCAV+KYrjQS6N2iD6RWHbwyFpWR8FUKvQFj0QZW0SZAIuDrCM
VF6mdhnoOG8J5sx2TGMbjdY0X14DYi7VcL7Lp6qzrsE6MtjbyOmCwfFrYMY+8JFuTt7y0iVj6RIq
4Q8T6Ye6BsJa4kPBCw7ZqB7v6rM5mRdgvVGBL04jbUd8QeVdfKBSPN7/wNr0o/gVSFFdRvhBEJSZ
fQPrbmmRI39pRdowugxa9JlYL70mBnICLYqoaIwTiTfBLmpQEpABQCR/WZm9z1F0PsTUmW+7+tBQ
BswbudwbkRgB5fnF7MlSs9lA3d4YIM5sqcq3/Z06Fa56xyWvgjkYq8wWhVzPdwX0vgTibHOZWF9E
ReeeFqvHZiU6qjNSMIF/AEfq6Lmvw2p6O+Mk79pkwyE5Mf5DVXj7mhdH1gEJfRV7kIpelCW4ym63
UiRowkpyF/zYONuYJt5xrlcTj21M2DGG9mWgciJLmdTb2wOrtub3xA1qeqnjHYgCOCI1JmGayiU3
J5TnH5LDUYwYkJduedGWpSVxpA1Xv3r4q1czveHcePTu5FYdtyuSwunTy39w/tsjs8HzhHYBY3S0
7J4B2JHK3d4Sc5FIFMxsPkGXSbKh8rGzC4M0odGrg+1XWB5+W+7PsYfjtu9MpJX4l19btAb5sLsp
+7jwRsQu1S26DqsgV7M6CXFlWQ/6gFROgh+7NycHU8pzFN7FnwySg2Asz6qLINSuy+AWshE9JqMp
sIlX7Zbu5KWJDvUwtAffvslJmjN/PuNFZ4bSiJ6UP4PtSXOlPq5/Rf2Yk5YoRXrScdtWE6iHcDQs
ZUNkAxHrE53YOnxVwS1MoVJXr/YLmLg3yx2zJemQtyMEGf3ZHAQTwBGA6avReSq2ul1simguqcvQ
tKvQtEFZ7SQ3aP89eb6lL9PS9lGjWL0hqusjBd/NI5WbvTNGb6qy+42dyUlr+82RNaf1zyx5kY4T
5JY9M3kGWfz9sigOviuY8RTbQu8KwqeUGnYsGjA8brFVm50p+VtZQ24XDXAmY22b1mE4WXIXwgwe
6i45izRJ5cDlX8zCGzN8nEAZi+9mbFwpSM8VycPlbLBF41euHK3XA5dX5RBGar63+8gURvi9sYn7
CVB3EfGAYtw93R8rCgq1LH7avlea+cjWXl6d0s4jNmts9p0vAjftyJc7qMdSkZ7aE/0Ndgx/lg54
hgZMnwDiirUMQttxGRT4TkwM8U/kXo9m1ew2BvCEqoMn9F8Y6zkijC5AH5Ee/EBgPgGDxcB/PXJO
WyGy30NvEhREvfCI/cMdMucV456X02HxueituuD77uQkhWwepor5sd8K7PpzHUu5Op19RTv7yBpB
l80PIpyXekVLCyTsOcl7oltr6+MUJsf0UuNJexEiXLrr0jflm6VRgsEYTLREdI/1c6cXEYHXghcB
ECNPzLcUkZQvTxR6M1Y52Vz76SqByGEFy9L55DW8axofJBEEVTUrfWK+khs3vQblufXkClDL66CZ
u1wk1D35hPOP3nYWYsz91ALeQb5CKHo+ffESDtHQ7zl+YSB/25sR8DvgJ/S2WhfL5UQ18CXV/WEO
KAWh+sMk26bAbE0KgUuGFBdHGt93wA2ufNbU9YpxLyGKQz95enQQklPM/5Mte5cwXoUiCgoghw+R
CU7OBlevL59VW7Dcdb5+JlHC8EBOb/zFG/2zfAWFKgbI5F+H7OaogYVZD1FKqYhEK2T30B3KkNOJ
W9z57woPTOD1sZepzOJow3qI2tqjKaWWaERKq9OO9dOQXIswaLy4HyZE/hJ/hYW8iCGBcEB+2K4J
dohNA7xRFWXDT9bi7WqZt+6M42yNA9csZYMkjsi6rqiIARU/tmvhiEHMbz7rAeHUBS6PJuFDyKpU
p8sCzkbPVd/9a4nr4kbcN4h8pePfKAledFkWKlyC/d9Osr2kb+7KauZ3cA+eslRa2ckXVWOIUqT1
kjt0XS4p2RSum9ttM7jZTeUWyGlwNzvdwi2u5WP1I2ys3XFWCM9NNTy2o5hVcidLvgUgA/gQpG6h
XlWuVJGjGJA//hq5hU3PTBS+pC1ez7FZKn//nDrn1Vw+cEyTbyqP1IYVr8Yv6rqqebt2GkZsSdA4
/QcpDC5ic+pF1EY9uhxRWJTU7A3pXBJq5qbH+0Js1opLWN//b8y3k5Zdw8ihHB3kNLKp2JL+aYGs
A8+Bs9aoX5Sov6RUEGyUdtSFzoAbjSCK01FnVvobAyTXNoNjcuVEvJhG4udsttHsNbOb5Did4Ng3
N+NdXpib7GNIoIbWFt+lpjvraH6GWMZlHSdXnIXtb7OuyB2qP9tDb/S1UaT3+zA5bBZ6gnZqCAlF
6hlLDsqYfD3j1YCUFAhAbph4htG7meWVoSw5Ioq7ufF/I5Psq5a5jBGhJ1FXenJ8KY2qgPF7xzw+
38d6Rgxu/TeyzZTdSKPrIePRUY6DGqTKr/NVhGwLf2cCeWZZhOXtg692zJbvQ7PeZ/FpzruHRPTs
0gThPUuidSGDYbIs2l88n8w13d3D7ms+iF8PBTnv6rWIkrO3SZyyL4eTwOQzKVMKcP8Afdmu0qN1
9FFe4vII9JJst1aJBovdI4LbMoNG0FqaTykyMGA80V1YIEv4DjdRDGhWJIi/aXFDZYc5fp2UL/TG
BnDrwFYZpQDmunFsMSKNcpzhCM9ll2t1Ej2/WNQebJXiYgZKOlBkO5ucR4iybWERRTt9L6wPBX4F
ttPigaMaJuKWSduqt6wSLmdJ7uZ40Ra3HDEuqvUcWLk4SinQMg6J0I63x0Kw8w7U7+uq21qSJp5P
OMA2Epnz056fv8vlPinHSHJIORZY77mUzACbB5oFZ+6ffE5v1E5DDXZN+51LZn4fm3DnnJkqCI6Q
7aXkTkTUzHXvX1wbYD+TzZZtNDSatE3hD8FJ3XOLLxmB2srcH3vuRPsRVJyiqbsE2H7oYCvpiKOy
acpNukiVIqmWs6FTK0F8FveEXBBkQxym4xWt0qjGpdrnaNuDeVkFAfw9vuhLT7NZALjDN1mlIa0F
bPIExnWBa9+yqU3gWVgKcFWBqA3jVMAvUESLe9H4B/TyahY9hhXgi0RzEwCTuDaQ/ymNvRs9X2sL
JyMlDTgaPBhyzFkGcFMJEU0K3tHzbNlaXUNULS2Y3hMvCH8AQXM8acV4AqBut76X+wgbaTtmmcJd
Rxa7j85PqlflWCzbkMR/1OltOFme21p/syFvQdhs2mGJc7CI/++QonFOa9WGxaU6H20vIVLq6fGp
SipkBWYfqtgHyKzqS6eUFvVkCa8I0Sz8NOR06ULC8taKZMCfsiFXf879lxL1uF9431tE0ddUMLMF
gXF8RtH9HmdZFNlFAN3gxhxeBzfPDfaVpHaQcSx4G25bRygjSihvumv0ePBdo4fGxLDs5boTUTGK
NeG+sEKPkQubXUhwkEZyRz/UOL3CBgtodX0MhoMyk9vPS28ZUz6519h2nbw4KTC9xxN4CQO1nfvX
ti1M/m+Pft9qVCFrbvnenVF5iqnsusl0WRy5D6vAMdfLdJhJ3bWUFQMQSCMsJ9O8LgZQZ1cDIssX
T/Aw3Mt63VWwuleKhdwzsfr5HA4PDCeH8M8JrES2ZdlL3pkgAQgpBN15U0applLPkiuVgSYZJxwG
sd3PX3siVGjRu+tDpIt4T9Bn0ToUBhIHh8BIuiRmL8JmQ5v+mWTlec+oRSvDwtl9+af5P3JFcDFD
PmkWIf1z/dY/ZN72KzYsRrdTB/igRwQzsdI+uoA/o0eMm95KsAoGNadSPC8SXbhHk2tA7HWaTTYB
kg8RW+fqasRITyQEyhea2PUDn3lwLfrbWqr/KY7HffCiq+yXgLiHM4K61X/22Q2gKPDDjrKTTa6N
+MVa6PxADgnBwKRzxxbrWxk8WgOQCOe1YaIxLV3BgxKfIOCWtK0Jj8qYnZsA37Xs2MI0MgokIabW
qQfmQb6MX6O5W6hyH/Qz08qWP/hplQfAOJmjyAw+LCzQRtGsrqVx4dl1EZXdcTrrJDQIuBRdZLPy
QNVWcJuqWLInSH/DpciHQWqWKSXSQ2k3BbyeMCq4/QYBpdDLoSnP+bFlHIgA0TSOcsKruh4Nm/Aw
OX7FgOxFg6s98fnSWXkGreCj59sVbuD/92O84PIUJlUoohF1iN1MZxwkzIeIkp/23f4FGietqZCB
A/2xbLiSbICoQfwCC778U1J4ETfexigBPLkNI3+LqNyZSOoJoRUjDGyvGuEx5oUCVKfhBxIIpZC6
suw6p4G6jEfa/som8ekSXt6VZ5aCjpiPTPyr6BqK7CqjzG2brbo0dQbjr9WmuG2I9PghpNYeE10I
CnjwRV2gIfiaOonqhui3JjPInnz4HCE4KoKXVTTsidJZgyfzYgQy0Ktxk3W3frStU45MHXhzpJom
1mDx2w3zOQ29IOBZ17k8J5nk57SZRBoZDLpRo1RHIqYUGOrP6/KmdleogEDe84qm9rWnhsSimG3o
T2ILTs15B8TWMIEKzFd8B7cRE//8cSMaKTNva2hCGoz7k47NPMsgEGB4tmjXaUihW/fkVITdkA9q
Ng8Jy8lHzg26IgE8EU89r+RV7/a+vqzIW9y00kwWML94/U7L80j0ikLdbsBVU0ol9RTdmnFcOONk
3K1lq58OoJlgC3B1fU/2uAK2+BxZ/vWn8txXRTHpQKWDkbzG58aS7rh2FxqGwFrvahkWKu8fL1IG
Qce8K/Gamyth+0ABgeCpchhkuRpEyP4lFl00SAGgspg47q04gygk8TGNkrkOE76ZtKvwzdJLmREa
E5iXteNVuVXcVQpzce0EOseCxYwVcwQsmP434ttuNUYK62JYICZGaml4IcUjYEYT6CkZ3KvgbAN1
MFz8sA74XhC7iIEvrrBxMy6uSFWj1OaiWwDDOroyfopSZS3K1SnZPvnbpz3YVHvNRH+Jnzp5gQfM
bGEIon5aEgxDyTUpoGbr7Awc2YS/ercucy9zS0L9cwe48GiPmdxBaOkvrHvkveGIBuhQhgPNz6aZ
WMBPr3KnQlLvDCloAyVauQV6e0LHX92ZCwlgoV4pPbhHBiJXjWlctDzYgpX5NeXw2g5gjLpgAEh3
PFL4Cmqx1cOfeRBH0qZSMpSdWhs9UDCrH34kXqNmcnC+hVVmAbzBZ/lrzXOou8RRckyY+F1e5RFD
GR1iPHacOg9zZi0wU4QFCFAVJr/MFf+crOrcnpjBeIryT6JTjuB2TQxlYl0az3LkkjBHAgsgb4d+
YUuASoMx4pht1QzwFllYIlWEh/iBa6XOK9Oc48KDEKAvPqt9YtW4PYGrct/l//ffG0L4NPvedG8C
XVjz8e2GTjOdky1lwq2+KPYuSG5dTFWYybulSFCZ58SAwg8C6Lh36FtrLjAGEWQVWnmbgOqpRFvP
VxZkR8oX1tDYhRFrMkG05YDHnwx0BcocmShZ/onDm8gUEFsfvfHV0eiS23oFEfYev1j2nh4BxnWQ
+7gzEbtthll/pdmGeyWrPQpy5zxqGsAEf1nOsoHCKonKh5VZ0/ft1F31/yktS60UwA8O7R/Aj6sq
bLQPWzy7dU8LZoakAbNWklImAukbHTt7Qdlt5qcfXhcU38J7Bwg3WOVZbONHh95m7nwX7fd8KlTx
hr4i273gUuD2+lfXnfUvb1CwjhfpOIm3sMrUJJnjLBNisuUUyqLB/QkapxAs/iRBaW+fpob4fScG
W38rUVLggN80iFzWxAfPsadZk+uzbNpmwWkDBwFk/Rk6/WhP2vZcxtF65WKD1y/5PdsP2ML5jS08
1XcsRMpHkixGFmYcWF3kzzl4MqaDoDmB6+MNY2fgMhjUJKP/gxwGD9TgCTKK0lj7SAdUzMxHkK84
pLVu4jm25Xux2Z82wEXVzjn7MC+pjABmEnMAmoGIYSa+h1rms+ZGCTtf7KLkt+NH8HiVAHoAe2nw
eF3JqV7Cy182pRPJIHqNU8SZEOnBbsakBpi/VLlzyT5R7SjBvDBXXLsdYMiYU2ed/9SRfsGAfWnj
haZMvZy2Fx0rkNre1t842Jq25GHavCDRPXmRt0i8QFnP64hHurGzpbk/wYIat2lUwE9EUoNSOK+e
oHGffD/yCQQyueBXYh+qbhShx5hGIqqyMLxnGzYnA6Nl6N/57lxtUtKmfDLdVnZbGFyDKgO60wqk
U/XdcNoxyq8sm+uSxGN4hh5ZAry2Hi/tNfaH1nwI2sjiDlu7gH6JIRmtR1zpftZ+QWoIkF54thzI
lmBpLt+9dPddqurjtLXqrJuNToAz1ynLd7fon6ZTnkAArwGW1hsZlUN/Aur3uZRkNcwrswIZZfAT
gVox6N1geWMfjbUYJf4QK7/llCs5EXe391VwVWhVeaVPFuDCddmKWke3fONwpV+bJX43fu9dAPfQ
asHDusToRvDpAo20VLbZhPa8xwLfH9lIu+dvn+Y2kCSdWNdqoVYmYM8om6CFQRkYlR8y7GdU/mAo
4EZIjdaRh3TIiCmLcb3dW/8chM/Ucizj7fFmjcBfuccmQS9Bn8g2eNE6fNOFudLP+IUtwar/PV9m
d/dzEl4EYGA/51YrS1aMKzlEaVGmqwcKXRc4SSgYF6N5bHT/yywS1djVBtVVNlH6ODafo1s5fEsA
bhwK82IS2RixkS8Sz+VvP/6bYnZEi0McD9ggV2yxFG3j/u7XnQR7xQ9Q/RTdc0IzRNuCCgHONsCz
cAoatH+0LA41wwgsaRx0G5dT3v+C3Ut7py6im4drQhxDJLDC0TAm0gz8ZUthITbPZVhJDznmr3vo
WjEkcOlwv5ag1XQSIjnn9fiahNpO5UfoFYFM5U+XVhlK0NM/HuaaRHIUL+DshYSzQJwy0pLa0JVh
zuTphkcW6jfJBLVy9eujA83vesMlsufZlzo57nUYNr5r5yHgcYlU3JFBiqzjoM3M6NKyIbLnYEfx
WFtK4U3B8H4y+HaTcf4ibP3nggkDV620pUvnmv3z3hupBNJ24VVh1k1Q0X+wQPNmOAuNz50eR2ST
hSFmdrut1MrwQwX2f/pm+DvAKqB+n90EvKluKKpamvt7B0kgJbjfTCHUJcrP2MtU3GEVEb/84CSd
gwSBaqr863hFc25u39AK35iUKeYY+A512odD0zrd5UYcf+KxLpS5gASmR+c3WtnAU+9jWe1Fld9K
YYhBPAxnRqWehrsCb+3aFHVwjo9LwHDfUq3pQnUAOTuMlD3jsynnOsMlhwIv3NP35R76Ej5msULA
XyMS1QYy13dpW4I8kbSe5RTgiJl+NpKNVgzle+Lht9kGVQwpNgrtNrZDrAinTLjqDjzM7b5R1YCG
KkuGSJoEaaVs+pKZ0zp+1AtsyYpDtRRY8E0s97CEIeMQCz7UPwLyML049nJgyxBdvqhF7iiPZwYT
zqPVmrYwww6t9T/YGh0YzonM8uO3r8NsVjrtJQ3j2V4q7S0XvpJUfc1qsbvGZU1wT/E9PPIT4Oyv
SypDnAHRc1+abEX7L9+gMy9xYG49TYXySVIpmHwR9j29qwJkmxUPwrZa08/XsjWCA8UYagWa9moM
ejIfCdNkOHz+z8wracXi45U0phTALAMhdczSA2pk3Bx3DwgNIl0VCmh93tQXz35gLSYiSyK0lMP/
N/CK3z0jNovEG88YhKyt8U+ox7+ubd3rxscuFDlDOQ84VatyJ0EK/PPN6XI5HiY/JWRAIPgjm3eB
x0LbRyU/usBXgZEwppreZxUGcm0cLH9ldNRVeOySiLs05V9g+BRHJQe/qCSIDinvvSA5XnV/miix
CRyfPIPKUPwc9UaifMK8/26UT4tgYIwTVOhvDWL3eXF6evsJSiusSYv5sFrqE+Lqh2tR5wZKKYKs
9kMsn3EaoI9wwRbC+rmxvdegPrLPX7MQL1/3nN4BuZu5aBQWoH48+42yd+fMDR8NghVc6Riq2o+2
aP4xftfYOehVgPUlBUm3ff8bJh0DP+md/X7/8SYqJEg3iEnXvin+CQYI9cbyYkjT0uNo/3fzBWFm
0Wo8YeOLaA/P+Liq8tdn+8OxrJfXD9pApfj/GqQok568LmpS/+3yqWiK1KypFWImdNoIJ7Ll/HvQ
76ZVz+zMz0ldq8d2/RKDQx3WtuIm2YprDpggezwkeC0w2Y1zZeyfeWtF9hJGD3zRnAr1AY97u/eJ
omLPbXLUrUXVDe7D/LP+IKg8VFbhKPRHVSgTMFooNXGsvB6Awrw8ZYzA4hydqAUzwUUzu6gKzrF9
CeC6R6xVzbWwOMWVT0epJpoGqb7diw2Gc3XdBOrget3pH8T2Up8O/UMrAksX/arP4X58vO+54P+f
axSEdkUf1Us0oJqOil3HVgrcq5MBXFNVOUP/mJCNfzOkB6xa1SFHybLPJuPkNZ8UJv9KLIdTyDoY
wZ+Pq50EinDIQ43L5SauJDj/35ggcZXi/4muk8uXahAJWPEDjU91nVMU3XFz+bppwWYLNzxh995H
N8S3sKIsf/5qkvnPtSlCMlzW6gztyMfrj9OMdSfwt2L3qvCeP/JD9K5OM5g/nAM5Z4twIshfI6Pv
+4LxS1JNZBIGLgjqyY6G0qxbMjsOq1m5fp/csiY6uUCYUGJ6qMzddOOY4ELTws+/doTE/9WlrcFs
ceOhraxBWEPQN6bVBUfefYy59WAU9WIdnfDC486RztTA9zXnuIHVCMI8yhrfyhpI0Ue8uREmAXIk
N0bPUNRrmp6ZTu6bGx7mglYhoRJF2IMkqLVK0wl2ACwJVXs54jVzUhhuDrZ3JySy/as4bMvZVvr0
FMK9gsex+YrSTfK3VQJzm3K5xrDhF0+5lE2kUiYkH+zR6CQBqfjA2U+7ukaoVQhkLWkgZ7DBq7sy
j8Id8FJO2PHb+YhQk/u7I+y/hPMkVluh/aYg6Fmy/9FdbH5bXp/4NjEMDXdeWrqu2iyg1QfgNstM
w0u7ewcoAWGleh+p3jt1zXUgx27NK+2tO48OD9Lc/13wOUPxVmtxJKs0cOhdOUX4wvujonBObVD6
BUMvu67cwE3o8Q0jK693M1xSO2wl9502twgiDgYGHeB5Gdm1uHAWpYDCnVUdmQmJNkBPSAuxDM6M
clkTSfrggnuOAI5p/n9PreBHFdeeQj7LgDqa/ugu1YJ5Ij1fC0Ue8nYSIb+t2GFX0nclYfq6/tjo
/ClyNGjoZdXz/LRFXXFti4VhXfloSckWkuMbOVUTis4mi+Py7qQlcZ5fysyd1QXyFvcvKhiKQO3I
XqR4SpKi+ou10/DJVVchDDzUdEW66DxKAiDAIxhXq6L4OMdwpQWqNQP10MMbD5qRNLoCWD0PKdym
sv0Oe4uCfdcir3+2oFVV+3EF3NbPhimdrTsqtyICGgty8gqQAYpDaiTFAL/Z8CDlt+okMhQFqw6P
4dFgjc090Ards/RndWAI277UFS1vJHqZXUsjp2MJSL38xuf/LPg9ScUC/z9ttTdayzlBITSu8lld
7WsqRM8aP6il1gXuqvvpjpYb/bkYXyH1FzWWS5WCOixPAZcmS4XcxrJPFvLFaWu8/9Egj7n5Ut7F
6Kk3tTeSI0JvBgye60Huk4lmjpl3iA5nqqCYP2itJK9jUC2pH4MkaVb72gT/aWrhyCtSf/XnK0uj
MW4CeaMHgNXBhXXqcb7u4q7ZTs60TNdiD+YQRU+ZOMiDyiL3+ZRvAG+GTyCQjKCHV3iqBPu8dHr0
SxYaUms1Ld3bMEIs3n86fxSUaEYGrEc8a2dGoMFnJ/G+3mBTSIjJomEHpz3cUFNELfYteO+3gfI3
sBPwvPrZrbEBknE+ZhZhsC5lO+/zL2mOjcLG01Xe+nFv98E3XOa2yBdjbeHjHtVLYOb6KdT5Jaoc
/JKKED80EbO9fYD3zSfPz+GTwVBcmuZf/+H90mCJz3ASTM9ojly230EpN64smzR1kP4sEQ1jpnP3
mmolvcDq/1uCXNvPkeGcJoCniviGpQmx1YHPH6QXUyUqoAJ0Eg0YZo0Gl6Kg4JgS1rn7dOXfMCpc
y6Qxom/mTfRCrpnxgyUL3XkyvHPXgv4UatvJ1dA2xE0vAj6B3qlif9tnemG8yZOLq9Rz8FCjURxR
3E4gLTp7/m0/PYn9WI7FvU3AHXMwXqve92XIBA1ssJB8ybdDxrjP4U4/cnDn4tvf45F/JVDw+xYr
vG33WWLUlNi3mzB6YAmfP8uIl+yRg/eSjujwDC6el2ROdRMwoEo3TNVv3ZfIGOM4TTN+x5qGPEGk
sQ3Dy5X9uwqXk2ZUe8kAMq/wUHeQtXVJTXnIGqdhzAhCgYg6LOsLdWSttfYSdvGWRnsnIL+uzlri
xBFczqoLCJn1Dll7h2bdefMKPDnDacF9kKjHiuRA8u2uzf3SnIrBgULhRls2WawXzovDmXtZj4GE
MgQ+CVSM4jfAqXV/eKYT2RcWEkfgJqMJRw+BhjjioADDGy+2j8yCLMNhnfRo517XSxzHmX9Y4jK9
gSDoaJXd4yT2wyKYkCNO9ehlTgeM/iPOa6YASrRH7VHCU1sWvyq4/HlvwaYl9silKQ3pLcdvMohE
mBWdVylXKIgV7WpGRZFMjnrm+dFMG17RFQpzxSeAI6nmvoK0xke297pkn7xl59G5jcTkxJP9z2g8
7VJDRqHSpGgC6HI5D2GD4XIIZ4FjrWh1DgPpMjWTdtDvJY+3dOimI5aYhcgr7tKiyHtQ6LSHsFKe
8XG9PWumQWxgjsJi8q2yj5sOut3S39rp7cl0xhechK0ELChP4KkNYOQoev5c162tuIVw5E2XlrdR
okuU7C5I2hz8cD54n/+sjxhiJDtJ4CAJ9URoK5v8+Lh26kDmDemUEPQ0bE7pg4c9+4BPIZgaunRk
ZMDO31Vq5ZEeN0nFVPSLTMTy/jnjLnEMl19Ln/Yms2afqcR5cTukXk2Z3ZWyK+L3olRc18lmrHma
XiSScGruHqIX3dLPG3HHhYQs1aMceIlOw3s6+Ddo21OpGMZIwgzTcIg5doiFUPEYZaALTqJE7PxQ
htnsqrE2qFxyr/4EAefbiQ5hpCmZtmiYniV4xVps3jQUik6gh9eBLPxT1QtXzQ0lAbLP83AtiJWj
AcqmoNdYTi3AKWHbq5fJkRwF3ruiH1FyvI9tQ3LNSfgm5uL2FvWC1XnVZ/2oBysIPzGZTiO/ynXv
MK2wZeWhBZ7PXpV73K23ZdAToKY42fmU7WjhzeT0UBHl2PAN8TU7+fQnlgkLcIRBcw1WQ38KvmzZ
RkYeE5FhKgd+Y6dcMdKEU9gh7qfGVazTvUMWlqYkdnTsuWzW4P82Xb9T2vXOchfuvm58j5nFubsp
AAjUwIwDmFlI7r6JFp45o+4W8vHgZolNJ9rjiYL6uJGC4/qvdCY+ECof13i7N83gq4+n3nGK+t8N
JhvzYdNup1BOwgLba6o3kZZevCN93fxN5fJVai2OTI1r2foH89xo87KL90jDAmW2E+hmX2eJxxh2
foVhKqCQgDtOiAD+tKchPAoqKG3NTqrajeVwB6kgdgWV2HntUbUac+cnvkf7tWKk6P5yBxtZO2Zl
tuznTJ4c12N2CUXxLC9VxvaaH5sa8R9LqTZF++htSzUDooLNIuxaUEL9d6mxDXXtdjc9Ntw3ulwY
9V9Y4S3JM132y0BFbm7LrL9Tva+j7q/eEmtFfi9cEqBHWQJqy+MHdSmkcO4eOMqcyyo9BXeZKgqE
WGwmFp4wjsYqRxDQhzhtvTQswUMSgmySXxfx6j3Rh8kGlqyG7AwFPnsG0mWFNTrbYQTc6a1VTXfx
nGtv0TU1pM/YdumBGyooRi1C8vRQZ9cW5m7qbxtrd2xHsutP7CQofJWl7dVPyP0IvDjf43dWcgCs
OoUQXtBL2FBVJ+fszZUuAcB0VyNdLB1/VJ/KHjY2NBMnIvmXTgXEP9cPXYQ5N5DxO6Y3P3ALAdGs
kFOOnSa++02tIxLe48QFQBNlE0th8oYOo4PsOQ4iKcuTCHTFv7hNCIHBwcYFp4pky4xbf5GzsVJX
Y5M+KnQ3Nb/2TsDTIGfIPBicPmSKbrtKRsqY8Xbx6KGAoFhZ4YHmTBxWMbjx6dmy3H4/abR7+xlm
KbDhvtIoDXWjmCoaU0qnGeEfCr/jAxZDH6xTs77YfyzJu8JC0fr7FAq9SyPYUolp0BiK/6k2eYQX
cNC39h+YeD5Jute0boQtnIBEsCvw3WwR+U6Nz6wl9tPy9s81u4RsH8XHhlz75lDuMFo5k6nRzSZY
eUH4bCjX2hgu+sbsU25X/W+GKNnpuE7OIfJxTrxSrs9FAmWkwzRu8mSBQW7giCjhUx8F1PQluMpo
TTwSN/RaP64gNZv465fAOuS3TYDVX594hwlUbfFA84Nzal8544NaxNTy7U68LfPT979vtGoMv+if
xIbWcg2yWzvrNBujjn+ZOO4s62CRn8RnmKCcVB0tn93kjUgy8TWJXKi7sKVRXubfTHkayEPwcrZ2
ba8zoii2u3MzpqrkjvFIsoLs9f6YYtIPhf/bXil+t6LwvwP5B+olVrijwx+N6dI4ot105Roy/lgl
P/RqZRvWkCuLl5g+8BIsMK0KNYVL5QphtLQAyUM7cQeqzeFixgOLqquOj5ajNhOcFp/PtkYVlmQl
/X3RVSXJePQwqE5dYAp8CUjjMDmNg6E6GllOJ4GK8leLpdCTDRZrSHWF6H6HblIysvWxP4PNjT5H
KwPOQQDZRnRH5lvrHifAIG2dwAsx6IhxGnf9jkuQaRFDoB0m/wzuCvhhvwf6wFdJK2+94KxlwhIS
4DKxEErACVMBN7u2hyookEO/uCTQKOKSqIxa6NHTdleP+leIu9yPg0rMEpDlfHzaXdCUj28vThXI
7pjAW1qCCmoJxW0xBYInzFaJ3IDL+GXXzq3uaJzlA1IWbL4pack1FOrDqUfg0ZGuhBA5ACLGd2z2
cxVJ0/3aRNVfwYd34uo77LnKnlTZVbsOFSMhAt4BoSRv2CdBcG2kcURaTVfHyrhvjKmUc+QDdyhp
qsVAljxJT1iPSQXjvhzcnbpLSJJNWg5Boh9qrbGmhbz91nunHrrwuEs5aN9LTGxmxdP4LbWefqSt
C3aDQ6Crrn5P4XrnLTOhVSzIHp5hnjsxi8XpEYT3GHlrWgR6X3m4z6CQxx5xtQ4ktHeFvgaCgACH
UHsx1bDHpu5G7yDsTQPVSGb/aLMzHJYVGidCJigqB98N0FKb5MMoiBPw3hqOz1e2kQtDuDfMLH7Z
oAvdq4mRydev3Gy3+SlKUyxKrNwjfHqYFHP65+tYkZgbYrVnVyb1IBPPevw20gQr0OYU1hLrt2Wm
qLk6n6N9dz6/PtqyH4/EFci70KsTbhTycTYJ7Bkcdu2KMYjNZcTiIZV+cYgeSGOQwIHSLxBW2ULQ
8P7wiwTvE5Q6W+Kbabhz59a8LkKAe5vMucQ8O+QDPCEhg5C7qy9uLRhzj9/5HFEy4CHw8hkTpYwb
mVor+M7/jUo6uZS70n7AWZLwTasj6PndelHr/oVbsEj+5VapEGSZ6E2kNDcBXQEV1yK8HwUXGTzI
P8taK9Sz8oCFAVWD6twK34y/D/r2+1Uo3tacLb6vtYyLz9ZZiZr2ylRplfP6mrCt3L/oMUT0hBg5
NcT+l5Up7iO1LRoRIZ3nOkVceIocEZSye3PiRnPHOAOsUqFzhOaZ6Igli2ueCxwjwp91EFtMnZlS
Zj+fsf1rxHFaKXQLeCBn3InTzWo9EuXxOM/zMyqJ6fc5r4+W3fDDcQw203Nxni+H9tZzmtUzPNNh
tK5enm1aA+cPIC3YBw1G8dAwRJsVWc1hvHfT5xn5sWX0riZe6AzFjyiLJbuhdTaUnV4KszqRYp8v
W9AN3faWCaRBh00mXI6M5xoO+B3CTZ7vp4SDFjV57r/QiTRHh30OutsvMMFhwkgyW1DceSRSNNSi
bhPiqb3cgC/hApdtON1p6ka2PEK8Wcin/uqEgt7xHGfvNeGsEIrqTTr9Ehq8wLkt+VPBcmQO2vGk
U20T0lF/5+glc6sI33Oupocr1izKykoPMb6hwps311KQWXjkEmiADp7t8FXsmJRUXuFnWvF+CaSy
jPSfowCYWD8qncjNmsjY9UM9Dh/m2zUi3CH3/fYuJSN4pFXjxC0B2M+C9UQXOrySIclwDiWRP41k
08NNHk4qDlA2JJ2/N6TxQVmDqltOXZJljmKCWH1M1ZFqalA+FYrTByWnREbLXGUirVqbRhhPtAHN
AFdzcJl1jqFVyOIyCoWgNmJArzT3jfZK4UwRldN5TiCkx8Hbtb5iZ7eZE7UqBaJUKLQ5//UKtwpl
sbMjmvYZzpcncot1JtKfbf7zL5O4Va5OXrjKZ2mTOw2yvJGEUBH8aKA3P7lqO288WGdWsEFQ8wT4
i8s2xZb5pwZrnCgXraBvsSbQNQacvegj76Wtyys9C4haoCnzVGa00M+bRz88MZgqSaPEIxIoO8ea
F4Z71BnaqU/G4WgWPBUXFSJ/ORaI7wZekqtBCIWpCHP/yTRD4uPV8gzcI5HSHMfBXrhgrZnwNIff
SmL+/71SpvtzkWX9huBFtWXnS/0cSUp38wtyCi+MNZISGmoJ6clU/z1jz4MDendZcCtoh816RwXH
CSUzOIyh6wPOataytE8fKKfT7JgEKRkLLextt0iC5W/K618ULCGLUakWNXJv9oWHL+GcuEX892Tk
sepQimBdbKwW0yQFAwnrzEF+CzRKKqwIFt6HzT5UMw4zKnVBNpleTSjIXmfFlNEHWjHrdinbk3GJ
yjFGMERUH03A7aFECy2X+oyiJFgFMnPfGqpEfZN7yqgO41nbhlsECzBl7B45dPu+RV7Sx7sUsmVL
YxmJTc66w9GLx7521qfNVd+ZmPx/FAXxxqR2L0fcvUFqHXysXCpK+W9THR6D9FSsnYVPzl/hk2ZX
UpexJBZOVJSL3Lt4eBGwltOWptOSVeuPefLqYoOVccBUzZFKwNo8DprAz84FdQp+Pq6G6tXOSw+i
BIOq5QDkTy9+EJ5ebeWR4FmLlO8T7FeyVK+Yupyzk+eQL2sQlYTSMm9gkUXbCh9BkoFFzt2ijqVh
MtApbRJkt7Qj9BWIy+pL7o96SiNDx0CvW0iHAs1dplMn6CuYQveBXcHTNVXvks3qV4GVpSlTijf4
u2L4dZMIuHbIz9lhHtU72GdZxh4ZGmvl5dmD2rFibQ5MqoSkT8vmtRValuwW+IqLenCSYOAA9a6s
mFzq853Fszo28iutEkiPomQo4Ds1uIOWwGsYSWXK/DCOSI/3b4KGHd+0x6lQEmiFgENDx7j/IFOo
BINMMcWooPK6wzDyadHLg7KTYz18BrSqUWSJKBN5xEAkdWIewjZvNo3lOEw02sDwWCbxU2Y0nHBc
TEEndE8hJEFVB8oMWOv6Z9MxKT+lvTrs03a1ABHeOxHRmsgt2RsqmVqgZ2N68DnMWjdNB86bdPVM
E+pwV/4JNUGbltIk8Zp/70tMtH7mxfaggu/ITYDuL8wslZukAq28xYlUPE1h9X+2aIQApElgrmwu
o3jDIOe+Mqxumx4/EoG1pMSVgzNeVxhojf0GA7ZWIuI0CjRl1BchHgArInvKiVPejahxa5xzMmIt
Yab3iLKCm+HBAqSzXuaF674rdwsDQEVij7uIKnNJH1Gs29RYO3T6DX4sGqcKFdfrmTKLe+CAgG0v
8e3PRzpBjEelMHB2LVtYGTg6Z2e7udXnmR8xbB5K8ln5JFD90Mathf/LotK6G6DjP8nZayUbZpq/
rankKvpHS/e6HtgNbFtVkjpi/e/w9YnLW4ws7njARpjXW4mROCeVYZ2A2fPEW8va6t5nmq6XBCU4
wOtCun/IllQE30TIwSYWnFHSEA6E/eG/W9GNejwqwXO2NzCnnmr/06F/WFO1lmOGJe/CNpDDxRK3
yyWqIsGJZL4i9KNC8NXINRwZUAfMmpBUiCIdMMK6FYYajOxc2SNw72D4a88+rxxyGvhcHmU0S10i
yuuoi+uT9FxDYmhI6mqkBaHyGx3ptFeTkA/scw0cz/OfgTG30neEcsDEexhrEui4rCCDNO1q0HTy
pTqeFHYSiYLyGQ8Pl/hbT38MDZvWu0/11/8zDbyR6XYhsjGgN8CaiC/vYmfiEK20T4gAvvoHHfEs
GJ+70hOrN2XIiBoMZpUyGjHH8YBBjUjGzBRLHRs/qv+t/0Tf5nOQWi93GJ3HieY77sGdEInbSucs
6BWSIW533aNaiCsj+Zhg5ebFeR73gun7pYTO2BP/qfFd+V68gQIokHn3OSBLX2nRqDW9klD8FMkH
sfhqShHff+Q+DgDGRYzWuAz81eGs47Y1NDaQMiwklRvb+NC627ai1QI8Nlt4SIwlQZvvZGz5+6Ck
6WKs3+aK2BQ8dyxPau3zNglqYBnek9Xkr/DNZLojvta+eYHe4zhMZQ1rHHvVesm47Dvc8lgCW7eh
ANXdZXroMRic/k5P5Imfy65Y2zszQ3bXn/YHeoFXj7oGiEnTGuT/DDQz2/kPicQ3MQtSYCB7gygT
B4i82dWnx1Bl0sEFRXhJ/8ewyV3Kt3BpsiDbXAZbPjlQd2LmIoKPPG/2fz7hGXGu6s6B9pOA8j8E
4sbg75sOCsaAQEJsYnXl6sUe1UEkQ07MIs8zzIzUmrfwCkl2f3yCg0C672suU1+sDXJiBStwpHVz
D4WlvPUjA2o6hiuDeQSp3FVcCgA72CeulT+oWs2YjeksKPS8aM9vkh6E/XMoQfX8CpPLq3zsoVGW
qJTnY7reQtZ/urtADMSherIOAatMa8kYat09UXd8Ma983CTxi9XkTyk03iH51k0WamxumoY7hppe
7phfGPkPAluHmUbtSxWKEqC/qvSYxlKPXDQEM+bkE/yEjD1Ett3rPTcyidEtPnnHnnL7JrYMlsIf
gGgwThdQAA4QV4I4XY96dRE9pP2KgDkoeUhN4qCRSxcv7+bIr4qTpBu0IFb55F/P9YKD7LRY2Zts
jabkLdI5RG4ftT7E7oC9tfWzYoO2yAGIvwnQdNRvMNpIDsErt/HT3Qw1rn4jpV3cYoNF/+oj8ToV
QFeHVJaOPWLihg1ekVtz+iJ2tU9xAM5/Md5HxFQ6hkfqy9LIoDjG9KvnbfepaQ4PMSnf/JoX84RU
bxdQOP5M2UScZpF5GZ2oi1qwLXx3E88BAKOIaEnUvpRNouLUz4HXS+da6jX+EoayuJ7UaDJkirIF
aC8oalfjIdRAGedMOth3J1oquwH2tRrepSM27YabwsFosARv6IV7XEH+kqb+umqrUmNH7HCx2cAs
TngcnFNv97MblD692/9vWl6UuPu7pNlP48azqJ1vw4wTFC9pFvSvLQI5Ar7YxdBxWzGma6+oAWfv
+UN17+TMvnINUmLKzKg8lhMa+CA+FxbpnSnExaZwm6GqeAvWRlYf6Lxhok3+HXSRXGXpe5FplEa3
4DkZIeLeh0isaP9Fib03a4GnP+U6bcRomOhar8UyKyDPFbbe368DGnJ9AB1ikhhULVnzlC6z7z7q
nnMWazjpKUIn4CLJvwGkFfw2bUDj5TsnVs9GI9ExiD4Hitvs3QFR39NVE0oilE5cUuD2O+RwZ/bD
RoM0s/DeqkuatFOLJ+xwlYvfd2sYy5RMZiX9U6h4A7bOrEjC71dXm5HLIPYBynifi2QJnKKXF0zm
DWIAFArhhGo9/Hhji/llIJSdLCNnm+DOX8PiFQkY9Otkvk/Twpkpl6Jh5Us01Au5f/sqg4gOwagC
1QsDtkRY6UOscMnp44RGPaY1IN1PQs0nreEgx0552jgnB02TaupUe9IjGqt4SGsQk8zdpDYm9rdQ
DTgL2eDRBXOrUNnfiUK1ZVWvE4jV45h1acBFRZSmSMIJCLxTyY5KTgHD/DB6Tz0K6hO9jltx+l/j
ylQB0uwpLC/49o75BE2quHKjwTL4cBe9e8i3QFATACZaSh7IQye+AnYpXOC1roQYmPHymLCehKpC
P9FXW0FLugNVqeDrDYos17Ez6qr+xr1++dM2EIJawzY1BUd7YKsijyuyrpmdvLSXxeBkYX9Kus4v
p54SmDClm3zFSoTwneY7qMpnR7OpsdwsmMOTWWgK6l3R2Dv8wOKTSPKZP5JGrslKouQsFari+dvh
Mxfai7Dj7d2cuGzvvdWf6p/hGzfhpGvobCVwmH5vVuXGMi2yXpcQw8ECbfbNxXKaTv27upK9TL04
zlzJT7kPqeqk1SW/gd3ag6bMxjX3B+vmv7EXII436+6IGFz/8CMTGQMWoI0R4+kiSWtHSgTbeTud
CWNWPCoZLPzYPsjM4kW+l7YH+/oB4kmmuy/IpueQnKr7x2NjCocHpamfVqjIzGe1+11zGpvQpSLG
S+14SO5tGztTmMbh+f6wLzupHeYVmeLYM+qlpeFi/WN/qh6hbxoJEh9c0dWDai6xsN2CAKRYJZBf
dPLl1lXjW2glOVqcYKSrmBFAgEOC0vk/NdasS9QXjzJHDwgPxQ8KMF0gbzVR1I4tin4RsN8NAP7m
DOjpe6JOW9DNQOzAl2aK9n1Hr/zodqLJc7OStPPjaRX/1EX8IsShtge/2xbaahGh9/YkzopPsqpK
IwD3QKfJdvmeXZswB4/bAVTCAxPGbkTrxEsAaVUNGo0lUdoIt4S4jfjHCWqr8X/4AVqyJTfXavKo
s5yQ4rwlELdHZNQ16+D/yyuNaD3Gik3x3qCS7qORfcYITk8Osj0cPiGVhen1GGyLvVGcjmnZ6vMw
PNz72/2oHhvE1brUy/zDXk0RdITc1GD2R11HD3SwCWI4TkKzKZOFQ9A2ikghF9nvBP3AiU4cjypH
2U7ZICt4sMqbpnzhiEtiIsCIk55qidnd7Y8bzAhkVRj5d2jXTLi4mfV+jFV+spUyNf45fwG3SRj3
rqkDmsaVX0GideDOBuUX71TZXF62gxmEalwKIBkOdzThS7kmQQrM98/EY+mIowjQZXBTS1sJWJo7
HK3YvMk/tQqnXBid1VTF+Nhvj5rO6MnevIHEfAxk4pVi2cLhNUA5l3y4GfBYhJDJeY/fJbYuo15b
Kuai7v6RXjKSi/8WIrHDBdEbVCz9IqjAJu/h3iMrpMHewANKTfbXCYjegwkVIR/xi4zrVVLdo9w1
jkhq3yXqqGrr8RibGUyMNa8htvRwFKS4l3GfKOm5ArlJuz1ym0tG45AVv4L57365hWZY7tY538Ju
qIJ94B3hKxVoMHiiHqWIQS+eLI+0Cf+G+5CkROUVyMXFw4z4mSeNdFgDXfCicK5lWwbPc9QAH9Vg
CX+rG2x0/g32pnsdEG8dNezCGjd3L7KlZqSpCBOAxoZgNcmnDgYA7geydKjIZ2trWEM4KfM/2+HG
r9cU1PtQXDUgHxA4iAMdNud+lvzJwBrODRlLFIbeakh3vYPmHCJrQSNLD1qEkKVLaDcm4QXHH1os
HE3EKRlN03RwSeytDJlzNSFQ0tCc0Rlj8wUaRZHY6tvg4gsKrD9DSOjSl5lD9ty/bZ1vneKjwKrn
pc+LmMdYC6hqLqpupds0eFPA40td2LU1fpF2+jkvvKo0BJdwvg3nDp7sYzhiAQz0fwJGoWchQK5l
83eJPSFBgKNg5oXWmzqSgauBwkBmxde3jaZKnC3ku8pJYe0uZxcTA55RJUWZFZur0vuoSEYAPpL2
FRdTSTPWrFkbgUwc4QP9asmlXFY8eQlAAtCH1Y3UTHLKECCRE7UevVSdmHvVqqd/r0y/EDc9QsXP
cBb7d0cRv31RE4IBbh3ZkCNVRPRQUqk8eN17iwkL51aqZpyuc9HPn/DlDQcB9P2dwZaO0dUOaBwI
k3PDQ9pew/PhV1RxTeJN8BoORRRT5XpYOL6DYpD2MXF5+x65YvecBeesNJgVTtU8d5TY1toEW+/q
y70p2KaDq6nq09gbG5p9aT+wB3ZpIH2NZVXWyltYWbOvY7LRsmLmTL3SiwE9elYXCR6gK7iWy9OQ
4z+Qh+MA3Z+s/23QI13BZKVjALCgBpX9w77wHJOudl8DZCU7sGovGlzIMFdHbZdZTuTK5OtYeLUB
Lg6X/ymtoEjBOAwgN26KxNrOTu7SSX6mXGi0CbBzWc4uTZKRGNsDqLn8jSyAvnSPEWL1g/gdEbLj
AQdQ+cSKGEWBlhYwUIPxKmblvHiSgsMjt6AKJJaxW3GNpmee/CiROokp8VXTxqoWKZnuFNmO3Ci1
W3dWwqzhqANocEDy7u6oUCIZxmHML0NHvnSgByHvC+fCC0M3Y4MARX2Lrwel1zazf2wSUDbN6OtB
iQ29rMZTwpZqvMAIzeu9PVRKyl+MsmoIvLqVVD++qgUNJ68fefDFlo9KR7ENXIquzBZwNMiiwgj+
i8ODMLa6uG7cGfqrNxIh1Hw3FD2UM2GnPWqiFPad2mfaByvWhGMxklPjNNa/IfK2oJQqFsPN4OPh
rrcZtWlACaunJJEHxN01gYD8/ySw8pJiqso6gH5Dw1FUhickNZbgD/ED+bt/Mga+DdPJQvbBR3Hp
188FuJRMd/QCXF19wWrI4sXtbCGRR2a5mhDmJFnFN9IttlacRnhxzfi+AEut7sS+aIQdgWlM2b0K
CDPoXRiNJ7U3Oq/RjcBqheQEfBgrCusT+04h1CWl9ikKhZDLBziF7I+NgXpmtv7stozCrzqBYjve
1anj+/QWI6xTJuTwv1vjfutcJvd2o3luklFikKBCEzPiuguOT900CzNzsXfnHhwMt6C/b9vv7bKb
BsxuMwKHtGj4jEIkuo28YYVODLt597WEhXBAA3IEeFGBOH1o4icz4EGNHq9XxhI4lW/6JjFyzV8j
KrRbHe9gZ0M0x64LaOhEzU0MDuA4c+y/ZiTwY3K8k9Kg3Tvmlj+RaycXm0+kWwzvuw/XGugBIZqY
mh2yOI2APTEgoYZpnV5gpEhXd2C0gUj2Y2u8ndv56enPjjgcKa8/Yon9wTc2S88Te07T+5l26Oys
kDjjYcatyfO0hYohkqyATnXjL/ieh+S3/zSqZV5T3MFQ5QXvZh0OAqeLR0Bp9uQHt9b22+noGTAA
hz6YjraPoQ4wvhhezjYWlq84IR2cAdbau7BNiUJVw0uHjUSsbz++nPBvGVwxDO4jvrUp4iBRK9aT
SbXmnsFrkr5FNvqQPJfh/cos6yywqyjcissYVVkBZjC2JtD9eRd7/M50VjAkC3meQd9j0S8NBpyg
gC7FVbnrGQF2N817L3zsZSrEo7TU5iaN9zgGYJjw/+gDkHJcHmUr/GlmCK2+cOn+5txvieEtSS2w
9tg1oEMSCF70gKVfq31nbg5+zUv/b4s0aeNec6SirqvX8nvAAr0WkxOyaW3aQF/TobVCd1hVeBAg
hsgwjp+tvhhfE2CzLUmArtdiFIsfBt6xiwDfnZDSMbXOVBUY6LndA22CO1++0868d3fzMEt1a70G
7WvuzjH5SSPZGqyDcIB93K1sDsfFWUzp9sAsyHRUBOS0AeBkphI30M9PdKepGMrexZd6783kXHRb
auNUE/LMUjTfplTbyHKNFDaWxb9jT70+oATOHCGW0VaXhDb7TEX0PskIEFNlsRM2sQ2VdjS/iPTF
YON1howh2iZTlwxSt9ZX7P2atM/B8+Daih3v5HfFp2uMbG+Pg86lSOmcjnaJe2fDioQ1Q4nVPJvR
mZz7U1MVfWXwW9gNqASE+hNGPIdYKX9YdTQTHAY3SqY00ANRrMjXvDuf9t0WMI2hFLoKo4sc4zop
29UbL8i+0mqe7K0ixMPHlvXyFnnjE4tsv9Nsa2yqNpeBK7nR6WfB/GoPjaVLeU0L3DaJ2peMSzDu
ou+NfiBKKu6YVr1oz1QRDgQwwc8P5NjyEnYbrlmeqKuQWQBiOQTEoVPAjJlUcKzdpeM60hPhQLiD
wm5bvqTxiS4ujjDO0XOLT4T81uqUVyrtf9vK8QZL+ANHpeqC1q2G/RdjbS/RXZW4ukimZaK4a1Fe
/VW0/q9CLmq/a7pTlwnglLvlPASEnJgi6viot2NvyExWHHJvBiX4+f4+3NpEnGusugUZhbUUn/2I
0Jm2aIDI/wnqJJDuTDAV+VYCAqViS3KXzmrgHpcan3gfqBGCPHaLOdPVS0X77sL7/9p9K4xTXu/R
LqTFnQxOelUdi0zu70vPN1K/JxsWkJ+5l1oFXX92cbHEa/a2I74KaRAnHqIFHIhiPa8e3QMAK3Jq
tlzIMXDsg7yUvB79f7DQZvqBwFnyhfg5Zin2Xp0AO1nr4a3R0tTXuX3TCS1sb9bjJZQ4mkXCIGpl
1P60A8CSRAhzhwCnUe2U4NLjeGFqJna+HIPgsNHJRb3E79tNKnHQ1OcE9Ud3ph5kSWEtKgpcUm6A
zoH5nltEbMmqhYYEenw3qW0h4yLO94CFkvnf9KLk7xSifXsIfiBdJGFUKcCeW93VFgJbpkzi2TD0
2jKtcggV2VO/W0HLFoU/ITCpUlxNmBqq7O3KGpDkBUncsiJrCEeubKUjOAqyI5/3NTcPR9kzB2W4
sRlfwZBTlubYAQJ+Cs1bccKsbZQQFAd7NYTvO/aOinXiWXjTiIh6AglyWV4Vc/dnM3i1BfdKwB+r
odFo+rPm13XMPWpJR0qmiGl09yOVWhl6PQmmRQ4RKlED1kV30CDWW6T1cUt23f8BePrmdiSIlHpL
TrBBiudr1JnSVuho8g/43fVV/tAHRUHV5KXoKewSwJWqJNd2VVW+evAEd08ic+DFA0MrpKAcn76M
VjKeRvrDU7ng0cmrooW7kqub3oAJw74LqPg3TBIcqWIxU8VUosMnrUxsZUOc6ip50m4pWg20BxZV
r4rutuuounEDJpHoRLhbn7ERMFFDGRlBenlpJ6egRq3jZ8dJQJpc1q82+U2Hxf519j7av18mXqSX
kqaxg/i/c/gTP0eW/Hu7YCcrZuVx+8Ml3foGF2gVqcK7wfJS8g4i/HD++ql5ANY9ljrdLuRPFGqZ
hlkXKSDK7njX5/IELs23maf/cPexQILDKgLLmqSV1wr8TpFWZbVa+HcPVb0U5qKsmb/Nyrr+YyxP
go9sU6QHoiKU7TV9peMLL91ufNQhft20ebHQ6fPIFvjXOMmiIAxd9jyW+b36O1O5rPkwTYlSz3tt
53WuOaK9idIDVh8zOiUftNkBa1ZP7kw57l4+S4NxC+7hGpDX/IJjEikJ41iyqIhG5zF+OEw4tJQd
G/qymwNZCbdkYm8viS/KWqP6McJ6v1owOIRmNQGQXQ/yu/jQcsmUqwYXSx3MgGEGxPglhRQ8sS1b
7nfiAf4ihZi3B69d0liKI8AFMbA056r/gVxkQ6brfvgGKP0qCpyXzQTSnsz6Cllw532FqCNegt3w
//V6Jq5YX97ClX0xYjx6IogFXIfTNeqcR4RrBr7uQUHK9knM3P8F7pUyv94W8D1aXI6hAMlUmOoW
wgJAdXTqxWHAZe3fhhJy7lv4vhl7B3ix89gmznil4uicTFZoTF06r83eqhWIUPbn1k0dm4n/dO90
NPTooubu5U3g7vTQeqyYYV6tq7VtI4FueMS1atq9LaeC5ZNigcb+hOjOI2oecDQvgLwzVaYV1Prc
uoF9L30p/5rphRk67UdjUhI0ZZCVdW7HzOvDjs0Bhnupj01u7nhd93kvKhgtkk1o+cpyrDtJmuxj
XSkwPxIhTdX/t9wQWfj9Jj/lo0GV/YCag+MEqMttMxtAf/+RS34tWbtVa3fG/Mr2zuuqVThD9BPR
PR5xP78TLWZLXPWnorCJAD9VFcMjYzvMkYgutLPnjbapclTh+yrrqcq2/ld2c6g2Lgwvo6HSggpv
al+HhkHznxDptYp7mxT7WvERVrO7d0Vf2eZeBIMhZh19nwzWuCAoH5+GhqnRa6fQhCSOfCUqdCuh
9yhZJWVI1AH6YksmXC6qbxEq5R7KUyU9s7Ly6ugwMNCyZwREHttvb/UmWJllbgfU9fDnncqZxjJ8
n4DpgINmaKWvGlnojLkriC2kegrY6zjbTN3uvg/YDazhqAQfADi3o4PTl4Mg777zVn+NX6saSPTX
gBuu/SP5umLpsLu/npSbYQQjlS4SJ/R58HBWL35aOA33KC7/flc11Zw6e4I5BT5IXp4w0EnXN2eF
TXNCwm+Q/TKCgjudF9xY9og8I3U4IMFh3MjRq7jomUfMv6YqlermZCiacOf4TTpXYffTPB1dSNMn
2VJO/Wh4CeeMgK/5XVEq6osMgJK9Db8+XjCNAyCc+pxMGLkV1haA9691y5qufeBkudp80sDVIKTs
1ZIkQFMESofmtwDWKeOaMuxALH1EATwBUS4WGjVx25paD7sjch9FXcbK5z/WptRFqp+z+B7B37El
NlbXzijBnnj2aimLK4KKwGObnUw6Mt1eTH4uu1f8hvhDFkj+KIs87xSIstRWmzdx7ugXqk2w+l0w
SkDv5tcUb4AsyKiABx0pUm90JPrA+M9nUn8qGg6DqgUUV1eX/eakta9AYraR3FUh0+G3ick/RNLk
fSs9wPzLjUCHfZ5AAQaYJjLV7BLD+wv4ENRvHIDnWrXHHEhy0HWiszDrqktYllraZHE/o6uFK5by
BX1IgqbL2k4YAeeV3BWpmHnkVC86M4fsI8CMtAtpUYU8rq1N74bj9pNWv5M4ph9kfw3cEhMk5iwF
2/KmYKvczRnWT6QPKm5o/OKNSiF8bKgS/pyFwaemCZB38GBFwoxmR9kkSRZHeqHlg1b7ivNrg+WL
gkZBDQnx+3xeVExDlEqrTVIOOE+Mwwusd/AgHMiQYGQyrfT7EglgwmCZmriDuzWt2f1eBroRADMX
wuaU57YelsjjMNQ6qRHswQoZu+2xUYT0JMooPZobYE4BO0tocEvYk3unfvFiBba1TPfAQTm4UtbW
hosJcW4OkVts7cSmiwTBxwmDEZbVck761U2S8650PI/Al/TIDiDxBhiqWveMu4ao0tgXIdkXr9Mj
UUlm2p47X/t7s7oEfa0jHmzJpWQ5f3HYvchVbUue7uSTSJqhDi9njRuyOItUOYLu8WFXEo+Z8J/d
yOo+ZEOMdeTHjKOc8ESMrknV9r19P4aT55QVFhmjQdvChVdkSZeQqKDAQFGl+11bimbkVL6nNwOj
vacKe7RnqvAYQNqv7LxNg4qMnshj+z7+0ne+Ro07gRpjl8ZQEkroPmEfKDRcGKNDTleYg9yr/1qd
mHKHJ4aBtaNTq5dnsdJd83LQn8+r/yMqQgQ5//gdkPqvNduYC+7EtE5R+AkfpGH4ZS+HpimoxWvq
DoGvAweQ831tcAiLHGmSVxhg3B/NNd2djxwxc6v+boVEE0h0tJNYNs9xzAjKtxPrrkT1nei39I3Z
EuYN7Pj7j15FG/RNxhUv2IjWEcOCvQ8DdTtRN+VExu0WiKeY53aFTS2VfSWmMJlLFpCcaPW/mE+H
iFhMncYuQEqOQtDkjVKXV8Vk4BLffUGf2RUvV6WhL5MoQIm4Or3mEEO24L/mQ6Q/KP72KoGGa7Me
rEcIorqvvy2txO3lZQoLr6DwW9LAezborxzHP5T6N7xk46/DV9vkKjpbEeiyYiiE6XVODFBkYxp2
vrOOvTiApT+ZRDC/94HgKvW5rHvKzbZ8Q41HHB8r7c0mLbI8TlbwND9pdXbQCQapIGkZJHApQ3lH
of7Vi0iZB9JKEDttQXnws/Oghur6kEAGI1ac7eAJJq3Yi0HHigfjrWkJCAMFpakPcocmdL9F6wXh
4lv51BTm6cwgGK+yX6i5lRWO4BGx5ApAB3mQsn1a/0T6bhR+8W3zXCWZNSjbd//1MzrNhO4sDOwO
qmxU6mMzVxOpoyhnQLSvmcIVK2LekAowi0RzKCR9AsOvP1SVKiBdSjcbpEKNZ0VFFgYebgvscWaC
4WifxOdYgEjoVsy3cRLA26X0lj6DUs2wb5SxnZrFYVWCuhHVzZCQ2rY6MR38IIcrXqPCm6eK8CA8
gd8qNj4orNV2w5iohLr2jO7fjnmcJE5MR3p1GT4eXwRDc00NF6YEBhm9+fT+xJ0xOJk3WNTzdGv8
HskCXqTi0IdmI8Wci70OYZOsgsezWdk2RYkx2+pDfTqAfcDGVXCLtq74KWwq/uIkebpSq2OrmnQN
J236gDU9ZxdDUZvld49gkh4gWuY/IxXldAwsZ6H8zxh5bheZFFk5oitHRBE+WI6zsKCbfTHlUrJ3
4VRk5Hrd+1ED7XNx0bU4vxNpax2qvoyJdhRHnLQqSYMTnEqm/2LAdlvq7z3pZ84QnIPTKQ4lfE4o
cvyu/qlR630yqskoXY6DiMlgMCgvHqjx/ggS/nacYivQdbFXhsAZUShaublSheQRlM1pZ1x/Ay9l
lp8BQfuRjxNEImkqFX3PRa/HCcNUFrVjlJ0Z6ADYebZVxIzyaEGMjZoKz5bg4OyA+s50ibOxjQGm
IBjmxf88noCht21GcCQJXY1Qys90IXn7ZgtxHCExCrsmMx+1lPL/5KMN2klkNcVOynr2sCYGXwUH
k3ZTaScpMQlUErV0P2DzZ/7p08mVaQ24M/SRwH0CS9KXGKU5zdtsIPip8aZVT79XiEG0F8txpTJx
VkTmKymdtuLZ/MlxP7VxcrwAV7K12ELP+sKGZO3nHvFEbMBHgdIPgidSI6hRITKUAMpD2sDC9IMJ
11kwDF8bPy07zbdTy0lvZrw9v8DIWkVPdoA3wdQnrQ38A7Nl4pE2qWz/T6hAczzs12JXZd7QpECt
PF9+lxxcwxR8crdiXwEtYTxq4gOW6AGB/kiKG4zKMyl7jGIeuJU7SKFpoCsqIF4hTEGsyavsJiTy
qjP6GCtAMqDBSkkth2oDHBMH3nYSjbVtNnxEg++jceNO4PqJonqXD6d/K0Fjh2mKCKAzfyM+JhIR
TIj3HdvC+nJZ3oUfzOAi2Twuic8TNQR93AmWJAPN6hEyM3jRG083ixwme9rVOhX4CDjqffvY3Ff1
3NQIm3NIiybXu3V9bUP1rFh8Zk7U/ilDFXGnDUeBFIQ9yV/QjYn9veD5E24L3v0+VbvSbyti/dHY
yMeRfpgsEVkhgbEjd7caN+GZ51M0BNc/BuvbUf+OOpwTiJDhd7MVuBEZooiSE3sqJgPy617K4tIV
F6PtDfUV2ZRvjHhJqWCOsCHTJww8aeDU6B1fE2uQCEQO61VLYbiBZfjh9+bo8jCdC7iFknompYdz
Pj82MdqEUcJyBnPZ4HjKoR9pssGaY8TBthHRS69VPaZo753oo687LGB3SRsjMMGD2qqMFMHWDdeV
SczywOrd/v9175rXqDz25+v0NZaiHwdLA3cdd260nvaSa+YLzQJaQsnQM+us8/4HwqwPJPFQtTMy
kv9EJ/ypPflynScURfus8wllWsbh/2zL6ub7afVF+qWmuA9XPs3g5soR3XmkmOR9MfDd+YuXiVKT
ZNISZuTnGPYL6EJsBhIlaXA9tsaM6JMM6Bt8cwaSHvBNd50yJYHHEg5hBVHKdLTBiL8jJSplsPsL
vkoF442YnDgwnRTcGyaGfaBAfI04zh7llTwiiBBOa4xG/9glsLTT5h3Jv0GvcLQjL+M1mDs7R5iR
TqHUYjzBnuNU66gKCMGzk3uZfW/cZDL9+n50pW64Es1O4Mv1sHf3AovKdFHS3WqzL4MG3lHXryGu
Y5o71t91LTvaeFRvwhjzGXCPmLJ0UukZB6vZaBIeJ67hcQb0APAkjPxJtNUnodkwvguRQuYZBysq
M+E1eUOh0UBW7ZV1kE8kI4X6HqS2KK0yM5SkkCrWJUQ2h0tE6p7QtqQP/YnQAhv+VaLr0rPA2rg2
DC8HZpTJFad9KtgFLTDTsdPBo636hhstAORnXWp+Mvdlcpj8/Hz3zvf1QvWVKuBNul5ab8oyI9fY
yxowgeoh4OhvV+dOZnl3SZMQpZp3SI+thR6ySSbZ9CubSDvRSuyKSe7WaI4SPeQNwPtTHsJsz1xg
E60dd3+ATBJrTQ6lAidwHlbQTwrm620VwcSGNEA+H1+wu8EoxhBxOF2zfdRMUPYd1lE9oq2QzV2J
gShsVkmsocz1TS3EM8h2MNOtRSiqO4kOKJ5BPyV806/TI3SYNeaDBrN0tcMA1OlbSFV3WmJa5mKE
I4b5ufkU63f5Ca6+B46DQo3SoOccyHwrtPvz58N4bJDnKDRQYCJ86HWsDqQ6PlGoU9Lct6C7r9YW
gpS6B/7JtOeU4eSSVyed7Zp4OB16U6KBP4aUSwDhRkEhlG2kJAroN5cSstVvNwLgkdpEng+9+0vx
KNpQYWRUIjTA1G0xhPa1g8//3Pn2FxOqTlI4zxfR/btjFFxLqlexU1XjapO7biFuNJeCaGziaKMK
Z3/7zeU+7LqAgX79vaUYqGwPR3aggpHHtyL9d7bz+C7gk4dijACtzZoZrrBmedTIKcjYYSJhoBRe
WWAFQ+k/tQ7fF52UpX4LKPJPNCzBnLK8AIYHH7zkE7IzPWPr2JOah21T88GYdx/ohtAOqPKw0NlQ
z/44JGDGNBfbnzshVdmGZGMB9tnir0kH107Wn7RAJqZcI2rotKDILtvtN9WUoIFPODxIm3J64Z+7
m40FPt0mHsNlh4eL0VPrT5cxL3IaNKeYeCopFmY0sj50cerf8Kfh7IXO9Ofpt4LWAolHpwNM1Hdm
0FwtMD+lcbugPiRzkULA1JAEAWr0/iVAAoPpSpIgQqdfNTqXvVvxRK8xPna/tV8kny35vvV6Cuf/
mmvyJMxf3PCwrh4llZAUDCzD5n65gvkY9tNW48lYjEAOFjpDpRRYR4amESgRar/vWHO69qHOZ8w3
DwvbYod3oKXOVhXQ4Bx9/PNK3h5R27+sdWCOEPJr+nXSDlEIZxEevXfmfKiXaiqTsXyu1/68WqPa
I+UCpEa4NOV1APiIvK6hD0gWqCq572xZMsyDT2mW4LzsVppy1ZLeDHxMYOrXspIKjoHeZiFbwp8J
nKvqDVHxsdrwMdq6DzaMBJXUoRO++eHJbB07wRbFbifdw1eoCs7a7ePjoL0PsodJ3lAqXXl4xMZY
SBQXlBix7ES5iY+dcN96s0GCFYmncP1WPtV2e1hYD0WmDMyOsRphjGJOWY/nfXcjq4rQHEHjb3xb
nnMVsEdQw3MgMIYuR4hV23nTlL2pEsFY1KiiDTLamccPX0XjH9y2DOWbh1hw8BDoJFUyx7FPjUEP
bpw5JGoBBw+No+M4tQQOWrQSvPH7biZ307jxHXw7TiB+ctdyfpQw1rTh/f+xp1R2gX8x151rOETo
C860rsVM1asXZiuZzR4xuykaBy9AtIzrYiDr6JcJm1zY2ySTX+VpjgOLwv06L5tAI5uLp2y/4mO7
CnQjJhv8EyDYUctM5U2keP86I+CZdtUTUN8eTjWALFoe8l/egxnqSSks3rlPb8+jmTDrrAfdEveK
inrKWqSM3RRVVv1+Qrp3ZX5d54jyWkZoW1H4rmouXyhwSLmQi6+KV2uKTkzTRHv7VQHco/24SdR5
H3j3u/JeWGp0dBLyVbDxEV/qYgUiL8p5wxQ7+vi5ZTwz8QLR5sOd5CZTIdpAzb1tbdDF2cJYjONa
6I4zMckb12lbNKBs3lt/zkk1jJdVeOLLUTdVaz26lGhs0EqibR23Qb4MWzblbOCa0kRf22cGbwVz
QOYbAMjoogcUCaZfCH0H8ZVZAX2XQhCkFbGs9pvE8N5tB1iufCT3tW4JGUDBWmShQ8f7oGWUPkEs
MdXN9GcCZPYSVirVt55WFTZx7u5uorgzPK5jdrZRWwRx/qgC10GW/1vG4wF8RzllOBShppw2fQXC
Eks1gfx8LZUmSrQ9DsM2nzaE77h+mLuC9WwemTjmZO6iIIs3UaQVO9Un52OBzHko+QGbETdkr5Lc
VA7xvvcjBY0bhvYurzuXHHOj3t+He4Ghhix8I58kZtf8PIWMuLZ3bJFUUley0uv0XF38Iux/Sn4Z
MxFSndcd6HYh/HUiCURa0brPkHsyvzyyffWhmK7FjI5fzHEtL1R7wgYafC/sQJpdwRr7m5ZtUQvK
fWlydjlZQz7UZRvvuEwUaqQs0jcuof+mOfcon17eZZ7EBFZ72AK8/cWx1U4XtXfrdwzJER/FWZyR
7KrT4v6DYM0YDbn8TtSrT9GQA7Be2kI9muw7R/WMPKx+2wYsJULwmJACv4iWNYyXZAszfQuektEt
QjOeZrEEB6RdNLRxJNdQzuuWfBRj83ZbeCsquW/3/L0j9DiuoL4OAZK5fDnnY48t/E3n51QLNsxP
OQJVY0n8Ay64UfFmiTC5+prhM0Ens+gKgVF3VpUNpPpZptwlHh8TvQCp9YPsfgRnCyJBNuKaxHeC
wUe3RP2LIXxv0NBYbPl9+7xbI9FXHPWODZGrxdHbqdHL9lEmSHRa0LHH9/0JGdBmYFL6Wt9CFmfW
KjKkU3JOFGZQu5uqx1xZx8O00mbM38Jx5z4fnbJZ6CIMTOIr/vg+M0DcoLLw6dIDlNottuiiq7h3
c9WEM2cbjCfroL3AUEkLarmucOXPKKm8QSh4zj/LP1aKFiRQM681ex2xmGLiRQXwppYPZdopb0IE
nha67sBa07cdUOCUod+jRoVHChNDptaXRmOo0kz2ESt4EXoPq5VEEvE3R93K5LceOddesc0gzLfj
fabq3RgYQLwhvW8ArMBvmt/VnQj2C26AYsxy/VBfEEBNoYxQmDH7OqWnAlf/2ZmlSuKlnfVOweWB
7rXMRANTaWERIfOhTr17wjJvHDiPXL1aVHB9eRAl7r/h3LNNUsrXXPReKCLIIBsmOXLDd0Js4q3l
jqQZGL4QnnqH3//qoVG14Bd6pgE7SVbB6dKk2P4zupqbwaGaqI/tbpKhty30QsGGpqIX/xbHUv1b
+BcmhRsqqnoI2vDXCtUYGO8B0kw1xxYFbxaO2iClzMq4UHdFDV2P2xp1AjvEmV1cfWdfNj+vxvH3
eAou9IJDTkzp7V8GNPpfBYOuQMKtJCiVgapgBf1PvOXySzNg7EJt2lLQC+/ZYxPqGyuZg+Oagyju
LKbFqORIBaSR/2SKNhbXXfORqSYLAe5sMEzpoFkvXX1YBp+50+6VhC4/ikccqkmlO+UUNPmPAXTi
PRPgsyVt1bZ74bjLff0JrJpguavPxYs5HoVjVnBWLsFm/JCSsiLJxpzoEvrTcrMCPsadRczR52iP
SE+rHKemEV0M1e0utWI10j629sg1lXI/k9yxDIplF9gyQLWf7IkZH/WBYWrRIZsqOH6jdSkMiGrt
UonY6sr9cpF+6YxPRkEyvLT41ElYMvxvpKBOGbE3irzdkLcBorRbH5zDve2fQZ65eIQ+86vFH1qx
9IdGgxm2rWfoEpD7++NKs3V/8vvRqfEQl1oRNDkuDdG5zUUG7wo+q3GewZwzEDO/X1sf9MFfUz9x
N6vLO85GZuU2IFsg0KVN3UFgScF/pvZ4ZWoH5tIXw8b5bqD7nQnJc/mHwNl8b0XKRgtPRfUGck3c
TTicXgJL2rAlRYwuxWiczReXAFKXJx6XeBTC1CABFWxSTDcKdr7BYKPpMernuQtpz/MfdluM/1Sf
paFge/LpN+RTKMIF62ialqqiATFdkgaXD71Qxe9lGzTe00VepdBSBPuRDuvDRjq+QmBgfXWCFJhN
nDDpFFsHQ6nKeN8DRJ4sndlJpHejF+kvGhZCAooWhNAbqi09XARG2t6hpX34V00AdSi23VRJ+ceU
a6OuIstb3y4dUDWUJOhl9EGDU/8Ec3SjSQsFiO/kKyMx8BiyyN8JRx4qidWTGg/x3QHp/8ToepVr
SGEFNv4byxltsLXPnFYiRoBASB2BhhRm5fYQazKzBi39vP88kppp41IHeI2VJlfKPIXOXDI3vbNx
Sbi/ES10Px8hhQySJMtuSOX193v0dnndYLYDQn0qanSnTk2kvJS+dWOlX64U0NV+F5/2yqshebHe
zVbG5ZGmHwAY3JUvmQJJCkXaYlsWLUhKJm51lGA/OFHws8fhxzb6bBOJnwi3wrRf4pIuxHY6dlOf
7R5uygRffY3I5hz13I+8fQsccnSHLKoeS3bDsA/kfY/9xQ4qXU9szZzh9yvdoq36ZPTPbQ0YI6bS
GlaPjSY+h4TcB+O291uH94hTL7TBYNikaLyJDSIWIhX0CYiRS05bITRuQNeAoe+fDejFMDdZA3nj
eOiHF34P0WuKOhr9Za5IRhog0N6Iynmy7vJJ89Qf0WXW/lB3UdRNrEiWNJMvEVNjOSb+8QSkJxl2
NOJ/UXeMqrZkcCn7GZ1pzCCqeRihhmSnJxePu+w+O6aPkX+LxffvKBryW9ZjsoUNKX9Ut6GPwQ5m
DV0A0Zhz/WpIkcK+Znzpvrka1AMoCFChUl3xEr5+HbRzT967yRU1JimnUq98RLtVwTVusXc3HVv9
09PJ7yKMUY0v4ji7lToUGqqeMlXQ3/2yN6chvLpijlEOmfMGP2XSMt7uLzcVj4u+lC4g0c6QbS5f
i/rKJkkI8AmHIW180qL3Eb34q1XDOh9uGZE5tnKwRKHgu4OWjc98ERU58YnZ80iG0mh84Kg9llSq
M56oxXe/UoO7CebEFLl0zeioGY924V7If3yAMnYUvvG3Kxxo7layU4IQ6NYjQcRWxNLg4oyaSMDF
dQZ8LXaW2tcMpmXAo89UoRHRhiHJIoZGTDRxLs4tDMjHLzNcznk5vTBjhMBkK8ugKkOr5Owoof1Y
O5mYTeZ4+f84R9iGzBHDxb39fgon6VzFDoce7zR45LJs3xvg7tF2ddXNnUABB9cx4P+80puzue6B
wyxyDBL/Gq3F7P92ITyr+523ZXOotqLvO/leJa6pl+YY9d2juWeqIYJ7qhmTjamIgVuVzkMhcsMG
si0h2h66TOPOFVvaHDJjhsYDGCP9RmLH26PuBF8VxX8CgNiLB6s7yUutI168EMCqdeYxnrrGgMd+
Dd9/+OTQX8743fqUEhi4kKan6ARqn501JHug3fbPeB36FB8SjFSHfUdD/PC7IwNZS4LICydObdjZ
6nIc4bMcyMdmVbZlYlP0wGdllaeKVtDwQGjX9+i4jmbzE1Nqhvqikg9r8ahrORGAoug5YNSt8QRL
Iyz0s7BHP0gO8Movw9oVFL0nDMr4pERgPdSeLF0WB3cGlZ1D3Rg/zTvT4dOC+3JV272LHylAY9Cy
YO1JE4v5DmHZ9Af982ArJSzhPCLHcap8xwz+aBdvIKGnueLl4LNjsJTXi9HzYANDjT6qzU6k7QNR
v885o1eW+IrybKptwsxnwJefW/wmciwiubTVYaKWPAPSmRlHYyI1m1luzkoG7uxjSF7aqDz4VjAs
D9sKolxiqCWHwVKx9F4hinWLLPG3LnYJAu22so02GzOotLIgQW8FDVbpqEc+LIn2JQ0rA390mg42
szbNajVtizrGhWcIdfI00l9Go4J5H+jR4eOFdK5xDSMCoAU0eBdEyLVoIeXXYU2h0DqWrPVhd37x
+yQDLB/wgZrxenbW2xvjqPxqc/zA/UTaZlXVIP7e/+JB3USjj9YEvl6tdmnU9U7oBMrWBFqPTimY
iLvChxgWYPKk5qpxkc6nyYJUT3vg0MMtSA+8g+tIbQMplQtRFC34xmlj+aPOWCgeG/9VNVoXiGUj
MKNKjNMeym2i6T24MqWdsLKvxYRR7vo+XVLHKJ9948/GgzVJJfj/QHDQbQvsAkC2kdfsIimV5XiN
b3eDAq712JXZQ7NNIlsQjjXVbKN62U7YWh894mEOrR94NCfdJAXIOI8cpYDo9zkGxc26oPpzn0oV
r2TPNIx41aB0An8pc9VvfIsRarozQ+xdCJ0JyWcDsmu3TVUqSsq4zFCViJ+H0lyntvys+GlfexWD
q7EfVHAZZmNAjHe6m3ECyGHooZOZtAjpvyMoQsrHMGYA8vxQbUXrvj5aSn5zgcqnr2ToEf/mmWPA
X3GlvhDlW5Q5AdEio2xFj8iNzQDxSXDdzh4Pk3+TpK+1qU9nHEmYQ3ZwDf52XxNb9xFlU61hQj4i
DOE42sbEqn5eAHVFmqzvS6+ujv/fwlGb1mYlC2PxHGOeCcJ3bIldYpQh9mxhfGQJFwDP8kTY0XdH
e5c3Tedn1FQod0FZkDTmNvwYIUaMst3CfDXahgn+TU7U5klUYlFzd5bw3E3bg2+7M+o0IvCEnWTh
6goYz3BxJ3vXUDxFAZsuxa/U4AW5fX2E4ZbT2Z0eWsds2+1UKnJfsZF57pLKw2zb+JOsURwt+ETD
MRoOtj5ajuZ/zU1DQ5rLloOx3yxSq7qQ2ta/lvrm9LdtMvyxIdbLiYxGSAqfqkV7qQyQbhwT+aIn
7pPduGuTdGQiTKTWqTfHkZPq+oQhsNEFDQ1sst9t1+s/rmYI0VXHpFG5FoUrsFk//d+Qqima50Me
02H4/FrrvawfMoSKG5j2IgTyMqi7bdX5Tz4XJdWxA67vutuL7694bG6nUm029xqIAhvV0EIOns90
IOMF60C8sqDCVoeJAlUKGo7tOKau2Lnrv3zTjbKpyngsUJ9k6RhIJXrFhuPJEkgGqD52bu8L8Czh
gs5RxnNaqlGn0EqNH+CmgGqD19ElP/j3cZrXiqrjxpOjYvyuKnr07N3ttFrMWJSZ30loP9la+4FA
oTKOPIfhvZXTCZ7KfutqUBjDTni2woirgU3rL9o+GWmN8konONDi90vcCnSSLH7zbFlUkfYYdNhe
x9CjghTQArX7Yl5tqmpjp54uGKrYakaYTWqKsvREY3H8TgYtLBXV6Eb8IfzNv7uzRMo9Om6Z97Z4
yXJ9lWuIZvbACFwfoSjGV0cON5TFcxHw0Uop+hi2KvxaaTIC8MVZn9R4UmxqLIHk0sRcLpY2m9yI
8mYuOrf/DkNF78nd6LeeXKfgmZXIPIcCC2NI/biXvyiLcMCAe1Q8Yo/0FWXkEfIwo/HAYsd8WU1N
5GXELPS3jg8RqKie3yw8CtPK9FoREZi5moTwYuDAoOK52WhSjyXVylzMhz/MVrXWR/vt1gZ30IVc
Nv2nGy0PxEC2ZOXzj7rJ8dz17XdD9kBHK8wrX90Sl05YmSLRvZUfag7/6OacrIWUMzTyPYZB4Tk/
7wovVAd/dyl6Zl3sjcnf774Ad6HADDDfPe/3ZoZdGxyGrw5MBEDrBSNiTNx4AU2VhnhYVPswAxS7
htCArNoJO5rD4zQS6N1QBNVwCE1NivzI9fma+dL8Xmar+/X/dilzy9aR3NYqjXQvyAStyOjHkzdp
wFWmtkmrcp/2zqHoYf73rxVrXo+NDL2trDYwMGRF9E/eNVW0tbD1xwa90vmjh25XVBsu0IoIR8Qj
Z/hGyPwI87I5is3a9nJp0YsfUSsOdDCOTiNkm1mkRaOj3fgzirPHHO7QhsgT+B+i/9IP6UqSQ1T3
RRaA9Y5YRKjoXCWn2eOHGi49o6r02htuO1WZ4RktSC3gsGv8yqVounFTLctKnjM1vUvAeB9kURKx
YJPc6lmNVAbMWe0s6EM1zYByXOcS6eFc6AWhCa6ITxwE+YYPVfufOfJLthvxSkmrUo8C4cxXxtVG
o8fRtQMrYuCbJ+iqglSkT/lutuU4x/c8oqTv0sSBBoLgsZvMUqH57PwaXkCeG/nt6u8JgwQs2QOY
GatWtZQ3/RsrD7h4c3qb0wBR6h57ZU6P2ihJKNVjrxBXg9RgqgP+ZQe53TIAmywEi2f7Wil3vX1Z
wmbhOF5IrzrrX08CUKFcZm1nn7He18YS9feAIHzXmkWPyvROCpv2oE3eukeEWatkcGMT8wKRv1/A
ruXWyQPtSh5gZQeT7zrJzaGqj5lJJIgJxOp12Nc3wOZ6M5PPm3QcuGMx0eOG0Wp0nZ/27f7iukbH
LLVc9JyFvuKrcivjt1ck/0LrenpjeMqVCoK6vhzYkcHEWhROW1H/+qMxWRuZdel6UCOUpv703M6e
GQ0AzT9wO39Owv47yAErXSqPWsd+7v4keHXa2JUucqLF8xv5uAIAJGLHl0LbwsvXmArlTBLZUst5
raPQbfObg8j8zyo4TZh4U3DtJaY5RgTHDzxyExrUSiz1v8IrIVfb/BEgQJdTiQpvbYImpGIm8lQW
FjAgFqKIeVhpM8KsMFl5WXtYb5QOZVqdi3gViyp9FkrUshr5pZfCYAirOO0WJKm2s13sFKpcrT6i
SQZgHFYlnXJNkVjZalOT1eqHXI3/G7a8NFhtzSAerZJp8YGMnybVi0DN5gm6h//DQOUuCkcMiZOY
CFSLm3i6eYRIqFBCvqylJpuC8LIF69AgH5Bm9lg/ptq6uMPPhKQ3LJ1hjHC+ZQ5Uc9aVSherLhrN
v/0gaA6BkWcSEwViawC0/WfLGziWwZwvylnOYeydnMGXmTwSFeNaPsUPClPeZqD/S0rRzmC6bb6L
lZKMDEtBM1UUPtLBcWh93yhWfXx9Iof6zgfE+5SMW0Wu1DiP2GM1ENVmd0R5SEN3K/muJa3zkqP/
k9azYHWASzI181kmmomdsGSBdD0MmbmsFkcPvuzuymqwN8BT12E1HkrtPBDa1R5a/V2UovC5gzBk
rxxSG8Tuufe68RJm0f0b1WUO+Tj44FGLWtIXxEZA6Av7QuHT++xT4NuJ6sO6bBzdHywi8VtkjmOI
bRdes7wUfd9a/wPaglwlyrmMgdvpf135RdrRWdxU89v+PeIUAAFECNNaUPgALJZcJPFksrETplUy
iL/qYAnB9d5O7gsLqnAc4tyeiYabRNrkAcC+/w4X+sjdmSIKuVw0ZgpKR7Jlt1yGFzXLtsm40Nms
wXsAqXgln9lrs9E6/rEXwdZH+tfkRV0e/Ke6MrG2IvLI0Mm2F79Dp/7BVXJi76mFEF29GIrmsOM6
ArDoQA+GMV/Hbr3QMcPYeC3JMiXVyVOfQCpYvSRdvSIqY9I4WTpUv1mtlR8Sr182OjBroIXapHsV
Dryz6NnUi5WdGdoU5fUJ5JsLbUhCqoOedo0VGY9u/IPi4inHZ+op9mtT17jwopzELg61uGgqIZmr
D9icEbgXLVwMZf3xosbt/hFYPDsoGSeKUeyxF15Ne6tmhxB3dJv7wvxjkQGoYi++DBYeQoVMnHp7
vr6TeNAHbHTF2UELqPJGA+tHAn3FbzQ1vCq4L5cyvLQgBNd0i0btOluVjYt0nI+9hAygGDlc3Nqp
ymT4yEQyDWCIybJILFwwN2TlJVZiAfeEkZWtbe31jCNd4q6y6Pcth4PJeygD5US8IhuOuEqBC7h+
IHqNPeo7GsDlq8AMfMt6BXkaWRgl20ube+IqBD6s6xfF/070vGgO/tZ92SfBBx/HHEWD/yoD/f1p
GijsGy1NjZNdInMSlzRo5Dx/DRD5YcBEGF0KjIDy/IFCFlNloReFRNQu2cEni/1QivFL0nZkw3ET
kQcI4UzfZ3IvjODMIelGRTAwuSOmCP6dus62EAzpVSdMLKxlMdUD3RxekveWh5XNsrKeoKtrXoFv
snfXxJk1xc+nqCr9+rjw1JcNR1YZJdLTiA7lay5P+gPwNUJlkrXEj/nvsuZvuTpnMnRI1Sz3tiK3
EaoqKc4E1qoy4goVwk4Ro0CgKGD5n4khhn2WASgk7nkYAGMBtpBZ1+mxvBU24K0kj4ViGWPZvwi1
Z5Ow2cudwDbsMmpdxNUYmrvhYJov9Uc+3yRg92IAbrAL3TceLm2G2ycF9xuknxH3VVMpuFFDOpyP
GMHUNQlkr4M79VrSdcuf+iwy6eQUmF0r+m8puRhQLNnxfX6EsSweW8/nVQAFOe1V8g9mzUzXJx8l
BY45gkbfWis09KL44OFbIfvrS2UbBTkcL4Gjl9d41UoznVqyS6z1nRn2ASN3qieCy/lcIi6wmoPv
oKKW18yc6CCAeOt991EbwDcHsPaOGa7bOunHJyEViCd+2gqx6/CM3e+P4xioT1x94kY1Mp6p6/OB
RlrB162KhyEqZRlLMcEL3SA1sfNEI36mvQZEYTDt14Mgv5QMjZfOxHJqdvJXJLwM0P7PdrvOoBBp
aI3y3K+3Cl8gHsgkTyPIn92lAA/PU8+8qncYuKiJxwUdsZ2HbWQawqqcUTqBuyNQ8YzvIuQeDmmN
45/dygi5onDmaBH4ggYr7/audjuo3cgdt9bYjYybdhmk9OTg3cAEMl3Mmuhgo3Vts+OIBs5N2xYN
+aN+hw+zs6KgQe+pIud5LZzqzCUnsp16q9tsqQbgUeV9pKf+YaxTDw71qZVQbzxU3s87jE3NT03p
CreRgQ/9LSNg5Y3O7ANoYtoEW8E1nce19GnYO1Dfat5X1DpbfaUqH+EJrqRZozwRki219hUNZDSD
vCewzpcDdMxBaHx8dsgobds5H/snhlCuMZ7RbJPeyV3IDI7F2IbjlnxJuG+u6Znpfh8w690KtvMJ
AtTV2n/486lARPhv6XDriKrxX2p/l45WVC/03kK3k5l63dYqbMlvuUjaRJPUTV9ZldWZ91/SF6b7
mguYBYmH/2SeYxWkcB6ujrkeXEH9vrRTBeCZBhgJzj+UAA25/xOSsQUyFaYRa1ueJFeBIALWbn2z
f6nznVnAbxno6TFeIT/sXdqKPsbV7hoZT9rADZAxMIvhPD014KibImyhovj1PWXA5i9N2hUA1kFg
j3kXcZzyJgW0A8u33ajgrQX5NnsmxWt8ixHuhnD6ZCIenVolsUnYsijhsf5ynGFxjXHQhnCPBysx
e0TwZp7lnRcM+RvzBhttt/iWGIy6J1RgHwFwd/abc8EZRe4Hftt2EP9WshBH5b8nhb+2UqG9gHTU
s/EOuOmluXBvSdNgSnhvV0w9rhkFCCILwijUqjcTEjmX66Q7cVhvmktp8MxFWv7O7zWL3CpsRbST
oXrM9KRqRcthrpvW7UIjaXnx8G6Vb7wfu7VW7Jjaq7jD8dikUW/02UEFBAgQ3zvWaIxKOsKXb6jo
K7MP+IaDbut8EgNyDmr3OZxrJ2Kkd3yDLTTyk+B2dfTft5K376oFx7QeXZ1S3ABYuva0IANYIvtK
HziDJHT85DLhSCxtGYAlE+whs1f7I9j3ARzx2wW37c34/oRUoHqrDVnUc816NjYopNFL3TiQop+0
OlbgCgzGh0xArkWKB+bhHkfMFq6yEftjtZpJzRr4E5XZXEVxAS3bOu++mEbhWEV7fJyvIEFCTyDt
lhRLoyjT+jD+mB6Bjo+naFq/vWF3Flx5dXpCgUvePtmNsmqQuiSMxE2m+4+UIuX+0UcFwZvmAlp2
JHTFDfC353J728PmZYqbSZ6RUvd4BcF7YQoAA64Eb8qlHiFLFOzys7qAGC9ocPRQ7KB0d/E6pX8l
CEUkUz1e5KsQFQ5kiiC7notWJsyPeHNUDiu7s/+HmETOXLQPLc2D+s3sY7lA5PHttHoRNTNLniev
DETceo3wQP3ynuxmorTU4/dbXYmdoZnGAkZbpTmCEMHPnOkqN7UwgY8xlFEEDXPQjffqnnKRfC3L
ml0iRqzl2AbnS7UqMh1tV/czW2PQ97kWEAi2+68+4MBMuTnJwy8rLZuBqwAlY81r73Ou7Bx0cFec
fiyvoS6ZKB2rAx73Npzd3kS+n4ErJ2sogAWl3Vy6Mcp7ke31wYrtZo2LIhQ9ENJK/fkrpyD97fnN
wtBhls/ENw3w3MVmfJmA8KhS1e+EFtoaEkEOtCGIyb8Dl8nDxad+DvliHPVCMa59ntQNiIxDpaoW
qSwiBVSG6e9gX0m7dGXgy3elMPuH3kmcBd2Ki1ElIW88tdK8F/V7BLp27EyQHmOpoMFOxm6o22qc
mCCQNpgKfDd5YiXSIJ+I6U7nCYGM9Swio5Gs9CmgvdlgS33ZOOTA/8ghQIpOMswgAlM/Y/vGEYVm
rPsq2B5ib5j+ffiTInnsd3gS7TdAhz1VdzIgqovvFgBOEZIHwL8wBcAFbSVponwJ8vCxAReXvsTu
aPsf39O2JKOBsCdSVNlSqoXYJSowVFBkrhebB5ZifbaGFHrF6Iz8woYF4vZBRk/qxKF0p7tiiI7h
v4ROILiqixVNuLcX4CV9BAT+WV8FSDNW0ygCEn5xZ7mtIfkNFmEdZFPXrDXrENoB1MSdbEFrrrx5
SeOijAijWT3fnR5mQkCJMopT7ckMp5CIHT6RGvJRkl8u9qztqis/TuLUCfMO/898oxHMJUPekChr
qTYVIYon5b9feElDmiX7CZMRhurWPvp6Bpmx9wHaIUa0b7qBM3HfacCe7dF+Fqfh0HRyeX0uNF/W
4SUhnE8fZgnhjbNYRzbdW73KB0NoSakIPKJIh2fuDcUgtyshRYgOmaNZISNGDV1u6v1OerCX99U1
0wrG4JyNfp2R/xtynvcggI5QuV5tz5r766qwieWqhbC2fnUzqvi/9Z7k5bz4IKVPccK6kPTPcC22
oqX8T+bcxpL0ByYbSzhbkwCeDIA5l4TfS29cAD4I4V0myoiTgbGTSw9RQvo/qYdTL9X2aH89eT+m
X8O2CSphmrLUYO2g8kQvrogA9CPfUETI5FG5p2wD3/PPz77gcFID6uzUm7B/yse1wmGBK0H43p2c
XMkJm7cKAHL78e+C60SHYTS2fYu9TGygbQ7gQ93fMbnQyQYjx79uYZjp87EgFfPlAF2Sqn3MLtAc
iAzYsskORJtWG6+J4jxoDaclzJjAv8C+Urj6Zav0LrOZvgtY8CEAZtmhilChrX+hOyLm1s1Dd+X8
FlvflaD0AF7C5jdsgm0mEuY8jMOfk4bbP6trTYL1YKqdejPBF+D1XgtouWslTvKU/xmfvOJ4BvPz
XoggM+bCTwQx1xE0UX2SnkvZSAmdCEFBbTRJpyxKtuTm2WkTlrMkJCjA7Fami35wgbcoxYfbAMZo
MXVegThGtqZKAnplrQMaQZ2tP7gkgLdvnYzghIesp8KOdAHjPz9fYzFO8u+rYC39ITggt+t98IXu
ORgEnUaISvRzrM0qOTS14EBLV1HSfkKCE6IBxTwKfb2tuffwCS4Jo1Ch+wLgdI6AHZ05ItXkyDKn
KsH7uuzE76l/nprsku1fw1ru8JpIvg/qE6pXxP0JxTEF9HYbgBqj+v+5N43K+FuydSh4rrHYgiGm
++FJoGxXc6G8o182Itjrz45jTibSR+O4TRbCXURwJ2TOlrfbNFjWjyQ6l7cDWXopeCkA/fFDxlbt
IXe6cDJ61nZ+Wgv29I1KsFgAdyQjkxPxVGos8yxY9jVSWIxivHMFxxwiujUiTaVsB7b+7mFrgdEs
cecbEHKoEW6zyo2R0aV19WRCDqNcUhdwADnaQM3d2lC00xk3KLwH0qEdMttFIwWPiGvRrJb4umJx
dSdcsTM3CyYsT2w/jE3zjZwp3n59RRGhSdTkrvoIR8ATZ8zNQKJGSFKpIBDDK9rfpbyJMQoXcqqr
rWMlKwgPrJmR3iyNIJk3J+2MGS7ZayCaWBUnGUhBaDFLlSz7ekkecepQ5qa8mhTAh98u12XDTENW
VtVbMoG2PRAR4K6aPH6+zufXzxNCk0f8TW/i6ftBcsBTE2eFNJNQ+VemtmlS5omGlGHblZG7BlzF
avt9y1fcv0MXFl2CrgMqtxYvZwMBJXNOd+zkP/z10X+qz01dafYmK3fXPPcyigk4rpixWr4kw1az
643lhrdJEqPIMEhDYiByNBEYB5qSs4pS5+0c12LFX4aU9ETYJksDmYKvDe9GAbfc763apU+A15BQ
d5wopcOgx7R37g13C5OZESP55XAVVHzPglClok8OmO3v5m4JTctKh3JUEPgI77I8AoMt3+l/RepY
KVV9I9rDH7iy/nVlW3gsJMFgjVyT/CuaaHmsIurRluuojwA6Xmq+wElxTAZ9qmWSSIjuYJ7f4QPv
fBJkGnLfdpc9CNdNCCPLV2t7wdDASg6SsvgQ8mWSOeDojLg3DeH0oAv8N8dYIh1xXjw/NGNATMGs
GLo7r81NCvlmQmfTrnTw+q0DvVhDF7NkiTNbgFpV9oLp/ZykMi1kmt14gfKA061VX4WaRbDdHKHT
lK/vgrfHOjxOQdxn326KVtulUwuZT8tyAchkPOL2+Qfoqd4GTizXG0k/gyei7R6TRiBxB+E9AT61
5TjrFvnGiGD5vpvjqWLJhuaA1Idxq+et5s3jXEda8+pWO5vvmxfLlrjp8QPq/7boOroEH1/Ce5yp
sUlyK5qz5cv/tTIXPn1Om/Fg9gVf15/5loHUW4Z3YTE8HwFpsnI9TXnbOm9BiFREQaCtnXgGYKVr
mN1QVeRBk6NduRyjQD58971b8X4MX5QB5hmkU6Oz/bfTVAmNAJxUDn4t+4r3Cm8YzV8NlMR/AtKZ
T2gCa2RSDeBquFy4V2CNHgRDr87yldVJ8AX0MHB9d7vmTJzAyYpMk2IlfkSPxOnS2pV0nHB42XtF
sM+xeTFwPWvdfbVnTL5149UyIlIdWwWuW0wcUsSHv9od/hjcRjd3DLoLSMiK+RLv5RxQNZQha/rk
8qqAi5dC9PglFn30/8qCUfbdum5pFupUmT+m2KLYOrtNTlOSu0SDyh/0kcTnxFOehhWkyYJaNCQo
OtyvB9rZ8lSVkY+j3tpeexfzZ2AWKgpJ7Xp8TXb2BtQbPFRPrY6UdXXOOhySAvk8ydkj6c+VuTEj
7g8JcwrICRPgoQWLp+rGkBRqbaXt03muheZzkxq2nt0fAmJNNbEY2EEMKMKRdr9DpffdW8kNZSzq
qQQ+PP8ACVffrhT3c1A6sWiLVkc6zxi2c8PtEQngTPfmthKxbNyXV/dbfT7hN776cbLuoTsv1ndt
rUA8t2IT2iligrSX4Rb0LRRqFcwNV/NwCofcknKRBTweB7Z3jF7d6s8SsYYEjDvl/HCNhMHyYzAu
9E0mQ0Zk+yz3M15SjESp+C7vexYR4Qem0LMTtHkppT3IYz0AJfhJJdalD0K8tCD/wbjjaU5knToh
tgGgkHR3547i9le5y0UGWpFiuKgPiOYJ5mv/Floc4l0YWUEgq0w8V0KYOKkSPpDVAZWuz0EIrP6m
a95YQJdrl4GphYBWbR7+TCnX7VJrCuVUdMgEtcD6TAA3kM6v88hTp1iih4bVq184QHd8x70Mh/qR
9Pb+lFF+pFxANs8dHdnBMabAeH2uacezA189c0KjTIV5KuT+50pzedS+uBxm7V42/7WDTZ625eBV
yioM+wBjUfLr9vbU0bSWZ7wjONSRt/El/5iLPrjgHJ0LqYFT9yj3UFAQVg9dkNWpE/DQEs/Mzhoy
H0509kEL/RIytKELaIdlO8Vl5zD8EOvztAOX+7tjvyqfN+JDZIU0WXCcZA7ZQ0ESlKzTyVRyYDVC
kJJH4tCViK2KV+Jpg0rHg4FYZP38v47bAKKV/O7f/S71ErFntbApWqKbzJ6g2+7AWNSSrHbFmL8g
HjWuhbNsHz5qd+39DOnNt/Zv7iQjFJFl/BPYp1wm9AatfKoL4dd2YbAnxm87vNBmtQaTygFZOTiX
Ux4wMhE3W4yHbVLQCMAebUFaTBWgPm7Qi+/Xck2G90AaJEZ2A5ByBNKwnd0ZHs+HpBYSu007rm3K
4ZWYuRj8KWbHJiy7qEwM+tz0FW3FE11/x4eTci8mJTDyqcrm2u5Z0wYdsgAX5fURFz9SpKaVXzwX
rEWtj3e8aezQS91z2wt0YFREe+msbOk5jhJ9Sva51Gc/ZMFHALW2MiecY6BKEGs3pVYVy3y19Z90
0ItqTZUIGfCjvpFdVzUdaz8xf0G2wgfdeKsa0vPKN8TvewtClHHCypHwCdEkl3RF/6inUgSEIQag
X9tLk7QxoT1Bcjus0w+Gjhs5cIyYomhzvaSR+HDQZyicnaUAEUR1TvEcoxKCxZ39DS0DBos0CaBD
MKiGC3/6PCaStz2o1ToMB4m2pGqmml7WCtIxL+y0horvzm5HfMJRJyq2ZWEDj24l2AmbfGBM3yoM
AMTC2v10tV7LKkl461efm468IvfEJBZbjNN/29kJ/3VHeWFrEWjUNzcAhHNq42mdSX4LKdS8FZfY
vFIT6K+4mZ6wQtW94w99JifsJ/uXrxcP2W3VDNtSuZ0+eUSzZlzNZtfP1RvHALS97lbeTK0Z45ws
4cuHUnGtfeqJ3GwCSUv6BfqOK0HX0qzvLMTWOg4+/RLBo07/aHfZXqADA7xJthWbIPZrEoopGcDY
o6tyv/fcMlsRNI6Mxwmj4wEZ2t7/caS8A+KwmgKZYL/5h4xUTFb7dB0ybR2QnJa3zcBXY45v+N30
JVnQhBPtPU0bxmvrPMiXZ2YwRZe6X0gIG2I7tl83qpTckpy6purL5FCB+fM71dfsmtItcK0Yv2ZV
0Ebxwt2pnLN09f102At/lqEFMJQ0PXoHGzwPTF+u+W6h0qen7WKdanNQh4cF8tAHhlOk188uR51p
kbg+a1feuYJtlcNRB+SJ5O32sAfcrjklrNSmHQob2CB6XhMqelQ6S+8zces0HaY9sJMR12PyMjp8
vAy4bHy3AajRvWjOzdV3AfhvbtL5qoyZgUqh5Zfuqb8xZWFnCZz1PKFBNp+gUo0yQdn+fP4bVbe8
AO4pd+tATC+bNg0pdHMLmYlnUm9xkEyEHWBmSflkrflvLFNuEf7m7pP4NW3MLOzdrF2WNYJhj4oZ
q7Y8mdnYek5OH9b0JMl8NLItB8wyjowkgEWwb56YqzmomnIZXFgIjK60bdC4+na5cDdt5pmQdBR8
ESYnatWBBzSfUS3oXVthA6OpmUkZvydv4iIhHNkKoIKtBpSfwFkDMLvMOGr1c4oQdb2TKt7u2TDQ
3RpjZfFSRp+f2CFK220cv7mMG8uwnlejAEkSoCafTZw1j8xbLa2ucQ3J07T8jTy196nHHLzJw1Bv
BihagNIBGckQ+h5oBwF2OdZRggy4rOavYr6U2HtQSgiIcWFjGbxImMqwd9SVzDygEuIivATmE9la
tP4c7tkcFGmXxuhPhjCaVDR/V382wzWKPTzUDDDTcDan3aAmwXjjp19/CS7jyMPSFrhRvmgm/iGy
I7rH3W2cjnJGLAJjXXaEDnI51kIE+pqDGRalpKvQl5CfaCi0vMpm1eQDaPrQQ/EMT9xdRXdAxYCs
fRG6shNztM89BsaHw+9vG1bfATYmMFJdjV5cJEz8mFQ3gbBTP/T0E82H7NikyGfR2ugODZLi8kSr
K5EgeqwmUIAtDO8/SPNn2HmTRNVUPuMS8ALDs7ldG4AvOBWdgbhys+SYuMYgAltCI8bwUKKuU52R
NyBxGOAeKuyzLRmYTA0ZOApNQSFul9Dl1PHnGRuJaNe2gp+g10YNrPLrpzgDDLDb0o+8i9U6dyyh
mxm7gQDnjScDtIMHN9n9PoTWwTixEE2COcmAdoCiGe139iYs2jdqQmlt/Manm6o88tvpShP+L401
gMzBnARwm91ssfLxE+ECbnkOg83BPNr/cFeK6npG5/O2GJBuFRQZOo0yEv8hZOVtDPut5cLvNVVL
8ojqgI11u3nVoQkrVwjD48WhL7GAUdFPTZC9/H8mEmcXicoJ1JLAlAgnNBMhrJBmOrlSz+lACmkm
J+Ou+RNA3hqfi8RuMC2Xaz1laNnRvF38qWx2EoI0qZxZCCfXgvg/cBCYshmdLz+1dUBfAfpH+bQ1
s8GZJRy+xhXLQiyKNM+tiol2Y+lJfLRwqYtI0/Z5FlwAFrT85N8sV04WY2UWrYmdXyZ4CMhn8ieb
uC8qFchyW0gGKzgloxZPwsUgFsaZzjiKGYiDjqqaICgb84+Gnsp+MPLCOOiEXLL3WzGy8P820gtO
bdvTRM9rwO7REDsbVl+rqNwqM1WuFSA2Ny9jtIwDMCNosW3J4SSG9oF8F0E1+Z2tMqtY2NhoL3Ps
rSxEds7vg0EEmz0ECOYokfO3x8Bs+wvAJ8hOa51qxJ54h5mvRO9B0nlgGIoUNAtxqNUMaiJMuS+o
poLIRu8WSEAmX6KXRiDZNgHcY35q+6uTjbv3mGnh5MXiPX7jShb5LBULl5Vt+VsTdPRDq54SVSyM
Mv4L8jHzIc4rVLLOGaQlWXbEYq8rJrYNYooK5mCNvNGz3FqcfAJCWzvsZjdmJ0Nmc/wQcaqleTAa
dc8mryuZBI1tCkIxr7d7yyQEY+eSwhcIlYhiwZFG4WqbxxGpmgUH7EnDo7iZ8K4J6rsl6ENPbn8X
Zk8cRvz0zcosBA9DiNOjGF28Mxsoj/M9ysRLzx4ckQatiSMWWIXtYlwHZxkH5JS5xyYHf9tEsVlg
BNJbI7YZBmZMA4rH98ctlhKGoR1rXyi0Ct3bRA6LffSxj3TIn2VR+DWCjRCLWpjCSSQqUC3QaiXZ
Ec8DA5kGbou57zzfdqi7t7AVNripMKWatVEqWsUNcXZNaRWfhJmHQbZfhO2Y7RQizMLpumdKMx50
n2h16Vlxtg9wzOb0/1uU9+s5TkbtMhyHMTeo6c+ht/KJtz/5kl8TDMeIAxSCQexK3YL/X2jg098K
i/1uJQiMVuSOGvOviWpm7HaxX23FDaXpHy3EvN2HuQtXsuxGhvjPmvTCdV7iNAShQ1HYqlO2SsBQ
f3NyEjjYra0GK3x/hD9LUBZ/TU3c5ruY7KQAtV5JbijFzj0b/r5x7IBqMEvl3An6ohd7J7RvbRPE
vDeetItkh75bGwxTj3kTKYr7X8I8XY5xD5pftsFTc9ZxXO7NEE1atQMgcWs+ZKuNbXdBd7zSJvOz
IUCA0m68aN/GlMwBxNG4L35m2PZW8RL1rX699plAtHT4vNkdEmbI+mqNyzbg+mkimu6sZ4Otc0ss
t6IS16PgTIThX7ee6zoA7h/eiJ82kl62PROwyhZUZTrv3AJVpBzSTecd/1rVkxhYEz1VKQf+uUWQ
805c5wbE0+vnale0AtZAWML0p2gyp9JD+5kkOUXJuk0xVHVNbMqlvDzTDKR0OPKiGcT9hkeRqMOI
fsoFoe5o35vakERB6SXKQpi5lFJ1teawNV9DqURgDAKQzg3D2rWfC7wIj/9PO+HLQT+47t0tLzet
ukBtt9U6b99ku0sZ7fvqcp1NHQ6W0Cebg7LaGh92Ui6j1qf8vxWO9hqNVkZCokIOYoTwJsbrwE0Z
sqatk3LTMx+BYYzALzPKhjT/W2YLynQ+3IYVXxgjuW0/ysu62UbYSG0Fn8aeU3+j8udV9yaVo7rU
ppRkDpi5AJ1RGeYI+VVz03omGCQt4qooT0bHVTA3IrtRhGS/VOUE6VkkEralajyQWfWW/WmISy82
FnKsvnrCh/rajFmAmn/cyPdDTteB4lq6qv1Bq8Dpy7uL/Qwj5emMv5Q1SuU96HakZbLO72gVRYER
gZcDdfQpEaA/cxiS9mCdTPpaS6xeRHIQaELgfN7woFv8rMgtK8xyABkTtqeMYALTiKfSpGXWvpxS
wLIpdfZ7QefLaXj3DphD2z723GVCH1JdFlrK0QlksAlPwNsSDzPfNQY62Mv8eHG0G6X4+uqMUkHV
joVagbrffpxEakvb8TB1CrLomiq+wTaSR9fCVZ8iLwko58OtfBQCOdIpnbCovJqAz5n3Lp3xcChh
2mlqpZtzbVpuqXoiHVC/nnBnu21a8/KBtYxcpr6yHRkX5yPa1P5p4svf51Izfq6Nv+6noSspyfXe
T+26jRyaJRpg4euTd9XaE8LbOTzcrhHEtlbyU1wiyOHVMiooPd4r6pf6HLXiFoGpTRfKolLzvZgu
lg6dj/isq9XLfyjY1VXP+q8UvxevJVwzJ+1xIdjB7K4udCPwYm1YWSQo7uTgwVYkExDruI6lMNmI
JJ9d3jsGXxlNRR0QfwoXjbL7plA6BHg5jcnD9tjJqmk/zYF14VvVr1xXvCizFeaFThFjg2flf07Z
S5rFWgqU189vFFQSI+y4KeRj5d0loKAku2lK2u/c5pIthfBxTrv4BkWOorunAHc0m+fp9XO3x0zE
DDjbNm8qgqYVssNGW+Y+R9npp6QiT7DWwQNcnYritYkCz1N52iSBfwGFJ4EMnOaNxXAqmvkXh5A5
1yuL0QWoET7eYtdqgbvKNmpOg0a3qEtOF8R9CPIvL7xGtyNp2NCPV4hTfv/4oQM/rTfbU+iFehQU
NQwJddNmYX+HkPaqtORjG/HO5/POhqojCjIeb+S6hvyDl5OfAxu3fXBF9rIUK0HBfAIPFy4l2LKJ
ad91JvU223fi2AnKOR1VCOEo/E/6bk4/YOh7g3oD6j6tTtcdKXCSEhTNsBjJlpHqJORhizMz6vsR
UsohrRc8AI8IP4wVUNdWwk16o6MBYCOOKpHDblYaIFf/WhgETdGdtVwYfu+fj4zmwmSGtIQk4o43
0CPsxLiu25vbFXFvvaX/RkdLFhIUghVeXJ280M73Ri2XldwcnuBGi6E6/f9NPEjZ+So/kKbw+yDC
FkfPOmcQi/aj35XNBKozEQI3hNJnnOHGFFUGA1F0W5hbG549rX5+cAriv29PoJxH+0p6LVNHXLq4
dALN6JrpWKLeWXpVooNVD+2zeDYG+QEOMKWIu00bpIrzK3+zDc15s3JkIirKvenibiiQ2yAuHA2y
fzMDUpo47GGVKlkEU6X3xbPXuj04GVW3pUX0YDYYVzMvW0z6d6p08Pdke7kMuW+QQUoBU/OkHegc
XW8/tBqSKpeu/24ZecU5extTwAIc/1CA+60nQqfxvInha/uhBHbabsykwirrFStCwm9FMPDwP3Bs
ZSVWmJ8bj9aAYSv839f0FVgcftvltH65+7MbpRJOq+B7AMNZ7SLSSKZaQRe80Bjt7ML1O4JrlhMM
JBx+BBRlxq+enhUtPEa+p/279bdbCk6pKFVQ2+gjjIRXpNYwBcY0I9CR3rzdyadk/PdrUMBD/Qjn
rvAlKd4ri+NaVEXcLntqaf8EL/OqGE/aJISlu31hqfi0NJgH+ujM/msJ2Ee/rid73Ns4qsWYGh8j
rQzhthdMZdUYAGn92bnscjQbTC28tp63JV8P8d2a6cijCR6yymlegdtgjEOn83Xza1dK1ILkVAXB
cfxuH0JgA4h3UHfFdYQN5c4BkDjHmzpF8d84kZSFVfHWd/KhUZo2C41Tpp6wtUeTXdpwN25mj9ob
4O6iSP3L+TMd/UpMrp/P36234pZzMixxUr2RmkuRjBTsqTE8fYGp7ytRuXRYlHxTsSqnld0LU5CA
dkxv/bBqdYniLW96aOl5Rbo8mj3s8UVDm0JurRffNxfwCXpK4gSS5+O3Eu90N1goVqpFnepOopKo
fHo6oGYhjiVYr8gA/IC1Y8KvPVyUUdO6+Y7FRUHx4IfiLZmBl0WLkHnmNzbgJQINOHwaAZ9YSVwj
fm1urRn5YjJD22QhRTIKUc57cQ7LwHnUJ5DBksc4y0IdCzMfsE++jj9G2izV49uFF8P1pe7ikWy2
3TAohXVEJ2wMTwXoY/NXafgIoXyhKDX6aXnSV8HHuSfGyS9N/UTJrAFHXBm9S3ZiKaw8cYtE30zz
+2a8lKX+DSufATbzYY8cf45e1W/PHUa4utzCP9RvgzD8MUmL0rzhXI09EW3zJpen/XdjvBWiqBTj
nPnZJTQjBhTzg/1Of/agFw40gKziPIr4O6Ipr65+gwOwgRdiZazV8VSTb8PNpSCaZXzTn+FoUsT9
H5vcKzw2uZVtppZGhb7gdziINUUcQOm5OUh70ASwtkoKcGTjU6MDsLCuyzUmntFER/bLU8Tc/EhX
A+Q9qml+ZO8j3U+T64VXSY4kHMBI69XtX5cYbk1tq5FL/YkCJ0YbksR210dnhC0HmuElfgd7QNVQ
FhTxJGxeEujvTQq9Vmpo/ToreUP/L1JRWuMq95sdp033g7HUpvXZkJtApapv2CQ9Mg7zGD7fF0ul
tY7+vl0FaXcrHs03TouuGm3TZ4BucDmdiel8KrMu7ottgeadVa3EAdrCWGOdvUyc9RxzwWXjUd07
C9J8QBrB5G6fhWlo/RVWpbDk3f4Rki0gQ8H8xgFKUFw8wXi097WtJcEas2JD8Xw6TSJWlNnNz4B+
ZR/CotdERgKJ4qTpZ+1P4gtMl4/YW5Vi5uwkcQagCk82ivHsjCw9S4vOFPcfZZH5P39YUnypYNcB
J7fRZAxmD8BCOi76QJ2MzyCRUj19cB40fJWcR2occk7Rh3y+H5cE7UJi3f1NNadCQqvORklcWH5B
mPbYDRvs4wPqpypcic5fEBU/f7UzAam+YGgGAKweYPTSKCZnyLNmx6pYEzDW2VZIkSHsWcrJe8NL
PzrdcRM4ZYRLg6/2Mk78JoQ7sJ2yhtCBqRHS5KlT0Wvi0Uq2aot699apv5vH4rydahR+kUylSDEJ
01s2NaWKU3a+CCWywivniPS1sskqPJrJKGvw33lFV8UXzsTHYzsJBs1MCmoF1DxoVFscmZnBKAaS
Rz0y6j06ggtEmiWWd7xpf6kMjtqSHZ6M98lk8J5ZjM5AndX5hIwLJKx55avypTDy4hQEog5qBCz6
0WVGP1WQhtkcW/re6G4uz4v3x2wK9kNE79TE8i7Ip/v4H02OUJ6mvVZv+680GTMCGgCe2Zh5GnpM
v2rEvWq9vKAqu8SPUSf7Z+qn5zv2lIxYh22UxUNYmfTdYM1vMTydtbzQswgQw5w97gVYYQonvi3A
5xO+rbTsgtGmXAXX68OQe9y13un7AiKsLRIz//BKwp9Igahn6owfevue6SjEmMrKVpup029v3YpO
2rHXaoZeIvjUj2Wp4tfukZeig7qYpyEWKr4Otom9jUUbdK0faL/WVEhXt2//GjdXbbPl4HdPxJ3g
56U2u5Ibmh26KHb+ncpUE5w2iS+qZiS0+yUN0EGkks2AEvdc+RhKVtcFL9JtXybnR+vFpQkQkfcv
DmhQczP38I1i4wUu7FvsXif8qWKjZnW3Yv5XXnKZcDUElvBOsk1oxTmuEENy+eIq53q8cXMOsg+2
ZiaeUnxwihBjmuWD6i5d+pFyHXE7UzMDlLiCtN+lMPg0Gt4/neV8RWZsVMRtNoil5Aeh4tnXB7Sn
sj9hzp2Jmv0UxKn8ac3UOGmRQIFnaL+MVEM05PRpa5/1X/lJVpjxd+LfdlXsZ6RuQdUTTuCgE19X
exyy0zIvyEU7MrWtEONVJcedPI84YwROBnmNU8TRK5+KFt0yOD+/2MFQ30zWR03xG6RO7oQggXt/
q/7YrUttQGzm3kS2S7DfvzA46fhPV3mZnFnkok6rkmRyP6JtvasH1LlFQy/SR2njOvHPDeZBPvaG
7jJF7QOYL49q5MWLXuex4pgZFDe7q5cOTll1ClAcd9IsnDcaY4G91gv/pyR68WTsD0IqsPG3sTzp
nzI5mA1YrDWi1XD3R+6ZJyTLw6SSvp/ZXzzYxQ769Ua0fErpu4FhrbvGaYcFuTORDMzvLRNoMz+p
1AJ3xB5ioW/bFZkQyE/lRdxjsSZUVDHZLhUdu7pVkcEGdRn1v7KvxM8jz2zM0HNQwmiEUap4lO6X
r9/cKcjC9ufQ02UcDVRf5ON4nwxQidzgg9gU1ClGSR/hg4UgUz3YQDnReE4mglxWIA0S2dYQFXmv
ls3BwWFNcwBp0Yp1SU8VvvRdlUeSTQnD2VVutD5aa2LX87eL4DGBnzw+qIxcArZ2s5r84FKUXULi
6ce/Mny84xPnYe735ugWlrOMQsHgGQOnUHqxHX3RS6lwS2brZv7wOPWrzpFgHy0uefLLaB8lknBb
OQXYfHtW9QdA3YGX/A8XF4ocUF4psyYfrmLYoU3EZLd7do0E7UwBdfX+hTTlTjVnyXCxHOGMRCZb
nBcgLaTeAODoFxWPPruvL200zGApNQ5lDNnwmURvcTYAydgNNfkIvSkQe4zjMs3cpw3j1F3vnpjk
+m2IN7YK+Y1Uu51bgLb3Vfir2v0Wn6pXqLwdsGiSVSIMbY5IQWXOZchHG6gUQ4/ArcgeeGq1jSNX
2NVTzYYvUMMtqtoPUSo5phBFtS69kz22+gNAVLhyInc4uGc6vjSGZzEV0e6hPCbazDA+GbgQuweP
f15KjY/bkqezNRc8/yCvdHHaDa2dH+SDpew8UHEBXk8hwYui6RAduhvIjnHKMaUu7uw5uwvWOnoj
7KXztjdawqVK2Xi60h+kXqiFQqOKHGzdIKYpj6XCQptginyN4bblYndbTyDXy6dFBy4lN5L7C7fe
FN5TbMN+9DBnz1VeIXqFxFVP6cZK79TJKghJ1XV/0B2VaBMs5AawDw8ee+dlm6nOLrElkIbqV2qR
4BOz5ZOuH/fmsJHtvQnez7KZ4C4eB3qLJzZtCFDpsGPmkyzkDV5T7k9TNmCZbz47o5bB87Vogl/w
N7eL40qo/GK8jkIkVXqJuG2ON/QEOBaFnHdf7IraL6/uCJkL7wXfGPFVa/C5uOY1s/oEZI1nv0Mx
bJ6hcA1zeViJMFNz/wdLqHjL7n6RXW/Th9usHhxaKjjCHg3U14Pul8TN4OsomrTeymcIf/kywXCU
67839Ckc6w50ccyzcymIH3+Yty8Qp/HI2MwwUnBlNoolzLpfHrm+K+oRarUU9HduwvEPxIEhkKLV
IMCJprb1ObE+1PcNV6PigU3VB590+LQ2uYIlbktD5R7l1asXLkKq8shByBp+td9755Fn5Ky9JPCg
iw2Cm398UjHkEOqy4oUadgV7fJyMbrsV63o9qZbATWmisciab1H8qFmJoPxPUsunonzakXXebleq
apjelOHeqKfLcgAhKvF5ColSXs65tyjDwT2EJSm0H5OjSiyrVPstc/AY463kV+rgl/OCmoKY3nkf
63iwzR/BwvlQTlI7F77KnO9lzK6Ve4R5/s4JsZtZ8kNTmLxQ2JMj8yfNIo+ELIBZOa5NuhmT0Wai
InpHEUx905t1eXS8pKGQPG7QN57Z8V2xrZj2h12a6yLm0UkAy1E4/VTusKJICtRgvEJg2Kff9Em1
rn3tiemTu/h/NHFoT9TYRBb+sLn9/yb67xwA5EHLZe1C2s92blwcUCTUn65X5ICHgof5IxdLfsDM
tt16KXohrYBMHHWfk9Q32CQ7f4ylD/llWkCmsuc1IMUtoywmWxGY885YKARI2Ym3FsNmrFQEv/J0
pkQVwsjob+WaovtwwvHdNSGEssJI42pmMJyyuAFRClekS8hEkzOpLdQ2Am8R3U0MPB70NFHWIRF8
66D++7pme0rVGhvpEy30Xc2kXjQ92Sxufva0BhYx2csjZ/IdelQvJsCvOZePG32I/XRfdgZh0HzP
Lc+qQngB5usTUKTk+Oz3oFguO0Lc6dKLcROMQ+0G711OqTWTogXOHU3JODjsAD0SV6loyK7f37op
+HsCF2mH8PI3TeaVHMPn/wSfxYMuoRlZ/NGPH7kpPq+eyvSQnYo/zGqKx1jWe5VnDn7nlxdFUtDE
D1Hn3zJYdnRlvkbFDCD0pP1aQJEBZaSNy0JQhZ3qPmrZjT1CPZf0O/pPYmDkPIlVCYey/aKvMZSI
+NJAF/kiyQEqq11T52kFHI/n/rTuRWYRSKwTQLDOLgt593njPQUjYlqNy7LMCytaIc1yIrtFsciz
ly5+/IWrzFzIha9gPhzL0duXVgBbtslqaEcgGU6TsQUoqLcXtv1zAG2SdHc16EywRFwWnspg37Je
PbNG2UMsRpiif5lPLcgRz0+agKslOFGYGCSg7EVk2haQzn9McJeUzAFbf0ASynLy7fdu2IE+ss1o
vQpXfacLLkdX+cKKg49zn1U7qdG5AxL4u/XiVWrot1A/E/8hmLiLGWkM8XcgWOQt3h8ubsQeL1x+
JpyCiKWjBPGzjFNUFM/2tMTiYmYItbSRhQ27KSZ6oKBjpF8bdZdq7O4uDBEHQvwvk0mo0W6lBEyE
rHARhGOfE31j8K8Vj8nQ5IIOQF+bVi31D4qAr1CLBsSFY5FoQYpJMJvFzb7yy7gIAkyUkFIL7mjh
TJvmFqCG7N+KD/haC0B/74MJgz95AjveK3eJj6sQd/eWBiQbTBY7IIHPJmxZV6e+cLY1S3lkQkVr
gdOLbPNVp4gjnAnIry1ZxfllXqsY6OXFeWKqKmKqIfLRFwNy+ES3M+n4sZ1Ww0mWZ7gAUrFYuOk1
cz2Ql1SsznmHcOHnElXHjZ2cvpJs2DhAc+pIb5O1IjJAIEHOjuCOIBM7wKz144z/R8gfWRiW4XoZ
YEbC/HwIqjXRoIOPDuNWU5kxpnesP1go1TuzZQMkPotDLGfGN3lUykrKDDPtDP0tb8hh5o8YlG1S
nIHg2QVkh9XlMgBP1Swq4jV4Vpp0AfcYM7K0X+pVD2dTW1oCJNv2ay7nsMOJ54hXffiFNl39nOTq
y4Z80qoPMp9DimqW2vBk1pUdSypVrfHyNm1t+WAaNUeCLe8BNo34cOVZmdjEU3upGstUnGLqF/IR
ELtuenBDSNnUQ4qdCsRAP4VD+2TxuKt5VcRE4RWNjSW46WwOb5r97kVnFZ+AMikrBnccZBOJYeV6
8b8GfoOfCbIkCF5cz0K+xOMfvWErLoqvYvMYyvL4xviXq6HyD/ry95qr5zBfdy8dZkEY5ijfmyLd
Tfo6bRt1QFPfU+SGWN6Qic+r4Oic+WDQ8PSc7CncAM7mZE/F2LuHZpk35nQjyAw8Wz6PhZq59QNE
oqNeORXDtKAiuji78mmreGqrcrd67tFnpNSDBWG4aqeqS+Y0QVRu1RItIy39y9KfATLko6aKta/x
xF9JffMYqxqnbhS8IXCAi8jW/Yqoi4IMj1kFeeKatEEoFfDXRY9IV8a+Xcc/3MkEg/MxFj0iipAQ
u7bvYMRyMwB2Q87W+v7WbBaGOuUjOv3sGOAwqtaom5LepSNLLZMMLXrPggiZnG/R4AGzv7DK26S6
9xC6IWPAiTy4kl8923mgtGLFNhKuMa+DGBS8Z42kaT9+8YYucD8A5f/9CZZmf7cW/eqqWeUTJPZz
qtHiRoILSDWwzlzMZcbhgY3jgcN2D50Nq/UKWam3iG0U+5xHvSRLoZ/WJ3HnIfCUDziRWVRuedGo
PGBi414SvTvOVYzN7CwG1qSnJQOvo2ICHZr8YpBtgbIgisd2lw3l+lbjkkF5ZT8CR3qW2tTyjc88
SCwfAzHD0BWdgbjnXlZIfhpp4RoD119iinL5CHWaK7ngQ8q31ACEThDtUjaOC97SVWTHDKUVkUZB
GavuVEnXKRMwifJYhGJgdj8is1guGSNVsRj7cWkhfE1A0A45YlYpYXOJsixR17TBltoIAr/dJ4P+
YAuhjMWGWYuTcnw5is2tZv5HSfdwPCl/gZkxVpMNNA1Cig5FLdBHGmv7SXljkfpQgM1rR7RlcQhx
2tvqzijBngzdsPae1zkpmeSpYfvMWf6djeWtgZofWOFxeWb6cbyfxuvTx1IqslNa3kIwjOqrs7zy
LYv60AV4niIUaDaNistdUk//aYnV9SpW+q9CK94Ro+zaznJWIcVKpkr0BEjQ//5k0Zhp1SzN41P7
TQgInQsLq9UR2fipCsa2n2HAaExKIM6DKft7RWuG9LUBCOSTIfWwsBHzOiWkE1O8JD7EnO1Ms4D9
HkOcgnUix1Q+TYAqb9c0N4MbiONgDrdTocblRIwevTzF0tFcM8b9emy6fzSSljGrqkt5IsXlnH6x
mmGMfDWyDWF5EaXapFVwJNAS7ons73Qv0GJ2HThVrqXpwlnIGTiyj/9k+m3SA7QnR6QG/DjzSZ6H
z2HqjC7Ij5f0uVzoogTKE8VnwoRmrMfrtjzw3YW5un6lTUDCEfBcX6zeLCYVoZdqCmq+xb6aJ2qx
7AM8OpmGKDxCu+y5X9oFRoqGUgLQPELVONZqqfLoObDusmGTmeXbXlkaSpC06OkOHk1J1yOt10rK
rdcuLPCkVhBv43P9x1IqXKrYgq8mBppcfO0OP4MGFfGjNuG54EP8jdPb4dPCI5Orcj3SEjwHu11/
jJGTfqPXdXkNMnnT7EuekAFbwCPO//GQ3oz4lYwe81nudsJI0NeBdEQ1+KYwn/SRSXy9Gsk8UoDt
RCuflgttZOInIbr9jP5vDqcv5Si6VUYjh+x6lA0+EcE8ispuyYQ1vXC3fu/+DmaPikwp31h9v0jW
bMbeZHe10LKnw6MSUqvRKTkm3Z+gxP+llFLF7mPhQ6M0w8j/5yHxhl+YNN40p/W8YH20JZmmahhZ
4NQTwlwxhkCV8so4tUXuammNxIetTq3avKNDSG0dKUaaMvnivB2B4oX9ftjt2YyqxCf5OTcP8y4z
7wPKMOh2YV4rG+Tw9fxO0QPNKdYGEesYDfoP6pYlfqc+Eo525Wl9RPPmk7ERK8uPct8biWUJUpbD
4zJy1VNA180LlDUZBTFtta3xjg2tjN2tUmmF6VFg/PAESYEhIL7HSLf7q5wmJXSiXQoZBE9CPjMg
JjUs+a266mX4S16UWuD5uUWpER/9ezWMakOzIJQVlrENCmv0huW3NOHOGSbT9f19+a13qcjmsGt/
Nbe6APQh6HySZ55SKSZIYvJaH9pGZg6fTY4SWg21uESU73+cI37gezFwUQUhxFfzoM98YkPk8oej
0DtOGgb/Y4VDI1ajE3qn7Hq2iKQcI+igWYP8MEc56Ib5hRe+hYJBm8A0o6hEv4bpH4ibx2G8EFXw
lgQ2iXtJZFOGNxq8Dhj+aPF6sLwyc87PfCG5/xa+fhToOvXPmfrWfCH+VA4T4F3twSdJMSx7z4X+
drPhn4HsIkKQ+iNQXXcn0jC0iCoz6XobE3k6NhprU/wrp+wCEw2df5x6jWHRW8ZZTAFyUCi76nw+
P+wvO7iyIXR+i88s/yMzFUAWT8KhRg1e2CEIjeEhygzCykNRojBBINak0mdaE/CwSBiGJNn2iPwF
eqjEWkXbr1xX2dzPKRqtXgloKG1MeZaZdxJzk+h8resq3D7KlV9z39WXKD6vAdipFR3mLbRqe7a7
iYKjqRh5zU6I92uHc1tzFZvE7xu73++5xCzhZ9m/cRA8Nb+pZrnUvr7smuixdTcLEEKRibXqXenL
fZ9Pl0Fy71KCuIcnQlPpEN1z6t6S0foGEmwj7UwiyJJCJFI2BcW2a7hubp+fQmwxt4sBn/dEVYEa
WfaJJ2Tc0Edr2LYPBZTMB5hQZlAIUH96PKx93Loe4jmTpf+PKX2R/RjD0r4nO/5Zb83ln3WLvDcG
UofYuf8aKL0NLrQvQOwJDJiMNgRIEUGSFSo1GUlM7/DL2vfU758X9fkQBrFMqEOJG58IclGaDsFQ
Gh4tt6E9VhVf+LACK+swsfjrS5EIYBhn5cMKh25c6UHD3Nm8ZYkUo3lbZnVkvRydpg0vnVS2lSgt
9veJaGXbICxSDdY3VScDr+xWcQ2EN1xnjpHjZIGGXdsxL/QcLoan4nFOG/iS5FWtidzEVaEqppzh
++ub3WLm/s/InghY6s/MEdVMMmc+yEPBn3XyxgJgxtu89la0Z9ei8AwArSmxNoYFJF/ooWaUB7xw
8v8N0rUQ2sJPHW5k8x6aBtg8qGjIWwYijjzQrjFwG2LynERX7ARc+3RKV3oXENTLQxoWJE08AhLf
VPyTi8NjPcHl16PSCeI/wDssPtgBmHbGh7xUGCotagnoA90WpukbYrhuz/cP4xkJDRGKlPk2WoDq
yHV8m+UacfBDikH/xkvbxTTkeHQT7lNMG0yP4J+lyumrqbsXEQARKfFqnQMECMmOtcwzyfmVw6qF
LCzuo/xiPeCH4+geF1UrRqhKvLjjIThcuqFKUTDQ5V4Mkm1mNt1ZG8lwysLUN3ody5AyAILWbWZK
Vjps9yLpw+iQZKaAce8tHZCJHkJPHINN2mvN46do1dvcifUEkMaLq3mj44KPHLtx94Rs+2KSWWPL
WAt8BL9xS3oD9/EtrKDHFs7zrW0j93H8m3lGRcPOmPgNBRocXeBTMcOFBF/vkMw2d5S89OtZlmm5
LASjotZzKweq1j7hKmcTGxeykv6T/d1TlZtCsQuRsMSLN8qlLgta1aJvhPJjxSrtvZOAiC9R31SL
GKAJ8Es43epOYTqF/hBMUgKIlf0jPJPLGd7j+lxLR/ODyD59TciYdVCVwQVi/S+PaOL6qw2MAnzU
VkJO7HBvm1C2EMJ7DW7VuNhCnApA7lSDD+I7HX3C5z25KEa6qvg5yMVjlx59FL6sTbfdowcjSVDZ
9Y15gPHOz32ofABKC/wxFF+kDIyc3wUgzyegnxwYKp6nx0I16+Cf27nqNMe90R6TEZaevDnhqnwv
DJPpNXGb6+gQYU1LEnF1XSxiqt1gLzmz2hQ83BsCnt41RRLClizTED1gGlQuEoOg/JqLarNU4B4h
lqNmhZj8quplwQzmFXpAcxZhc7urA5vQluFf8p0ROBhhatlVD8vT0TzYTfp+0rzqT/YnVpqx1NYH
5fv5AoA17kKegvvbIVLCO4Zvk7Qm2au1vFNI0kc2uNftux44LHQna6CbAqs+AR2Aq7t4WPz5Mw9e
zdZZaSQQd7JxCoPt7fN7H+/Po/BnliTKpHghkWf4a2rrSdpJs+V7szKH9RwtJX+WvEPLCmHsTzkj
BNTDftUl8OTWCufwzlLTJWBTJfuoikzheF+dYK2xbVmT4uY3L6T0E9f2gaSfpWBTAklzq/jukRag
QwTsu5eaMR++awqpzV3Kc686lpnUr5cEssk9i6mynm8BFIpsQuneAr7tOVVpfrVySuzwXYlG+B9k
cA/qLjmU7pPtS9yJ3ltoPW5igqKFmj0MsNOgdVXN01qrQA/L9SP28xAQ1dpSI0zoZqgLUxwYtPRm
8FFvbc5D/UNLV2TJtlVXOK+qUFYW5GcVQkWqdVgQBGnYIUVjL+FBqKugUrc9sUPvt9o+yhIJpqWa
krlN+EQApNhUaJkqqKtGHPteTyaghpR5TpyAGLl7luq4CvN/Nc0yY3JwqDWrG5uZCnbzPlmy93Zv
Ec2fGnnmnnt9Dx0C+KOT6y0+h5xL7Zi0NRio6IRoNRwoxdSQRttwsyexkSR8D86FFLjoAMMObfDN
Z5yV3lG8+ctLEAO5GHXuSQSDCFOS9VdfvDLovr1MuW6SFFq7ygqvMRkk4vYCYkzDZTJt+1FXJsl+
hYDhC0fvboZXXlh+nfg3rcatmaCiJrxigL60CPyq0MyqBjjBRclv0UZliSvePRllAS41m/1/dPsm
xTk1MGvKmL/q3UtW6X1C/0pbagYTa78pf34Fn9F/YQ3HPH/T2ZKhxjUmbZY3FuN5+qJ15UIKgysx
8EXbRGpMGtBHkDn9KHLRn2h5qCck1D+R+bJK4aLhBz9Kcie1gdjhygZrKBIloOI+enwBRuo1nMmJ
NSu0VR0oYzmFbqL2XeUeJesp52F9VHu/GPhmC39ymq16x4AM/TlfCAj3UvNEZ0YUCt6WkRnjZIZp
ezUE/Mm8ecBzQRxfS6IrOLDMcx8bERQNOQq7sWkrENAAYsmTDBgBDg4yWIz2YIzJeHvxcMSBm+zr
95Ns0rGwyEuaA77oOMi1YGrv/HSoFIAxVutQNs231K5plH7B/fK874cG6ZS1QN+IUPnl1MH+u+em
wu5nA3s83X7f30TesCOHWpLV6nfjVNrwC4eKXwLsX+p6XJok6kSHbSItqr48Gs3A6CiJqx9XEIvv
Pn49l7+RV+vV01PI4HhYYdrrPwkXsBJHSdFLae1Q0sCPhPxPd1oVRoQg42JxVgdBTxm3m1skh6N+
wCXjAoFia5X6o5ZLTAqxsAPLhm0lIXFdGS0wWidibO2/75ICI0V7Y04T0ue/95QyqY9NiEqMiXgl
Yxsv46dYKwE/t+kJI+0zrWK2OT4ZKNDTBiPqYSciVyobNL0vG4NGdAnRoWR9cBcZyHXpKCtNb+VS
vwkY6dvGeUf16M+OFGICNo5L4xjyfbnm6AIfFkS5eSzxHhxU52YyV0+1r2GIsZrFgNLY2PHbU/Hv
GiLnjeqgth6a2RqATJZcNlZFuzfUhQ3Ljj6+/vx3TtIahpdRNDklwLbt9nuDKDS2jLaG83BWTbVc
69LluQoRJ8oRyg4zRk15WmzInvBwPpF3KvfOwR+obIvlg9Ur9WAhvNY/915t4yVLKozrvg+Y84zs
1ly9QOK1oMehijcVPv7vL6jYiIwlWVVuuSJFEXQ7Q1i9mInYoMYVe/2ztJsd9BsaTZ/uQTLKiHkn
CQuPEsbO5vbqGBNZ2uUWh+HA2lzuAJ+VEAomaDJ7YencX8yw9+chmfi8QE20yQeHqQJsuEZiAOsW
5PNc9KVntl3kKshLBdPNVDGfeGv+5alZxt7hDVGzU52zea3PiAZR5NiVICgnmG1wCL/zwEr+IJXl
vkBfYRr9hZRC0PSby/nktxj6vssQi52xFZrUpwDygfXq60H5+KdT0PBJwXBRjh1ry9gupNsyM9zR
ZaVCmgg5ed3mNGmJgpFcUhF5R9VSPK5hD6qs3K/16WdgRiNZi0t6uodMsaRdWPIc6hOn3kcsuy7D
FJSwIMmpNhFCAT871SnfQXXHIbgWO/3Ubkx+eOM34DneJMDT8Yj+2qdF8rmCKsryVMigoczA9rnG
GXeKIlSC+FZsA5G1TKQhfHHN5ryop3xw9k6MNdV8b1+XhYxSSJqXGqAf4qd9WtIYntx7wQVzhngg
awiGdWAhybTwrj0R0mEx0koW+2oJETlT/9EG2JDTHVL9L4xH9cGvoSpDfMgNJSIYkO7BIx6GVkoZ
L8Mmqm3YsM0nRQ5OQOJL7MD24f5FehU9VwX6IzxULvpZPCwDaKh3nX8fNqw2xPmF9iLqbbswO/d+
5ZhFF7YLwTOu0uc4kOcKsjt2yQx+rw/0iKtCW5etgougWVahmNVKX0u/oguhzuY/ouODu6EFlknL
K1pMssOGn8KBM70Okv/FCDGFgr8Gxrt2LwKctn4yDi5I7Vmd/HtV/Tgbq+I0LbyPTwK2tSwZFd4R
YxdwMcmuJGR/U6I+hZPWolwhmBL15u9Y/WrEmTS34qpfR6SS2nBQb5ZNCAMuANuN9TzHqeEKOhF8
8VM/XmzZ0iKlFTEPJvZiFsAmu5uiqptueCVhaX7OdA6QFe+CceOu3r9m6PmaLx0V7+e7WPXCBFYg
6UZKZe34SHN/QEXSLBhXJQldbRm9qqT+CK7dKylofLxWia/8GDNcKflh6LcaiuDoBv3tbv/gxInY
Jm0LS49ZzL+PW6eOApXo75fR1UmA/+XdVFdgjim0hfIWex5eKmdarn1kVd0DadxT6i7MCQ9FdGiA
mf9Gp1ueq84NVmi63ndLK/hbelkuGOJ9fwCpl1zhTDMfTcQMx6+j2eJByJ+uFeW+0gGzPE32ZsSQ
MISv9YOOIEz8RV/659HH6IfwJvCn51EVdRHY85OlKlNUWSbjKHMnW/5IfB+7feBWL1cqimeQ4DI1
L4+ANg6EUN0SyolbZY+oeIbyrpTw/EjCK/1akr7ZblbdyCsyUII/qwC4jeC9ED7CUMTvanVl7sKH
8RLDRRKVFZqm1F9PGSRwhzg8WcXIiFTSK5aTAiINPsCxfKjqDTX5RcNWBnVfOd6A+qT9TqS96y7Z
Pou9cUVSYl2rmb1RJD5THwXB7oyfK2ioGOhcxUqyVBzjIXh5P6Qyh/+ts8t8e2ddNnl1T71tbl3T
LIaXje0Rd+E39Dh2SvKoXSF3MJ+oeQIIhecrY0CEqrVrPD0CEWPixvmwXPO2aQ3TDP8xqKP44cvm
EdnmUk/3Pjiq09sY8sKTwR46K1MooIEpFgPEzdFF2n5AGXAlC3ftK9EevMDZqMAlWKzxnNTAexR9
O1FRC9O/SFCiRlMkwSdGI2rYvypzN9bop5Vz+eQS54z+Okag2qb4dEDK1NiKmKgCdL6tFOmo8Znp
mtzH3MFt7ZvM79k7FhWOkj3s/dkXKsvoUVmNmMVWiG2tN6k27A6p0I0aNTnQxmaCnm4NrbAkkeyw
lqjqPl2TWpY4r1B9WNVwUYLtpGTSakE1i+kivhRmTZxWiZmOHE3Uo0Fav6PYB4AWMXpE3fOCM5id
uH6oCAn/5ir0Dk41Y9hY3kzmyU709ZKYOgcBINCL6xeYw5T95TG4BAilMaT5d2IHKB9egv3C4HBF
Rh4ImTkXG2HUHvjJ7VNZTvme6ECSa+aexMYOPp00risvs7D3gjGgLEfpdJkLqr4NwzqfKKoFuHuC
JHmtEpyMfsfb6VUceIUaxvefmmj7EoQW4fKLWfqnLGPfElvmX96ZoxMSc/hhtP5PAtKHhz0B+kBX
mZBcMRGZSSpeVtEJ3kqXCwYUEt4nUW7utFKn7cdxxyRPxQUtlDE1GpDI8sPlJpEEDgt4spGvu/Er
EoQI/W+sS7JlwZ6kbLuAB/iOID+sLWfJnjbjMMAQy+a5RHzSOTJUe+eRcw4xDA1ZtQhvrBffFM2P
EeRWdya0AO7UNCPze2hXQzMcW0V/7VTxPfXg/0Nkmbg+IZVwmoGEKUIMK6UlVUzrtBGlVGPJ7W++
u0SRQNXh5GmbDFOIIDzFZR2npOd3L3avcbKe56OIncOsqjDKEi0+dUo5f1BesHGysqSZwYKG6UfY
IuImrjlny+R6Ct649RTOqUXFUuHOAFhJHO6iFqK3bgVHaaDBmisXDCSnNdXyWLG46KsJGZ74JygO
QQkoFXb/I9nLeKrFNYlxyQYJ0398O84z5tMHG7nD/Z0VbglQ7f9mBXQ9LQV5c4onRX3TttrRFDTl
UQHATK6HKWGlTys+YAPJ0YCVJvEY53pU72qRHqCK4XQu/TpajRo3GvAY3RzXLsW+P72oSBXz83Bt
pRUfug6DOZNFitd8tcb7ThOlZ7ha2tmkjfNHDoRv5sYAjXkgdpiLio+6mPJKX6hmOLurY2Hbo5kU
9+8j8gM2wqQ5R1VLlEanGa6FljVXsFCMVnndMenxwX4Xdk4kKN33X5KJCytTYvWUSmf52rplpz6m
qjU7Go7Y5EGXc/yPZ7WBCcNQxRajAxtIw7FChE9otK8dT/lshFGrtuo2Uxr/AcSqJVDqZSc0Rs7B
WaZdCSjZawbu/7rJPyOl5fK9rs1c1FJS9x2pPocj04r5EK770JYTNvgbXAoHE2JqS1WKSAuT0dvQ
NFCkBdEsJBzHGUasBRvnh4xf0eF0yN2tyVj1WVoort35hMlKvdEnCuzNy9aI3rl7zqMI7KulUhvq
DN0AlQU5zs5wIxDk9QDyO9l0mN423Xk8U9dhHG4f5tQQt4v0bJW8nOaKgQ6AQqO9idqqxpEp/S5j
VEYtFQSRg6iPNaZplpmwUiiKwQ0kQVM52j3N0iafBuy3edr7csy7UYt+GzDiQH7AFMF+MPRvh3eW
S60ScQiEeX3NwVgD8Eq38vw38wzkzdmlFd1GMC4bAItKHlIqNgkAzfJiOmtk22fJ5xwxwadaOGv0
rdGKo6oCH6D1oX3b0nRCsI0G4NvaWQVJs6Dpd8cH6dZzks8TJr3H9Du3PYhDKZuvsC0uITkimldt
AOXa8nBvFB01sUunetIpbufCwGR8+UeYQqKLfqXqQIYIRTh4RjhWq8CkOW3/uCKmbJp8Dr1hK5Tr
8i4NKPjWCpi6NpiGIED6/PYOrqSRrtUgAqfsvErW30Y5SRZLUdv3I3U4ZiWx/0oMuhukE1dhqKzD
wvDd064rpFSNkzWh64C/0EQVizr8z8GlE/PcxddSED4M1yqUSwThxQZ2ARrzKnHGGR0BkiFvnwM9
r8orsR2PnDFzWGTXqHeHY/yJcCIkLpD4N3Fem51PGwAKnfG0humPtLkI8GkIvnHHP+RppKEk2gsL
+PgNpiy3S/0AGdMKJdrM2KX+L+u7/JFAMJawfn8WCXwJk7Ht3cru94/H3mm9nhsGlq2curHcTCqA
tOOq0Ju/r0cFmoZbqKzqX0Lbx1c3S2uJH87Vh8zSND1BzyTLTi3sg3a3HkclJjf9GiCaTAEfwj12
+HH8a3ZmuF/llT3xASpopMgBV3mIKtENILoKDw1mm3nywf4m6xzygTP3pe29PwczH38xpHBp8Rfa
kNL/p4b75gNbscI43WGSDIlEwNHmW2wMZYGu1ycEDZwIg/2D9BUNevrHRHo7qJECSgloKKpjHkx1
SmtS1956d/erYJoE8xV0kwcsgCJ+UdvefrayhckgwFV2AtlF+y2M/jLz3vwCURNOUdE8cO08Gnd1
Nf5oBwgcj0tpfMxnO4tpHOtdl2xOKE/8PMXdMqd8Yss8Cz8bfNnThu2elwissvNyXqGuo1xAZ1Ol
fgxZ8hQAsgo8Rd/e64TWlqLXhgt5amHNme9xXl5zBXRfIfma0/jymdbhgOgjYqGjBdMBlkd9N8Ss
JpsLzj6lkU0GpT5ShIMdq1kQCvSCjyrUMCp43K8iklsmqaYXTgoxhcXyVvesr78t47pvqaa/OF+l
KnXdYGLqAbuIBWssFO8hZ2fknAcp2K5djHxGDjwQ/5myQddtq/9v4lzTNTX93+t76gksZrXNdVgP
8gmyrxAIEBL1vc6L9ny8qahJzeGxM7WTbh+nsldN+et7gkcSATgkjxFa6lnhgEOupW/OktYEHdRC
LUwxDvgdmTlHbGy9vWIide2yDz/AXUka+Vqo6mvIxt+U1ZEoGnLB4uFH4zw8C37OF9H9jcVKe48l
bW5qeR12BiEJgz8ITafLK8o2bHA1+Isw5e7Fqv8eokjwXyHC5iF39DOdLyMbiA2k2UUBnTCUFbCE
LY2L1q1CWErl/tG3Fqk/G+Y5OjOOPWtd5GWAz+DIaDDRGow/5kbYoLXBYxcSW7UbN51bAsNozEFd
VrM3g1zFj8lQZrU/+TSrCLXLeU0q1QBsioJ5gHcL2HffQfokXb6lNbLEuf5JDdwNodpv4lnEqf1F
/S7yvaGEQaPRroTDJKVQm7L4r+Fkd28olfmuu5Tkur5aAmej+Iz8v0RyCe6Kzcdc/ps+Hms4zfwd
lrWW29YAItv4XC4o3K/eeqkkCmBg+5r99kKt8XQIIzywvOCNWb7d6QKsvQq9ix77ucJzojazmW3d
0kZR3/4X3/Du8kGM2RrYIiSnHLWm+5zNsVDcT2mhbx6yCdPH7U/hlY8jJ1kdKsr+n+BKsUMnHBWz
L2h03IIaGN7z+ewUFsYhP+wnwyPwLyk++aRX8qUBMEDX3Ud7W0PcnyEJqULJ7fve/kXlNkbT6MBT
FwOOAZ2gsniGWiXQpLG5cS3KloA/qe4OUKOn+joaQlrjgILKvbKPpoeumUmy07d/DThGYcgO1pn1
4F82/rZ06LdshjMe4I6ei4EHeFo4eZgkUkKmiAJ2Q8l7RpcewjKr8fDvER2bHmWBhv8JzCEP/JeR
rqvotpXZsIw78mUIE25iUgNdSX37d3nC+s6VT1OqdGOtMj1x6Oetl8vrBxFR+Z9wOoHM38jwaIQl
fGUU6pC0As8soQXfrKbiJnLEJLSFob/abAn6gkTXcNh764Ljs5ig2Ph599jWAlIJZuOnBDEAAOgR
BBdnejAqUxd0UKR7yWZda1mV1oHHfiebiBhARyOVx2OZUadTjXrv8PcgcDBju3GNUwVk5WBHriHa
mDrw9a+Tb9lBM6GS6sSeYCqY0HMscILOFjiCBHvs03vAI48h84EUKoX1+gWkXbAh0Fx2dGvY471b
AurePa4LqHNX0RZZL7Ktjb71F2kLdx3HzUqyoCBf4saT/La27tOHyae34jkBPJ3SU7ouwBGmzd+E
3Ikx0fwzoNMzHYYdch7P3Ez2TB3YdDPYJgHdws2PEDthQHX8bgyPVtFuuKE/gIcc/QGu6auPyveJ
OgEhP5pMApPHQpP3/OWm3stIQxHVvOKclj8NCeIkdpEQkLKMbEbNJjrFaRqIgc5evUtvxGsApBcO
PgOYn3mm9MFnkmZpnVHIOgzFUtSFeig1DrC4IxrSLc5uv/SYS2RdYPZycJHSm/XARgOQFZSMjSL7
xwGr6lJXNEjWdtK/Dyld/S1Pi9um1DucVii73Bz7oVO+cVEJq64FbQnX1XrQtKKdAC5u+qDIPMd6
GYsRCJo7IZVJXU3x1zL2890bVDL2y7L2xvvA7f5w9WqpVWwHZP2PqrxeezAeAfZbsSgqZnzd5vqS
GIaKxYXhNcnEtKwhw99mS1AIBdX+jwkczhs+xwdBEFScdS/BJe+nwJYGJFHV5Ig/2KqNS1ywIDid
YOBkqZ43VgT9cfpbQjsP4IUZcCbfhGCzbZ2ZtVp92FqPr5XeSA4FInbX+JQ+Wc2JBjIiTz2nOJe/
jCTrCzK845pqLOYNMjBOXnaiJbf8EtAHc4JqJ4TmsAfpz79n6+qDla0PSgRV7NMUlm69eHNZTVEA
R3Ra6Jy8RyYv4OQ5R5ipiHX3dLrlWy6zkhf5q//zW2SCWEDlgb29eDJAPZYIfEiXJeDd/5qKdDfC
PBaKXHBcdkIlZts1OTDSKdwojSFLYFG3zET7jMmC+ekVC8g0u31hbanwZgkgh2jzlSoZVk08z13U
RS9LNt3pKcSkOcRzhfuzkE1tAjJgGGP3reaaiSwjge2Srqop4opRLr31U0saSODtJvxIpCfNYCrd
tHfMmZOW7fMSLDQrwYbAoiQBo21pYRQmvBnE/8qEo8LtuEzndgQxP9mIj9fNMK4X6viWIbo//F4D
uMVzWH6s51la5lZaju3K1H8mYseT0FQiV6vHUuoL0Tg900QSNdIY/sYmUfsxyZBHiBVWRHAZOtqq
VWSjJlWqLonx3KTzzWsH59UxsspBDLFSlKUapsegOXyuVWsRHqwo7BEjPPKL/rhR79e2TO1t1j3n
j8t9MN+nS+6/heVxQVLPb1++9s4myx0rtCBflOgylaSP/ksVmaz5wD3oIWrCHeM0eTTmBwzy1QO4
79aZZFb1DdiOx18T46/X18r2mpBZaV5zOrQvTyuTPHKkQiQe5vxb7RMqduarthGhpCXEd1aRXZPS
chMwN6uJh1FHuENKhUAHsh70ePLZsYEXFZOd4EaNCESg/gDEU/pk316ZMQ+PfiHdbD6zJhm2TRrv
087bRWrsNU2yHlKRCjCtVsabROaU23SWqFQfe0E72ajFnbtW3BifZJoLAywfyM2T6GyljdnaBvo/
19Q3wDonwZFmWXatdCFapUPMuaWucM4GlO/mC5huxJA4jn+vzRM2l3yfxO54fJph8sHUXeo94UUu
iZHegTKs8R0jz8Wc85/N1DOeLquXeClry4NQ6z+UKQ47yNGNkEzA2YI2q9E+p+JMUjyMucq0t7We
TPPimUkMy1Lfm6tYW5lK+hddruS60YuQhEFOwjZ59+IVHb7hIJEPmGMFPZlaU9q/xTXL/B/swlD0
G9Yy+Wn/tcxMLJpn1GexJNK9bfLPgA8hw3m1gGF10EtnzboG3mfTwCDdkLTM6jaBqUamL3HLb5s2
7e6Bw40Oku/4tdnMMUSUReOKNPAHdgCqW3A/GvZA62OTmVeJXYr5n2QTTvN8ZUGITF99pYzWbmug
GTvDZv3Meir/f2LsH6Xm7AcVc5CpgB4NTU782gBZJjkh9mkKtV/zsFZV7rtZt5jVNOB9L/6DIs6Z
QL+TssGKwes0Konju2wk68WEr3VwhdqNzyZpqCNpGuvr3wgM2avfu6A52SMlmyUV/CPoLeLn87Az
1Vsn7xl7FvYIDqHpsUWOuVA+9pi1w4w+25sSWAA1LmyBonbfAcFP4bucGVDENXldOoYyq1Xl4o5W
vcy+tg1fJInK/+GtwiPX/5XakrHt2v6TOP5klLf/I+uoKch+taTCj2r76tRzFxvJEdP/1awxl6hw
xjLHc56cYPxpeTlfKMpZysxlTPLpDGPO5JgbSnRzzHlqjcL+nkhOBJy6oQxByQ5xyaMUU5L9mHuM
CtFghCVq0CLUSDXIbjx7QVVTCLprPsEKG3Zy+yxWi2Yeaslgdm6zB1/UF5C+H3BTal/wbktEkYIY
HGvfdRpMFBED45P0YgRtnwmfN2un9z+DHSQNpwuuYyJcXZFUYk1ZqJYbDT+ssrR4BHtLOyy/khK2
8/C4woNzOksFX56LBquEoXQUPAHSYgb0Hek5f60L/biBk3Cp+SOGUtStb+r009QqGEH5Pd+h87N2
n8nnceAi2308yWwiQIWjrtPsq2zovVsvL5VH/P2QMbvSnI5wAwDKbFMqTgRH350xOoTq7NTNMOGo
z6oplx9YgiL51vqe/Hy0BVjW0UtMbyj4VwGZD0LxZTzV20NfPnJDphHeXf92iS978NifMV/liO6r
6+T3b/d2q/1sb/TlC82iYAWV4prRrTMExFuoiHGsGE4ZBZIYYbPViH1XweVoNMoOYKD8VXrIGGXM
DLFrGehG5r3AYSUEvO1NJxxqh/YKy1OcTXs02ULyMhMvz0qBF6s3hBZPSWSlC5uPk16Gn9EbWC8s
wp7amAMllINL95IW5f8fHWjLd3IFf/rCj06/nq4jccAigV10ykDlEZlHW27GtBMIr9RB8qVq6qfQ
5G02ikjtrdzOpGQBLcNP4KkGstyTPTPRcil7tIbg/KvGck6OKw0ByqBb/LmY6hE884kcW2WT2SHt
dBtXqq6O73EiMFJYig/G+zDKcW2Sh8ZzIaAvZ3aVuz6aHZPs96pFK7B9Uj8LfOPwYjj1vaylxIcd
c188LDym9eOEjd0Ow76fOpQguRY393lzA3pKWfJ3ORnD5XCwMQDZTxzLAV9AtiR6yk87ODT4RvBu
bDuRpQk3B8m0TmZQslmIeRA237ybKdfh/pdssLXJu6psGd4Mh4piPuxCMPaaN+8C/CYQ77Aw+wWD
wW7oMXAGUiW7YNN4hoAxxEW5/0N/1skNoUrrvTn8P+a+WzVdTYoRDu18ZDXXReKOF7HGEt25LrGZ
Ehp6WV8hcQA3VhQ5WmgbWHVStLoe+KMM79cbnjRHDehx7cePrHKAFHZVyCs04b+QwCkhnVvmwjtu
6K0BOfK7CcE3jpO5CcLQiAzDzJ4tJcdcFgVoxMSTtYMP46RhztPz4SkpaSj3KmrdWEc+OXYsovwP
6UnbOaqi347pI+fsDyApe8t1XN6VHG+HTg6ZTQnbswdq7T/HlReUbKUr7+XEn52fE7VexU4Hymd8
uwxfafkIcFQyyr93cv4LiqgortqfZtjkPtddSzqdTguLn3ycM3QyluqbijZpAkui7vh0LTNbqAJr
wLG9YHLYtYemVqFRnRlII8qxPixFEpFt2l5SqRhivao+Gove1fVAKzASFFFaQuAhKwa5wRwejw3u
qEYlAnSvTgkGcw76p0J0fWFk1sewJS6SzybPoqGskkGCvB89gwvJWUnTJrBCN69uTw0ddn7v01hv
Xi+yO8ZhYSpwETHtxIMtPRWsL8M+hRhzSWtlG5VkpVrbScCm6bd5wnZ1p3n8O12QK3XeCpU5VetQ
qKbVuFn1ZVTZWtISy9BfzRWBGHp4V0ZL3CYaGrnqn1ieLe8XjThETbcQy7/vaocH/17cE3euFtDg
akSahWBLcuG74RkTS1EgVfN+fwaogEaLocgkQASVPeJDyjwty2vN/TgAdenu0FBLl6iw4uwZkXzl
kRgCCHwB48UBWIJbpRUoFd34LgwiMRfdr8QXjMRHhD8UUfH3Fn6OwqTBOkv+1lBWrNBT8lyZo9Gh
GmhUTTXSMowCI7+ffCTV+eLj8JeZVYndlQJmHqTDgfHN9Q8FXmUpITe5UfvV3U6ihDEA5yN0NBde
b6MIZmfvff6Hs/bTtf0ZmvxAz7obQL2S2YBHGaQcJO3UjbdyxcNpylWWB6niHrGxYoSa5q34G7Z7
JKFHRuSGSQ/k7U2y9J/i2XyFzjrawA7CCbbgVTHyIEpYdcJBb1MEnbXBcK0V38XazaGXGe6GU3kh
3uoDvSe6zbAVcIyUu0pEmsDjEKHnEgvp9JzA7TxvylqPM4w/cIGhYYmTFs0uvMW5IYQqG9hYQlrw
+m633PTXNyBlmP9ioN5MNxPfSMqWUcV9CdMkTB0V9bW7bCD2VBmIxFGcHdE21Lsd0bG/lB3lhbZo
lcv3AUtJLxpC6/2RMq/dHEobUPrXIEMrTtDwSEmCL7tgoz7W2s1eXpQhvlKpkyI4YwlOPBYT6HQT
bB7ptFuP9vgtLTVhyhKCS7U7qGjilUhFw1HPVdRgyeyOZXz7USm29vB8IZUduLr7ICCA/0eV5MyO
zs2jX2BcqVNREBDuWTNqjRJyA76deQMn0/4qzQCdKTSNlOhen7FxZNQEDS1pX9dgBGS76KZ4iyoM
RuKMaHWDmnxbwQmaMwqh2Ar9IoGolMlNi4reoiR92CxAVX/mgM1BPkiuZ5oHBBSEripi+kei89xk
pWRwLwTkO883u4zs/Z9Pwop18olHocPFGsX8GvLpP8z/3KNtbyviPhmKwLUnW32nmyJUtX1M0a1S
nf1w3kfiSddQ5491MP60CGRwDBiPj0FAcgRnW+R6ihb4KXAkZ/bPEH39zFDoYpFefdEAbEPD9e8d
5lMyMLWAzU2dqkRsX9O1tKzCaRBQ1zdz0fjtq3VzRik/sLJOwPQoE233mB9IzkTGWdrfEU5RxEIE
TVfi0V/t83vTRBRqLwR0SwNOeqCGWL8oWcG4+uihlQqVddNxWxxKdmNpjWulUqw1gc7izrnAkM8o
J+3kwUQbLNqeO+e+2GSQMRavRviTeM06LcQkh+mRXW0Xf9Nkzh3Om72hWEhvvKf/jhs30yPGqw9l
LuEQfpUBnW9v4Rvi/YJSyWg7yFOHOsf3x1SkWF9KmIb2slZaWCy82mDT+hfOIADj0bMh8RGOFBCH
eDspe4sF88h2WZ+ZfF2Lqh1CH4p89wLFbBwPeQqFZuumc2UWqor/MuuvbBtYpXxohs8IrwbulMVD
/GjwAco67J1mqaBrLB5l13wgIZXjEOuq0bL9r2WaeRo3aG25ETAY9Ssutm9/jZw53Kq1bFXYNUy2
DCJ8QmXGyQcF1/IobDP76eDa4+B7o3hcVW5jDz81Osq+TtpwOgh8FkwQqXglfn3c+kCjY6jgoSL6
zgI8JKf9wQU0875sYxvDp2lRzalCy5WF/Vl4ecWa8FdsqAc4V5ocaSxnAya1d9EeIobkGBc81B0F
nVrckLdWhMAEfpAHU+IKSu5NK/IbnUMFaD9q9HAiy/9/y0Kp+ktuG6GPG2DdGtBXoG5cFmNkC+dL
u3W4o+Uuh+P7GK3vyAoemgAmqrKTuvSx7xSIzbzOMxGXVI7aXM0nhb52kr+oyGVez1EppGHyBi1q
kKAeg7J1XPkkz3hlNtxFdzJYfnulIJXD9nS07idmnt1g1doDUmNq9l7v86NLl+btl/iPT88aTP3h
qo+Vqwnn9i3KRfR4Ac9InM5BPh9oCXm84dHnZ8JU7sTe6MZutabOaVjNuBl8xwBUlJ7FKxzkuc1T
SnTm40L3QynI5NTqGAymo4CrtjCintKeWP5uefhZAlUELLi9TVn5fM6fVJSj6ihKcKPRS1mALnwR
pcq+mD6jX9WfkNn8tpnwNIwHpRL4D9mWJ4Q28xpcCOn+ugXdwU7C/4D99BXBZEJuoFaTISpURG0u
pYWVdOWt8pHvJsUepQqj2BvMYZUmXtm7HahDNP1cN+xNZvdMq+0PKl3PpKJk3aYWkj5Wn7xhn0vU
ADdTbTLSN6jc/HENeuIUhctEdLF0ueign5wGcvYVGr9cY0RpzKFaYywjODaIsIFs+qH3Hd3v16Tq
IMuR8ryqHiLga+wC2VXilfwChAP5icagGRWbI8Y3z6Nq0CcSiPmVbz4oYIhjPQEKTCPX/Yg/sffm
swZoM1ho++CCqycJsEzcZowF41Vvo5nGjNrYZ93yCVTJP2afg2FU7bldosoiN/FDy3JpC4+tvwN0
nLVC+JahpzYw1OJaTyetzmWGFSoAuKkkC8NGh8zslD5eypkzVgYgIzb5K7SLFfzHvTmBb8TvDUAW
SHo0tiP+QtHrDg/LoeW0B0nunn4oJDkpHAt8S3Mz5hliS8ifeg5RLCH9NJUyIfJT66sGeLPY9eKk
+qGS79dwyQnwMudk27SYc0HXBtV5K2KWIO58p7qlLkLptS2IRuu47dK+XmT0uGiLuZnvEZ9o2KRD
0/hwqEyduZY8MegeAMcxyJYQ+XN0Frsg83ZJHaoUQPC9kB+lNXeZsovPDjiEUBrf4XnIcr4sUvSc
IG83dS7PRDrDk0PQs980gRWumYA1MSZs0tCGOFA+GBe0aZkolSbstZmvod1DOkuxKHiQnkSUzPtU
wQGI2/Sf5EY+GOZo9YUw0ab1kHlZLkJnisY/klb4zBvJTiSpKatLA09qXXfXU2GBfWISo+RyX7/k
SxQpB5hkuXxYE5a2AcHt4/Y7OGXWYQXpaklSWtIsJ024in42+w7kp0caYQVL2M3oPzOjtVjLoxvB
rzlnnFWYZTrfMa3aLcvJmbwBSGVRugcs6Bia1XiJpqRAIMjUI0MUnAdxys80lqu5xAptRx3Y9Zqq
SgnCsXr6NJohIcmntZJm+/sZjPd+jSTM7dd23vDlk5vuUwk/WTIrak8KqXT7fP9BYpdPqoPn4XHe
epP9zjnyD20bL4WgjWiHY96QsoZGqZuGxmjyevAW8+mlhz/DE2SmTqQIZ88B69Ww027BlkXxX+Z0
cGJFOfwBsCiuaWXp4zYPBQ+LrkYqJrhp389heAAWNUbmAVJUA199f0PxlFvlP0K9oZeukExZtN9B
oDResORg5Vru75iF8hBEUM++zH0RuEDt+wCg1PC1F/PfS/Rr8P9Rz1dtGvPD628ofQwy/KoqFdpK
kkL/sNHss0+0N3hsXM2i1Sp0ZW+yugA22C0xTaRNbmSb8AkIv9TJUQEYB0DkSIGlhzBRvu9sHvjJ
RVfxl3OxzgWudTCuKc7Y54VAzRan7F4lbHFxFshBbKSZrf3Td3PlCE7Vl/33ue492e8ifwbn2xIQ
FJpiBNq3gu06uPfTm01z/4HQL6fqeMpC2e1n4PkDuUoDj5piBFhsnSFsZVYdk3/1zSf0lJgMl2jW
VzmHTJ9qS7mB8ufhInb6E3azLcQOdGAo0opevCpidvHZ82/E+HxnlcayoHJ3t6hWkV48l042xuQb
AGLGC4viwGdsvmExbg10m1a2zAxpEksEt+1XRtdFa+x2Qt/u4zZdS8SRuTigRr+LrcMKqSmqKgse
j/yK8HIzXba02POMXa2Obq3pBG4xPWgyYWGSCuEjOmSwyeXJkmJiTtY0X7gogOg5dXY3ma720cse
++0DmCS6tkdPqDOC1VcLWMYcE8cwAAVpult62YXSaKRktBe5FMnuprv3NdLRwP3rVPpf9lC7r3Me
82ttvhiqBsFVOOQsgmSnnneSKQJ2oDzsWLuceMXjYioQPAe/QCIFkp6zaZhDOGDJJzZe7RCmsNDB
77w/xxORoBXzlJIiwMDEP+Sz+nL9L1W+mNcbVFLY0d+fD1MFTYRhB99gCesxTtAHFaFJZCBgQvzF
p2E9vnm/7DJJRLzqjWcToln6ORXjOeizVR/4ezjUJKDHLP6GW1GPhlvbFDM0b+NY/kCz4SzqoGEC
qoWYXilwTC36XoAe4XGjaNdolnwgqSLn98wRs0akJ9HjRjhnTvlYgVODKpkELu81tfOGWPRH4t6y
dyMcSliPSE9T0ef6PIVruQWkZlbFCL6DEjuUq/mZJUAFf3j0k65iPfPR+W+unbOcklt2n0u+j/gi
J8uAFfQMBr58ak+1r4HDlVh1LQZa0XlUU0iOCO2EiNJ5HLp7bPQ3Ps3O5UwVJjldiYf8yuTKYxDK
bzytZSz2yGXdGLLe66clG/kvq91nC4TymmbSLjmcFJAe+Q79sszxwRo8iKbBo4DTT+vQng2adokY
+TdA0s/goc4dZ+4qQI1BVee3wNYjJUztjXTBfT6m+JyywVcBlWxWSzHaFLyDALFet9hyfRtG/frp
6FScE7L5scYLw5uQHkGaMlvW1gZ3DeyPFmp97b5t+4Ffl/AqrrS1Xz5uhgHuKWUBE5eVRG7PyQAY
H9J+xOiahPI4Nn96yO09Jh2u8XS8Hznxw9tOdO9PLf8UoUBkoTV4/MMPwCPO3fwNr5LeF6KC8xhp
vjI3LYT1juCUfgA7DsmF8cE6BXCZSOkoP5VaDh+54W2SsUTb1m4vcuk1npK0+NOgIasaVuP8SJi3
TSjRrbir5JdYa8s+4n9HN9mitKCatc4u3dPwD4htPBVxKTNfTBkV2ywDPH9VDYXxvOiVpetkXM4W
n/zryWPOaRXYfHhP/IbjHjZQOICtaKwXwj8vVZD8HpvB01iYjnjunQ24bGpPXknb2KTfk06GAw29
8VrtiNqUcAEvGBXjCubCwGmHdzaj0XPp+wYGXjSHdCb2uANGakns4L+QXymUPc9BGrEJjeeF17GA
UBsBvMLJbxE3x1gAuYA2sg+xXVFbOHzedK1GsbkpGL6xLvsqv6oWGdhhtevGm3KQ19XNeGQD0bHc
SykE7/cVRS7LB1+AXwghqA8dMtGCkM3Lfw/JI1nrBHpSc1y0M24Bsk+8K08PXWDXYVsV6+3dXMaJ
gSb5jaT5ApMBUtUhwtxqfst53TPjPiq4j8dJSSCKs0pIOgZTrTr/0yc0r0WfgSF4mXiOzYUDoKdw
uX/16ZvUjzxXpMV/wIWFVfPmjNUbOz7PNHteJrkLaldspewMSDHd44uIiBfdnKAqR8qkSiklknNI
UbnTUpQqmPbqdEZCP6wnJlWN2b4CkdR5YHToe5zo1kBM5yLeLe0bFDa81Gq5kkVSU4WD5o7YKcqL
jI7/gQDGxA2FudFpHDxNGiqm/V2Fp7FJuendULYpExPrsUEgnlUZl6vh77PkBdN8J1Pky+uWnWMr
aWtg64cxg09kCMab8pPsCoV40ma5lbunjPi1d68Ef/iyebWpgUdQA7OHZf9rPqnarVhpKFsx6mBb
NfterVQnmVZ19rcwUwAZzkhc0IxYoKK/HJO259qCkXFszLhRNNYH/jO4tU0r+hIO+duFLCA7NV11
mFugffe/6u7IiI8GfbZsf2nCXcuqfybOrjeJgp1Akn7rWyY5j8wtKBMywW6l1TrOkJ+Hca2UycRe
OcthG7IeyreC4bgyE3G/eZOWNEetitWUJ2Kzax0edkdSjCdACydkTz/fcVryBVAC7KOVe5RncfjP
Rnt9NCdhiS5fGo3MPjvYhRuerTqxd0CXhsp+xDadoD+Mxwl0K17+B9Q2+bmQoNMZhh9RNHhCuh9r
CW9/cBQyZN7QnGilXnN3E8de3Lupja8UMrq92XQkwxjHQy+mZuPYHVtTsvAZF3+Glblc7M7IHAl8
x7Ms4AiPV32x61zgRGDaLDtXCneem49U/ag66q7503tsh45/Jp93Ap8IJiyc1eUgvlP7XaMop7n9
K7+lNyU1k/6vX2yDmlbeRlZo/4WT9Kt8GEacB6SK6Veo4T2loxP9OLegmhj+d4B1MTHYC0ALVc9V
vTOkliD6+P4IIs6PfSgZN9Lti4fhGBMx+ndYNNzjVk3ASermzJNrlG6XjPCUC+nDUsv9tgbfULBA
dHsenFVtbJbWOpcWlHqTqB9UnlKYCL7//fXW58S7z+E0+LJ8qKY4LKuqjbl59T3384b3MEfEIDmm
2Aqg5XJOnzkJS6TaWxZ8nP8qLlZ53LP/vZsjLQJMnDysTf4HtRqm+p8RzmuAFUmItS/yec0rYmDu
cMHelWv0oOYfBxGB486xOXaDP6fwJgk+WoghfkD5ztWlwcmnD2qJSsNGrQI8KA4atVTsUUEavnfQ
Av24xbhfktLxtpbpJrGjL81e4MBfJ7Fv8MStqMOQWudrr1fd9J7tLW5bwbBTBGiJi2k+3xT7N2Zo
etJ/l9aCfFzioqSV4S3BpETrKrdu47ehnc0FZyrQw4dDZoHnzEH94qR0IYkY+w+KbOc8pkQjkagZ
pvuZ33h+QMvZ/rLY0PkXwPnQm0VoxKqmq61K14fjWE30hVR5J44dDwdxGD80xmK2bZ2i+Ir/9uZF
kSUE9d54xmb4SSdJZwOYIILKRM8GEZYvw1zxFBG0oWA+Yu9SIinvxtre3gNfXqz5BVmbreRFMFbT
m5ssCT/HnAafwCaQ2LAtw3hGYGBjKY8bG/vtAnp7xVDizrkcZB3vL078CrAsgim+LxHePUefnzwh
UDziQH1FuSdYGNpjeK7DnDHa8AZ7e/oQv6e/1DSLbHSNw5AgUYitsZ6+smaaxqBuInlTUJEVykI2
TuCVrVJ/9Uxed+zAEL9tv+B92fjLXJmxPyoiiieo159Vm3EYSUrIgY8QYgCp4whZtR8zgT5/DqsG
26z3t1h+7/ooa6DdD0IJqzabQt91mhBhlNtvAbrAx5AgIPTN3cqpN2sbN3ODM6OBFZa58CxHYYUS
3gszsqJ0KOjstwvJPlR/isOJ+n87434I6dU5HRditSFJ2LyNXB5D9sc6PaKHc5AqYeqAsmuQNJNh
LQXftGgYl1fPUlheRpxk2HEl+Aq4awjSWjmaqcdB9uwu0PHjJAdqmXW2UvWkgrsDlK6BZ0UEJlzS
G33wXgr3U6zoFtOv39yJAInyQtS2szsojCPtpt6zshvRGNvYloAfyiU4r+GqO/i9x1Vq7bB77Cuj
Os/crczQcJnGj7/kQV8lA8BYBEQMK/7y/F9oox5QKKjHXj12CepMGbbD00uYRXsIdY3hDPjzHkD9
Mqg56lGbw8o0QSJ5enu69Q7XRcX19rsPUG0TB98DOhA+K8GOMfAFwVdGtx7W8MzZ0slqgJT6d/ho
Kv2nbnIAyYnpCMPsritICO5jfU5xBqcnU4FdXjEa7q85BrBb7VkRUSikE4elx9F46xPAIsF9XdpT
tXH3eNW2krlKkubx55Tp2bjx9VqUcuUM5XZjhOUzefn6e65r7LNzCvRwJVH60cSganXIbbBPRB9z
P5UV5XvWLn9SP5mKOtlCnCdZhgo5tYKcuXSamelAySkQBfzA5F0oUqQmfqtTpYYcOYEjBD8oolco
hQq1u/IUzgGQJX4FPN5YP3wUsn/2YFncb1k9taYhLmY/EqASApFZxqcS8vDe7u2dT7Ui8mWB1VWP
hZvaL569Wh552HkhXMgIc0IGwDLLhcyJ9D+dWHIiIQJkuCMu+tVHMJMrHhCp7+iuRo5ZdSYfAazs
jnEocXCAGIlmkVm/D9Yp51boVhbgTTQy0cqZG82khLrkX6XnLuB5BEbkvnt6WW5mxEUZCvav+WM7
i2lxmhCt26oDSYfREZvkutZvqhAWyMcuh6kTGOEvQ3yAg2bGHUlkJHkcAJz8QDwHwON8qvXIKnbz
XX9zWONysP6s2pvCs63eDT/WreaMuQgV3FuX+pq54B/HEfDw0qmWdjLRvRJFxet4QaSwrGYA5QnM
ELtUbRXXOnwDDzpfetdmLQmxMB8hyDkLtjwlIAFlgrMb32Qz8wVTzH2Z0Zoqkb6DCsi/Spdgu5BO
dDtol54GU/EuOm16Fdi85c/B+khvLtvGaw2K2vrOjBRaQgnYX1BMP+mAr+cyzQ/Xi/XPA0DAx5xt
2WX/2B/8HqFX7g8LUm8W0Vtus2MG1FXfzd6sT2a1de6vQ5E3vP4oWfa7+IXK7qaQnFP2YpP8Rgpi
hqOLb0tmyZEwqT5eK/hWrN0mIh0gOUOJGWa2w+QrXEm+cd9biMx38qUaKrtDhKgjTRdzxydPhehf
FZQ0n4QIHVTCcA9yUDaJjNXDBIEH9J/otqVKhHIm5eQx9o8uIrPQdYhSIYksTT4xoeLKv6hSD9hW
Ao4YB9qiOmmy0sjhxu12OhmwTcadD5MUYkU/KVwnjE7n5L3QkLCMcCd8i2VrCyFgmmtNMsgt562c
BKgnySMEQr8LcnJnEEN3wUZc9L21oYmZr2ycEFGiGGvDnIdOTTJYnyiWhjompQQN7/09hTS12GkJ
ohG16lfNyNQfNcowFcaDw4q5Iz5jx06zDF0vkCJ1BlGdjj9etnhV04Mte+PXrrBwDiEu8DG9cqzZ
Fe8cx32PpXmAKH0WpCvyOa7fNsnclQMk+LiTp7+QyBlAGpc74J49iQ5ey+Oly3NEVeH2FOKzVzJo
FyUKSF5pPbLWtYtrPjyIywulJXNCOO1/EFAcQhJ5BBkIOEXUxIDCbgnuScGHv8LNsjQiF4aLb+lH
WphAJtyaud9YEImnnWQx2aBnFjB//Ss8DoviD+JnLCdsVIu+DygCXBw0P/hyUQtg7MdlM3AFt9+G
Lole+mju6kCInqeupYQvfako3WbP2alG3zf4aqH80Me3W9Sv8tAHnNxLEfw8TCA5tXMpcAG7hOCy
9grTSQoh9eGrCGHbGfeivEqt000rjPZFxC+MAU+6DCfHKJz7YeRNr26hJ7i2BMrsODm5PrRBsaTn
OUZa7xHedgI1Yvr2zFzDrR/Zs5hrcTGCTl8yP94Kpx/JJd7Ix6VupJ0/g6r5mrLVFvq+41VgHjnW
TPjg+bhb0FcfrBaaliA8iN0h/3FnpJSEtO2nSRXzHKCNle21gUN6JWSEZymOwt9/uANI6WoE37yT
H4rTiVA7B1YWMb9pOhbNGOMVFeq2CGlXIYwF3KB7FDXXCVUbStMCvAMeJ59FTTTAHNN2mbNl5/6Y
CH25DDWvbxZ58tsZEyhCtKBh688+S06obhhej/b93OF8dXIXxCpTd+/OeHDsGw61ujBmOk5tEc85
0UqpuTWiYMzow+nYJWUlCIk3KAgumNQc6tDYDxQpE2VieZHa2KULjGjN3+8hfnXnaaycrEqNas5F
RQoSxsNnEnc84TmmI+MmQ0rHUdCP4Z+alsgcuWLsvXK1VBcKSSnWnfX6ek3qNDi/LiHuwtmgpWlA
qzQOxBJJZyWjHPAbeDUIXQO9+5xDQbqvnKI+a+JIazQ4wOWY5w/FuVngbbs6RhtYw+yFG0KAFg8G
/8JlyAJLYMlgxDhtMGcugSGirQFA64MH2v6Gbya+JpmlX/ebvSCIaSRq9feFT8KHpG1pLTnmDMQk
E/EbM/t2XMVv14QhkIbObesNQ2sA+N8J4J+CqfrF0N+O+ypStJIvEU3ZrnaaokikkAE5BAXD8vTD
D9yeZtQv/MeqOO0Po5I/Csr0U0V6rAFkngJ5ideRtqKO+rvwHK5dBTER9Vhdt5QkwftBIsgZUj/q
iCMfPsYT1AmazjjxP3GYyLB79oS8uDL5/Yzw7R+Nn0bFoTxL/KhBmNp+PBA1LXruiMB+z2CPJmFF
Zxsa440kx0rRac6o8way+7CxUiyQbdW98op6f4ougi66OYF7d5+lbe/ePDHiqDuJYWuLJXIGAatk
oLWHwDq87s15Dd1NHmNj0KqKOU0Y3m6qliPP7Jn96zGpt+BiMa8hqp1HnnoePd9DGYxF7UKeyv0x
/4wfSKWwlGwBFI34KgZbD2fWVAg9XXv8bpCQ/CZZ0vU6WGq4G3OsMThR3g5dg5hfelHpi4oeIXaS
hliFpQdfe94+Lcb6Qu1jfnqsUTy2iv8jWYUARW+7VFha8do+khnbKdYQGFvtgLWBmr8m/32RlfMv
611cdT5AHVqIbGFtxGQ3VkxT+aBOoNJXdWsUG0AXP2xrEerJjyxBCHJXMTAH0nKPEWBpx5wlQwv9
PdF5/cKdRxxneDqJM3nCBeh3V9/L9c2N4tjR6vJaDSb0EkAOkURlGTWDpO2OFDXpJeCGNa3USehi
6Ctc26wCRGP1WlmmdyIcQH/KYj+idITRcHXypyoPThpzn1MQDRv3KVyz0bGiELvG9C/+pgWwfI6m
1o5ir8MV+zSM4QmLe82fsbUfmKr1vPUEzDiD8Wfri/S0RUYeyJ9nj02kG6zL2sQgGcw1wbcqsaK5
q6EP1uEen2+ddpuP8jQFcORRp2eW1QTnyou5nHn0zU22QicEgLTTiyv8PS4f+WNXD/SFdoM2/Rdj
Jzuf+jU7H52PdJzA2aNx4C/7zExhqDH5KqZLS2bzHfLxt3MbsBY+pfhkjQ0YdYg6tDZQnl+FOGCt
PFL1HLdHYydkmFnMKE4NDpDVsWOcTExJ9VpYHpvBXjbX/5VPjM3ViE2V7Hfpaw48EdkSjeyllWJD
wbR6TMfxAgcDagm89QW1a8M/lG7tUK3dGzSkCURw4wgkSfZ83p+ytEDRTiRweGFVo8fluvv4xFt5
xuiyrwomsLuD8228vt1cLIL+QEiFfBST25A9vcSHiHnv0TeoWs87p6pNXii8DndQmmm43ZONYb4a
7t8nLoBngCYagaYtx5iZ+bkri2sXdVXp2XWYzM9TH80QsQ9slDXcpasHCNkyN3nr54grTShhIRJL
oY1vEy+XkzLY4N1wqn0TuvAameBg4k6AF7BIbgT3v4JZjZevNMhSlhvrf0q9c667TBgTHfAgiKsw
pfscN2kNmMQ6ecT5oWgNwYfAlnzZMN7yWFYkQCOm7Aobk4wCfRoooFMBHDuyFqzantXs08lCOe5r
boWBE2smyJDUElNsClBj8gcfeClijdAV2Cli7bYxbBSQ8rvW+41W2QAALROM7QjOZysysnBOgpD5
hkTzxTyg/vgn4QN6zvSCWN68bkIJWBH9ZjmPkmTcnD3W+tDSCNZSYHifbhmJb6Ra01A+b3KPqTUx
CEkvHOYJy1untz7UnqqLn1GMJD3/izyHntcBzMuzbjW1+Jjzk23DWsZDrRTMKZ6ux1VO/+YvD+Az
TYwe6Kgod0nfTHcPFeybUdPcY8CTZhaxlBfzc4LAYkw6ClffS0pfqzJHi/xjt75w21DhuRwz9TK2
rxJN3DO8lnf9AvaIc0DYQxGitOie/hAW4SFeWBIXBJG2hjFPMdpqmniPUObyVXd+fDQ+rxXJWdRJ
Knjr23dCasCt5LxbhbQJAuZZzZMol+SL9MnFdDYkZO6MWnpuNyuNTPWLQePY11crJmgbVcrRwytH
kgG6qa2uWEmIIrQe9U1kPH4F5XnWOJ3k++vzNYdmxEGnq9dkKKqv98gBlSoH3kyVIWNFczUFXIdi
ggRWHxls+xCwVPYjaHK0m1hTT+lqWCZx8EjENfyZh6GC4QPhrBVIrSaCy9D3DWFhrp++IIAnbMMk
bX6vTXdcUzIb4kiGlDku6OOERtFLaLzT7VeuRubiQkLuor+fPjjMJ64bbGhB1lcUJ8L1+1N/o2Ea
85WlauNt66ECVfZ+u/QqGBSUomvBoLD7KNsWXSiSmaKINI1O6z3R8M6T4j3PPT0N+kxHuYlSiDyk
qMEEtqjcj2cchV5QMVldPlAjwRMnMVj8qpSPgsXrr/D2brXLi5AZvgIMWaaTYZi7DS9e925+kV7l
T5ry8DpG87gurPfgqC0hDyZWfR0zkqh1s04AlR4z18b6vbi6SvICgl9oma96WrfGwqhEDlqmMoPn
HB74CjRDnx4zRrnhna+FYfpeNpbjwaXU6dcEwRIhxPDX/YezZgDCdO5ESQPgGEeDBUXUxcU9JMOr
ljGAEEOqg+Tox3CBl9gGUrBtQurZbcb46MlaTsSYkTFLi8HHouNxGA9xf793of0Clfnb5DeSwi8d
uHuL4dK0y1gQrN/dv6j2hKf0WzR8idbLFMdieg7plvnUqKOEw/NJqTWi0HQmyfI3TquJ7ZoGOHag
PANKLcWeUbmDDD1ZnXTTiqlple49O2qC44RLFkU+sHy2hvZ+Z64NHqCBnzqdqZpM0CkOW0F88H5z
mNJIK97LFX5QiWrjIsFTfvMZ0Y0DTUtBT/PJ+RoITumzKfCGXS6wNIDaQUoW2ytVuHOELrNkvxdX
mJmM29HtVkCzLF4mULqyZVvq6G+H8e6+BuRx3YnzyJfdOldG/otjfsWHuRwE5rfy6Xz9YNiq/3rR
0wvs86zfis9FZqUbhspP8odefDi2+ZED0hyA1aIQKWNa27TaW27G9z4JmknF2NZqS/df4r+5zmcg
UvIQZDRBePHTE7xY4yMe9oi8TrdKEDOg2yUCDQ4Y3xZbrvQqZOQYH0f0wOOocS9Kh0wumjRvWz1J
TRZ9QfYjE8mv0BF/SDzIcNOLGbsitRaVs+y7+vLePJ7T3glWsPSc+P8Dzz/CGmaKw2PKW3d/nVWw
A3AJpCUx8VxYBLjKqwpbMeFT3vi+xKQ3Hvv9FxRKq9sh3VjAWG+R9GDds324sLT5FrktT3RdSHIy
pJX6wYAk7IokZBnxFPLBHZzE/osx23ZpQY/4WzVAUZ+B7UZdUO4CLHHcsl/cJbToFtdjcTZgYpKg
XRX3m2ZCZlHPdJEJdMlqZHTLQP0Nfgu5S2c16UJKmnwepveB4qqjJ0X2+BKCYZ5prBimTLNzGJJ7
XDZPGIg6y97J8LKx+ECt4HeJSXs7KmliUg761Wlok0sXY+WZ3OqL2Pp7rjbEsUoIjqgvJ9DJnOT8
usT1QRl/pPrRQ32cHaJgyGLKCsAmetiAX7wyEy8djLzWv/KsTEU3DR4pxoE6eICwNR57I+bZV3AY
wPO1pvcFNWs7DxUtZfLtBD9vXqBjmCVFIck5BO17yCEnkbhaRpTHUGe9CE9ebocAjTru/Yq6vMg/
/toknqQEO7amn+9JVWX2uoMChFxlGjsxfhXrVmENV2Pm1ouB+t9iyHMTzGMuUzR3QEOoNdOOVq6j
Y3Fv1RgSmHNfLul+OY05l69u8YDfyRu/aBISjvsnM0mi44LvKabyeJQwFylp0FvcmWxp1KlNmHnv
GeesJBgzRItBg7Kj6D+hN6PUriiokF+2Jx5dW7jZr6fpOFQO9jw078P9HGaQINaiD27ziUnJ3Mnr
oI2ODVnXSfaK7a2WdS1qXab/DKPImS/wegR6ovjDb+Y5tWCaZyZ9cc72RcdzxvEsq3/G3Jfgq3TX
tk9DKvObKtt4AONULfnV6wYaInQ70chBTELIC7JfXPcRZJyBuaPIHN89tkHLu5ZEMuzrKnPIKSdW
r+6jAMwOahfROpJxyhFxPeQd/aeD1mrESsWXs66VFMb/huK7cnxrd9m+xapHXYm9OP9MeSrIjGHe
FYayI6fUCbOMvka+3XsKCRBusc3Md5xj4rVdmZJMf5BDmCvaphm5vOnn76FCBqCkFjqo7accS7eo
TBMwJVF9w2sOXVhs/y0X9G32ol8s/ie+FoUrbapO7+FrXQP3wpz2oKkfMylfd6N5JlXLBtDyNIBl
wV3jPJ0VzWZsxJlD3xPf8kIVdRaqyLqvq94h/ti6vyPpxDibRos7qAeG+efzqYYJ0OzEADpvWBDv
u8CKFeswE0NYI9Z9RkFfF7BwfLpBP8v+z8VwB3idKKlMr+bo3AHy/yfOAE8Ytd+0ZzbA6BCKfmkh
DxbOCEoID6UKOcGmgSvccu/2+r0+6lUMF4ypUWuLzeKigE9IdQA6U7ke+9gudUTKX/Ay8j5VwR5V
Ypvzdz5GvhQWbLfWNV2ZWDJ/UFhLYispaLUuSuSY9aDATsc4lUuVnDriiI8zu1wHK3VaPaVfbmNp
MwKyU8cfSdwh4U3VplK5KOeEKKCW377MUWFoXlZ9xd5MobgA2UIyNv1PubomW11nhXSrrTOw039q
iJzJ45znnOFExPSTybxeBPDO5SMOWqucA5gdZApQHt/DpewLHogqRKGOzEtX23v6wFvVlwneNAV5
tuwpWYVhs2qzNBI0FRIgn50BSDr85XEyt0VmDbM2jQo8l/GLFZ/ZbUDmt1k05M4Miy9Ji8Afs2Xj
e+dZPQT9W4riJSt4z8S9lONma+cFzsNM0iHoiKqS4hiRhxBGqHCPbSTeiPlut1A0ctiAvXMSd3LB
CDh+X11EWETJOSn8EQa9gJr7ceXpBRwqnr9d7S4mB1Tp+rkN+iE2I8PYcv8H2AlSjWH1QHuYdYRz
+Y28l6vEMaoFaP5UYGI7U3M7PvjIf7+9ySVzghnUyGKDRvJkMpioOfUAIgdst1oBgZHCIOG2+p1A
70rVmib3cILQ4fuCmkddY/nSg7+7zbsCFq26iAEo5SkEcjlGuxw8Ub32zap5ieJYjqDYbgpXIBla
xyClwPCNeBAwNvHKdm99l1/7cy2GQGUF0r5NQTQh6Ga3lQjc7GvXsWhUb6jn/gkLn5dli2IEHQXN
K/QwXJ0O9BnSXRHhHRnNDPsOLBzGbUCfK55pOOFrFdQoyjZ2eVHZi2ZN9vtVWdGLoKD0bANSeHbO
TaN+tp/v+cajUq8Z+NwjxwNjSqbmJyJNEXngnhnxSUb+HzR5Eg5021+yMK5wGs5rHbXiDjN9NCxs
XRE+u07NX09kJP7w0SB3Lw7Yc8P7n6mDgWx9qB2+tOUzx2EhCCwVymHisSKRbfmnBvyOLRQludSo
3MeUEVGNbRvtT6bNc3VHxTF0qUhm+KlZ68+vFx/A9xiYzqZLITRr1+cfCWJBVveoiiYJri0z7CZ9
/B8uGBOvLF5jZbIfMPon89GR9o81XGwNjsKibZA9KpIFC5oxuC4a1aYxOWop8RNTIzT1z/Afd7bA
HQOAl6DbsBCLnZnrcG3fki6QeI0NUvo+VtZIAwGOyzleFX2aij+Metzs7HubKGmB2oJBEeXwL4CD
b2Fyt4w/kboJkCu4bd/yxhnRLnVz3emXKZwPHiWMxsGwb7BjQZqSp5P4rQAMZ1KTk0v9bdE8A8qz
mQCr0OX6CeWZwuNTOQr0NlVb69I0mf5oSZJ9XMHU3FQuyfqr6OJEQIrWOWwShj61GjkSnWD85/Gp
ULjiOOkUzbZ0hK/m85+aFHQ9YmW1uauXDl9k5AufiH1+kFHqWvIcmqoaBCD8YXy0e515hrWhRlnt
GKjcOsOvs7oLI8tXtwoQqexMx432yfpxc1nLsISRgk/Am8hhSaT5iIZWG5icuqFXcoNPdWn81Z4J
7+99xS4KvwiyM2IYp2jaMBoXzxYTXCmW+tNRlieS8mR3T6AGDdR1OAwNqa+Qxqc/1PBvaq0OvAz/
NKvYfSUaehe1nSFKewinROBkiiSzDCZ9aQ3yUOIL7NXuRAfFtoPRImN1vatK3E62KEFQOHZRYPi0
jpSPv4Jdoh9R8g1NP6raIXrzeE8dOPFgJsSeZ6A7pfMnkOcqZIV4yjMehyQn18wc865ZsKGpUZTI
5dVKwiXDk17gqMTKNhRQ123+rEEo1OuYJ4h1vqDy3RqzJd75f9lQGoO/ZzLV8lQ8dOfDnrrY7O0H
PbxDepZYXDLBPJBLCiogqaQUN9fHI/4uxhwTi1HsfyDiryUmHNSQvrBJ+uvzQ9qBmEZ1Z/EEMRmP
54yyNaaSUxTHwvs58ugtx+Adeb8yoSdZfzqsyRx3eVMOMaWbNqZfRzlsqvbERkCfl3AZEe4m4+Gw
bsiGsa5F6++w3SUYXd3voKJISMqoPv4zw9CjkR73cP/cKHmV/4Ajeh3/zHE7kgPR3Nac9sQlYIZ7
c8T4KmfhA23BD1BzDDsLVvYL6K6R3+3Wp6zojaZK0ZxSKt+vFaxaa3glmJke+2YjofyAHL3VCQDy
1878j28xowygFe/BEX8bSeiRVDrSZbbhMT5h92+O0eMIp9Eeq79Ydc5j8XLETFQIlDcVB9toijIN
dwGSZJBk5RiPdp/MKCzdwL/m0RBGHyjLqoIOsvnlpx5E6u5D9jz0Brh8yZwxWD+gP+UbV1qlWgGs
OsMsb76QWBFDe7904cp6OsPxAj5B3VwQhKSS/efLLp3YG0RvHX+0uvkTw8oq4OpwNtjatTRtgglK
QGi8/DjfWo/kL0RMH6/wH+yGsy+ml3XATbdIFTmZ6Lecm/4TlvPsaww2WGpN8sZlwT2aHdtNfA27
DRxcC2dkHGN2qDhsm+uLEuIbUMLoOB2WIvUoeLOx+kyQ8auwhHZJlvJqSNH1Az5YDOH6Cdgvn5Dh
24Nl7KH90wLQJav4r9ucbFItW6vniEKEkqJG8HBJN6uKfzolJopzK9UWGg+g7ZazfWvOFYo8Tk4s
q7gANQ4dC5DWtO0MS2XWHuw/dIo1vwUnZuHYInWmXrHq0VRMj3JUB2c8xjTlTwY5LLLoYLZTbar5
Zjj6E2G6aDprmgtXN6/sJnSPd1rbqgGAguSrhG0LjYby5pAwDHDAQFap2IbIzSbRNj8A4OWRqwQH
V1IQ/CEDhB0fSmyoKvXwZkYFLHCRVE1TorDIusGfFLACEbM85bNCnNa2+ZpivqEQr2DQQBZq7n8p
toAdJ5vECaFgTssg440BbTF+ymm0T1x0xGZuEEmCD5flPUwRzU5eWTpNOgsBv/TY/arwd2ziU79k
H3LI6cVA4HwzaZxFhfohFNo55nQKyDMBq4KPHuOtbIE/Kp8tsYtupCw2V9/+tppFXY5hzREGEONt
gqwk3+Er5RhgQReCXHwAh84L3TqMZVUIOzsQAw19npDnIZZL3yt9T/AdSDSX3Vl7U6/SoinEsJri
yFGtyFkv/UroHShmvsChoHGK7zLo8X6OcZ74hobuXjsLM/D4ByodousUzyowHSZdxLGCPaLTK8ce
Oky4njpCoUxrXWF/6VRrdIgOLN8vyPLht6LUdXRvPXv/JcaG4aW+UoESj2TNI1w+WcD9wv4uM44T
DlK9600XCpiKHBLHFOGI3bNVOrr/W6iwa2oY5D86M8ACqPVnUprKtDQW97owndqrPiBOp+TtH490
7CwnOdkG1bwo7C7JShrnC1U8V3F4TAvRYqG/ECEojlenoJ60zfpRdNBym4CaVos8BeWvzikmU5In
CKyeXnqEUy+8HvHL5w2aeQh0VhpMkgcVexoL5Vc0BWgYQ3A+TrfLzOI4t3tWBqEV262jGzKHWcTG
f0B6RkQ0bdms5JoInFqX7lDA2wtrJbWNtCvODF1JYvbzfB7VAsxrB0ZG4xHU8gc+KysrASUdH/Bp
m18ax5Q/aF8sLmOrD9iEzQLNHbdVTx0xN1OnI+Ai6P5QjVNk//KA5PFeGfDyRtNHWZ7aJbKhDM1/
rQ5vS/SvgELjmMrEPXhTRJkhsRU9AJNVj1e9qB7UVCF64gCHgFudRkLekFPS6421jWH/iapFH/++
BDVi3mRtc5d2Cs+8+h1kA7kuMgkqS0xsBJyB/F4P1AOxXFW3yQc0s4DKW/tlg+vFkrdxQ2u/SiIN
NW0gVvfJ8cIWa1FHyvbOU3NmCprjgGU0WnECym/H4mYO5Jut4QT9mBtm3rMWa9Q6UTXNlkroOJPq
SmXg314+eSANDsOrhxCkYonRiY1TnzbVjZzZnDDXc2T1vNq0Kag9lPE37U4T6FtGscO0+Y8F2ppO
3cXsdt5ZaUDYIuY99o1G1HcRVdl+a+gUw75szFwrz0j9008z9Ur8nvDxRZ0cj5oj/v99yE552g7V
4DTd1G+dFl4ibnDJJht4manvdi08uzIFerTz7RcXdJkkyrVk3Q9yGmgX2QIF81lCYusyJmIXhxtw
LaOm7jtTttkcg+ClLKdXrxgSCgtDvZRjhQxiiuG7BUMCB3zSAZEccsGb0tHCNCM2r7w34i1f1WWn
Raz23z9jiJcOZx5F7TTZzRIH7a/hy+t2kUDeFV6reGeVRkGjNvvMgCLOYOOd13R+JM7znZzFwyL1
jo/BfsncCNLRXSSoFOFdW999zdfdMdQQet7Ki3oxHLC3YKnMungQiWyGu92OVv+yCsH1fQXyxwuu
DBcPCXsSz9VjRMuoQtvhomKemIJHOfih1HlSfhdqur/XytCngXY7dBypRS7+MF34rwY0Jx+8t0fw
tfGXet/56QW3usA4MqMgLE2GChiR8pd9210TcQJEkRY16cXdcytGBRneSHHeYd4yNSCLbKqPCzpv
VJE8VlKARoBGVVoAYA3DETFHSEoGP28v2c4fNbyRCUHVAGzbnbIzxxxo/DSVGhrf8ydGbbrPKnS0
KVtfKTJ0VNpGMigkmapa/+Y7Z5+lcxq5G7c8be48pAnNQW24xzF/fSr7RJu4amRF5WjbkRgpEzvE
eBN5SECWUpkjGd+HBIYBuAUJvc0MpQdi1znecIfGi0RA59GGI3v6Rm6J+37VYrsS2Q4NYrrEBrz6
LS5hkyqqcnbf1xgOvri9fPXlYJW2kLqRFiqQ4rfosW8bxWA548hdORIpQMYHQXvdFxUemZWUNmVQ
gpEthCyv+NxUfcPXmN4sZePWJdJSFgwnArMx5vNyOZQIICabFqusdF5kHtqHks3N8xwm5lv2JhXJ
eM8x7woSQvHfxNHeLLHOaPdTXJ0MKd+JZ0I+Sv7RpYMtRGZbEQOq+olQJwY7oqPqxa6V81ZldLrf
zoZKRBRxfOGPZpkS91E1KbYjyBBEflrQK7ulocUat0WRUVBFlM0T2d3/dpNj4I0mEAfZ2ZxUaSOG
ajq9NaWBpwJ88S57qBIBFX9IVC8FxV8u4f/ise30n94Vf8To7Vn6Bw8dr/9u3274yLx/E4MarrzL
0FpsDCV4CZc+xx600cdDo0hOxW4AJQozcJlsGaBRDWqZ9FxwHyAHUjMMFw3I8g7SCdUZ1wFUtg9p
OY3xbdrDfjivEJF4MtCi55rNvcSclzXrxYkKxlT/XiNw8f+0yd8jbXWJbuW2xyMKzq2Bt2rIsDuM
WdZEeG/cRV6ZsKaQ31+dPqDzB2Iqd70q4fhn5Eqxr8RmqetiRDUIAjIYS9BRFZQCN611DUJPIwa5
6tq0Vj9hPYS+1oMmj4Lm5/4DMKWlZMBX+9gjOekI68Dop+qNY+ukNgGxNgtB4b3Y7yldZjReiJ4O
iIzzHYVxjpM9RV8q5+br5QSeKehoQ7ByNPbQ4AM1GT1Ens8SzFt7JuAzeyzRgxgdoMkwRiPkQwwP
l2JuEUxY4IqcQia2ZUUXvdi+yTEHM+aiSCx673D+VJmKmNVKPU3R0tx1BkJQh4qZYfC12mDH4u0t
41WAVp/DA0n5onSFLAfRxkhDUKlE1DmS6xcjkl/m1P7VEOGlYhYV0gTt0caj0zmjaF7g84S3oovM
A2AaYOnct+2mpra/fLM/549Mvj5YnqrbDJ35X3An3LIHUCoXzeLmcz78LHU47n/GoF5J34Vv8o9a
1M4x9w2znXXD6YAMObCGTnjHtULCnmulI++JQpMuf94FGiUMHJC3NFpSmf+fdp/F/S8iA9kdCsJi
zyKrtd6tsFuDAmSN2IoC7rZahA61yBQAwt8OixKpqfMhBQ8lquZSBpFEQhzTk9GRLyHa9qaaR91f
3UyIhn+F6pVCU3ieoQ5I+WTBk8Lt99yeAljAsA7DrS7GQ6xnma/xbwxeOZIACdjuwLOBsCBytL8n
NPHiFmfso1sh3EN6fiaIXAGC2iA8FcdrlCEUM5a/Cy61WNx1p8v9HrgVz2MQELrngp4zsjdENjYy
jqg5EvsZZw245QekXnmRRASz5FMe20yHnr5OlzP+Hy7CJS+4mpMOzCkBBOh1Jwa1FhWLln/baWP2
CII6HUA1b7nOUtaIQiUjHt67G1zOVEoNfYRMNtDlj9H2sZ+nQI/n4QL5QR8HZL2G3XQeDobrUs8U
CZcyqUeTm/cB+5/wPwn4cxTnNqKPCQND6j5T55e9D+nmAWOysYNBpBsJ4qBcqvej7KmvakH/WVyh
JWzLWnNPN85+7Gbk/RbtDur3VgUyZME9dPoawPpRlK/nm84GCGXX921U5VmwQTJ0Ak4OS7IFmG70
q+3jixd7wv+AHjFAk5pnDTiSrCIbzmpzJwjbiADTN9dB6SKLi/yCBO2OTxS6kO2v6ASw+yyfyrv+
SZlSpDl5F18078Ht6N9oUtE37BmpOFQTctF/rLyA/O/JCg23psVsIQsVY/ReUHKY4KppQpbvY9lD
N/fE1KN93U0UJG/f1kf9YlKTY1cR4NcakC7oToVG2e9XfBFKowZ+4S8UwDZZPklyZvbGH4VqdCZr
tiZCwSMD28R6Sqo4xU6fFvBJeA75lwbVbvDKNu8tzM6XYgHXMdW4hPsFU3lJ8QyNwiqm79Qsksbq
jJzbQMGEu7qzw2HnktXLgvDZkwCSuX2D1on8HWD29VWKkYfMnQUq3p+ERDk78zLIthbJOTDQsrq4
noL3L0HYf9w4X92g0tz9FxUxu9GEQxBm1Cd8zqUbTvf225s0mwzHch7f/o5hLLfRcxYqVuyh21dq
dLBAosrlvgv8VOvKn/HBtiRKatwzzDlVpuBkbIIRUeDF+MhhU/CApvLEhAYca+hJzAs+9yID1DXK
yLXPtTu3BZQRH7bkXgs+inqh0d75BzcjvQQdF2WwbJw3V/8d+PdMB78iOa/16HRjE/4KV01588Sd
tZChHH6xp5/yhY9QVPQanTxdWkKBpYnOkyrAhmnC79kYX/GYv1Hw2j4h6ZgfwW/ry02XP7BItpWb
nAmgpM39Fl2D9vgWwGLU08Ke4k3lFzMZFcxGJuAXFhWxpZNM854y3x6Y/3DjHxCgHtEiryCytRZJ
kcnLNnH1V6NjpG69lyF6SLcH5nKF3Ur7yCxIKl1spwJj9sXLjz5jKloTe8ov6PyHAKICE38LK/aG
bXvPlUvWywC61Xcn3pC2+wxgN1f7qnzJFLrAGG5z/H3nJ7paOC2eKFIuyGDKcEqR1DmtVLmWPg/m
VaDBLFKLQf0gxRpXUnlFkDe99cOJpK5ee1SRVMxxVjWjIOSdwz+z0aXXNQl/dCMUJMUoffmgaqRD
UuhQOL0qB0VpU3lXBNR8WzyxuGhj6XzyVyz8Fw23C0atgFQK5Nyv+FQ4UzNWDJwk3IiNYgaBoYuI
yyUzT0ZS3c/f+op+8Tg9wGtr6VQGhnqgDbbPdrM4zsAJ9ulSWkxLvz/4uD1j82lre7xL4zL1uZ56
tAHuaYyXrpcVq2/Ca0O4MKEmwafIZs5Ij+s7PkxKnuqcYI/Aw6+EKtSB+I1/abtbVfENf4dag4ht
8YRAGexXmcEGyzfTKyTGCR36UBsVBbyCnU64okTYjOYliGXQcdGkei8mLOWwpsPwqOIUlqUnwdhT
PDkeeX7M38G3ZMOvCMpxEGZ0qCnxvq/HL2QzFeSoOjmIn1rWVlf224+78++XuvllwYxNZYt9APJf
v2VQd57NakAEvPCPoqLaHrir636rrDCLf1qEZZrzQ3e0ffw54GZ5X1V6/RaQ4bJ14ChBQX0nMFJq
+FgJJDl3DOXvdM7v84q3kg2L3khBVfxOk2+vBDWl1mJzTu6utpLJDq4ZX6dxpj3+xCZxEEGyW7X3
xNfZINnbNVyNIN7ybH44XGDtXTi3ofEfqkqko32nY+OKydSOGzHYVnyUXQAspgtNhJOBWVY0lqdO
RtT2Aio4kCg+ge9s4bSf7BwLpIjOlykaAZNGDmplYLBeL6JryJNAUCLjM2/uHGxmDHNdUIgy0Jvp
lF5rPwXWxN+VavnUAsHByy0adhY/V1NT3vr5PjMwClImF8xGCasjIfErUv0Ax7O8LUrQiFHKVMCp
y5PDzR+OnWS+BUiz82+A8OzFMBGZuuvYlvETvf5+gSPolI2UZRKfzstNgB6rtvdIHcG4vrOi8/On
ZkTZmSZS55pg/3TEhc+YQILSdYkhEaurdPtSdUWMB5JpBvfBoqWWTQgi4uB8/SiwmZYbhaCfoZ1+
03Tz3bsOwN1+eX69gAMkhpnfmf88jpk2jTu9doyVsoZeR7mKv6savz+99NNPqMK8GHHcGdJn6Hyb
907nW7f2Nxs9beyQCz/q/g3iTKqA/IZU/cx7YDbg7KTv68DvGvJgEvAm/7c4sPKUAiDPhXXN5xLt
nnvoZMYbNZGR3n/ckNl7LSXhKWTHTXWbGGWBcSyC+O9TsYtjobbR4UNYRg0UMtSyvFBGESocWNH1
h06rgri1DE6pbo6geLXqihLcWlG1XJcyycmHjT7fhWI+SXdI6n/RxXKyDQK7JU/t6u5kPvtSyC+Q
s7A+ACrO9/UnxLshs5YfA+X6L6HoHT4lDYM+qCQS3tWZxgi42bHG8RkCqsfHqn6O/YrwDcNXHg/E
5N9EYKi0hwny3AgWKRvMrA3ZuH8iXH6sE+73S4SWiE2e++2nMiFg7vxrRPST5m/1fapokFEJW5Yy
sD9L6BUpLA9DnETMtes00Z93ol9SK5bkI5TUAx5dOzTYnrwbciImUyYRzO4w8TQLW0r+dSAO5UzJ
wXPh+YLvaH4RSXB/0aADiAAUUQ8CnW+FbTb6gAnwjzKEXX2/CUAKkcH56gbOjC/0BrgI+AFGttdD
72Ku3eSzt6Jcb5knH8WnBliqyc6J9GXEZy+6oNpqwrBnCkszG+wGT1jiYBnq6f3L9n+85Ji6IHkM
lKt5e0QutbjKXI7WRjP0v20ZcEbUnQdXZaBCrChRGSv6VexLixVEtjgsGk5qJrARXTGKE4KX/p5F
JU9PoQbqqqQJSEfy1wAYqIfQZ9OVh1L+7rUWrGN3FH6BxOnJO5xpE1iBzd4EHKdAgfzM2IB+laz/
EJNOBBHU0lOgojPyt6s6NY0JCAPd3DTATJyJ1Xeivsak+1aAEZnfXvdDv/K41OmT8UEFPS43SpPu
Kv8FEeLnswszaDyR6JD+Pw1il9VVLgEta7u/EOp2fjbPMqiwdxAQpdyjXAepYYFmyX5UX6AwNH5T
XEzIAk2OfZsaGtcKgzj1vAguIXC4UQD1voDUwKnJxrN1iLurxnlT6bexJB7v0uIru/a2S0JSXrfF
GkX+TTTgojLipU/6bp8Ai8nGRCl6EF/X/s8CTA2kbpjuJCJ/gDewZdP5xlXsPzbWas3dyvhuWMxi
Hal4HCD5XP8fd5/o4PIpbtuZ4siwzBHPtNwbV4IXUtMetBR8HpEdr9DoHegWxwh+UWVNPt+UydHj
oJI6wJaimgkMyqE12fbiPGYT6uU2Ir0j2pZKcmequOURboY+uzHCCF0wfPVtTpqX51Quz/Fa2KqW
5jz76NOC5e4CwJa2n4WHx2C1vt4pieiEPa4sDGY7D5L05JknHSp4lXRSuzoNLO89q2DoqK/1EOk3
bklXoYUDuhRvhllrIb+PS/V3sGaD7zPSxE0xRwxOCyqqs7yUiRrAIWQWzE67bMBOYKGTOSONjrJt
w2JTkEys2IyRANQ6usc6by8CgHlGg171XAohI98FkpXooUcRaxyI/IRhmrE5A9fQZidBHMLvdk1L
5fbZkynpty0jxIXdYH6d/G2kAPe11KXbZrD5o0dx6MdRMLWDpWvQocSNi7FJeGM6p+Eiim1s2feA
z1MA0sn24sBLMWALqO6RJ2mG1xqdiFmBPGu0YC7rIwEtYmCqABjE+hpFmjR2Rvi3yI46vtUMiibr
Y3HT6m6jZiC9cTyZWVB/OuvVrNEpt9abyzdsYtqHIiuHd2WMLMh2axnQwZPU+BeH6MO0H5jjLbpv
vqMSD6vTqqLB177xES906IQvsSWBh9Nh2cxpzWyB2XDAsVAeU2nDGRLJi40rBbe5ikgVS83OmdZf
K84e/pfqYdbjEamZDFbf2wJYLxG9nUDb58SK1wAPZqVWoISrpX0vJQkfP14TUn96Po/+ngTZtrie
ZR2xmOCHNBIjpqtq/RvjSytfl3cT49AA3T+6kcX/ww/gU24DkgeaIkIQOVt+n3cI8qWjhIh08ifD
lE2nb/BztfK5RYEtCFCKXGt+ImqjZlIkmMf16l96xRGZhb1hTwPaGfe6D9o/7tT7PSp2q2xNk2rZ
IfhC7Ohbjpghg9MCveS4/C1AB01b4bObUMsvxAu1isZmNsyxJVgsljTvfyUHGDEjjsF8qUWcGmES
1PkfzekCSwpDBR8sxN8RaIFKynZ3fbH4rOcMFtexFRRDTlDUgZc6KG4jveVOcERa8UI3OX2YPI5K
pw/2kVORLzxb1j6DGH7bmdSYQdRAHSgjqiaivcPOpDmPUR/xW2LNbXvFrRqLF6VPpbi4dIn2wP8M
A1c0PCNkafVgyY9g1T/6h2v7K+xsjZtqKFph7TMiVDm8MnEJ4j1dn4eOz/Q/IdIVPyDI+AR4S63+
PUA/RzNyu2m56NVL/ZRELrZVjdFV3MGBdyAIj3S8Uwl5IqyG1A5COm+7rd8Fvx5DsE4CpywpeF18
K36mLMVdyTB+Ggm/ZGXhxIpM2Yvlj8aXkfES2ofXF+tcTuQGFCe3GVhIklFchPfeNuV1mLnqPcZa
2+b+N0liVdWKcMymILEdwEhLAxeB6fPKo8R8YZk05KwAU3isD37cYlOBmzCBv/h9UrHECACAQ4Go
vGSCvHuuXY1GOJUR7IrR10CFnZ/c9dRqUGY6N58BwdOG+dH3s3IxTiFUInqeBlc1n/TMXvBrpKqs
zSYSmJw6I+4Qn3nof/eWBEqJOtTnrtomAE5F6KBirCQy7/ioHeuR9R5SPl7/V35bQYuZeR1E7FN5
+T+ZyeKZKBAYZGO19johGJGcx10y5gSpXglw7vrI3xknzKy4Yh4vlligq5zlB/IWN09G1uyPRQNl
X6PE/WwAqxv4wEQCyqyt/8uGdSH8F5Lhjk9OZeb8n7SajWkNJRZIKqpUtGkGA5T763gMlUoOlCqb
PrbYn3u/vAl/nb3fpbkEP3ecoNqrmi2sI6xAF5emfM23+ds0+fMNDkj6rfs8IgZL1dSlkLwxVHET
FKB9Hor3FxQM2GjSkOcPzKcHZ4QsKXXY54Y4XcL85A2tWnQQm8uDvabk/+yUZp9BCIruvnncRv1Q
lTdIPCuopwe/nkWBoUxePAo8O/crw8vPO4QO9NEcp4i+pynkCBA9hwj8wRL6CjR3FKbBsjLRgkZE
nfKl09f7R0jKJN29DK6wwsl4J5NwGXkB1jGWiG1yUgDh9rlPwcwKJW5ry1CfS6uFjPD/uH88wVAC
J8j3anA+A5vJr//txH5mNFb/X6yLxfARKM09NbqhazgWzixefXMnTZ40BCM/tKazZRtnuZZ0GwIF
B3wKuHJfF7NhdyygM/vg6CrOToa0kg+qVKwkDYdg2fGgWOKqppxHJ9yXQHV5ZvoXpNIgH0HdP3hj
ff5v4VtljhP9NN35RhFm2yxP0HCGPTa1awHMGQrBOan3lo8x6/1TfVE8bFWjc1Lo5pooOn5wDai3
hP3UAGFLQ/PlHzJkbUCFK7ixu1I2TvH/AFrjqCqHvfglLt8kphccipTcss2HSvtB2ZDVZH31DsRF
AFhJRgEIsq0/9+h2u62ZGFKIqkIdVbqQwfgOTxQzsVI1I8c1gDhdwSjDbnilUJHf7/+2FXCJ/I/G
xfG/CEfBetptPW83zkRCKvz28br5BVNGQFhlezpzefyzhGc6juE/CMXoyp7o+vmYLU9j9pD/5FIf
hH0i6ctmarUt9bb10OwfTqkcnt7ep//YVnUOqBZm6GRZMJ1nuIJJu5zBouO1Gp5RSMMhXLWJ0/dC
LuxoKr23CecT3nUuuAI9VLjl8G3xv0+2p2rqbqcYcTaKu2A+Du083RS5LL5U4Kh2y7NDCX005zzI
QCUB2vfQ+llP6u1UaPqJ8ywDCAZIGJn6pHddHvvEQGtPyofHarOR7DfeP+ByUNg4fniiGiXZl9yT
DVnk3MRPBjemNZyNuln5de9YX68u/guLL+l1YIUyOj0YUGs2qCzjK/xc4Y2xiingVNmGxH2Q82CL
TbwLpHKM3RzP3gQXsLlpRv8yVndWChF+lH2yzAH0XHhpdAgCfCx0KibRprPaVK12/UKgtpdRwpZw
qlLEVP/l+DdUJJJH9hrqD9IGNyO8gMmexf8GAzD/q33t77liDO+yxGLbFTOdT07NCKyGZpVGvD3F
sqVFEEmCodXHy25SNp7tN5leRlXP2t7ZyHzfjUbV3ux3LxPbqocUESEG4vIBiptEzj2+17ig2LmI
gt1j6+5yRSznOeNiaDfNOS8gwd1nnbB3Mb/u5xel3fah3iwDIogYIQ+wLhsmWSoIJ+Odfrkh801I
9cnhqhJwUlwVjXz11cS6AwUkfx5v/1mRmp7Qo1XuDz3AdzU+4wm6h8siYDIPdfmgoEniZAA2VNO5
+j5HhR+OFct4vvoS26PbipBsw2pMC1F1kRvXTONJRqrAQzWGV8GiaBCvSiA2UTrbASkCbAMLGBXd
WgpIN0yZMu3B963bZDTRT2Ivl0eQL3xNHCazZyclCEAmvUew2LbtV1kjzfZkeqkvMDKv+wwXTVCm
a33uT1QIV8jbblrtxDUC6WxiogfUhTgv1FWZlxq+tprg7f74/9HvcGcXYfIGVAwbj/N4BdahW2uj
LYGMv7CYEbzfFDsGN6he6BfyP6wW0bXWKhwAYNiINx282dncDaempMVRW8VkQcf8bizBGJuOhmzk
kQv9rccNUjlPt94zncRWNob63rIuD469rgVJ9w4ht8SM0f+l511Th3iLdqIUDWX6zoKB2Zwco8Mb
b+WNcNdORw7xINCVohL+uIrfWxjpp+BKHyWDCxMA46Frgt0rfjv3Mix8NBvyPxx3KdWE0ckVTDmK
8l/2BN7u0PvAJQBuXv5J/aByvufZeoxH8ajX7JQ3e7zXzjD6dKQexOlVw48Hh7+6sHoVp7a+p6X/
kkzjpcQFdeTDskXYj3t4EhJefj/6IVeo2wy8/UioyHM/baweBSOGCNxxYc0AFbJ5dMlV7pY5Lh/2
tvQ6T5Lt5MPatNz3tHm45dcn+W/sGjp67baVuf3wV0MUVS8fqAr7jbwIJUZgLxlWiWkh4QRNE1mH
pG8/d5KhrnNfj60ZBzhW67tYRZ1eI/zgIdrPoixKYchIEfGoy+BxZv+Ai9FttQ0j0+ve5xWV4NhF
DvRk86PY5Ntd3aqwGxeLvAp0l4htAaAVMs5HlcYzViKFiNffqsCN+xGZrBngz6HwhGXDA8gMySof
ZRvm3cWJpl7dLu+TNeKBXj5KC+VmElEcOs82Jo8Q4eM/IwJMeo95lTFLU90VUvcvR81r7g9Va+2o
F8MydCDIs6b1oDuoVj+4r9qt2B8KerUywW5upJcQg4KlbG4osi4N76CAz7SwB6FkoMkrbmb5kVH+
lluv+8Xc0rMebHpOaxfrDeRmvMsYH6l+HhcC5RWnjXgCNQOOejeRwhiUgn3fKtn+yoHDb4f2BpA3
tWBP7YuPuxGuhdOLx6L2cXZLrMH2YvZtYfkxTPLjQ93ghfHMRfEyBZ7jp/25lJlhNls1AcR4JQCV
I7t4Xg2dPupk4Jcw6S4vFfPPUhgghtv3EZU9QJTDAsPFv9IjxngdCqC4KtgOJhc1cTuF2v0YxRa3
/SGvSlsYqYKga+AcoXmmuSiwXEf/Ks5qLB3jWZeekgtu2++Ld+HtXWjkiNyTmYGuwqTbKcIlRUet
B3rogYovbtvNZ0p/0mSWMBM3V/QKamQzrhyRhwUycP7xB5qmdejZmGwhhQs7qp+luURHUpafBm8V
VojjYgnEgcaHiCqeQiKJt76kGXGgfkFGAWd1fHeuYvCl4OAK9UtMjv4JeNonzPwdW7R//exg8jmE
/i30NJNh6NBt50U11EDZyar1GP6wYn/88oT4oBP3kOcCqJwo4WTQ3YVyArxcGi8Ozhk5ARYWGimu
TjUpyMqsRvInDt54UKVN0VtIz3poB6UVcRl1nRQPw+wVdHixA8WSjjqzXtvsq2375tWUUiGyxV6m
u46KGT9KKkcaKFND9U1XL4c6Qd4mTMH0LVOxVLZneB6E9lbuWGRdnLusX0Th3I0Rq9E6YEUnxbvg
Z3k1ZM/O8E+BpMusTJlPnLijPMoWCw7clLtACkvDwWkOQclnWYEHoNWl4f4H65BGPOg2pkPh3L8b
7JQn5dfvrszrUjIAM8SSyZFk3GKWudPl5FxUApwvOYM/9hpat4G+5qsPhf2W3D3EwJUEqEdgNAjH
OVJLA6PLuSWhJ9ciB/RhcQL3oj9ZxWpGLw8LhXoH+5pR+zC6DNaRIGugP5w5v4gSKD4PTqFhm1ml
7/S8gAxSp3EQ0U+MR6tdowFlJPJkbvZQc9ydmzLWhGzggOcYdFiy7sQVvTn8WuDe0rGuasBcWu3v
SSw7AJDYGY18IlKCcSE6Wnx96LxGCKbpK51uoevFPoT5md4FcmH5QPQ/Rer831kLJa6bvMKWwdw4
w6UkGjI0CFK0xc/Indqwjtn1u0mgd8HCJiXHRwf7hpMRFd848UQ5zQXN0013Y1nB2n9XhuWaqKFF
18ieQY9n0/ooBk/Q5P2KWf5+8xJ3uiomoCGOftzyDsVZ22gP3YTJB9/ujL34ibFotY8tNQhoQMRM
L8FEwJq3GKQV1qORwdrk2Gr3iMkAzfnpH3ct22DOKGcYV5EehgR+6Ha91wVoWP0Sfd3ZadSk2Y7l
zxdHFtgldbqP0jgYqv7H74pxXHqSgY3r5TpzlFt96aqoufV9alkmw93ovRn+2CtDJMCgFv9BKq14
VufsCcKNkHmx9YZumAqEcXzyRACim8Pw3h9c0X9ZE+BNzkgmtCTztkdfnLCZULhjfRnxC/mwIpfa
XtvYGBjOUvRqxHcZe+XSdLKsZuZ3ky+OpEYjIMOoRKskVqVf7NN60XVlIo6lJ6Y/Z/dbA9qKzAIu
An8FEj0L9NCt/P6UZ3BpaNJl6owv4eH34imUUZWhN4BzLuvZfvo3IlFyousJW4Ns0SP/Nkj2AUhi
SUXzPFgAA6NUATX3s5ailA2ABOphxsUgOYVV04KD5Z14Ho6Uwbq3pebZ5BVFZUPFWQ8ovbhZLCyo
koe1n8VHhbJE8BZZluEZrAVV94NDAJmtYFzUuWH9tBQBOHfOFovX5Pzc8kOkNpU3f8+q74gm511f
S9V+NjdDYKXJIfylJEmcGDfkURPKMktszY86fnsGXsCRB9fB235DQewGwDXSmE4fPkmKD5J0hjUI
yPnfpRIgH/d7IkA5+gRKyfzobM5KfBH+U0+K85OjeDHwdKTblgF+zofW3dKT+COBduWVXzUqV1lG
ALPybmcEODS/7lTSnWmpl3W7F5XQ5b3BTVIvjzpQuKXogu4LzjDZZN7q34zf//tR7j2/b4aVcKMP
/w3dX8K8RJyAyApgXxCbfbyX0urPpECQS4EEcI96CwJHQXDxDhp+rHaHSwmwNJCA53QvT2+mcrUv
mhDxfBonGdZALNWzzb+KCR/GpdEps4Pip4sb7t1H/AsrQY4yiJYbPV5alL05w1Ekn9/1rSA7mt0P
defKy0HiObe6SSj9eFwLh5ADYJ4gXmma3GYJfU2vLDE7/VIYAcNPSOZwc2RbD3dY0LPsyNIECZR8
GcyAFYfcSQM98WZKIBJOEUVPFm9ppMnPLZ5g7L6hJEBMr1zyiCTScD6ttaCHSphRuE0dilWnVLxi
4QjLeBFMxDidixtKCqARdg1syZELiX/M0FyUS05EkdiKkH6bEWm6Er7z1LXYPSSR5lcFfXadVtI5
fuEti11qnDAmyG6Xr4XtmFyVOVHdHXU3CV5sjyT1YkkyP/knHkxPz8w12TYgPYgd6EkB5ie3QNJ0
MYCEM0WksA0X4G0bLKa2QE9IUWBA0mIV6PaZj9Pga2MTS9RfztY13GZoba/59UmeQcDtiISvd9sN
2XkUT6x8xZ8M0Z9f250nR9IWDOSgCy+y6XoyJILS6JyHXGsQ92yWWb9kJpn5afPTSUmfSydykzC8
KBal5mROq1HIt0H72mhirMsPSU8TIi/8+BzxWKDDkv7lp0vGfX5uxnOrQ9YuRtWGIvIxYjSPBWBF
i24UmsrncHCMNMhGegP1F7SqPgj69Z3lo/2SUl6GhYOcflzEZ9LFX/IwcCDyawNNxgLUC0zTSQZA
UfwJDR4aIoqNB9+F0ensGHpxkqlSiAzM1PLIIn1KIozmlu3J7+LDNKFw71DrPgRxtP2ENSYzvXgO
WftP5i9lt6MiYIbywr+61Yfm3ismM1n0ya/emC0W212CpYQpWLjN0t7jznA70pxQwUvOVCts3ApC
u1/mzMf/kOW6E3iKVvtAj5D+pwx6iQB5BPWgN7jMnttI9tFXcoymYmjwKb0ffxNQ5Dzr0W5noT6n
0nCmEWHMMmEH3H2nuaOa/qsa5+Od0nl6EI20E5yhKjeeKhaENch5MRb/N2fZS0ly7Fwn7oOcKAMT
JtXbPWr9XxhPTpmFUeWzr5gS2/via0qx+fNoMs0OtPJDTbaUSTvzVNtKDzr7Nbh1tNXym+0lirAP
TGT/gTPSdy9rrfEjaeYIZewuCQW9RZxbO3aGYuwuHBWL9KIKJlswizWtueopMWxzeXdNqUVDKwXB
hTgtZ4EhWipIr989Ry98beDV3w6q6NuPTaFRb2vEvkd+xx5/fYJoZb3/u7O1UtJyo60DRzupfOdX
y4cxzWI47qIo6smFI2rkIVxbcPi1F2NENjIfOnjA6yASZxTEpgANQPUIZLda7rnf0MqW0mbOGNyz
CSa1xoCDIBgqLt96mtGFA7jexPsHPCiPW17hnMSjU3OhkeodhgOEndErC0k20dKlIw5C/rEskQkW
fnyJVxJuFa0QIHBwIxThD8L5kZbAVM6jIcPu3+laiJVEtOrsDt8Ba0XhupJx58Q1mJoaNxQPurcV
+95LRT5B/F3K4/nGW1xGhf/NjNxXxSOm+501SnJFYWnvr9lFMVRlzGaeZ3UMaPQAFep0PlGFIbN3
uQ+1nrq1nDjAFJTYboWWR9aMKOBiEsawO5JjY42IUBXMF6zA0Nga1wgUYMY1GRu7LneLVg210mmW
s8yaeejiDLhC3vJ8nBS0m/DUoTTngVNt+fjJLQagVJw9V6GCzN4Iv1qsKeapI6snpYKTP1v42j+T
QphFzNA0jazkMlJ13egnteUnkn+RLREb1u5kC3M9/KhH4UFbo+m8du33kzSl+75Zl/qhtwFBizlh
rg2m4ape56qyhdkUk2/fRjr1Cy8eNAHiu4mwhSOdCgjkZDk2X1bFCcEimjzKZswhx0ol29AXE7vx
0t+ZVnAn2cbOSqwll3gJc2+nq5ARZFEblbUv9nr4rFw1LxrvBH+nIquS0uyPnPaBAkt9npo7PKP3
IoQIh+ac3KiaaCRZeqIAl1JwCxrbxPh3ZGfXUEBngMfEcjBNvtlaoDRDzUAC893h9rXAIWmo9PVp
FA3OQwasSzL4KL6YCeNM1eqftqt02R8NrX6Z0CjqD6vdsBYjeHUGRNRMWDRoyuS8lq6DDbli+NiY
g28PQY+UTh2GNqO+oALOz6phRr1SOOjTk4ZoYOHR0IaLe+pbOkF2WcbtNhB+UQsZkV/kvKNxSZ8j
ZULle7IvlcDVDez6YoZ3bT8ebo2QfWpWkgIIoxByBXsNHnkzfS1qGvXTLzNaVWhfT2sr03glmYCZ
yD57rujeKIloM7yrqkqkJarBNUdGBsJKIlv/jXfI2C6O2OgpXM0q6SFwrgplENa+b1731qx0lMld
w7/6NQSAY9l1TxhBfRylwXAKTtuZKWWbHzPparOgWAtJzuIgNBG0nbpXDODgzVOfC98mJHwAPRR5
Cjpwv2UkaNz0AjyX5IKo51b9RypaDizVN4/nIJSCx153KbiRvl8cmcil0VVVNfSw0vvGVsypGnAq
xENNFJtYSnkgo5JuIvNd4ayatZ9QOkktz1T667ZU0/DAtMqImLdOVvc9pWwG+N2rAxFBRSG07l+q
sbv49heEKgXffNN650jZUhZdkBSaqxgDE7ZQMlImhdmEvaCmFGocPNxVcgWxfWO8D+xvoBPY7f6P
J4H/3ukAFTB4uOlAp4I2WfiMG9XpJKWlOoOQjg7bYeaCCalCYeK36AljwOesC/RlGWbJl6FMmJ4y
7AV6siFo/wb+jp9gYh7Mwi5Q3Hgjbq+8oRhBiGPmwVXbmhOMAHI7RrmuK5UiuNEaTQgCdY76zYod
d7ddoEhYms8S4o8X/GNT3EnWbH0LuQ+GF7nL3TxpIcoAx1ehzovHB6iFJbVSQveGf2zA/O4wsIUl
LnIQBBZL06jxVu1yyVwiFvu0Ut9gCbtFqPn7q28lLYIR2/tGKPPOZTtXatlCGV08We9PlzlKvu/F
6FdYhhcR2qUYXyYAX4VRDdti+N4xCR5Yob2tAydf1M2uQoTb1m2o0W9RN5UEzqMQILtBFL8bRddl
NhTC1GdGdSSALQTGaK5nqc/ryqRsy9TlGaCbobCmxXwzjQoTAptCujDC35VR5ARGI8Pvkwt+JYcP
mkslhZa2Z9x7N7snY4ulq7lZOIf6z6hQtRyqtpPNljtaF03eFhWkPW/rkHqhGE8Eh/Kxq10xzjcq
17/t6RnNpCrqvlNHmqsqC90ptVuM/UQ3ET0hb8sZAglYi7kz2UFRr0CW1F8sGobhFDotQG1zJIAo
yZ/bT6QWY0kC1TQ685eJGLcv7mjIbGI58jMIztEYLnLX1oxQP/y6KTpJVq2B7/paoWfqXdNPqU9j
CqoDnWDGbmT+bwgEU79eK6xPJPrSx7GdDub2L67FPMguqjWzSBtlk07IfXga+NzSoVlFMZ4BUhjp
sW3gUAtDC2QgBg3tUDL7Y2zCk3RdWduBA7qkLn3orMJDWddo6RlelKX/sPzfB/TQXu7dRXOk4TCV
gt9T8FBo2aTB6Rus5LmHjOw4YX0Sb2voRQuEg4jXem+Nl+CvhYSllQ2DghAWpvdxhCVoozTEvBTE
wRv8MNOK2Zlk+1gN4QMSOtOUIfL+vVDz7pxbBJ5Iizd0aYNTJ5qvlz6m9kMWKu/LLkIw5AoL7GdS
AufeyBiUTAIEkFfz2b6t07icBH0KLfUcPvPYYt+qx7M+KmOiZ4EhsBv8bOC5teX6Yk/fymmfjEaH
bH9318DvYd6DpPfuSCr99zEdKm3MXUs+N6k2h+CWQ9iyeODPr9f+fegH49LPQAkRXdSgdHSjgeEY
Iyokjt8b1lEn2v9uLzyTjlIOqFHThxxqush6jobLJW/WNL1QaebvQ+6nwCiMqmWvG43aGPSOxdRb
oyyJpclwemDipytnNdsHT7OGdaCMSy4YzoeadDRU4cemlEHzDHCZJ/iSmFu9VOAajMjNOb+R1RhI
GXZBKE5uylOiKvG+nbdDmX+61jGQJHo2P+NiLSQyKqBL0F4VArKAJbh4uNVx+4DSYLd4la174zta
/vxcjoow0LJa3SQZBMnio56gxKGXZKS4aNW9Gi2AbsbjenC9uMOUHavRgcMHQTDhF+jmgzBfWKFK
wy11axWUAJQyuXLCiCqY+LCn9o4ZRPSJXUjHAsSQAi5mw6mP1QKNkw89kC5HFtIDyFzkLq218c+a
r6TboKk7DCv/vzEryGo0vVJZO8sPoSzIC7U3UtC8glkKkMeic5ZVtoBVjfXRg6Naf7Is/z5PDR4H
7dDssvfjDgG5YDhgHkULvuqi3W9EMH4Is3MNsRK5FpkhD5gJaIR1U3Elo56geOJSD1YTI8JiqTPK
Ujs+zq+3EK4iceR8rp6dLBAYwOXJ1c8dPDNxC4By8IQhsCqpbdt9AJKDqdSvpYOQrIXZvQUky/NC
oXEVYV6kLqRfoER8FMIkdWe6mWD6xGBW08d0sWtykVEUl+K46SNl4f/uWqgvJ4u/Ars66O5wZiSL
oE03uNd7elF1lSiE/Bo7iWpOZBanza8OjcEugL3d5bTdjVf63TQ28B5Y9Omdshxz06PcfMNTV069
0OPp+wTqAPefrl0m0/WxJtln77dzK40OK54VMf25hlPSBy0wdki/8vKHnKsSdsDDRYeioycUL7MT
szj5/mWBmkz74DcO7eKBi1JoxlIPiHmdpVOy/Rbqtin2nie5FB+wiLCEcSYylomj6x2PjR2tMUMt
mDQRMEy9/0Y5SmRwnsZG71yAVw5D5XLQ6gmk6KxgW9jQmXeFDvmPwcRhNyGp4Zk+Pk67ByhwePSr
vXiHYbx4Mtb74o1U4yW5Nj1WflnoJ7cFtdA2+rPXRc3BDAHPJRbF4NXsOf4jNTVsnJIGu4RW3kzc
wC9jP7HSh6KSC+DdjPhOxB69WjNL97Zk3IIKReaZoFWD8cbDXVh7YvkVToEsX0G9MIceZ/lMuMTQ
vpwuMTtfvYf9vZQovuX9BduNS8ESJlPkwiVHYrdDRXR8Tno1wk6hTr4XsfbV6e4F9eKg6JlQ71pD
uoP43JlMhNKiJm6hWd8tLDMGutGj4ilNruwSgWtZ12kRYplcJA0GELwExwEpeOXRLGuWk0cp11X4
E5KJfPuqTuwHw+JZWPS6UVzenuiFsZQx3PP2MhsvGxmXVStAzAJ25DEm8nofSnIxL4PR4vD+Io7Q
Xt2noYGW0bAHQxdtGDiTH5J1bd2LXpOM4mm1S9EsJzOEwnMszoJoHLtRKEZZuBB/6Pj45KF9xduS
pb+gvmhXJ1D2UB5RHuzXMApNofDWiXVQNN3yJdpatQVl8IWeay3yHvPYzmQMWstO9/PmGyFFIccs
ZzGcXKMi9ouocDg00lUJysUiuKdTDZqtUkzXBxYHC7Qbv+wx4c3zI0T5R0PQxbx3lssqC9vgRYwk
ct78305P1jsdwyvyybGxBIdm/A44l8SXN8CcOUA8UkVlAazmbfpxhVHqkvTJS/wnpDDb9ZVVO489
FKz5r7mm+V09VQWyz1PdC3ipXa1cAOjC1E7cn4hbaxIGvGv5vpgRKxSmY5mZodkRX4HCuI6KGlKg
TfPr93CK4bkAcEBbS+wh4RgJKNceMtvWbbHSvOGKNCN/NI5/rZjY5hpAJ7F/jOQlDhwnweUnEPwQ
NEjeZ53jwNhOftYpxDz5weM9sOIc4GpMa3FAqVLuW31/H7xJoWKty2ojpOs3byntNCW0DM4LxY8X
JzSNiSAzpj7W/IHX991SgZS4Crf4ujtsLcx29fDwUYATJ5efznm++0rMZqHBgKLqbOsDzJcC7h1Y
tJW0I7qIscu5mpfa9G4n8apUNL2YK21r6hUB37GDFbDqB7ABRjxaTYfDqXNIVuPiB8C2R6Ptd4+N
zTKRbam3htlZMwfOeV6BekgVuhZigRBBbD+ujJbH8mLrEbuOMGI/pNAS5Y/UY5SFOGFo5OFr3yiE
BXOyvEB3xxyaNkLFeWcyRgvtyfMOcr38N+siXNrBOryIsLIepXi1dtXXW8hlBmAtpm1C0CQCqGPE
qBHFylcD5ykFCt8vQ/bWt7d1cQFRzOM6Kj3UkCk1b1/H84e3iHZUcuBcacyoD2uIc6R8oTk1BmIs
3iZH7xLvQm7GLRjlsZ3c7z/ccwaUpn45UmRylZYEk53JpRhCI8guwofgkMSgw8OxQJgGt52Fz1EH
hphvLdM7O/ZMlxA4PzzSgezN/OdHQRddLBVg//fRQhyuXdMF4kguuHfy0E1aI3E1xUD3j/5+CQQq
uIrVTgc2FQEbUciNFePTU5kGEMaYW3RZrjmXa9aaIeee+hnEQt3QR3w2xu3moBo5Xf2eL1V6TICN
vSRuLFjiU1itBrrGdk2k91X1jUplNM3vC5SxrfvT/ovB8uZyKUDz3L97bV5hUT0i2UDC36hA89Vj
jLkvEkfewCy9fPBREamPz9LK+ySy8vGPbcbc0HpnOqQ7tw+mb6pdL5JSI24YCE/E5+Y3oQcPWAiv
6oWsPzyyNU4s5xH2rjyrjLxMupO6v8PsvSaLZT9X405y3xhLLGe7lPeoJ351zWImWZYRVTwSaK1T
bpvHHuWAAimHZ3hcs0YMeyNvWD3jjUchyC2cQB2nv6j9PljZ7YDU9EHuqP7Pi9fuqynfuIeilEFG
uY7vkhoKS878FX7o/8yi9nQdSiBVtMLAg2taw7mlKgUbHLUtUZEadqlCRWVfAdO5D0fSgnbmav70
xdRdw5askxxal32nPB/dUuzvPi3NTMwrkSkP75JDDSmT5RDZM5Pw+8cUmRgQ7ZRbwpEoV4FjJq5f
+F1KoIE71RofXedLx++Ht6c77sYWS6JPBU5uSRPlwzgyhqWk4IU5E30r78dUXFSq+YNtX3D9v7at
PQNQRO/BVsxDhMiNCVTwaZXkpO7V8pwKC69YagoeJLX6tauXxozhMn4Us1fn/N4nEZepjBb+NkZV
HFyRYx5CJ12J4gFjmjXtkoy88hKFq/61UYRvUVu4Rw0NA3RWjQRhF4VDhZgR1lcCBN/THcttAeV0
QsKM3B6ooY8J/vgyZlihVTmm08P4KBL2xdsWtUHKZVojVKWN19NipDzz4if4yWxHeViQfqNta963
9USKPRKwogkgonamaOPiMRbWDfo0Fm4LOyG4tHmqyzBgFcAOPHLLKZ/AivhFsgiNT1vNisbFtOLq
DqlebMtaRngk5Nk7MB4UPKsPn1YLTt5PrCLp+gwwYNpKvop3CTuhfJ3mXU84sBTaEibQL7lFnTdX
5uoaV0fwCXsGcxX20fiLSkGDlrD1bPMTzCqII4KVR/tact96T8agCZ8WTNOaCWuZOrpFP4Nuu1zZ
CC3nMMYE2n5qAgkautawbXexgIySfcWIENspKOqJB2a8DNB1ecq+J9luvFIFUidIYYuUh4BtN/CJ
ElAdcDpohUGOoQHC9gP+8EAVUApOTFasQqm4XMLehRlfckogTemxTRM8ZUcwsgeziR7PRe/u7d8f
0z2UEeJmc+wUukpozLkUbb/6qCUhjN8pCZHLBpZQN0sXzWCMqP55rTCe39d7CfLBr16/33zIkjIR
pJH0vrObz84jJA8sDd3HqfOGlS0BYlcM5caV56ixM8DikVuTP5Ra3ADtAJhjz4SjYk+N0269IBXv
VN03RKCUhlNlo9tzBs2GzQW2YJwGBLjiktdvOOvlWFWRe940E8/H5IJhoaXUBvCNuvI5XQZVsAmh
IFhKd9U5O8e11P8Dw4ajLS92kFU4fUv/39RxTBlRPUF78pl5+swQWHy08pHXVK0pRbvAnmhmOkzo
y8x1W15+gKK2sQp6whRrRVPJO2tMa+PAtUHdU1P4nm5mWTfj4S2kv/sWQNrE6ermJ5nKQPwzlRbS
AD02JoUjD6nNqhSHjiNNzHSGYZmHZMKCjQsvWQa0kAc6+59prtV0U28DsAgGOlm6fYaIOgKkW9+F
b+lhrjJvvgloT4hypbuzOcuqpIIlCdL/onsyzEePqPg3wfF8Mfb6zt1mjZwLeU0/hZ75m7H57f7w
4hwMrwDZgNpKgHRYJrVz6keotylIUysk0UFqppJCEjZYy0yQPgD8XcnhsgfUfHK60xDQ04cMGwop
r78x7CrURFet3/JXdA9L8avlVunp/leaRDGE2cyTL/ueqXYG6kojgl+iwZ5uM9O3uTSriC6dFLkn
cX2iZi/l2mHXchTq+F6B3ofItDvtMLXLV/LqXkYBRXMCLSXzZ0QACYqG6sLtrt/y527Py++M48lr
EfDxD+j3DXOKYR3kDVS5kkqapc9yze6AhpFXt8RVYNn1OBUGjH+rJ9AZRRK8cxZIMW1pbEfPzbh7
Rw/DQ1/OxFobP6DwAe2AgxzAGnJXE0T5ILZVYfuxf+rmg9jdypcnlJqb4NVaHfQTZaRQeJf25dpT
xVKfmv25re8coKBl6MorhT73QJsVRYGcMYihVVsACdEFkPB1gxxws9ThpcAqeGNgbfGSgU7U0MH9
jK8ftg271XtNrmUu+KiXUkKCVPoCAOQTS0yFpzlzdC+65VN2OOKQyjLOJg5qTD5bcdXYr2N9KIoP
Ji6++JXTj3f/o04NxDnYQa4W0erUcE/h/+L2HIjGsZwQ5Xq8G+Vh2Gtg5K5euUDwJj1vfaQwJl5T
npKVMJRSLKzEIW3EOyCSNAYWX4Hkb/s9GEm8GC8rOmi777r5nGX5a+ZhRKGUr27Kz2vFb6CupnUC
FhP+qfCZ2SHeDxFq/g5nnakIhIkaUwSBI6dZFEXFDlutoAohUIT7keTGe5U6/MptmqpfKTK/LmU7
bBZBBuyWymUNSUoXOl9uvVRcqkMOPXgj45dU2HVz3O6pdokL7auES2O7oS+xJmPq+EqeI7sFr4Px
d1wvlKw+x35uILuXmOTSw3xFU4Elw93ab7NtySFM91KDsXaWon+DmsAg1Scv+LXMnvr13jnPomv/
VMAj7vZzRZttukTGjnIi4czy7zR8pYTPIrOumLruq6VtfRM7EVBknFbfTEJTyD8zOMX2UWF9SFpb
Xb12nJdpIwIkGmxKxvQavIS9juEt5T2CEEjM+6WgAL7OuD8qHmLEOYk8+1KDqzI5lfDtOXMMh6Uc
sHNHy5xMZH88I5SpP3+z3ZFySSFoTP+7C0LZvAb87Wzttq1rRYkGOYBO6Q32eLnaCsnvGaSISZ2m
u1Th9iDz6wAWzTYdxlNhjszV8e+GKbfgPY2ZhUuNu+aii/NISOLw66qm6pQm3Rc4raWylYBlkj0O
anRTSzlrFt79AC1XhE1R/PgbNwXC8DM088+HLZqw3esGKWLw6as2z/VeSm9XPIMwoJXGW2PCTb9Z
0VTo+Tgtblw14108uFeJ8BwknT2NNiWRtxiAhbJ+mc5OIruoVJKj35X5W6CMWYejHWxXF5CQ2VKO
iJ7SFMCpC1vaa9+L05n69uY3AdSF3yPwlWT0393Z5lMRf9qChIC3kPR9Ll8XOQ2tbYuWneADszQp
tbx1xj3gf3ZSqiBgaGh7TkdFtNq1tDHLjHWNwocmonhwJneQepVMxjeZum56P56HtWdzQt7X8mBm
uzT4kUAZOqm3T9GAf2N8YkNzvN6VMa4h7+0MRLUWtRgEAi+KAdutjm/buFKZUJgIH/aHZdOT95d1
6kSkN1Vq/yKquDTpmHdTafduHI0DZxwWCNAMOgH09nFX+FFr81graYARuUmjv6liuE+CO8KeHpR4
ZoPythgG2HVJOLfFhETAqtCCnoxN183ZcI0TItw8R7lDen+Zh4POUaBacmXNqzhnMesKyflUW6/U
ev+Jj03vVpviJvQ9lJKZv0Wm6RCkBcNtIL5xg87sYTAP2Kspg3WpHurQVeiR/Vz1381ESCBq6T1s
ST7accxJ+4sztJTWpfCOmhZJSYAYOfE1Mg1vPjTrRmeQ7Le2tnyhbHAYT/MUsb4Zm2SNkFpZwYzN
nNuwqAAwihx7o1twy5QZojprhTcV0PeYNeJDp5SVFAT0UTYqW/ibV/lF6CgglVSiCjcRhOwCKDal
bgm9NJx/xJGVUi5QGDd/FuOqm5Eh3g2PFmB9V95zauTyoMb2cmIbUn/vQJfkXnlQzdjjt6v/pUey
C/Kfan5XtCeM3HZqu4ikLJsWL1QyW9wB8H1RM+pFAZuXYCwqh3K79ayrwO1+yGu3bSWZmvJJuhtN
RHKjpgZ3aUcGSLJ2oMLGxGtINqzKNl+Ht2JPsB+5IvJEUNeeonDIlWthnDRUhxsagHONUdb/hdZm
aVV7/ZpeHPrVdqNTJmjNMmmL0zu5f0xm+RKggtqE1LHtjlCdXaKBxHOL1rWsImq+QZ9eTGi2RGmF
KeXOUwe9K6/YvA1yAlAEcS5C0jeNf/qTWvtVAGHymOrmnvAQE6vQINUJpIh8bDCQekzfxnntDArH
FKPRyC0LZHmut1p/bUtQeqEd6O11pcM4D3q3H6btSvEMYChf4ShHT8NTFdiOm8a8SOTeuShpbb3X
vKTkeuYesYGJbb4PvfJjCnNc+pHG0bMLgbAsXYTJo2CCg4hzZ4VpfLtJ7M1xSJrIpKJa6p205l6S
2aMjLCoNt/nBqqBrwIJFkLI1Lzp2OaB0nKb61bZlXuLZv+2x3gJNUqBb8aSg9l9gDm1aopuJPQkg
yJJDLRy5BkGVQ7TvAdhcmI6EGvdgAdTH1utPRgVj+69uBdK2YoO8xgzT95qeuxP4vZDGZfPODLHW
/LTfzp7FmZV0tKTfPv7Ccd7kiDLP5dUeSvCDtC+Mq110y2odiOo1JshBYYsXDlo09mIKp/ONSGnW
Esd07w+5g8oK45qZJW/nXctIx8fsisbhtAKB4tmsmax3rB0k6UYInYhkIV+Dv/htZhvaMvFr8Ao+
1F+0UEcrA8OJrd1rNOwDHJmV9QxtWE8fTa2ZcN/9E2B/tmszYLfd9BaASGk4zskGSBykCOlwqBTU
YOl6aCbkheX33LcpkgN8JgrBRIE5SnNgsupKw+AEW1v8U//YnBPdLQmWAXKqAOPpLrxxgGyhfqKS
8EL1iPEKLVwmmRp69H9BBTaUnt3WMIG/B3h52gEkmZJoYdgmSHtsoTorgRjpgOfJQl4EYbCd6bjW
6/F568CRsmoXN2D2fNW8XhwPwP27ork1TqLmefu9BAZ8gcS0LjMblQbsVaVNF2WP8id/Cc7mlDnb
6tSCq0C2jXBVePS+dCDEN6zWcOP9BNqdKEbik6ElkcNm/EtN9FfsMoEBbz9FlG9eTgckolclfuK4
KAqqaEfyGLhxOXxlf8FFaPkvCVkgrLJbsKS/ORyf2Lasm7iBYKyney2EkhaaZoXl6xUn2fGr7Ryi
nQukgzwfkzM6ks239A9ctcoeycakLC6AXBVIihPsjwf+qSoJsj7E7hMMzxzloFb8JPg8nn7hmBXR
v6dWaipTdX0ZP81BQsig6o9374XLYiVVaeu+RYre3bl3sqyCW/6fCCG1lQpLaZYWiIYUjO32t4Ct
Ke2gWhqh5M/aOe8DkXuPhV7lz5/N1q8ngwo8Ht8ePEgLE/80uBVXWozDGUlARboljpZ7dC3LE99f
9g0m4KZnEhjAMeSXv/BuJSJyYg2k+VEfqv/LIrSiEjAqgKcvIIq/KXzI4EI4LDlmTYTJlkyPbqAm
eOH8pMAtCb4hDGD7itaq8/J4QLA6oxmJgx/FYk+snxEYkWWVRVmQAaMskGSbYyFO9dd5qMSD/TTS
OwaKanqrKVtyJ6kNOWihBnGOQtt8xUOaw6mpcHCcOZUz7vcCyx9OzOZQ3h9d6M6my3ZflmSAsAm8
oEBYSQuFjAPgHfmrw9T21bLJaIiFni7FEO1etprE087OZT+1Nel8KkBpDF7vgnpxeNemCElh9FzT
3phUSCxfwUxZ70FQSW6uicgBFHpL3ERncXxlIPDiXzrSMISY8CSuhl0nzdlzqcNa1GZyU1SCkU/m
UeVNfbpZcZ2IdusoC3/gW1u2RtFNCvIEbMB5f2xO0yhKNwXxt2OXNP1q6ienrYpZalNjUPgq5+Sp
Kbhbb95wO5rqcW7d6O58g/21RN5RnWP9m5q+YRaRkIqFdOI+jku8KrR990qj89cQgZJpBpOgjx8O
Zocdhg+nh4/lVW3NVPS9IL/O7u3Vn8Xt4pMqSrTCtfzVQi6oVckLUv0qEMDxx4zqWM4ZJzhsgdKq
WfRZlTO6vZU/+3qIjjqjtbHFKHSu0Jlp6dM867c7zQk31m76WQ+BWRQPktJ1gcnBVzxWDXMgd8SC
I4b7cqOLUg0r6jeluXNtU82Zk5W2gWNBECoYDbHuB8Rcord0XV9A9ykzhGvoezt0UgK7kS3uUfhL
a3vX3ABpAyg9g9M1coFQL/U6WukL2OeyikpqhTdZG2kWjDA4kczloMyscYodl1agTi+Lo8cM1izI
I++BoV1x/D1RxqZ+KARay0/p2yqsK83a/OEfkfk0rIufCmNhoeqVzeswCWZAz0EmnGPB5oI8oKYE
GLBQhE6d6gM3tgmss173+r7tF68TJ4ROmDSeN3Qk0HfsvYgzs0HhKgsdxET2Ajad7WjcA5bTsBb9
ahvneyT9PyHBpfzRQ5TOdX2jbaCUi7AD/J+O22Pf1yvepY8q3jXpiV0RPDUdXw49TzMBEA744+F5
c0tJEBX1WOF/HU4vPAYE6A7aTphMVM0FIn6nisRzDefOYPKv1AGkcugz/dxUxBi7HEMwrVRhCyRa
AVQRU6x7fPYGWjyaOXTmUfpK0KWKr84Xt5xOqs9m8rBJBVwaoQEziIjQVUrkMeFW/OG2HJ7XyucP
h5Y+8Eb4Dm59Z/vzSkfCfEK5eq8N3InzANfnduLChQOx/hJDJBcazondg8LHddIyj0e7acsz4pNN
0tSvPC+S1zH4di4zVgJmPzi4MIoN3uM/Z7qehF5eaB+XEqpBafaM3z2feWD/VilB0Gz1cIWjf8ei
GEfUzQ0sKg3XUXk7SrMFN/qa2WcS6j4nBZOlM1gpPU3Ht7Mqr/c5eFSr44F0Z9e4VRGGp0I5KxwD
2I0EGX7Tr+cW1X+7kzxewkOylPQu4oRp2Ag23GMw+5SIjpUZWWpbc9182LMSOrFfSnXHXm2ZrXAo
7mpTKZ5CRGEQ3ZLkmT972eFEg92yMWmHd7rph/UKLN4TLGlvs70UayjOQNaY3DZ+ZN1ObwFc/ngz
mqniA3XiivYP+7XaiYzVs1C0/us5N2aTEuoEu2/L6s2T6Ul36xxVs2u3akjBT47+xXHvl8n/7q6W
GTa2KMESzhoFa/por0At0ZJwp5tk2Mqs7CT82hFKZfPoBbAkhwA+CoJ3Z602I/NPxh38CnQW3F97
uQR3ZBA8mIdIaWLmrhuLMuHs4YAar/HVPwtfH50v0b+O293/vYkdQoYl6RthG1U5GhikeiQbhYQB
o5dZJuRVegwH4UpeoH2Ga5RdMBx6j9X/wxe6R5cODtBc6Ul/BvsrG3BRjbMcZOlJh4vnp7h+Hjqx
k3LKBDh3Vt4kDAZZdsEUACvU2hwJ4piAGywFkFTucsPGVyiUabETCUM07r+/Vm+bZRUGRaf0mTy8
RKtV3bhXtDMWgfB6JhOPrsvtuKEsGALCRAX4Ai6V4mRt9BKM0zu+9VzP5EWVHDMjxwzzyrIu+Te7
nbNy06HrgTIojSMpZ48Ep6+0MjnNQk0Q0uwDb/W8VU0e2ih9QSqyQ3TxDFyNh2ev9HRzdQr4NE2s
7ZLH+gULN2BILheFtk9/LPtzWxaHGuvSx1plLmGkp6lv5OpS4zu9ADVHgxzev5rJi3NTHy4H5u2A
TkvzOJK04zMorKmYDBiA/v8vX4zFZfui2Se03Z9+wEEwVLe0WOalJ/mP9ExBomkmoSMLgG0ossvR
uwUG0ddmf8FlyTUbvpecQCYPxBplDlpdpsCc7KYZNV/8bycxQbWW67UfL97cz22QP3jieaKkAzID
wdn0CwPdUzvPoz+/cpHSCWOzTFtWoRAFXZZ9JKomcQ+dYfClTTFSF2UOwdhM2jxTlJNwarGB6sjS
x7m3a4Z0DWJSPicp2v3Slg+6l5+Npo2ePbnMA+lcVaEgm5DBch8dYJT8d8hedXd4Bgz5POxXN0sf
LyUdGY4rvIUop8uJe4HO7nF9UmRPivgwYhUDdBydBlGw1ujZ+mn6MmGRbq5wmTTCsfpDkJtVZC+W
XdkYyG0McIPBW80KRZpDwJtKbbStrrao/h/kknrTYVO6XzLwz1kQDRH/iPFluVBGVkkRPNcY4GtT
v562daGjt5k0UAKh4iw+P/v0zlOWRnCX0PS85UknLXHhJZLnMySOnGXHqhpRJwZ+GYS8Ic6Hm0gR
KsFYVz9Fv05gPbwqwFwOJtj8J0gWLdGzBaQWOghjSh/qNin44Qkc3EZrE2NvHlGKSnZunqfwd6fz
HEbdlqvEYOYGdEjSQjDdOctreNAQ611Cqnd6kkB7lka8NSsCconU0CMRg3ZAYwZOv9HZ5CvbmAyx
xqwb+BVtUyP6cbWr/rQeYU+DDX1zsw6j3OwhMjEYiAPWkxDNd0CPRRehxWpwgyKADcDtbjImdc2k
KoLakhZ8PGW9bdhoq/ApEMA2NrVa6f+4UpuXpRqhnBnYw62ZVd5lZ4DEvWrjkjWGrZkK1RC34cGW
4LrP4HEVXZ7byzJwxWTE5SqprDN2Lol/jnZIbuMigKB1Ssqavqlg3Iob+gXosCNAfZkaFp2mUOwH
wWy1rul323ec5By/VVMFtSAb3U2rT1GDDBbHd94alLt7V/pRDnZ3Vsfv9mgjv5iKgeIuzaU7FvY3
ml7nW1nXmfQhavxcrZ1rGoKM2Ov4+CMnVZAABRm/U7Dp6yN/pvnF+90wTHfhKKepkTJd4Ad4EoAW
1tdUaMo/xtIiQTXkSXWFkPurX9KdIWYHf/xiFIJpBORKzcSxjHgkzG7UeIASeZzjgwo1pzQe9Zro
4dpmRvw/53vJ88/2rAFCW4BQaguvB330nU42Vpwjp8hSeuBu53IbJ75oLhFPSaRwr+mLe5Q2UsRu
2kvhr/8f2cmw6yd5/LH28VuTMy3UN6aGi/uVYiXUtv8zZrW4DLWftccw2tW+iHhiiuuUnE3Tz2oS
UPPsih6BbBKyy8fc7LmY8NRTva5VCzfPcqXBOUy05RjOrGTeKMoq20IV0MUqHdEthzqDzqLvKE6m
TyAb9I0Iai8ImkndFNOx7cQDLdeSv5h5SCtpqlzqIhHisVu1Db8IEoYyoSGXLQOFj5CVrxPLBfXC
tpHFmINpFjEfZNnHVh14uLOWEuMY1ZfDKd0ESleCtzSpfDeRvOVsLZBL/99z6Fjkr5h95ATNCAAv
oexenJPy1CnIjmJqJXDT8ladWz2cJ5Hn9asMni34LK0RZiUV27O2fZMoeyMIKkSh4yBz3mUyOHvB
74oNLI52Q0ATGjRt8F4xQHZYdsLym7ggYqYwhI0N/zOvXx0CU0elp27IAj3/oQXRPZpNebxxREF6
rRcTZEb/IRwUXXu/hD9lpvF/L7OuMunCjpGMgaZcF0R3Of0KpepltQrDzc1zGHtm4qzl+HkK5rO4
P+unzkBr4dBBdnZRpoOGtsa6wuM1+E1Nvsr5Gkjruk63LWMLnEVrc3VfH3yqeB+vOQVdhIY/yyN8
1S5yuMYxhwuzk+ntFJzepORRRn79WfDIig/zqYdgSd81AKdKg6nAW9gGxMGd6/GS0ng/uV6CfzZ1
uUf/JtTIIk5Ixc9hvQOA2POcjhJYFvvYs/qvOacnW4OWEUiwcu5vMLydgxyw17zBaHTC5RtVY2EZ
ayG11jIHGxTGnyoJRmAYgSXVK8wFHvs5rX5YK5s/bH2kRmhfAigFKpO28UONvMQ8BGwfmHXekkjs
5cIJsX8OOWnfnPDO3tsc6mnTTtyUU3HsE8IzGhg/dGQjsbkK9bibaMdhVcAH6RvB8mFH9oTz3JWB
BSXgZ3kuS3KmZcbpSwYdNVY2JAwtB1J0c8NMwc33L65TuoiTL+Vz0oSd8Cp9m5nF2o/yAaVZzB6F
dHVdaAX0hlEBDKAnr361Talw3spzHZQifTNRK9y6SyJ1vQHRVHV/jVWFWtum4Gz/qcPrwTrzyiaR
Ly7umgU9irWH0HSKhRPklw0ER6xRM/ZTKy4ir9MJPSl8kY7LVQO9WFCaM2+tIMSK94xAQouVcSjU
x4yluCgIi7RDkTUEh9SOup6q66r7xiX1/N62aDw/uqONo9tV2bV/cVPSQvTBz+R+eJMNSOnEco1T
+sjka1wGVEU3lx1brG3grx/kUBGwzDoY9AdZ5P0XCj/ND/7ZxCQQah00XbDvI+YIDkU9wykZGnoV
+YTp5y7yqKm75sXqY5YPolrw8omSlQk1zxE2YJPzDDlNQFawf5KXvG75VT8rFYScsF7OGpCoCKNM
ycXc6bwdf3bj7m3eotFJiM+/Ow3ryaDJTmapHMsc8lqm725vGsjEjv5DH5Ehef10OusEXR1DwyjL
BeBQX86Ylf0LUpaQ370QhRgxBuw5qFoYaxGa9ku7bDjvFzo2FvTioGS3y+av0k1LS+LvA4qPpMSq
OcTGox6lyVW9oxr0lX1lTwZcdHw2vwNraZHKsDiZVIEAz25mdK6FLpTKRgPb8tYehTqgt2iRTv/t
ywZyVFNu+eJLR+LePAIuL2T6Np3XlxpzbDg0Gnwiv/GVNp+pQOJwR35qmGrg5WVjG+m+e1c6A/lx
FTZ5V15D9rc+uX2gIdwKR4EcI1k0hYHzqKMRPcOvbeHkGoiOgOLIUwpE32sJ+AJGts+xtI0zE6Y7
jDAQqolNEaSfJP5YznRdbMIvyFMMAVcl7/58b37/TR5160xPQPxl8TbNGro5jBenFj5YJZ1alnHE
TbC1/C5oCgb4HNAUvKbgTIwIKy6Ap3CgpNtTPf7207guP5TcKO8QVUVcixFElIkCEoSsoHkq1Gh0
MkETyQSg7FI94uw/NoJ4hJeDBcbqoja+RynWCszlJz8aKym5ROD/MZy2UJQY3/67qjUxMj0Zjuif
QYSJfv1kwTfov5lfL9jCBTZTqazT5RiuujCY11upL3A3kX25gOlYO4cKAPi2uAoCUha3XKeqSWnq
E7fdqV6DMAVsTP4TjMANr1mJKNCF6IbB3FHGTUtMVg5aNaSPqYGxP8cUbAsRmklBJONRAR5VFqx+
OQPLM6T5wCFPvlV4dejY48rfocXXbrbk7/ZGQzcroWn0Qx0x2kfbIlqB1Y1MOC+wm6sX3ufTEpP2
uSzr+n8ZzfpTn4TkE3HsfWO6ocZ7A4CCZGQ4k/LzMyzf7FKd2aooEFlM+up9TCADYFx6NdDTAuRQ
Mo81YSXRKRgCOQQHqsZF05VEVU8IbGctm5+74gB3FE9SsCQeA/bNAfFb+sEkkRqPW6ktfAzI8ItM
YkNCgNzqBQh7X6BxVKHhllicbHrss0v5/usDJ8Y/V6p2tlPE20a9ccJPqiNawZwLxT1SjhUKvfZa
PcYRJYBR2JTRWFk25iNkcRopOZ95bgPUcWXlFtwJog14GWetxS7z3+QQIp6k85kPgUIwdNq8hhlY
KP5sOh2uMwo9kEtNA8vEuhlOIVYvfU7OsrJdKvbvxExud5ox8Pd/16uAF7GPKgobfuBiWcgx4vmE
OeZAZSX8hHS463RCLPgzyk0WgzVHlkbha8uduCznX/rOf0z5keKINEjzbwR/+019u3aGQidWZCtK
YkCkKY63c9YcBpWQAwFZG/rwyctfITxHGAHijJ4SiK964J5fcjCdEUuuG5y4hvcWyUNQimrXBU46
NzMHrHJwEsxjqMlDV1yps7IwzarY4iKc4se9AtLs147CjTHheItzu54/bdZ+ePa3PmCWMLdXzo3A
18wWTt8Tewzc9PppA8JJUKEyauxhOow4RUUW6ZTGX+9gc97GK6iFM7iXAL3+sHd8UYdFwAqtRFJs
ppk0aXVSv3I0Z0txYnUz4z+cVAk75YCwqkhi90qdy/9yEtD2A/7YgwecjGWcwBuSzFzAUGOpqLOE
tNj4gNVjg1t731fglGge37ibrkIU6VhtOXpPEkpUk46qKA+mxuSxiS/5F5qGzMSrtU3Lx4dJmkVE
z0HjqA97R+vcCn9go5elqSvCYLagox4JigKbwmgRbPYdVEJ0grN/qer+pGjbFp9W49sTXKwn2GKH
hmUIxj6EMvaJn+xUfUV3DUY8XpbQmOSbL0Y3asspvhTK1QAdAeUVLilzlPjnWbrC3mJ1KdTq+rWs
kjApytVf5FlAlUap+8DImZa4VoHOTlDtjqD4oipY7QHlVVZBXXpidJ5QCcRjS3GSyAky4oN+zCwG
8ZqA4gHlWSgHDtbGYb/rsXQxOzzHFdb6M9FXkJRcJXjDvHmWOIbckCi+sRk4u7x+fi/KFN2h1uaq
IXQnKCvL6XHo+QY04WawehNZTp4rlI/A7FA6mT+/ekjDynebE41xPREGwRqvJYTEq9wfYFS4RfrL
nevASg+b2xYatP4KMgo/9brMIuq0VdUtmB0533KgCFiPtT/PZXp2uBSD4fYLhB4wtwNiYUkLbTFu
SpOm3j2ocBVc3ySeicXWwf0oV32hNR0iO6fGR0hIwKpxyE5xkVrExKpg/zc+TwUqn+DMcH2vnUpy
GSmFAH65yQ1A8dBwfoHTS8mfU9LyQQEO7PSLGKann8e8nE58TlgQXniEixfiQPgG4Wg4p2BqbttN
L3SRXtYLYk79Wd/Ut+iaN84qb3RdJIlZGz/gQZUcph26AWgzcXuCmG1QJjE3fpXl+vZDXcYvnyjK
0aZLpngImyLLTQi1G4xThUsqfg+bzzF+rfkWYqhv3gPqqQjXOYxtLuMVl3OJmkjUcQ4ZoT10thSw
ZCDktzMziyw/Q4Guu5XYP/0voPDVTbhwGzGjc/OFF+1eJ7H3sw4vG9z3awzrG+OkV0jatdyn2Lk9
j3AkCyLllXAevJF8Pqs/Ue1KUWnYWIqNsdFTP/eltrxefPBLJNH47+38GwGdY4J30Bj2Sx9/DqFS
EVT+pz9XucpY23HNq0rExr4rV+NABCFX/TTUNIjRTnTwlAB8a4nkCwB8KLxKU3GJgKYl50g9lDvH
mb6oDj1jBPwGcT8Uu2YZlatDG2nq3PJ3b8zikYreatmzMMF8AmHCs8DP5f0g9BA/J52xLqK7ceSn
nqVwCMDcSjkNa5tK/W3a3Arc3G/7cGd3QMMXGAAmifDKhsDY/RE+/I5WI00Rc6vVwkB/dY26kvrG
FVpLbPoTIcjy6SLP1Ls6wQL1yyYuvixnStkSVc8dJMbQ+FuH02TLRWvXSWLYkC39v0z531tSqxgC
2hDjpncKdBVykR+Qayg6MFKlnG1e5vzsaTSzii9Hl2o6r/Z4nMzKA6EsNB7M1TcBGjR0A3/6N369
UvEWVFBmWEMcL2DNGIADMb44BZBLDnsXn82C8nYdPOXoI7KKHy6o7xP1rQO/eoPA8vDkcYozr17/
Nt+Aa8u2HAGGHH9/+z2aDEghV1NHLiYDamKE9e4sHzAOWOdcuXWE4pH9GIk+kmvZVDZ9oIl59pVE
mRHPe52JMpwu18CAi6Zb2luh9deDimlfzY9NchTdsWXZB562uqJSSniJRqn7q7qSOOHcgnoqoS8y
5BAUkKYxtiSTdX7ddxiiIxy1JA1SB53sv/EITkD0RtwhSQ9cYxl4NDpFDmKzu1sv+4V8MYZ5jFA/
hDQsKlfde47ZFQVaPDVIL0/QHoO1rYAO0szwzsr1lXTgyY2JkEyZxQgaFazH6aEQqhiaykg+KiFc
p6O4v6woD+THjoZNcCSrR34XEutY3S4PCwSDupHt3U0Sspy4GanFFCYmPac/afN25kXOWHybSCv2
0bHP+qohkF5pMnB+57/WlUHLaH7NM/RtUPOvQ9dOk8tMLV1iFtt75P5VgolbMpKZorCqJ9sTZW4V
dWRLfETYYidmni7dwBg9kGaY7R/3EFrEBeaLw0nKTqNfxZbUIz52WZcRqgNnBhGe12NtLX52E0DR
5yYVJbuU1eTDqFl/0Bywkqyq/HYRpP9Na1SHV4AZtEGAglSSTgk/hin9f70sda1CKPjCuaUwpYpB
PQwQs6lbIsy80gof3KUEsXYDCkZiz/2s46m5dNQfp1bCd9JtWTi7+HtxJzKnx1Tkdrhr6Z+9Aee8
l40L4aZxaoS1uLic9zt8kHkCLXti0L3WcQ1PpyViBw4b1F8DJkeOG1lHCEtwCPrtnRJFsH+VL4V7
UuzvlY4VR0cBL6XvlHgjDYoOXFxXEQY+8LmYllywhE/DyUdMe0a1gZXjnNSpxRSF76xz7sUZqku/
RYf3sUPeTOEcpjZWsCvyijpthFqz5o+VIiMM9k+MII/nHuNESG4Xe812nAQ6YZUBOEKEnHToeQW3
5ku9c3CpV6v9j2JNQo5sZN2XctLwysD+dPjWcDR6+j7PihzrToJkWQoB/38lfXaCqqo9zR2RuXWy
VZzqjt9GEMuXwf4UEtZ6xoDRAFBUL+AFogt7XNHsSl/2KjJ1BOs+frJz/m0ULctsmv4LcjZg+vdT
XYgz+HiUmOxfergOhOYfz72+WwfiYgd8VL4uIqlbHY9KdFy/AD5UQ0G9oO+YzP7iRqnwydY85uvH
mETsGFCy8w8RcILWI1EL71yWvLlEnBDJTqA1zv19OdqYThRlQrmSEHfWenOSWM/eykwhY/XzJGUX
b+Bm2flhfSGExIbxK8C3IuzTkie782PRrGBCl38xazfw57lntywpMBeUGVpagoOf00h1/54vMoUm
ydkRLGxL2uAr7fWljzcpyFA/dxzysGGLhG6lQuCvnxua1WPlvHM/y8sXQpCCwrmJsf+r9gIeQfzW
y+HxfyObf1S7vgKLpGLq//8CTdx0NEbNUtoO3FDByI2lx23bFIC02y2ClkCdd2PgqYWtC3vNH2zp
TtA0i37vww6Go66guFMsbnFzTSuMJIMz4xgQvs8GUeY0J4SQkTKOXWMrr+Vv772HDNnFBXY6veCA
I9crbiMl6LccKLBnHwEl74WmXGFje1jTr5eVcIkxqeV4useI0lJM4fWC7fE03ufCs3/M9yE3Qe7L
agGmok6Sql5D9matzM/CdNQWXUcxor6J2QJvNcQw0ZGlu0ReOR/2sbbZ7EtV6U9wBjtoa12magBH
+S8TWra/kU6hhaN0d+kwVf9O8RI6hXubwckDR5aEqJnz6yucBZAGbdI0NWf/pAIwCz6HJY4vA7nv
Xcykja+2+YcuZ+3RnaMZexTkv9LgH4qq2kztbDyQbUstkNQAQMHshNnI86JC8iLRlq1uOisoSkyB
nc/x0KeYKYwa6CaIqmBeqVkpOi28O21H74wPjUrLCy4dDNY5458HKDD8yGGeOxTwnp4QcPlsmDm5
QVHItZfLfMZedFoRyhwCKWGCYuFFS+BUCuko/+4cy3p/XmrEXzIeEr9JXH+7EDGjAGE1CjLktLyu
8xCJ52rwYyjZjmgt9tps+bsnAVVsAWbQ/amKx9bqNo4DRMtRatcDoS0beVFX+JTgeQfnxkoeuoyq
YO6yugchSl+Z1+OSK5SzgE82J98qVstyC6DTnSNKPnPD7val0ZNNk8DIsESD/JEzXQRM0C5GfVOa
x89huzVELoNU6zC6n+/XB7Mh4UlDuEqi8psLLO/XR7T7nSdEBzfKsCpEIkrl2E8ywPXMOIxyHNWx
5HJQ/lAa0npDPidHmPDOul2PUgEwR4Et1AGP99G2Udo0Gyu5oafBdaR2UXv/FfpwGkGpgMYORSD8
EcI9MMvzY8WCbcwBv4rLhOG3hHPpl5hVm+umMwWqXl1u1oO3kdy6YbtpmyK19jdmSrTHtY9qO4fR
i7KYUZ0+Yj7c0jSpju0tMZ2a/yJ1mz5nsLKMvxz5RM/nQcs5k1m9KdjVga+WDMepx5/LgJ7n5aTB
P06HjANAls6oKJuf9tFYps4D8mAObC7WQSPh3tZtwcPl5gxNx/DCwQWhtD7Mf0FSyQO4bvW4wJRt
+laM3MkUBRkmFPhm2WcR6zFfzLcH2BBOoCbNNrgIj3L0Tdcr0j6cWDN9IoDPvnuIssH09spcHWMw
xfZBsD+U3yfDio3TuBMbAWjB7L8T8s4wm8JKUqF1YFpqCNUOxTz1EM5pc505nvapiPKwgSNFe39C
8bcy5LBLVy0ga1n8fEjv4JwMXihscCsf0fdmw269adHKD9ODGg64Uyxz3DmwRpnIvQHYFDNLKpK/
KzZ74q/QWJw+otFk8EPae2c2FnYDQlC2WOmV+76/+TIhOTB4euK7/pChcroF5e9crQdfYF4QtljN
ZkOfzerTI4baqnVOcWHwyGrNhN+oEORdhTG8lMlHETG8XRyM4GQAez7JWL68DZIwT7g5SF7T36+Q
G/xJZAsfTEB6C9wn4UeXCTexoRhTY3OpNSaQjixKdHqyOlT3yw3tjZQIDUoeRD+v8icBLrH8segl
womzIig0Oyyihmvs6oERRGlw7bE6JFIFntDjQRb4pHuLa2f3YeorLndnqPtWLxHph21MFnz7hMQV
ddG7rweRGaF86JEQw7HtHDeBfMlAygqB+eR3q68TGP6i/lpEbjNxbXnAUV7fW64Hz2kojXdsv8KI
SHBVnYLT8idcEMnC+EM7uunusqZNr0iCpcOzGA5vJKg/9P/JurwX+WisNNuWeiLZUZ9noa2u0ooJ
6O737+QcE5AF6wuzP0EG8TLl5mNfgj5NjgK8M8z4mLmesizHqNBVsFs8t9p3mjdmGphUXKW44jeu
DhSoY/TrkHLJ0YzQ0fsaAQ+ahmnT0DMPlOCxo+nrQVCVLBlNKbsDLRZWVTvbn9wX3b0NY98fnWkc
G6JihT9eT6+s2pwOyq4KxLteQJLVtpl7lecnaGK1LwQ71ofcfHnyMCCSAjh7Yj4wBQ0gHxvEm5YN
huupBVTExN5kdOJ6qhJPLq87CEuBslXIPr4x9vI9dTyJP2ZFZW+l10KfPEIBe8Aei12Ly/wtPNGq
yEknqqmYph7exBS5i8KJm0OqbPjh6DTOeIBHwFlt1IUaVgb8l179h4dP+/HqYt0a56seGqjp7+Qb
mCD6zGE0h1NcBrJCD0V99MpAV2URLqL4Y32IwfebqZ9pqNZKPUfN7ioNG8l1wprtMrs+L7uMj3Y2
N/C8Ot0DWPhTgbyGMUPGVae/WBy0eL0ikr2cyTiXBuYLp5fz9r6PXNiTSgF8PH4DAMiRWrind1p7
TN+mmaHf/qbZqpjIzGX0u4hvjEkciFnXayUezIJTpAH4unvQoqFTpsq8XLnATKx5aWiGu9v6Kb9H
txO79sz94L4VR9kh6Y5cmeEeS0lB97FzWJdkW2IRIrCTA6KI85W6ugS6sFtzdVNhA/4g4rxOlBQ3
CywYR0fZQ+1VAzCPSgwkaBcA9DZGnX0izuNJCWEs7p6ytcBu1Qj9AmhlqbDqyQzkU8/LJ/oPCp+W
YJxHy4EBwCINbD+AEeaymRgf1ntq0JGLlfN621F84j/FEXzDTIc7VwlKwUqa6pXdNwVv9BOWI1+j
Jx1oC0LBt5nl3cj2AxxPZy5fOsFDX0AwSaKHZnxSs04fgl/yPmpb/zwM7vGIE2k/t0HZOcMK77sU
jL+11WmPvXTn8hD8nwqwH7K6wZv0EG/6ewjH15hfTWLAIwYQrR4KKylCEDy0L49GGd1jEAvJvGkn
NU8p/WmHMxXCto+6CySj3b4nxmhTLOPn7daiHcnYLn6aOfHVLgDFWw7jwLgkXEq7w5QpZFqqBua5
gJfdmn9TILEVNx7+tmrwJNgDIulOkFstSbqKKLrIOEJ7hoOS0EWskRxq5mPBpIf3NMqZ9fs1Tsxh
WTtdrAZ6v7Ua26y3CzrpUaJ2mLNl9OtmP9MbOXc2csnq4yyVC7GKc5770ZEByoEhSH/ZnoWF6pZt
SL16O2M+AqK3s7n0c4qg7IZCHhRMmkyiFQZtYn7c6NO5NJOtJA4SQ69httz/6cTdWCppNM5r7AU+
Nkvu5+jauJ5ua7sdOsE8CngCGfaxFL3TXKus5mrC3V32vA7ifiu1jV/SOy4/VAhZm3OY8Mty0WXT
o0a0X+6CLgYB8jsygnE255nwshuXnMAh8SXblshjbRxV5crdBFjdPVtr0nTw97V17QCpIfDJ2FU4
8q9WGtL/0NdYKYwb0sShfker9MG2mFfrkxag3JiUhpc5FtJLPZA7Nab+2IhTcysz1dO7TAvTwVBn
/LcS2gLR65UK7Yalgzj3vJB8IaVQwkjdr/vCHAUEgfB+PUbOQzgbNLPm4Da0Me38uqzg0emU53/4
cj00m2MJdmJWdZEhi6jWaLJjug86wlU/0kh+yy1hAz46e6yuzVhMlryWOTG/mwKgzxbngTr8M0li
+usniLXCxp1aoGZy34tDdeWDr2PEx9gYb3IfQWt2iK1VFuY2mDv2fIY8IabCOYVgb0DMGTdLNYlf
S5dLPnxW7MT/JHljFr3VYaXeTCTZKxyn1Ph1Sw1JGWuxmHO/Dq1LIbsto3B2fPuHIy8Vmz3o7UBp
/HgEDnTBzgGRdOPlFfh4jFyW0bKwp/s9S13m59Ai0U/pYQVRwukvI/zbvKVPSWsixePO1A/8ug+F
3LxWNPta3OE/avdiohuHkJA37+a2kWVI17cxXeBc1J5jPGTn9h3kosBg0RSm81joG/a4f1o8fMAB
0DWYA8tUv3tyaqLjzbdqLlAKgeq9DXeVXJ2v6xVdPukPxvaDEBMLoITS8s5JL10toFfFZzqPY82s
9lVBhKE6V5/vPz11T5jRyd+Y+ZOcT+TwdhP1weEljhTDSPXEOgIFMukOKprPRXojyBg5Ke3URbtx
3D2AJyEzDnEVfkDRPvCBijhaIG6Y0Mro77Ffe16T3GVzjd8dzrmrRgYRod66RlRlI9J4zKPOL4fE
TNOkuzrGxSXr5RVwF2JkgVYGsqPz+bySpWSlI4ClFzEtNYP3W2INuQjCkNUKWQ5TawQhN3ZrryN+
l0qaEXUUON10xkQxLB/8QzZ+TrFUpn4BEwfs2cmi8PAiKcp701D3gAYXWABGZmUYGcvrHWbIFw0r
CZROF0ZY83sE+zwowCy2jPN3mveMooPMA7Dr2dZgVhzrOATLsMucaFm8snjPOBzYRe0NyU678o3V
bsYFfcjUk4P1hdqL42ZQb1Ro2ktEN4fG65+BZI7tgCnHyI0atxP+O1sUbyh/cdJsLYcwL6jp7TUS
U07ew/hy4Z2RI9kx1JS6Vm2mNYgNtmSYFii+Ja2u2Kz0wzy2TEcjWVhuMrfiuZv+k2XSq3slh+g7
oTQGTCCzwb/v5KP532qo6EVSI74SalPMpIUBd8AouGSyVRatKd0M8SbIh88jGlHRVxDPcrTwqlmV
Gmso324ReliF7/L00Q52bdwN15xEq5M/c6qKMejkOVvXnDO2sZMx5bcOaPOLSieO7cCitHJif7uV
hBR0tkBvwmYJ11Hy4t6jMneOeOhKsaSN4FGX8FbBY7jYahKJqgtn9mgbY+ojVMQ1pqakC4QDak3x
m5xmElE5qU7XfN/Mg1H/Nf0q82UKycxIs/RrvBaqV9RKUNnpT9VJEV1KSua+hV9rjH+UhmVZX7AE
Bdv6MUKBMkDA43OjA9ufTVj9P7ap/Bw6KePlPhj0c6e0tzmxrNtZEV1UvXYb+AZTTTYnt6bC+pLa
4UeDsAJWxFwA14Pws0ws6diPpILzQfoLvC+dYtbJIhMR5p5L4BRq/YcDnFK+ZNLOK29NYyQ4tZiy
zo+1QOxcgAT5L34nedfCa1BXz5n71Vv1rDqXCrjlu0GWia8yzJfcCl8GMX4DrQKcAKl1r+pDrfrh
ENXw5jk68hqACklbRFBboJUTApx2jliXskP7wrRKzhrWLdnqlcJuNLmz6HIhyP/7h8dnsShRXrXZ
o8Kw8AruFShKx7b9pFqKAcpIPKphGup4TpDLejTTxJAzEyTYOwPfVjHR3TOXp0H8SRhSlGgVV80r
nlRb2S0vCU8b7OdtPEdlUlS5cWH3pqcTlsElpT8Z5WBdFlgIt9D+e3j7jtgDbRQt8vHwJuiWBnCP
oJNmfdB/u9fGhs35U81mXh1iY3pmvFGYZY5nKZA4h4a/GeHaiuKTcr9EXz1BzoW72GHkQHADf11N
wFgbRJNN1C61/tDX3mOsOC6K+9DXmxRJ6eM7/z43PI8acRW4thQbpOF+TUIQXUUyskwd13PElOlS
9ZQxWv5mHtoTKd8fwyRm6PbcRD6ZWFecR7u2jD58mQAfqSyYkwiHSHONc91LjnlIjuucHb583Yts
AUd/OBgQA44TgYcaQZ1QoOpAvXpPtS6cRlLY4BbTRX7erFVSDHOA9I0GuyYb3MywvrbNPCC/6J+H
40goVM7A2+dIXdcTyAhJOhX6EfzaJkUihAt76LfRmMia1rNojF2eZi2zHBhe/B6zdALYRXOluCo2
KsMRSZD9rupWT8q6aQlosy2WfabB1kqzKYMT8NKkeBBuoYeOQ/r2upJi0Hk8wzmkZxI8SKjcCTOl
BLpqemzJGD3OHEqKalXckaFma6uHWWcHvdwHfN2RAYRvg7mp4QGEED7l2yy5yD6fV5PE6Cd/igDQ
cyKz8XBeK1YoXs9+tHDEl5Nr0qjehvWNuryymhf0PqOKLksZHYU/sEKKES25QkJChiUqSPkffDDU
KcE/2yGOZtQnf0CBaSG14ZSt3lE6FSBOptIPP8uJ/Rkf2tgnZulqQ7Ca+K4RLf6BbACQeXaA3AjE
V5V29pHw6HKFbcv7v5l5/a4dJ5MnsAHaVzIrdxGlCd+66eZ5oZZk5ukAu7f3FPZzH8Y5QhV1Fe7L
gP07uaM5yhSU9yGc9tAXIYCwLqpUNWk+6zShPkuJdgxP+RCtkCG+KaTCY5P0awt1FesDglXGvMLd
vfgAfA1QdjE3SyPxApyZHg9IR8rMJqGxD8Xg1sgjdyK9QPchDl+jcZrqZIUzoYV8DdyMxJ1uDXYW
jw/2imrKe4SKeBAMGHYfsKoOsYmdKnsnWpVg5v2gBGPwYk1pSZGrOXf5fkZRhCpUjWiWMImypLth
Ie1wjAUgiw9t5KZMwv5V/fFzjsYMHGk629lu+gHEBt8mfxXQWSIDyKMDYM1w7y3N39i8uBrfVdIr
i7PoSEFmmkLTTNuuTTqDo3TBJiQExkHfWIfisu4sHh3VAg/93IUgibBApDzoKCaqHUoohzaiJ4Hw
GVHE/eJEpl/pRP9xU9Xhf+oBOHKH5XXAW2hw92fmIpWY8vceaOGgmtp85b3rDTAibt6Z3NR2sDRu
ACynJrDXZNYXS+SPWiEi2uXak1XcDUQC6b/7QNswWfTXte+nib8wGy43dOh7dcCkaEytRKh3N3yY
g773JebbUpJoqC5SG+hamC0ivtJ8Rf9tLmHLtW8SWEoKBoffMNjH2B01DitK5WMTvPejVTEGS3TZ
wiR+QPx/ADeg9J4Wy0/o5GOljLycgDfXOWjGgOPgbxWQ70cZh03JFGkjHzsRU1uXwI5YT7qtv1YB
TmPW/5ZhCISrubn3vWTPKx64E4PfWsfuPokMTJb1xKT1BXciNdtOySgCjhklJBXiAkB5YqhICOlU
aTDtQuUMtyXvM3K2eXvpwGkazjxsJ3Onw6nKMdz70iNW+Y6DpUvjDVgw5/6Z2DOCX4ayv5XGZmV5
oY0ptsIjazo3gcYxkp9KKfcmdtkuS/WBGRkrM65z+klxytx6EKul1Q9chNUN+L6On0GjYC/IZ2F5
FydpS0/RnazDhqTcO3xnairjAal8ClqQUhYMjcmDo2osDn5jHR03CmkpA5KzX9ReGNIhhqiKYt2I
7L8Ci12dSl5zZuzhQUE/Gc+wnBBYDi0SrXCuawY1BBrwzUOlyxFG+SZir4vdgFZCB+1IaVWX7etz
0slgIy6zP21gZTAKrnV5BfncR3zmPR8kt2pgZg2DD1ODfDipqtd3ym5kKdCZF+Xfo0ACdaK0kfbO
1MiHys81muVZe9PNNWjW6S1hnxU85FtNTNbGg2A7XlwADfYynURQSqthvWudlcK2+quv6EuhCrHf
drqhzx7iDogASfUshHnBP+xs6c1Ch/OpSn9daolMZuUxkEEoyiajCiapCeEyNAXZYvW24H5ZnPZ/
H9toZFYRf6cQDcqHiBCQF6slLB9XA7Hu/5ybBVY0NzPQyZw+VxdfMu0z+ywfk/7NFhtHHx+1nW7u
0DI7bSQtyvB3PgCFHjBIXJEGZL3aRZid6QRScPKkSjmIES+2QSWHDx0/14czZkFkCMNFT3gbtvt/
S4K3qLNV0SFy4IEh+EF0G5npnpJqkmQYDHEnup1C1VHAfwwgzAjouoJ4Er000vfX3RT/BkMkMArB
gDlgwHwz60dihSbH3CgZo2Di36+hSL+YvARKrY68tJouo1198jlMkSXaCh/2sRInYXK1VpFFbxbk
Bn37IZmLfHYkXreIAvg463cvrHwpkPQdKJ7xf4AcjVPdVJJ92FFkmsIgY+jTUHS4f7wY4ZaxdTuH
SusGLs1qxTGZq+bdv44ruV3UNWCuNW/kAKef8mFIi15c4AA09PITZLAzskeVExfn7juCeXcFgRAX
g5nGuTdE5u6ac7lm8uITnmv13DOibMPwtX+gtwndMikJ3gTfxQKoIOKFww67VxYiy0wyXLTuLfjc
6KhC6u5y8hSdzvrnbmKWk6/mYd6n+/7M9SG9gMUJgDZ5xEthwvqC3foWOpDq4dQJCb1YHJ+tHj5r
UAF65wYRws6NZzaaX2tOX9Yze62zBGr6z5+cedjlnjOSMT7g2WJ2U8xq6qhXYS8jUijn7n88386T
oMEN0OIRtY1Dql9fnmcyt+L/7oyLWecz3t9NK3WcE/91R5FF6uqiqWjd+I8XqSUEBCq4/ga51TG6
1ekQWoWPybONPx9uSp7rW65D3Yd4lRR8IFRFrIDHgsgpja/AVMo2a9rD59k1I1WgwKz4O1EAMmUV
PTG87AQuitJlBDpNZWpQ2hvkwq6IUnzTwykosr4bT9dVct3lNcrIqbxm7wnRg7CJrmHM07xp5jDE
850cGs+mkX1VrEQD3MfLXBMhD5jiO2bEbJuJxarueUhzfgqhpmNaRrAxJtvwDZ+f1ao2mbUWbvyl
sxKB3fwVTwQizyH8kppAz63l+ZN7UqtxkqWUt+lDs3sKJgp2GSDGqNeziDV1foYAv+8D34UXNAVZ
3PxFBqwJPqWXV7hAQX5Dbli0bQPchEsvg+gCVmPKDvDnZpBBHwT8j1cBgdwSJSQn0RRH7e8JhnfL
vb5kPxmkikSXH7D7tdDc9X3o6yLTvL/72p7OMt+jHm33MgagjfivxjMdF3Otg3iTV8d7SUfYKz+0
wEajEMtupOM9DTigYGDzxgmU1wF4nB3BFAYRzhcwUgFDcQVuKsaZXvgswbM4crt7CrNvIjw8Yy8u
9asQw4PfYNWvMYNvn513WrM0EnVj1jQ9CrpisSZ9LQFOwM3aIxa3rCPKLvCIcw5GIttqctS0GeAF
Ekl7hOVobbwlYuXGZD1Veu1LJ83BzeF5MYgAiyWTOaU2DOK/mRzRcLE+gVAL1dri9LfuSd1TMdun
i3kccNwxt6iztrmoiKX0xntJoKHYC3QMyYtxatPwX1ZWq6yWR2Gu8ubkaJYfmbwDsqCUQry1+BSB
5UUC3SHIJsUhos+JJQyZ6xJo5jUvBF5cFMYACLbOumKzQllFgsnk5UB0Qw5xp2FVa6BQtzEODlc3
NrdkYJxgCXVPMZ27P0WPnO7DK3eo5VFthtPSeIaryOuEh/uw6+INjQbukq9k2Or4kacvSNMrZbTz
sghakajsdYvWj/I3HofGLw4yFTNjQ7m33ti+AxjSsdPeJz0hzipkci/mA71Z2cC8HOfh1tYDSmp7
IoNRkroBJqA17G45D3qj0PNFiRctIfPW+qWOKSigUhG3VHTO49tyVjN6PyXR0E9Mqdsin51G5AJH
Nj4r0aQqYi3OXvWFshtwtJif405t7PldCGQ2LGt1TkOwpVoHEGq5Q0WIiV1CNDCF+w2CHMmrdTZh
fGBJXE4s5Zo3vnOwpz/fkOJYSkVWmtPuxbKU6UkEVCQViU/CSCxu8d/Srcr19A5GA7AmSaRFECCY
RRHmqiGyhBb5D8bFojHg648By/8HQ7neNx7s4Z7rKSYOEXQqmoGWeSHBUVksmCDmeBeu1EHNgHeP
U+wXwL6sqsh3JBVmhznVoY7nR9Idtgwf5HU/+4Eduaeu0IG7xw67CZr/ZwHs9uyYmhI2HtPWc4Le
Bvg5Bfrr57m8TukFoKnlleLjhuyva8BR7tSlRQm6PiJmyZu3NcSL68zMe9jA+Q7m9uRoaw4OE1oi
zldeWtf8IwSTQayUZrTEUlzybQ44DiihIth4/OH8JwGsU8X+AlDSDaQLvlJSAREkTMG3aBpu6WsF
OpiAlwSZ7ucr+uyl+0W376X/fpNPOmz5ojvzHnZP8gsoFjNDcwv+1/PP6jYbvBDXj9d1rm6VrZd9
mpfM4MH0dGA97h8BaD4OyEHcmHjhe0qsAq/S8WnGCYTyJWPblZtvdvQWktRikWRdB57TzaCFwvY9
L1MeKeKPPbDFFCxo5tiek+xf5lmYV8mPk7yKWPDsLCwB0ahUdzHaXrKblyZNZV+K1aiFPdzMYv4h
poOAGAi9O8UppvegPS+rscuRQ1vS3nFS8FQu6TT1RyEBAAfaaNq1yBtWlqKnf6oIYKw0rIBx0eU9
mPoV+QIQ/l0oO0N/ZCcv+GpGxc1QPqPNhBxGzNPoSqnhiJtaMaCkUpmOY1xc7ZWuWKEs6AtNoTQt
8VZoY+lf5Tf/lyMhuKLeJZe3BAIog5ucISSdQbIPM9ELYdCCSgECOM9PEm1kHIMQlHz+iiQf38BR
f7xU6zY1OnwgHHAsU6k+viFM9861y6Xue/yyDegfPicpAWSNx7cWpLeAYOGYdAV49HQRlqHYFV2x
EWFppUZEXnuoSpRemkJIHBFQdkngGk3ZUjimLuYX503UPGYbuTTgqTGeWc+wetTlb4N4JWVBCkKJ
zShkj2Y0FWXYKKYcsjar/H/Shly80VxSOfxg/o+ivOT9KxzaN2PEnLjqEGUq4qxy1EkgKq+kS03O
HESw5w9YyvLHgywqsVXMUhUpKFBWUMOfW0YQ+/RXgyydn4Xs69rMTh5ocApoSLXvjh13F/PIxN4M
4jgdp/Jni7SVXZv9mP2DeQ8h7Lc8v3R3uASLVu54J/bM85IEI/+D3UiXL46GPDWc+wKyku+yEYx0
FQoM5c27vr+aTlKwntLJJIYBT0OP2rhKqwybChl+eGRJm9zXbed1kFVyojFgKtd+DSAKIKIl1RI2
WLlJbH8s/LZ/ftAZcl1onz2gl+zx4lEZUOnOZe+yChhS6KW06rg+aZ6ttme/Kw4OhBuyXCE7d6cF
O5OKAaQCc5lGtvwIp43SQi4tODAQ2qDxd77K7ZNZAyUqVxorLlWn9lPpz+3OFbRs+VHyK2sP8RlF
Ybinbj8uqLJZLvA2rPRNO/ZsdLEn0sPi9jCq/ICd0Kb17Wfh/POSy+PntgX2VSCT2mhpowvogBPP
ko8QIvix3ur1Im2g0sO1g3fAMEQqgBXt+THEcj/CwoCnzNN3ELVmpXr3y0x6p/HD2ZlNj48XCOzN
Ns3Jkat8qKM17CM4DVpJX3XzDzZK+3BnIaV64xxR9+h0vicuJTlaFYzLLam2KNsLnCtxoS71qFrh
pSYXX9BSBGwPCYgQcIinWn65c2bY3czNbGzJT/GUOBvYKigrpSDEEjbErJfmyv+4jq6Ucni+ope0
ZizS5hd+k/9Xj9oXveLDmIDm16qO5VBJY+khZOiRtUp9jxLZVCSsaqKLxT8iOB0HbZ8eBfhHCACQ
EckPo8YvVvYvMTb5RTrobu/OJTm9JwLhM+tCy1F2nIWms51PfzEqZO8IxWc2k+6HS7Wa2kiCZGmE
3D6oYpaVMHYo5HwsFARmuRWZmK3p5gRZG0RUxpGi4Z+T6AG/SkzDSwirX5gKk5JBVToh3EgOXwZR
gUn9Mn+X4Cb0oIsy5UsalzAn+EJyy2sKShIO1w6dYn9vSKcDKHoEtHyY3dz5rVgiM6/SkRswVR2l
nNsojZtWn/qddcXUwRJZhQnQoJ70AcmC5gDyM+d6i4gFWHC9QZ8UpVFPopbvog7kfOW68dz18E15
0eE30F7hwEdC9PDugBKwOQS2jC64oGG/s1ETYSez1KTy0zqzuX4TRhxJyiGUMsV1LHEZ6MxSIyc5
6dbzkPumU3ZRbyfOx8At6GxkYJLmAelFaqze1zyHbHBPAHw+UZbXIbYrNsk0TqtOswjIovDjx7g1
7Eux4dGw7A9F5/E5Cu+uJ6BsJe9lZ7ghw2jgGAMcqs0eC/Ox5BhQVWRU1UNpqMistK487wM9EHBp
v2lSKmbWyfntnqvvyihMttw4y33OLwvajS/S72tgx14S2K+QxGDdwsHkmJaHrv6Vs696NyqtRh+s
9v4a5rlirRAjsvtrp4G/TM/bEciJInj14L6NswA4VbElz7/vRGpxIpOVIQAbkTAsAIbO1NIDsKzQ
VYB5v/GMIWW1SvbGHAvFzqLaQazpyGJFr90svlyO7EgyHLgD9I9J4Hn8C2zTI/9HrWnEovxaJybD
0vj/kQTGE7DXP64TARWIImL7PYqfrtFdYFAnZ3N3+EhSQe8TVvRHhKoTRayGFVUmBSP6TJjnUGGM
PxuoNYgmjqpHe4KroKwMWsGfHccX8fY186jhZE9U0nfI9M+sFmn+5U6j/wbePWvxVGalTSqU672u
xST255SRhDUxzmTp562rl2L/ZT02mTF2yQAxwzuYFi7GOYgntLPJwFQO9WSB4VILzJBwnnvyulIN
uETMWfpktPd0jUF8SkQB+IaonqG67+Vv+kAO0lwFW+XOfiqExgemIP4rnUDikM3k29eZsZOXwU1L
lm/y1YVzA2AYpMDEFfIvakZVyI+E+QHhLWtdzK8GSjH5wo8g52G7uAuVNvdka4kQ9TnrY+t2vhC8
T0Jq1HWwaeTtzLOW/0S1bly2SZvFj0/HEwy1pTpzUqqBGSRtuk10HzdLWyA38iEkn2wHLe/fkzQl
bS+8gWxjjLN8TSlGQl16TGXbX6aB0lpJ4P6xI/ByUurdV1iKMet3limmBAdycLPbC1B9It3ju9d+
0JDS4ufIw659ihDyUr8FY77ISBlmmZFvYBt7UfuTT8rFU/5dUCnQdk73SlPLGQqz3lmtfvcnlbAW
X6wh3n2DcaefCCyu/M0T1uSLOWnfAg9c3Laq/5mkOwFzmW/0jJg0EDaWDTD16jGQ/GnxIPbBBN44
P2MYE6x0SemUwRteG1USi6LuyjVjbPqm7giZyijN4n599S/rBYJo9eON7EXWZ+3YS9RUhlnMv2CP
Kk26llKQl1mBbIYnLTUoNkyraRVMJgBxnI7PYgbAX6jNziPNcBMXsdQ/Tisbg/ac3J6Vqihx3asW
yMHcaiBVQRTorec0rVF5NNXJHc5i2X8TgMFyKTbwynIfaqTkcXv2gJMOX0bTQJaLLpbebJjRHM/Y
zo1OwG9qzxcHrGaWJJVFNgLhBMF6Uv9g4KPm5C3nio4U74E4Cf4TUj+EeZ2WEYx/a92ndR0FIR0y
ZaUeibKBEYRgrpaI5flENck5Hf0t7booalgPp8RDMKs2+nTJAkULtlQAbSwhEbl1yTAGKER3vjr+
QWVMEufydC0SEKuiXF6K9Cet2QCQ1WFpkWC8vBoTI5tJYm6UYs9t91sOc63rI1U90Afw5nHpQGCR
tneqyOLwnDPyvA/+Qf4tQ8jJSnoK03R8Bicbamztf190Dl79Lz3mjayONTbY02B88uNF8LeYtG8L
eX+403UCF9coREJXTJHolCjUEUz0O9YFY+jzMPlzmXu5x74tgKSbEf3zoiuhnyokx6XrR6KrW+g4
pAFfOUhj7GKLFIgIE3eR9XCguyG58LVvZ8Y/FiMyMGMt5LJhq9osHl1ZQpgHSL4YdOS9uHoelnuJ
7B0qJLV7jAhzZwuPD2FW/UmzqEeQY0NrvUD2arzQ3mi0V0NVXtXy6y5zTDDPVSXFNO+cwZQ0w8UU
v/WF4lZ8mnNzvX9mtzU9Sf8bavl6BVmdatI4GeS8WHhXklvCuQjxYYZWD/I9zQTnZD5wZ2AFU9Re
mGwceuW2tk6tvTdeo1vfECeVUqhOcwyhrWe2OBApLMUqmz+ZpChPsMaj2B2w0McKbY9uk1GWL4F7
jPt/694JAaeLDuWD3X3m7zqPQx/uhfv7bnoiyf6W2Y/JEKIp5zz54Mm7aZnK0BhV6oc3r6uxs62q
WWHQFlMJnxRz+428NZXZDJVHww8YEESGWGropmgFF3nHjOq+Qys6Xrm83xiayFrWXgQ/86wWl92r
dCK+hnxnX7QxtlAnXQ+RjEcYVamTrKzyhD3upolYPq+xUZ/nxYGhdWAssL4yqBK4dGUKZrOqLRB3
LrInuDEkhLJzAg+nfgxt5/k8SW9NYEwfP2hOimkluyWoszdQrZE8pnmKSS4i5VY+pJmh36QMCMs8
GcOXe4kYMu6f8+sjgfzi3kGAJU5uF5io3ZXXGkD7asiN5++SMJ2bPcWJtKpYQL3YuyW8mCo7ncA+
4jsTlQZnSKemUWRSVXrWWBvm9TlochK/5vgOsnp3/aznXdfuYd89xFvQveYr+kDzk5MRdd+/2wzh
gwUMrgnryFpVSPqo9FjM6gl/FkfSal7FBal+M/ePKRpechyKc0bkKZnvCRlursk6GnBn9vaJ/Ptj
cmITF9feiq3+MCLfXex02NXmV5MGjD/x00Zwg94M/qxjDI3usQ3Kzis7QvXFnhG5n3bqWxdcu7uD
85jWv8BJ9mNahbcOSLTQJM3PYybDQFmyH2dxyv5SEMDZgann9UEqEkaeIg96rkKSht39H7b1/QDh
AQzBRGnZbH9pPxSAGq/Y+AzWUNuWYztnqgkS25g4aRtF69ko9xDn9jLZxQgAKgroblmxOYPrz2FB
GlOTuYTSmgZ1y7aC8bcHPN94QOgoNjn261b09kyVvIL9pqbXYaq3ApiNowD9owt4Ty+lknJu1kMq
Pt7ElyQyiCDZTLkUQDSSMnsoDhg/KQwlfglLxIm23J0GGNWKDy7xWjm5dfHEamOftT0qJHIbvyQz
+ShMz2O+rujmz4/Bn8kOsaElPL3wfF/XjG3k9mTIsp1Y9PtkD0vjMyCcvNPk9Y1kJNcJ2HLdhLWO
17QYXbrGYw5CO+gjG/nPf3rDaRRif0GUTzSuTtgEAZssKtnXPiMK5+HpCRuxaBgf2TicVZIAqj3G
J4YsN1DC5/KHXXocPAWh3b/jOTReh4moDsrnMeolgpm+mEnrjuObLk2lYFqFYxnQ+R1Loo/EsSqe
nUZb7HDTwFjAOtY4uKwg9ApVbJPCJBd9DdNjoXWP5nX/Koe85YCpiWGoQAWnttDztp1MtgMfTy+u
tcOjhvx+tZouGvhcIUpIfKkra373woXpZ48Cy04oqx32CZPhpHKmlej59jHb7diai0gr1247k/xJ
6/SZTNdwsc3K6n+t4ZxkT4RuM1EezFb2QbccLNg0jK6nTQpVdXjZzLW9OuqPMoAHo6TBz1EdPyci
WTJ/5CCRW6vWG12yrhtzeuPYRGRRO6xpJJY2tyUIpWI676f009xtZVMsAt9zJWRJ+G2xs7amtPSo
IpGjhgOer90RQmChnJSMq0bloSEOwpa2NIuGItRgIedQPMdFO3YTDdztVY33BZkbQJ7ZVzi+KFtO
BnFH88cy72IImbtcum5qCbzIvyMuwxdKPg/nGG/zgBv3YKdWJoMqjbf5N9iRN5xpyUYBon+61sgq
GMfS8FSaVvposZk1Lduae6dXO5B7SFVQcmtrySSVeG0EFUeqaKXnwgoEjPhl5X/fj2lH6ih9l7uq
oHKqJFs3v10PPGh546DAFcCernTbpyottKvOp6VMBdKZ9QwaSJ2grvUOYOj0QWNP7rpHVVnHbouP
CBKwmM3T5jXrbYWigmR0SIUB5IEY9KxZPjhDbIFJw/qwO7/Gl84euQcKlceh00DHbPYWzu/W1g0y
YRJBU5+uPEEo8nqbr8lWK3rCEg5ds3iFRbG71pMpjsmq4Rz1xceorNv8rutIGvmg8vTjk7UQ2eXi
oOn+c+qzYZCY+hlfzLbUN0PYhaEB6uzFXCSJgWuwJRC+lfK83eVAbp5awRWmDyCDBwHCIqqw+K89
z7k8VqRHbNWp3UoAI0xTjhA0Htovglojlj1xSaYoefB7dIkC2aoGuQTrktSIlDolqwUK/t9W9L/W
bsz+nnOI+MhSzJLnhl6z77vzHIxUDimD/3/18F01Z4k2J0EsMfaw4LMEeS4SPaofveQxv+Wer3Ks
PCbU0+L9Ds38ekI82etYQmjubbM/hy4QvhiLg6v9A0k1faeFplL18EVoXe5cdpRuk8UmRM9esplV
le4WpZtIhS1f8Dvh0DP/sLhfeHMCXSv1W894TNsaxKZNEuCPLaromN0T57LkHoUI98DjCPN0yevS
+B24ArljdkDePk9cwNGc3lTXdQCgvfmKVsx+GDl9GgVp2pK7knNs1oajXlBWpQuzTQa9xIj6paAR
g8LCPBPEiM4diV5+WhP0u7IR3M3he8sJ/u7Nv+/pCirl7XZc2MKspfQ9aypI/cNZRr63+iQl7wt/
/CAPo0FBvtHLVM9tuCGimeeWbPe3qYM3RNzygd4JZPP7dgL8AuRG3L0+xtByIuhz3j5WH7qhxS1k
RrJEzpnfgoaWVHuxIvutX6G0RDJ90JzU75oQmmRehJncnxgmmpllqULdgoFtKF309sBaEwtnleJ+
oMrrMFjKTETqqdTomfotmZy5Clhx6Vaq/V1TkBK/jGHutUhfHUsfMfXYiiqpTbfMvpWLjQf3omtC
QubIWYsWqSdlA3KynppZxbsmEOjMvYlXTCegZxwbpHGvbZEPuaAkK+CBrvIPIZS3G3As2YKooSe3
AtHBBNhkH7anPhsD5davtdvzjos4CEMLplLPm3o+SZWtTKhrj+8m1Jwkz5HBY/PVagyTF0C3WB5+
7aejLU5nIghfsCjZwdOGsCHJPopwu3j3Y1w71HgwGFSzPmxN5TKhBFpZpciSvKPQOq5x2EEV5j3x
48Gb/nz5lK01wt79r80A0uB0jXRHLHUwJzLzkSz3Pu7bFKeh2HOfE9ZWOC476DGhPeWzbsC3XsNJ
kE8Iq5eoYobr6dA7xU4w9MirVbI/XdohdvVR9NijXcaSwC2stlKxn3soaPrNSlrE2bhZz9JODh0f
eaAdzQOtThiSqZYH+lWKs6w1fG2LdU3Tm4FntO7NgWEo6OJMHa48/rQXOhO6np6Y779kc3ISolmQ
V1XxYrNAyqLbII1OE8V8oTdfAqhEwe/z4+Mfc5OrdgaSSOLgMUFxPLGuOSQHaaVuuXxt+SgLSlBk
c2kezM+Rk5HgFx5+xFR0NmXL310srgTGmnzSX9sjftkuueo7JG6RJYEWZ33Hx1z9guxjLF1yuXmk
A7ADTO6Q9RY6LssOzeIUMt9Q5yp5EvtupRoKrRjEbPPSOQBnbES/rCbW2XUQm8ydjjbc+jAAOSOs
76NEtVAgx/NZTK0Hso/hGoZihvFyWytuZX6Y4RbnP3OqdzBxSfU1+JycmkD0HY42cej9LYqwM9vj
q6EbHN6DoLNRBfYBRH6j7C+LsV9Tu3pCNJIq01Eu6lJfvZtWVTUDAOEwlfzozheObOSUS6DB5Wxm
bPpxDwLWKSHbEUroI2rf0VG9wezORS/SkTaaeeQi1tqHx3ZCJzB4m+0ONQfD9Zp7EKchjVpy9Tos
/xq/fyb1DtSIgdi6ETA91ForEavyPIckEoyWj5R4XXhQ1b+itlL3WbvS94sHejNVjI3vsUos+Cuv
b9d3tw/qtTmxzoXzB2JUlsLatG5iudzRtxesSGm2bnw6ipH6J+Y3bG6JjAspQbgNXZ1Ujta+bTOY
8x354JgyhQ+4jDSjilFUopoC/yodNkNjzTa+BJTHgeKFStxcIH0oWQ5yUFRXSrcNWmBwFsJ7+BFa
b3HuxY6ike3Tt0aNXL+QKGteFRAI4bmuMTtTN5XrNnk8H7h1XHBivCNbYWhNl4n/uqN35MI4yGBL
9b1BcXGmWZfLnyElpFdurzw+XvwA9oqlgrxsIoO+vN9CFimW/qCDeDli1qMOSIldAqZkJiQYyw/1
NNqzoX2YpFfnoQyU7538EEBZA2i6FF+ERHOutSCjt7I5eZ/jcVBryPXrv0ebprdItUFZ+qm9Jd/p
sAHeK1NF45V0FGOr6+Sn1PVzUxvf+dYiEzo97fU3Wux6ZwzP4Wvymyvri8INJk9VhGwhd7qYnsQH
Ffx6uTez6sdFh0RYS8SCQjyAjMomXnC5fjnToQ8sBHntF+ZgRbHGWLMrq1OO/2a6EkZXoTsoIOuo
Vejn5ryT5fANF5QvtsC93EozqShoSHxqyredZne33uqajfRS4uHYQZ1ob/98Uhk35jIWl7evfEy0
GMcOH11nPtkGNqOWEBrvX+LtoJoKPx5BeZWhk8vhs5WGXuZXh1PeNcSIRERK45XtngwQErKrEDNH
LsW90sqgbswPgwLYMXj0180CbnZ1SnjcwqZSiS746U0NOObLyrF4OX9WulY9b2tvmef6QjMzWHgU
gb9C2osfeDajz+5n3g1kYY6beR2RYR+D/U5/PV0yzqkxYOV+TzAZ/1uL9qy3J0JTryWAqv4mFQ/k
iQ21yifBcj43GIbVpwsQQ5nE65Oaxz6j9Y4pISgPkhbIYIL+/WtqhCVJDhciXT/tBO90Bsxzywz1
s8/QJnhajqBu3sY9S+MFpcAcuHxnqUJJoe/uob9C9cZB4edJm72P0sltwdiagwS+ksGDt5wJUH4n
D91AWFvizgbLWsmCU1m9Tv6Gsi0FiA1CVZj7L1wPlnFKkQt+HqtdF8S9PE8IHtuBGCYUGGKRFm0Z
QgZ4H1cw4skzjHI09fhfegFH8+wQLc1+k+0o+tFtRDB6zyjqud6+xtQCRZNJf0yem3iCdFPzVZGe
Ca46blSWLbyH4gYj45+AzLGTd4r01GsVun1ZAaLcOYrqyoS+G08sOJtu12hw/99L1QTPNK/6UuiH
VLgj0S/iLra9ajUJbFZSKE4sQG4xUuN0aTzQccJGStr2wayDY4P0YbPkS356zsQbpNwOtmzwtfdJ
OWkcgKD/BxTB/k9491gsC26MlDCN229jzKDQ/Q/4zO/f5gHNBXfEDmnI9p6aXAmdV23vzDMTNMxc
ZPcnSxponXoqXKXo22QjRNLLBqDduFt9BJnB6/mYRjunsdsVbjkQlv5jp6V9dVhvOTsyVSpjXbVa
J57keKV0aJXRgjZy++AmGQG28nVl9ntF4I4g3RYIVv4mGXkx5UartFHbjoMQic8Mt5pLt9r0TzcK
013TcvInp8xssTXiVCweQXmsiA4HVqbjO6zu66Sz11mNSRhdAtqK8Uz+t60obK8iyxxpkEb4aMr1
I939lizb6+H3GkgrrLl7wS9/kLdXflaR7ECnicEbbMKHm+yUnPVw8l7w1YGEya0awPH9BT+CuLY3
OmleqTIObMy0D3/cyKpiZHkAwZiAj3LeZhU1sumOY3+oaM+Dtw7gANg4DUURCOSMieIdiNdX/x5t
kOwPPP2SJJEZWAfX+g3qejhfaXLfdaCewlvLtsvxIcmBAGQvB101jSMJ2gfb9SkEUAKoimaOcYmy
vF+UfkiC/6KSnyko/EpZwFtt8c0a/c0k/qJjtcfR3tczlaOBQG/Sdcg35uUk6hLX/eRHxjzUcMY0
DeGg8egbvJN6nry3J37xAB85uOsR/iUBunU3tiaXJF0BsggXlwjrvkypEMInrNtlVD9ndvJqc1KO
S2LXygXm3TEFfKo6UJrkQLE+33yPGMq+mDMbXVz2qi22KeMRdOANo/j3yOKpcJjcSPv9dR38JrF/
6iTVm4Xx7ocrizIns96CsEq4cU+d2V6RRyigqjoxFjH31FNykEabfmFIwebNIcs2Rfn7hhGOKceR
xIXvpjtqs6eTXEZ+1ivw+CV6DoBDvzw1VHefhLLMTZDWk4kmz4TcsP5aon7Jek35gisfv3Qp/MBh
24JWYEAiBaKhRQkMldMN5W6gTR80BtEwWVFabmxuw/KJI82e4xednoiBIFZqf0+78nkLEHWDOErP
fr5u4MPy/6AbSDGXS5Y34LKGYS/xucNr2wUAqQSAxRjjuLPp4jM/rSAS8Q14Bj5pFNCE8/CVH+Mr
er4+Qu66RrI3Z5vf+F2X6D39mGOCgonXCkix3ct4YXrJjwESu6tBp5ks2b3IA6ILxktxWoJ+soVu
lbcYZMGKjgL5rkmlKk0c6yDmeT0u+ngV078ElEg6Q0ffRYzdLEAavgpR18kgxxO7V78pHKmOECui
gFeOQhxZ7vg5gKENehqMHUn90zQAb/+NP81QEwsXhHwthgN5vJ6rR5RMr4OZmmo8t3mGkv1P9b8S
Ut3iOgEUdq9x1y/LTnbeYTkEl30x3rmFyblMm/N4j7YvgjPlE8fckdkokcVkRjgdbFdvVgAxyeUu
pY0T/SdEkTGwdqq4xBPy270M14UVQYpkPWlQs3BuW6A0gXG5tBX4ApqZ/b9sri8mLI1wVN1b28PT
pQrJ6PpnB8GqEc31JjWFRkOqnbrJkyyqGuBnbWy0vIbjPk8WI8L8MnKELKY5Eqec1TCnEyM68oeI
rTwKgiq2ZKMcrn1tZzNNqn2f0ftHyF+ZqkUVJ7U3LnlffuBwt9UKrqAdl6n0AZMFNhg+mo+XXtvz
rLu+zJ7mgJiCamgPRHQ++w+zsHDN1nchbwA65wso6DKUX83lra//uvVj7WLnGgfntEtNzcQdxB++
k6G117nWohxJhZHgwZuDNm45Udqh7IRwGYSpJYjz/+nCsRiX6+RRHtoDzN/+acm9JXDapEPQHo+I
6j7xmz3vKfHYZfoEk7WnTDtVgHVtFtPTBMeGAY7BC/O4auVzTT4h2PT7z3wFYmVrNJQ9nyzRfAoQ
d41ce4t4ujnQaVLs17Fm0dKBmDH41yhd7mSo8FpcTgnHq/1zrvi1QV2ugcQfrFDmnJ4ElLv1gfUz
DGgTAYZ+z+pbk/hQ2ISfgDXaL97+uoauBabrLeoZJPngYaxyc2gIJpxC8RC4hoxto9Xp1bfMN2J/
G57Q8UmEnwx7w+NZOBtkFVxrQzGxyZboYkGy11zuAXM4J7DRIJ5A7nCTPH/RNcuUIGJqVQ7UUhXE
BydO2Wn6+60Yv2chV9XIcOLMX4nBBNcrM3W9Xp0k3eFEOiFYbgd7VNhgT8FiTVZJAzkrJTV8My1c
2FKCcthFcUy8uxZ2k0IoVABfztFR0POtjXwbrSML9yUoKKb9tZm7ME2l5wtJd/jgl0ErUQNRCcZ5
i7jpb0Mr41jp56VZ9sPmEOA8dCoVBJzgbJTi6i2IpbS+reckfpX+MXB6gd1ipLK72GTPWJtC3akG
XczoxmuT28kx9FFnZIBJc1Jk4yylFX+ALMDhM4cyv57x3M/UBDB8E9H5dCyGi0BK6xuZhDJ7lspV
PYctuXk5q67i7kjstNtGYKcokH5SY4LxSiTn2M3QqQNA+HQcknNvfUanzfMUBnxnEGnV8GoirxHl
klTKmnJSpqbbvY5VxIry/ZIiQFozxxPUcQ4ft4UAvNLPXETu8eqQuVt6G+aZ0xI4yqqDeMnFYvdF
axoQu3L7RBdMjSe0gVZdjbk7WlAtKshwa+jJse6IewSKcq6R0PLrUUl2QYP2jPvQrYfz27aO1cmg
g24WDnoi7F5WcGPV2g8DsygwVB3L9RasTkKZgzpyzXfvXstonoSCt87TRbpuqCcb6SGryrvhrqtN
O6n0Ggl/mLUN/+OhrfV0uzz+kwvHBViSAHetrWEj5hHAHAsvoE3mMmLoEj//Dapdf2aMxItZAMNK
ObU6ulkQOLOwpPFQvI4hBstlO8N72hDJtgg2KJwHwAORU+cb3kCH/XCw4+mkRl6b686ZRiVCr2V0
jjsEMd6zQZSKDLdcE5mvesm/baIGUw9NT14Ap6Yl+yGquIPipduPHtWBIEcdFZeGlYyRlVbk49SL
NJLpUtvuMRji4FcOTorvpWPyq/moIiOpWbR8GQMXW0FffiG+S/045UJ+mkCrNpDiWQHmVVjZ/X6i
HEM+tT4QFDgNwt5HIGVzsegqNltWECujzrkXscrRqOB6+eYWtlJmkm0zPKuGMCj/L4W59uqs2gGY
/+YYMdbtbDUmjkJpoujqvlRVc2EqgxgqGF0NwJgeZsPA5voBiODPpDTBtq52SBdvEGFLeDELLdkG
Hnlksd+0bzyLnHNxXnKvz+jG6C9ZIzdg8HMyaONEsfMVvVi+qM+Yhh4TO3JzeF1GFmavZTo7iSzs
cus1znRrEN5YpJjlHeCk6xI2jM8ci7GJWlBTMQOysz7gT+0EJJQpl6DUOY8fjFrTGGY2MAM2Ga3P
Sbc+gYJhTLXEJnAx40afw6x9IgiFEvrfLSAdy6M/E75+vCjoMXQFGQkIzE4f7zlzQaJ9lpEAkArj
+BVQjh5UuaO5OsrKYfAwOZ2BZHjDityFhx4vcsEIxObDeNZwVT66kvGtBJ43OCze6wFfHWh5e+HM
24iPKBQ/FVvP2AfckNpz9BIEGG6iTdpkq89GWIhVz4Qsl4JOYZbSm5d8ur/kYsuNGekNoQZDgE4T
uyP513QP0AwIfw7pbGz5N7CGqZQceaSagEaMzD7lmFd+jKUjt+XJQuIOS+LKsgGRKpWEEretAAyg
IIg+wZ/PtL5A6iraUokBMQCN3OtMzXsSXoy1s5FsAY4Zy74bvDWbOABL/LSie2ELuEZMHg/B0rg+
NtqHqQ11FP0whYwBuGvLzXrnnBg/iq7B+IhvwJV0HAbpcrPrN/l0ukZU0y1xC+qthg8UTk1zh9HK
q7FKeW4qxQ7YNlVwC9xTY0fS/3Pn0UNvyxs//UFEhG4ekHACdPRDCYhkXY2GdwejbJa9e8HqUsO/
WCfF0x2NKqczpnqqWG6YqSzXEft+uy3TAUfmvFbEB46p0Ko0+Y2dUkPDrpU5skPdy3KfUuXxU1Wt
DRx+dg4ibf1K8YshLissQQ6AQixPrOO6oWxT/cKnxHOTTE6SpREqRrJ6ls+2Iib9odpAyhv0U5fG
c1g4GJmcDhBAMotIcpizwb1rqO0wz47mnXdbZqFzyVa44UycKNL1DxfYZByYlCQWwankKuENJYFj
zo+nkDS0xg/85oOM2k21Hv+OVIbjVpfPYcNJL0eqsVfw+tW+eOyur2Nk8FAxZDcuILsIHZAaQWV4
BkcaU1jWXfIy2HZZwUoI9fWh3Xq3LZRhauZy9Yr2V99mUtDVgj/c/bYM+THl6HBa83r/XSfoUHaC
aG5flI4iPG+oUf3XRO7sn78bTfGOkW/mQG+ho3BzbFrMx6QobZOqtd5HSjxcHoYbY35+3miSb6P0
xNW6eeZxw3W5oyQWmuPalmOFD8fKfjK4PXJDVkyXUfplJ4haldn4J4pNbuUjlNBOh3afvDx9z98J
QQSoRnnwahKNl3rEyUC1jctxCDGriXHk+HbOBhkoUXXPe9SP96bATAp7mNVOqHZ60lh1HJw3ERP7
zn3yBwPF2Px/Edr0q97QhDKxhhl6duT33UFcHiLoGlNWKpPrOejng2G6Tt7jLfJvncLheAvDcBCN
kYGvE1/lWuklsyaKHdZ1K3guS4ZyFV3P3gNXo/IUGQzxmpFXIksQiK+Dsz9mZtKfXnusFwL4vMTg
CHSX8URL+mPwRAnhE4FRyTSsuY4bKlULh5fRUZ6yaM0q3juG5ioIwElgJyGvPVitt5homvy7gmiY
pTTOhkDDbitFinKQfdaJiwnm7wQvS6r+F1OAwMujXaW/OtVOuMvlujngEWnN30XCUXi7ASaBVGeO
fVJplmO+1OOzP3U4GrNymW9BYPU5wOvBahOEIIGDotehTrboLHs1kfUwAiSI4tXMTRLB4A/jVigV
H98F1WV+XDFFj/IY5hes0Fp/1JEDrHP8zGY7OUDsEc+NekvJUzPlCu15CPdsS6FN7goCH9lY/TEv
A9iZnehqYkCGy8ZJStOSjZBnp+3pj0cfO9irHuARNpsC3FhPJKccmX6ALZwb4wcIo0yX83D+o1RP
QMdsOrYZ1WDfouOBLsWZkWkFDsHVQwZkEZKZf/eHxlizEQ7m96cZs5IwBN5WVD1/sI42P6r4C/Hq
27/cqdtiNsjRetdt+WCzAYhLC/C0YbleUDf6Qr+w6YKtNnoM11yUtNs/UuGpYOKVSWgWd3HDZVnl
oLKygKdt4/3Yyg11Eopug4XvbUKSQ5hPIbMjXP2YW0wYwi5XRlvn2A3uN9DMymZwgaTPiPwTiAGi
TTU0/PjZwdJFRphuuXIqqPiYrb7vQqZMDWexKRJaq+0m+3QUIj7pdTUEXZ7TjyUbOHYM5TYnjX7t
650lhOCAdYTL93XY2pH/lIYAhrLyzaTbwRrySkhSpv1Ck0bx2mjzSNqHyIj8OJfcLIKkOOnP0UbM
l65P72R4cBm/06cL3M344zIBQ4aA3F4fqXygE2WiBxeLOWxdIfshEQcmKeo4dkVx04dfPTvuimhk
i2SmksRwBNmFplTguk94jwUPqRmgXZsw+J7xjlZNWayXy9pNCgUz7x7CW9gNwy7eMOYTzREuPbBL
Wl+HcTL1O9Q+XcXO+DM33jBHcyPos5CMGzKawMmwIdXUvOzNzxwzpxrmWbmXzG+xwNqF8y+Od0FR
lTa0u/m3mFtkmOkYyZI8udGIk/egs8vGLb+d72mYdeOIJtXQ/4V/H6QjGYJECb77yYzP9J+Q+86U
Ca+PBE/IadcGh15l+jL9zHflOeF+qU/AAxVTR4iITJ49vVhZqKQOe+MT7oylXLDozrrg911Q1onH
Lit/u4P4K5eIE6Fl7RdjTKlxitORL2G9QGw/+fhMnP+1ZopbCH8kjPDIFExsqzaW5MzK9Ccctj8N
GPQU2AVBLpepWdBjsDoFDstkuWVjcPPw3GzXLvqSiaPzCzZ4Sv467ZYhDIcCtDQhXB9zc+zGLT3K
9HAWV7StvHRjVb9xzX9d/LkFiX3EK1w8vBOfU60ugqb7bIrNqaVTt2wi63G+837MY0Wm9/T1Y8bG
qH1dNFSCsBcZtNTSStcVrudND1VsVQ54fOOfahf5F2AixTuYmVpo//pTA/03vnMD8rtU0/SNMNQ1
5dvsMbKlSqLNhb12+zPiUlVjHAaF8CKY/F6zoLy/61txS80BkTbsRytMEStHPy1KBjJ+89S8mnbM
D9Wg5GocLJaoN8ZUCEm/VrYb8XsIgbfTViCoIvgNkrl1ImpTXKJ3PffZ7pyiN3q7jfvdbqUtNRwH
70ajl275Xkz9u7mgRXqMw/WrXwlyR771T66FVeJrPgr4AWutgKSJnRGfITrsx81lSKMrBuvIL9c6
5cBoV2lNd9F3qcaAwpE6EvrND50gYlF56zG7nqvgtgBfCBLI+C7+C54+qmU5sk3WVmFo3LZ8iY/4
EJNPEl1IgwskiNSWuYPJn3Q9h81rjQIRB3LzUKYAdul16wmRcJQmWGpQa5J4cOHL6MuyvprLmHuo
stlgHrmeY7as30orf1FiVoWUze0O9Su9Qr/MsIwuTfvcPVaa7ut6vuv1oDB1ZkfSf9Oc2FsBXYCI
3CXftUGmuc9AqRe1FFbFqnsm/G1KzQBZEdadcnGw0PBYiurWhRhidUCQzNdHWGz4qvhtk4uN+m2Y
t3VQ7NLZTiaTUzh9tFSK8FySgC+ZZ3Z4ySyPimT/IzvlIqPZ+M5VcXOBcTGpSihQx82jedJeNYNr
TugQWh44SnXmJRWlGLJoqJr0TheBPG+YhYY8sigmkQNwNF2G/26XnzbhdkwEBL1N62XhWv1lsh2I
z/wVGRJn259tbxt3puhdkOkJ4hARY0LGn/B6m0GAN0YMPfm4atFx6R+45fz9Aw/Mn8kG5v1cAFuu
KLCWtGe0MQhz1pdk30qSBLZBLVPNgu7fwUb6ATn/tEK+cG0Ni6qmF6xsxm9J6SnA5Nr6WXqvQcfZ
Ugpkhxnpf3xbTP3PkcPL7nEwC19WfovaC2BPH9VKIgXwBqwaTEL3FF6M+gcJjtbb8YisugD24cDR
mfzItEeswG3K0ZB7Sdp2cGtxEMH4XvzEazEm05gwWIh3Viz+MiYZjy/HwoW5ej5pvpyhVo/GFMIZ
R2NaIsehJsCHoqljpIuUIyEBa8+UU/3mn0hoKapSBRL8LzLOkjXfsGsShTrDUw3sxzSP+HrFQ3mq
AqffFaXUVF2ujLu7z7Bk1c9V2WIN2VavENU0G+p6mfBZhKAqGL6cvS731oMkM+ZXFkGkf3BQG6gi
QCKzYZVWQUVxIC3VT4i1VDX4gUPZjGwWIEJVRTGSRUO8RWRkM8tEAIjHcBJEUQPVfhKkb/9S2JVQ
PDv2s0PzXwBnkUc+WsWJqzxlvfdyB53Mj3mHVMbmdFJhRWlUlSSMTqxS4rIvlt22BdShhCMd/p0k
m1VkArJVGAcH2OXy2JrblLtkHXBX5QBbrBSFlf7vERIzIOgc3kC1rmJngUBUEv9PEykQPIeai71P
593WkYRxuHEX2xFU8Ipvz+TQ7qGPyVHzlnFf8Nt5kTTbEDf6ZOwOT+XDq5FIxGNHPJT/vqSLkShb
TfjDIOicylpd0cSOaqjOEkbQJ68dT66cBz/oR9vnn+V3ApJU4aMRSQu7qT16zmWpzD92j+JJERIp
dZSCSPquUzVjGdcgLt5NxgYDdkq/Noe2jjyy1Sr7vIOcScwGrVbtE3jdut214O6+1HJaukNlfoel
tVz0btd6RZt+k9kx7OMm99C3NmxreiuLNsXL6dp5o/Ms18Ke9ML6isg9L3ovD7MrGrU6mc0/0gfD
FWCsYajaizJc0kzcaEmd9bvM24xHZtNnuAg43mgz0U7BvbOX3tK/y4supSdlpjsZb2fbMui3AGX1
wCJUIynfrE8LyRH7Qi5Cb5HoiS2fUajGWmnBzK69WGBK47Obg6lxGyiWQbuxPbg1hHMA55rUIawo
HQrkgyC0+TGJhF3RLdEiF1H/FF7RfGjHwk3wzfukuTQS0tIc6kHYPDxhzzrSCmDjJVCDFGlUepvr
I1tQ6aBHaawGu9TwoSopiYXF2IAlQPDKY69KHM5XvpM5Oh+kDrvPURSeCnPV18iNv72FEa4koyrU
DOliyddZRtPt6DPchOHXmbq0431q+ZOAdgYnoKDsc5raS/kr+6/H8wQFwchqXC6tOkGzsHwPWVKQ
N6jnWZ4ruQjn8BnDzrQ+8Mi5ZzDjVcZ9Xc8aWnLRueOzHr05Iuy00g7QgLYMJOBNa1sBxe/S+VPa
GOQwfHdNYbXgLKtLckPGbvnaUFHWcDvxPpg9Io6RrznitWYyzcpylAKmGCO7a6eJ/ZaCUSRz+55X
jVpp/ag3NcPkKB3mvHeszd+5g/JUIfdjofWzfJI2eIIH32GRf626JJXzfY1Kgl7Gvj0VoIzNTVIl
O1v6tL2oC8IQF29idcrNY/ILWMZpfaAYuNmbZ/BV4ALMhk+vGORlYBpe2g3NdAsIRMZ7EA6xACgz
SGioJijizI96SjX8LMV5Z6baWafS770w7/JrI34kMV0tr4H57y2SM+R+k+j8FwkdZM5GUo2ciLft
CD82n9Sl6DlPXzph0M/7Cf6NvSm2Ylry84Qe6mNlsAPjFdRygzpgPn0utuzVzcIubq+LboEI31Mq
qfUPQRvLvKpVrZ332Twuo7Z7QNdFYhu/C3xF20euUg2zlUzHV8MFQrsxZGa5gXPcZVn640vgCwhd
a9q0HMF5E5Suhfc7AyIn27duMqOOodC55e6sKNYCKK70PsDvSR7rOk+/AdZd6yuwiw2p8bvm8xKb
m1Fw6r32+M5OvhNIMKVNyOj4zrVT9j1qGh25GK2lZsz0dfMf/HF05Q+DOmImBoifBZRUBx5C4AW9
qf08LUQyz6g3A/eSoj1guyOBe4Lgs0VDOPv07JFJx7uF3IUHWyxyU+f0gDGO/k52r4cTvXL3pIHL
V6haZPtJ/eAg0gxx+PuPHgeTTBv6+0k9A/HE9+NaChS6pn1B/9UywmuJtwANsFRpMZXfXrNL89+d
bihMSHHgkKSe7Tf42PKom5hA8vuOrhizu5oDxYp4jwKSeOfe7KNqtaDFyaw5nMeng200SJw9Qrt/
kCbhWo0jhczPic9sf2XScf7KeL1BkSUFo+Sf6SNDq7KE9kFJSjkVo7N8oRFDXuTKG8ImhvvYUb7S
qwolL5rifIWgTKCIkPh/K1yxYve5y0QfT0yE4gVKW1x9Z9hVyIuIMyhrBYfHzvm92SGCSaQRN03T
FtsfOdbiNbbNkvCFyazk6BQsgKnbzVxVSHf5KJRsbu/AT2i8CV1jb8RKJZrrMTcXZMXQUDGz02sj
I6cc3dl8F/GZSi5FaDMooojTjo5c49ku7oAqOop29nMb7MRBLP3NdTolFc4AgBLmwvHXtirTWkhi
TN5ExvffK/cXneWjJKGwfk0NlPjfJp72To6G54MkmalxdXz+V3rIFWR8YG1zIU1pMBaXfAcRv7I8
V8xeeyLF5y48Gr2/3hng0v0051pswNOMULCBH7oUS/o+ykgrGUNhlnhcsPhPWW6fRoZHDU2Kwnfe
U0KHFZZfUKcCZY4/CODM4lqg6WahlpMw4JJHGonTrBNeRsjuunxdKRJ1biz+OJka7o8HcU1mGfVR
mLSeTNsymyKwqi4k5I9HDUWyM4jtcMVRCYukVldq4M4iaDZGIpBXuEctTc+0hltcdCYD8kKSCBDK
k8cUFejt1uZuxvVLUdlzGlQfzq4MjNmsZ7gwGwEJ5Scl5t3uGOCxFTughKtHsUVo59PrYF2ZphfN
CQir85izuWVHjtv5+LiSWLMQI1SefkbXH2S1bsapbhyqBdTEbtLrKIEy8/gGMKaWg1L/ZrXx+rHe
BVIikI5TF/sKhhNHVwbFebEnQFqUFjv9H1PsBzjIVTa/5aAtbupJSHdyIlThGN6GjMfACjwHvBef
QbOZZAL/cI3/ABHmjPBz/DWGPdq2AeaLp9npI1aiGicMxi63X9dTd4gGZZmX7LqcX3Yukj85H7nP
h8qABPxk4MdebnQeKyUy+BuxJCN1loNOiI72yGpltL0eeiZaVBS3LFz75foAgCCFp4aaUt2T5q2g
Vz1A/oTq7ERtA3L+XcJAYJ9Bj003qXOkR39qxaTk6pqSX595umbOLD2roRAb+QILkU/H2MT3MiYu
SINLHsjWjHVY7MFoOFBa8+sGcDNxGzxI6CIwMHlR5VclCb8oQBisBy2n18RUpXqAkv3ipuXMABXD
ldFxd9cxuQh2vZz+6BE6BhPmzSOQl0UyqIcwBCiav0xu0YPdnz9Ve0Q4ZC8dKL18IruUo9U/t4VW
eJFPsQVhuPkpN+ZhpUEWRe2cLCf+cAoF68G4afuhKTfQVOrZ9ONxDKCEr7a4tpbVWOUv7rPoLQBB
wQsfIToWGWnxzTetPcDLdqNzKX8qvYcGjBp1JxLWpaKQYEBk1nKh8s1SFxmx//YOaBwqYiGfLnO1
+qs3WXvo7BLVaVNOmXt+PsQdpjk0WPd9TDSGuQ+LvkRCNgeVtwwzWQ0lar0nyEe2aGdWKMICjR8b
l7mdarXDtfsNzVQ6sQpv3/h86Of6clRw1EvKQ6kGzZ97/Ook9Pydeq3RLbOredlbSwr/Lp1msZb3
ftbSFGn0UgyV4ZDyfO5+h4oFkt9gP3IoyOEJW8KsV8OBGyOaQnOk10r2dI7cFwfK1aB/oc9Y4Wuc
8ZAmN+lLfcBC4MC6L8cwbztkcfvw+DJqHvt1rVZI9R9OcSZRVko3wnJDanT7QOzOt4v27SoQ/m41
DI1LSnCRduG088kLsfMSYk3Fv7n7uDdqnZ9xB23tt9E0bD4LsM1srIOCDpDnGJ0Xudc/96vjVQLG
U9rjcHIy9NuiE5zpFx8PGoqarhv5IZgc9oUOHmiMfw/RHu1d6aw8+bBIi4gUFRtOZNDHBeMjjPva
BjKwgwH+u5z1gj390HoCUlunY68oYF0ntR52SppzyVpcLP3wShhrg6WV7YkeixoqtUphz+PJVw/v
o8qgyJL6uWwkkhjP1qdYYAJY4/cOLVD/SoEecQzGUTghRKUGUBAZpyhUsTM62nSSXPAPxpDajD9v
4A9m24t6GMzR6guk35k9IVACPYqVW9+y8dnl0ymwMahEOBG17jSKTrZuRLGfTWtfpBI+EsEGVtGe
9eRMR5ggJ+LP+4vbTQIn7Pe6B92ZofAIxO6triEZ8hIdtdj2sZIAsGOVRqalONzInMaiaLcHM/R9
8Nxq50+BZB1ZPSEqNHICWkxUWfmLFaYCx1JNEHeGXlYrXXsV4jXUMa+/Rm+SX6ysnkjnIaqy1XPd
bkqy/KoozayMe50pR+cl8+Ng83/bqRxHORH/56IvCrB2+Vxzw0/yxlTZNREwMypA9in+jE2Du4M4
XDea/vq0puJNyxzcaV/AAWO7x16zsemY8tRQ9g2dO7YSfWYM5lirzjaW9x9Ak7P1vD3oI8l73eqs
+arrfHcClUD/9JZHVariH7EpuD30MiR6bfYVW0NlKvw7Fm7Lx1vMUanu6z+Ww3dYQoZRCp0LrejT
m5pA3SzSk6qIpjbveFc0Wkt5m/VP7GdkiUFearpMkXFjRIyuAgd2PQcnLl6BU+VO2PSId8qvCuGO
3n5Y3k4wBDw8mIFwpGUEhsOVYWndQYEhe2/Y8Kf76Xl4hrwUj3sKSlpsPWc+HZ0YJhdP+SaMzjwZ
s9qQFlBnB2m6AfxUHR9C84hlyPgDIMG8pl2sB03qM7Zr7rukboOijS/p3oMHE3Al3sDU+ynEf6b9
eM1aW7nNUNHPMjVqHW9SudsneufG/Nwovn/dDgihLbkTKygkRYXQ8ExnbkC7NGYUVyIDc8/FrrsU
MVV6CUJ4jtD5zQd0iRQCeYM0kDFq6sbpHZ0ypTMurdpjYWTIiudKEEVpH26A9x8X7W0GlyjacdVs
Clz3/LdUwixrSwvhA8nxzzdKiBHdkN8nh6wMN8nm3UZPDhhEjtSr/cSvjUEFit0cTjOsI0i1ghKj
TvqwTuxIvKcqtIxs4btNQudD+rlcRMrKuynlTTOR889V8IRpkxguf6B6H51dyv22dxeBorX47ZQb
4KcBP+ZizZubbx31xGKnknQy1jbpSaVxhAi2rvkB4Ptu1l3J/2BUUkCJxU+GTV0f9FgWY4BUhCK8
VB/hlpB01UwUe0m4V6TxUJjTwud06PC0SEwz8ZzFrAtTHO5SAEATf+5sryzstxTMSAgrcz4En5lZ
GV0qk+xHRUNbj7jbb9CZDRFahQMhnovh22nvRgQIW0Ggd1LI88IBMS50rlyhoHnjJo44iTAPX9c+
YOicLiFoZYEk3iBZMDilqMiwsDZD2Tq3u4KzuM7LbCLOyIOMaJG5UGuuQnLAAAB/VZyEFCQiiAXV
zcZDC7f8Cbp3gEJNXRbWlJXixUbylJxLYTIcvChOuxHkvIBURyVQqqt8UxAOxJ+BLTXqBoMROZHa
khZYecr6IXl68uvAJm8mx0ADVfKzDelvxeHB5+qUNaCq6nrhBH+US8iHrizJQYW3MjMs8e0YNKWo
S6xI+w9zVniqwvz7oepT8YnvFfjlIkJ6zINRJHFj3S/4hjiOlHCKV1c7Yw9stRNlUtPuL6jk+PLH
B9mHVr0APVluprd5f581M5kxEKCgam/2iEle9MkXT+7pCuz1axJF1NxSvQNlC1NbmyQ5fuxj3SEt
RpiBNOFNBLtszHKLIJ80/9hYf3KM7c9lB7z1mnlG46NsuGKSrW/yQ4M+gez6GErX0t3BSvi/AjDm
VLIE8LfRQVKrfin/AkSmqMR3er9SSoASodA+iEcaKhrcePf0p0S5Fw07/Imj4PSnstI55FRW5fCb
/hiSICryz8wCBDehs8EshMJ8GWpm03nB37siGlPcKUq/XlRxtUC9PNNgqfwuKRBN3m8y31tKMfVZ
avT4bs2QrqYcMPvWh7JB0GjTesH+TodDOuPpXJVxkSnNN5QUWxVbSSQCbedf+OC87e+v/enxzSQF
3p6sZQn7t09x48PorKqa3c7XYERgF9uZjCrU6DhR/T+KgJmMS/7LtMLV/Mwidx7WRjQ90ZtL0fnY
lLtAqrcwq4umx/y5nHuqLp8A7f0JAvoP+/Lxz8kyForK9BtbEjje1Xz8w32fh5qcddsbmP7CqWJj
iMviF/Pi1r7piR2oizYIlH3qqmMf5B7NvD+EosLl9gwycecsKSIaKbIs99xYbeYyJ7v6LkbwgPV5
2l/sJdTURboKa+CDHKXQjQGanpYSHX3iovP1zFS9gjnUjFcGNfV8pkAkbMSudu1gIvj4vlNrmmeV
bqZ7Iks7i3/P9384FrRmqqvKKera1av6VAxR6+yiiA/6MVIlk40R6ZfMsmQtQKz3NP85diSArWqB
b5FDEBE4vNHSSSsfug96QAToAyc4+KhaPHRZfrJgrDIrbEYtARLY80oLg5Wh+AmlH4IwR68YKLBi
lhfuRZO+cbQ5MP9putGDf0/ul8/ddLQtJALpLxtALzZj7voggjLV+WIA1YvXISRHh8yeHAaKLW0O
XCrnpP84qCVLUnaPngYp8WOf4SCWWafVG1e8h3IeM01LgCroI242Nuu14On7Ju2vRIhePZxQSoWf
M3s+QArO1vFQUX34CcxczDYnAzLtds6A9lFgkrAp5SqmyHja9HDJhZfv5rM8mma97MIleXFXJ5Fj
wzJhRvMeNlfy8MDDDVP8N3N8GJEwnKULAc8d1OOu4yH7UCajpbWhG/c3/KKS2yeSX9rIvdChas0L
0G8vHw3C8F0U3RuxekYLpEXUJXpg5pa30HHGfertSTbBEUhTwOpQ5rneppUbURBCq/hu/J7HO/P5
h+q/K1ba1GcNTQkVZej8kgfpiD2D08FtR0V0dEYml9s83LQbp+KgcvtEUBP3w6P0mkhl39CCnQat
H5aBsTnLS24wqO4Yt1FR8WsMft3wD0kZRhGE6KtfmayLdfLjrXYZDiFgaB433TMpxzGamXxGmKES
K19rVITX1D12uxnAOjZX3B7vDOdr+Qj4ino+YK0f/ac8pmyexzAk5vYNlPxOSZdUX2SqD0mt3V84
RdtHv40VuZqAf4yEt0pR1W+vC6rgNHvvDOepFSbzVG0ho5bOGWvV8BnzjT8u5O7LYnArsad3gHbv
22SFms97Xr6SKML0QfKCJ4+NjKeCBEK7FeLhfZjp/KJuPtjSm2WPBdPlcYvPABgY0MXABi9HjORH
byvXi2GyIcNnBJ2PDN8RWk/TpEajgwDqr5X2End5NrQ/3/DN1yiLg77fzUT5fWqoJn7Wy/SFZckw
CLx4cZO0B8oZ85Iz87qiOTUEnQuTaEAUo12BstsUFvwZMBNrYCQsgzMJDGukogu/h/Go7qfMrulp
Jjk4qmf7G7GDIjVG88wFfyvmktHnY5s2DdA48NJIuvWiwp+yB9AkGCXb98xY9LCJ8R7RoHcCCYbP
1KeKSOAyrma+sSPailuPZp6c/Ds4KDt0PHK3U4jB1RjFGCQ9mWq686FsnOcTAzTS2kR6STPvKD1B
Qr/1eWrmz0mM4Ad6wP+gb49EAKEGYizxwhnKb4FbxavmoLeBhrnNlg8Qt0puexbXCsPcGCjEgWN0
B0z4v/eNWNxtTe2PJqbHICIIWTDn6ZtG2UJl15vlACx8xuqXcbyYgG/qWgSjSXUD6NCjjsJ5V1RU
+8jCM7nLFBVfQBYPoBMoGm51a6bMX/eDx5ZfwXL+BzCkRLCyNQqRMLdRCSUNJ7/cac8P6ZHE5W68
YX6yojWEC5frRG3t2olOo3yPw5BHDkTZEwUTLiGovA8QhH1N+V33yi6BdOhRkwmQ4X1pM/skAyCn
ItQ9J1C71OPIipLCifoQs5OEz8qh6I+SoEtdJlp2+asFJ7Nyh0I0Likr3BjFNIJBHRlWy2A+CrdV
ronzI8LmsSHWm5i1i/JvEtXwkUZcNcifhCF7ZAlNFBzIhd0QFAVybXtmWy2FKjKAhDplLtNbHXIi
cMJKh2Pw4yHokSWsA+PuCSQbp2SIikawhi3+Zj7E/0inTXbon3uUdo6ccoX5ooPvHTcrAHtFTN+q
S/arJ8aINiIVPWnKksR0xQ1lPWNZqZ/Hi2B/L+1UzHfjNaNZ/vppJ12Of88ygPNDLNdQz2AB6uPG
dMPSqCap6tOBGP7xdrc+zOzYCp/4tLktisE4X7eBfKDV/RTzB9ZOjoUyc3roQzJ0E9tPx0MIkhaI
oiKqFD3QuW3PJguOe1Wrc/OMUZ9QlfctPL00nuWILj/SME7emwTRebZ1ge17tjOqRYztZEZVy6DB
iXMaccQMM5JYd1HYk8yeDWirKloM3vpY1++cAabPv5Tfk/+034kZ4/XI7hV+kOm1iXpXRWynnUwY
SaIoUhIZ3zOQDs7hByyiRfZDCy++gIEye7Ru2ZISdjD2lju4+tCa0woj7npzFRpVdKL6Qra4Gl7k
ac9l6mLVX/irDITuh/CBbbRigut2Am1nSnQek3Skhl963UTUJsrJJ0rqp5iNLbV4pJU2XUYTeyiF
/0pKsSwy7fiSZOx7mgSEuDVjfnttP1h2shEco3SF22UJKg/MFoPWEe9qHdVVbvkHRRPy0dsdmPdh
QDSyomy8yIeb3JwIqyHPFfFSiNPMQ05+3j2f1XdDq/3IYir2SieENDCwT1KR7BdvID+HpBIJIlnG
m2cWxV5b+zqYaQidBt97caYtKjfBgaY9s82MneiGQ5Zo7ewZ82CTIu1cEWOt/gZARHTknySRikfm
+Xe82ndcrVy9rDjyhVi8eWczoWOLNoNlj6AaToM17CZivhvt7N30N5qifbDeeyi9B6Qeqil9/DEo
nPRNz8oL02T7svXnxgzTpnDBgZkum+BABhG3+euVmfzB+lAYK1O3xbMkwucCeCzmeDcOPYy8Q7NP
Fwzxn4SmTg93gKctGe3+zaz/be6FsKdtJMBdZonNLbRj6sO2UpxhPCk3EhZWwzrO9QnwiGsZz+Gj
+rlIKbaH/BVaKju/biC0g1UV6BdgKSmfLKyLY5fqH6aJyBcPvkZQZCeG00Vmtg/zp1MEyKUdDDAI
MSgB135JiEGx4s+vhbMm8kLLAGmFqNtCRA1YB1RpbxyzSDkdPa3DaCcShk62gqxiTsPQybNTmDf2
+/1D+yIlAxPhoEyP4ROYpfjdpx2Rin/oGZ3HVbwZ+WjV/hAFO/ndLtKgM/RrZfhidqdpzyzdogZL
ig7/XVQXJmZWfhRCR5F1HJ8w3gDWRLRWKdQ+ctka3sdKi8HuYUWVu6Jgp2PWrukcPk9u5dN7dIf5
lhb0qAfFV53ltO178HtucNBe+HgIwR0w1UJ97mFFABos6jDpGDh9EA4sGc3xrnO75YWB6Y91CjZz
v+lDAwPDOzbv8yODFYKTPo8K8GxiyoAeXbbk61LA3X9xsHVYNww+6GU3bZL6HGCeIxYxx7N0/CKS
yNCjowgr2NtOZ1e1el9OrI7fb1B8/UiUKymyvwjNC64GYt0J8PfiZ0IsWYbtdRfK5jVT63r0ajgk
dvd42TnAGFmyD9aDpGyh/ThuZkc5J5f5SRlNbezI1FlwXS7bDxZrMbUilaD/TV71tK2VDd+7iBQ9
jfYHPqNMMK6gB2AoUEd3mVzGDh1H4ZV8sCIxBS1hin0zKj5Lz+vV0GTUffSeSbNdvnSl6d/S2+1m
f/AhaegZiD2WAoRvIORf5zaknCw7a37rrDFRNXUyCa0WRREQ0dXTLRUxONZmO1c/uCObA2UvIYEE
lyBptX1qop/X5yWkfMTlamffU4gc1dQHheE3dFhEpANS/I0nRTEXr/9CsG5s8ChaIa4nKkp/QU5g
Mz4s/3BqAKxamRNYTupgFgIRNwQDYocnuffzXPhwYSPdsO5nQUYWMrINiDQdY6gD4jEe4ZIb7num
CMT3haLOo0i1nhvz/0gJxf4MVYxPJTvrv24lgkg7DUJJuPSKAax1vLGRY/WkrAnrKMT2LRquIHNt
DwHugmRYzr4l4shNvn3iJNwU7/KzWYRQ7F7kqlAZgeoMf/rdgpLVt1P2OnwdU2D3ki1Qj/K6EKwn
EyN73SHBhNZ7vamUQ2LGyttMwhfnzjhjTWKlP64wKDR/iztG7J0MFmlLRtRof+7HsCNhBORjMRLm
z+l3bFHOIow/9ZoBdCFE0jtlNqXPFJXusLhs158oiRbWU+FIJpwWVxCDUPY2hLP7YUD1jIYa+QZf
Ib9ggVVcjt+XMgPYlb/ooaWLjtIdvdgDvhxevq5MeKVGIddTxe3lQILaD7m38+xZxG5LAzhFqUs6
ZyKYVg6UYxhLTJ4sX+M7L01sZUpuonf6hMlqjng0UsasK7ik1129eogBe0qpA8wK0K03M6hmA24z
lhiI1+JF66POff4kxQjBfmRb0lCPef+htU8gmXB2mHBai8w+bBjjn8Mj4kdOjdc9v2PfRydAWuzi
KaubomCNnOM7U+ZIZh8YDVxuJ7wJAlN2XYj5gWvvGM1DdRf1kYWNbpVFQ/ygz9VHVld8VSrmVtz1
rR7oE3OcEVPPwbogvRNh07PhOGlYYiD0bEv+fynqyufNlHC62scoWdjKeumcs/v4uBxPkx2BzYni
x9TuITHFVvRceY0W4DK0eMjlk5bm563evo0wK33nWs91T2bz/8TQR0cLnKTawQFZe4egh1GrJw2m
IlQ8DCskJBbpeOZcSiZ3sbnj9XLxtTPUwmHSBOtqu+4fAAUyH7Jj84Cnvgh1aBcyxEBTX3xfgl34
I9fKCUH0HVMnMemweSeDl7eR31H7DS3fb5RdB+AzqOsb7t/BfE53Q02zZJ/KA/IAuZV8xaCSFZHx
rKB9dJ6y1t8Z5of5pziHOh46l+2RP68QPP4al3iGCrhedjNdzCzUEoHk7susTUp2K0QGj2CcdkOX
cFtMAHigxRssK7TY+XkKbmLZXFoa7ZWS8vpgp+sYDHfAheNkksHqUsLGiaC7y4wA1q7X4ldoeRbH
KuBEe6Y/8Jz4DcrDIL0SdQRJiq7/9KM8RWqIJXegOyucUAASWwvM6eqPZ+6biCGh73ykWUPOpGLE
taq1R8buw9fQK7PX3OHabXI3GYpReCtUkAa+R02be3+YyUFuoAK09oSgHCfwpipV9iTrPRVgeT3Y
TwRQTWqgR1hL2MJ6aQ/f3KpV5zfx8+C8hFCPiIW7/JhuS5K/fL0V7egJmXaM1ZCW1sZtE4hCH1TN
wKhsWVyxOjVtZVAlaQ3LGU3BG0YWYhI6xSsQPAoWIGaq+VCwQ57HuQniZgPxspFAJsmKnpMl3lPN
xgDKbSnMRXks1bRV8S4ZjMJmgieCAQvpHKxVG8NzHZP97B3o3C/3pJyt2Ozs2mNyTRsQlaVEjSbj
NkOI7fE64IZl6kL3cKtQ2mdo7A6+1V9WGyyG2N/w/itzPUySbuzNnLrpoAvYTQq68KsuTBT7SaDS
aBSK2k/hWjmspl+evafXT9lJIGaKzcWeeZLKGvSWz8354oqk/B7NNgvEnbiF+/KXYbG31+eqRpmw
adBe1wlITg7J0jerc9bxTlQDeTT3gvQ4/2AzOx9WoJqZ8v3IGwFNrTmQ/lRgslHsTSI3qMFm0Dhw
bqwquiiJSYkXmKv/TrKB7MS82lHE0Vji7cjLLQ6CdGS8+W6L63qmRavqOD9ErICzqy8jmpbJXSoA
aBcUI/r91TTD42moTZ9Ra3mNtKCjZb01kK/wdFRw4zT+v88AkHfOaxioiPn4Qal9DtwKxY88vsEu
bxMQZy+7LIgsub8Stus4Bslrjqrnrp1i5RM19B7ferkS2Z/Ukds0+UrhRV0/wSBcJxPmCjyAJbXO
c5Po+aOtuCF8SLj4Gi3vJUK7/Pl0HaswHu4FfdNGFG+s1P0kte0BwQpLnPJCMmc2fAab/pB9iQvy
BH6a32OwVOBb9rMRY4uXO+BTk42+wn3oEmnFl/Z6kGAygVO1f959fyfmWQ268xsFV7vkhbGI9I9n
bk3B+JwKbNjAamqQT7kjioVF0d5nWrdf3TnTEOcSEjcpFKBIY4k/iqNI4fk5At4cDqgqK123/Ko1
9PQVRuN7AUSQ/+DfKVCpnDx6DkijFNddQKjL2afu3NETWGR2w9hfiZqx9MITbSFW446VEWtddHRh
sMvodqn49pj5/baNL0lBm0mBikE/hB5KSGq8yMfzugnw4stM3DaGYMtKWx++SCqwWKWD1tpCHeOK
04dsEjTCGYxostYfILaW5MfLRdDdB9Y+mtGyv+08pumEtKFdQmPlyZ2kZ6RBC9DEz82j9yWD9Vsc
8Gw5lWnJF0+mozLMx2eRbonmb8qIx0QPwYZcYVBN0fVMoB3qwI7zZSmEvoZ17uU8EsQWM7K7YVM8
AhZJTJtec6h2YuO59uVzHYI2PPtPJ6Kiyoq9NDfNhAwnj0DuQBj1mjulRqN2Y0g9LA1JgjgNEQVq
ENXPj8oS61LamdWhrPrsVqIQF0dSzNrwgUa2kjlFJj5wwV2qp0Cvvy1z5PLrDhVf7k7nAX1AlWKJ
gY9LIYPC160lgmMf8zTcaqxRSQ9JFTW6eRZBJW8afvRhPALG5FPUr6xAefrMjlRR0/53CeDkMYNV
shrMCfOeKMejGtZuO7HM7BxOdAFI9DhZIg+Prrrm6irUN7yAs9rC0ddarQlrktERiROKF0r8aiv0
oALHnOv5GU4f8+PX5k0RqhsWIyoQ2hzQzLP8FabFGS5rLzhYE1x9r6jJQDmL3YprXODdCt2R4Aq4
H3nfrEAOX/COMPm0PWnaAUDqX3w9CGUXVub8SNZnkB0QiCWJvNN86UgLaZHOPnl70XOQ2U/Kzkwt
rED/4C1P7LFoyPQXg27plmRdlcDnKXjavRT6vem0/47HPDR4NRPrRUQokV0N79/DzIVsGukjxUjh
9aS6p/CJK6F+ux+zA3ReXQDvf6U3kalimmRT8EB1avMmEZYKohBCcCyryEWFeDUkC7ILZsrTXaN+
e2Gh/reUC+oRwi0g2tbB/Xn3kvD8+fhb0nwye6dj9O8Jd1VBD0kI7indT1Q38ZtOFPjmkAFgDorA
dURbqwXgdjqx/Xwh7Oie5zFN6qbx3qOBmCCmLs6RsMHzEtqAD6XyghTK5c0ZSzmiyubxJh+HEXRk
NSBo3h5WU4x0SK+UMjtD19LoO2zpjtQdbd4hWzgGHIjS7UHK7m28i8AepCVabHPpeeFELaPsz9kd
A04lcotwKbLo7q8XRVRFuaXifQzVbts5tbjFpdY6FnKAwiRG/pe56O+IQRihhfEeWx5kg01u4xKD
NbPl7GJAHVfddtBpKU8gSHGDR5EoQck8rpdevwQi3S7Fvg05hgERZ0xIrntOgvXeVqltbm6njnFO
pM2aDJWeALz21v+s47Vt2fKcAIHAQlkypthZSpKmQGTQ7wNygW3wyvs8dm6l7v6u8iImDT1ZGvK3
Ngki/23Y0nxwml9DdDCPFOzkjnYgB9YijHBnXAbhReTPGIGOVW/1+PCbOp3+fRgmk1GyV54zYw9l
5UaIO/5qwo501DxisWQkZzO2j6QhY9CKNmEL1VFyeL7OeylhPsObarDHR5+RF3vqUjikyISUwkPI
5swhp3JPEvMUF9u07Cb6gf+OwXTPo2H5c9mRaiQzen+WJJPluldok4wPk3SK8N/CpE/kfSRpH0kb
aAppldLYgdF7tuq4I0Jk7q+dtQnu/bgx1ZVnYY7oLVdo6to+el2u8kYPs73Fz4eJoqQzSP9OsUo8
Pt8toQ3k3y2npKRowG9+IBGS+sdn8p6GXnzmT2EK8SD3jn2BolVunkQ2ddpBJJUUJPGiYAXtehRG
tG33VHRCZhtTQVHQk9f5s9ihFrceazh16lzT1rEwczxRXQ6tFKn2eZHvK7UFsqP/HvfHk8+sMXdo
1XSkkOK1raB6qBbrbaI5+hBRfuQieVGWKi7cOzQGlnYBvWCcY9Pl9KaAPNDKkSBTMekVqd/vgkqH
cf87Mi7schURDlvAoW7VSvAneey2dpVD67txXvue+jz3F7hAN/dCahVea+z5Z2xrPoa5h6xS9RBM
Or+TnkIXq+ecOoGlTA11lizkRccLSgXOffh+1o14am7gyBQ2lblm2COAyoGioUMQr+LdpSWJ6GBA
nj0w1rV95B+2IZLvriWktW4gDXJyeFAOAFdKzEDMQsf9BGAgFaY2KfEhIJqWGoGospgl5HaJLIfH
1u0HbOChBX/PwKpsY6b+ax6swkzoXehs7Ellpf/taEmu6uwr0FJfY0DTXAv5KnCBiVchWgDTtq8o
6cepq1pFzxLHQgn1hyx7PCF4uoqV0cOEJ3yNL87PFhzQWzb60AN837yUj0lX9rdzqDqD4bzOt/dx
SBzODEyI/rmbYo/3pxOSVAm9H0JPIX2YRfTnQ1Ac4PvdEDFZUQCI9tpsSm00aq2mkItso5lMiwFD
3Itv4AEgFkA2rCWLHwcZVi1bp2VqpvFv7oGEYrmblj1Wq4YysfyVdLwMnMufuNETwueHRiMadciY
hP4JopRiELQGtKXD7Gn2LIdg7q119GaC19pfb/1FgnNMmEl0srn0zMqVQXCxCWay/UnN4k6rJEtL
uzujvwiaSlMhBl60H6yvDkxpg+yhICtj0NteyQncmTuebgX/aaFg03P7bawREVnBk89EsLMxGBjA
0ocw21cIPVEARAxf6/NyQM2nkPyxBBC+7eSDbdwOhg1R0Ku6dC9AUY1oOK5dDGsaIcg88yMh6aTk
o11p5PC9wKzPEq+F2cjUEqtiAwfr3Ipwrbjv5d8z0w9rzUf9kLid6Zaxr/Zw+sdScSvI6ro2Ft6p
stgFzAbnFqPqYNgNBpYeXOHctIb426cwscFQ6GWG01yye4L53v8yjBkK1urVKg5rJmizLyM9KNK8
9CFLD/OXhRgCbFKP2LhtE7nifsDRaUUIo5sEJA1Fyx+x1JLSX2kdBYJiA8L+ONtxLiPa07RE0jlZ
br52apVJjywK29v9+jfSIGPQ4uAC7vwucCQvpGMYcwGdGZgZLwvCkPy6HxIR4sex62XZ2QGzMhE+
syDIWAcs9EjhLw25PXFacJs8g6oN4k9ioY4f5fDQhyjapqEbj572A18MRJqia4W+9MPLP/eBL0/3
XjmBr9j4n6TcQJfeYGqz0oj+O8hFu1uHx14fMjmOXa2N0/qhw8on9a2/IeJzShKoU3PeMS9x7eAc
Z7sfspCzes0ESUlPwMnaigIbDMOOsrkNErvhFdWVZLfRK4onnkriosAC5ZOfYrVUFO+pEzLkskOl
Cs9pXUmUSNOOLyhoZ1db8F4Cwp0kTYEwyhYjpzanAS92WqYXKBM0dASGworgz/a+xyh/SO3EDqYq
uQT5ZOkflBDzgn57JM8n3OwBaVUSR8CisWCe11Bp5vziJvKWnVaIfOyqy0nn5AETXNbg7Suke9SS
hu4OUZYW9gi+cCm45H4sxPD8pAK3yHtiQ7I1upYbNVw5FNH+TeB9GK1VRJAHiskk/8tGzTajLLZ3
xMuJn/i4td8zOXPazkDWljAVqzihKbnGOHxSrXl2AFOAmZSuhqR7U3u6qeKaTHGOS+hLTnUDdf5k
P1od8mHeoGkvW7XDGMDE+IvQ4yiXdMNtw1nukDGnHLLkUMmCoy/MZUG8epC/PYlWApko97ByU5zg
CBtjj5h6iE0LKAdyH5CruHkLPS50x8+cYrdyVLPQE7fXoEaZxtdXX2XGeKC0dGVoDt/IyfRX3s2a
+BT1KPJmAcwqhbcGnuFP3gqjapRdjW1vJaIlQuchbUHvxswQal6YTBlYnV2FZ0rpvi52Vfel5xpk
ZJe16aQkBVgsXGgW5L1mk1f/RCq+RRwzPBsN4ujxOwRsMFL8ozK7iK/ZQwefmjesBXCL6tFprhDR
JLeK81SAwnzgrSPLwBGR+37osAKuar6y3QNQ0uXX/i74xrYWcng4apgvv2r4BoRWP7bOpXaccUnE
/en0wOdM00B0KXxTIhNsoQH//uUL6FOj6Urmx+1pY/uFpBQn2eNlDFD2K+cQv7lCM9sVgyVxclln
Yib7uoa7BkcrDiPw6HMnvuEt2mFZt3PdYRDDVah+ffXsnB/SyUcAy9/xvDYJk1kfPHnUaiTrNzmT
z25fFLVcMVQjmo/pibTUAa1R0KPqXhXxs9VsMl4eEK8vIQvrukuqWYdx35BgwRK1H0H8teK51SIK
JYIt6fSjtP8NVz0WFQfsvmVexE4nio3kn3vdWm9eG8qSU0mPCyIXe9c/8HigcJWSdTeAbSTHs8jh
6tOMn8dQoVjgk5zoPQWnC1e/wp+BGLb3KF/31Rf/JTME36zyL6ejFBP7Q9EciCBa6khcnVwr0yzo
OWFymqU3vA8QyDmbXoRL3ppqRCTYS8N5KVdfWqz+k4UaPBoDRW2+9lqHVzhW7au+lI5wk1xk+UGN
I0CtRNrJ6RGd8C6qVZERfgeVOyEytLN9VBkNBNBqGimnNiUKp4JAJiYDcyGDviUGGJsIdlcZwS1v
8miNv2LJQRZY9Yr8wyNMC6cUCv45nhLmYfIDUwG3MjBUIrxKB0egRNolsNKaFJjRsNcq3GzzWRjb
ANy8zyqzlXS5OVeiaCMA+mH7MJjSzQ72AgZhrFh65KuR6Iiy1mNaiXvDW1Dg51MKQyhluVngi2Ss
63F/kqr5H3XWI5v5FHHS3pQe8FTX5CHkETpOtoQKugi8Fntoh/Nafuutnh/gscuaRNTLx+hVMYCO
7GSGqF1XF1bcHB4Pa6TGDyWLNH8az7Cv9W9dVugUOWzkDXD67iyxjucdURZ5qSDrsGHB/pJz4Ge2
KyPDP1ysf3wje9mJSSakoTEDa4U47rHBH+A4j5pt1zWVJRxorz2oCeiW0raPMhfU+EYDUbGXnR1D
5wu9ajCZeUOnsPrnYoRHpvc3Vh9d8p2GN5ZmjHt/UzL0uMHvrp42SuOmmFWiQNKyEOx2/Q8Yd2Ic
DNPqFzznuTMifswDTI1HkBCMzeb+rQinOi66ysxJXAnTY00294gbcBI9cG6VXOmJv3lK9+iU24Wn
QK3dhhI/m+pcnFX6BxiVBQn2L9NFghyrzBucbTvX78RptW/ngrIAa4RN6X4NcnsugPQ5UNv7x+MF
jDWLpbau7edsfpusJuipVFYgWJwaD57eflyQKaYCXYLn3y5Q7rWGMXaiah++e9X+UoShLUkrPaym
nxljorc+veO1ldAFYImRzKSF6v4gTrHEWR/0oRwr5ICbfTIf9XvyUVrpDf1dGrKQM4xxvfFuS/Dd
VeOPBVr/QeauYBOAjAJSd5D0O6qgUqAwfWFmUdwyfefIECNGecqCaVar8k7GY77XbSui8Ci9Gm5C
+FzUppr/QIk5km6TER6wJYZ7rdlFlZYAhC/F2tEYsxT1X8aUPo3JE+eiAYAv/QTSW/d9eDrRazXr
ZZf3ikwjt40AjhTa8iaD6UqJn4RE/xphaGWFUozNKXEA/wkl8QKGwKgdUPtytkWmDwD0oEQ6249+
BY6WGe8DSk3NR7v5jP7czcJzXqrD2fYNKP9yZJa/osLTRLwc2lsslR4Wg74tbVcr1GP8Swiip1k6
3JeCrFq/n6Ta6pkMKaSpuwJpillk9AV7WFowZgm4bBf9Dj8oJfm8BI383KByHvv2rzKCAy9NNH5m
upjaet+6t9tJZRiOxPkh5J21M/ZSzMgRItDxnYcNtuQx0uWE+2MwLZm/dPlU2C6ajW35xlKNp1Kl
/fCqF0eRkRvFtotQ9I+p/YgCLaJUogri0/fwYZz2c0sitWlN33zOosdckkO0j03Gw/I8gCzmcAqn
qlxI4nyu49/fGcu5ZS/VmKoiNmy+HSbzxaCg6rVH/nPDF+tzsCwQG7hYISMQKWsv/yLMmJ8F1bWB
qPeOo8C5F1HnErSITucL/1bJwkzT9rMX+s/ks3eR82eQGneTcjpGsrG/Z2yV1MHuktEkOAIDOBXi
UqubhGgBaOBMBP2Q0l2QV2jvjia30Cmg7jPH8zVWIia/xI31yIK5N8ktc8wz+KxfbnRu4xU57qWz
uCrg9RA+O0PuywbqR5KYztCGLDxOeV6Vdssl/qrucNzyp6qntOHX8nYhj7Zyz1Aj2TiC6O3Ujh2s
mfzjpwfv6PPoO4JTgLpIrftHHHBFld4hjynVKYsLqJpem3fGw3+jtjiyBarB8FRj7lOl3IBtMv0l
A8lOBmBJvm4HZClmxIbDzBbHVGnKL2eolxxbdhovzMytChJbEwkiEBZA7oTZqIs2VTE1xvZbryj5
Xz5IgcC/byJyHKOhwExRGFHKq735LovMK9dB4PEn/j2cWfE08ZeKhbUjqWiw9IrWG640gzV4Jxdb
Gg0yRl+GQReMKZQDY+wChrvtceLwrh7Ptw0CDUeFe109DOOLb0Q2KYC2XsAl/JRJ8n86SZrmLFlT
rkDP7P4VdphMRP170VzJZl6sCj2ys2k7F6xPhpzjav+6JrMm1sDOOBt8eS+CxmN0FRedR/z/2mn0
WpcOscknNtm0HvSa3lsWDmAl9PVblbBzWCtRmFCe+7v33o5jHdHkFNCBzlLAWOH8KXaVgLSEcZJc
JPk76bieQwWvNsbdxE11x/htCsT+02Npt/9FCheBX+YFufKGnmxfLiji8dhhT0GxBy6mz6h+DOCj
LJLsPY5YRFkyaEKZcY2C68rlMIBSeR2K2kDfAeqxjf8HQ+qOihP6u+ZuiAsy4ih9RXNFKv7eWlxT
2JVam7XO+fCsD2PRF/vLB/zlfDlwp9invrJH/GwaAP807kG8XSLdN+vHXnmydYvsjwZIV7oQu6x6
/JkVCvuwLI17Kflz/A/TI5MjOIetzjCKU2i9fw5g+j5I13QC2lavE+m8pYyihNyOqRMWXue08EXY
Jq6OtGMa4T0P2vrXAAnpeydDo44ZHuvrSe9llgPXv5/A+ImZZ/KJyTIruQfhpdcv72mjZjGW6rWA
Z+TzL92EXUWw0ZEeJqVAxlo1OcGO7bABDQt4nf60QUw3X7B56DwYjGdNFYmeroaz+obxS/BgBhCA
YX47qwYlOf/O63Cfqay0dngyVhkZj61DwxIPQb6BFatAtoqvrOZy4kSniIzX2bd38JtajtmhI1vZ
jtko2DQ4k+iail5QYD0tWvlePU5159pLykwV2Ct4iXvHFRbQ8S981qpmrrjQlnE8BjzXRgx5r2hB
AEhQgleuqNHiXtZy4MomjlehTtSJojkhlg5LMp9crvFEsFOANITpUaOHTHICc8KatIMUcjgkhrQu
zZQl0oju5URTvBlZmwy40yzaWjf1fuMXIHmifDhkaShNfotGoTtrkWEBSDTQQU+G/cGGKJabRMSh
DpPfrR/iZ5sF7zwOfHSfNZfPUxZWvnwz9rn+pCTNrUDd/4C2wapwZ7xiYQhsatoBe4jxoimYrF6U
EwAciloMrYV4dl2gITVC4KrmQvVwEFNkNXGsq6v1obOZwhdwZHUFGxu192gBcElcegOG1lHMLcZf
dDf0arsGJ5ushJf0muMuRSRIlgWYForGZT3Y4TjCMUFpuOzVY1ex6gW+juItoBniFBtlkSbSvIOE
FhE4mO7TtIqnjiQQTNl7skNLPkHVbE7eioJZim2RZiGAE9V3s2jb1CEgLVkkbuisTWMLtYMnzrZ4
skasj/WSXggSx/W68lekSyJwRJH1BJRrdfezkDnzON5e3FeVm+BWlPYHJfMh3U0oJhcmlrwpV3c7
2TmqHoMzN/hkhmFZfsOBUf4iFePYzytDRcn6EaP5TkaMFgt2zWLxHGCrrL+VdtzAsck2DcMYafoz
C82ZVIikOZmqOA1iV99rExNKYq9AH/IKs8gXT9XzBPCBlj8XmKo9PxhWyO6R+1ts7epQ0RWxbC5R
CvrsOgrL8LVvtzy8GpGsoI+rZ/aYoiZ1Sw/IWteDsS427dF4iBsIxFXI+aHCsyYsp4Qj6MsiFSQs
KkPWHZKMeWbSgequ7lqjUIoK7bzGgrTj2l0OsbAmdKLLRZATwJSmnsJqPR0s1qCw4+9CrhQD8bwI
Vgic/MS1/evrLhz30x48PzqOYim4vSw2/jde8WDeGNLLdqbq/Z1uTW0GAI2rFR1rMCoL3njIumEy
rqxIuo9ZiKKlzy/0GMttra3jRALoT4O8Yk3P1DS7RNz9j/95+eYNzNc1p4iHP565rHh1JpiBF4f/
v9lfLceocErrVDQ4X+V8LoUJl2BoQCXvMZraOmbKaL6WgxvDdr9dyFAGL9+ghgzOuoMTs6Ybrp3k
oIAT4uHVlkUnBeQ0ayLGMEcQXXlYmeKz0o+bv2P0iAJ4thPVFf6o7bZnIfgzP8+knHPZUAHCqWVd
mV1oG7tjWcj66uU6dPIf37LD23j4kJXtmMh7UH/YLP0lswvsac0R2Q1a1pt8bwi4DZUKhu8+Y4Vl
3UEFdOv5ECT6ZBIGY2DB8VohWE84e3TbLZiZuV53GJ4DqG94sjt/IGUjwNTllQCVa5034fJhCY5E
7FN/X6+2ga8v+ge/yUuTjPbFytfV3GyjoswVgB2zc7raqVV2J6fuHw2FwvVSDZerfxEDsza51chn
noE/ctLPGQrfPI6oczJGNcMm2BqLzLKMF/vYZK/fEqhaH5HqEIQI2MizQI+gfO8Aj0LtNxR6Ykpq
U6D3g94IdkZZflGn8RrJ6G7+WXjQ4UG5/i6YCbXwpK1PxAZ/kxgDsBE5aQNbxlfTvtmDqQJT2+z3
ZTIEIy65cOSUUItN/fY5nsQIzdcEJLLZ4Ega0gaqAo3/JES43n08YHERXrvpvxrkw0Weh9YWMYej
jVT8vKU8zm9pMzq+nDydv6dR0YH3lE8jdUg3hsb5awPFsmWcM953jPj/Y7ygHCcpTD9XBpkOF4lp
8H9TXDrjU0vxHka5y963ZOSjt8NPEJQbg9ly5Iz19Bwp4Bs5nHYWsIJZDV0AOHTsUp0mO8RyMB+J
XN1QT9iMsaJJDFHXkdPl+Om1VMCv31dwLMkrZf1NQoojmMEKibUH/7h8aJl/NlnPFF7vIwrACmAZ
TUwjfyGDhlyERAZWy8kQkVR9701diJ9aeD+L9YCaozhOlo6HwQ9aysniu9sYo6xjBCUSfgLZNiz5
dubFTQ4Trpm3gXbsROG+HE4182YSJg4tXL34dqkgWR/dgpDqy28Xi6NhzCat+6eIxBJaJsvajUIK
N/Cnbn+AJvonKat4v7/PkdBxFqcztzFfntCD+nbuG5S8hcefpMB5vhyh8QtwH54nQEtQ5sr2+O08
EpNIcnUo1uyFdgFsrH31Yc3Y5APWkmDTQGOUk7eEq8v806/F/KJMuW58ljcR/mStYu72c61Ry8L0
byvsvI5TPzfLz8ArAofldyu21A71IHtXwpATAmQqmMyMv/OnnwC/PXE2/cxF4vtVbYa933o+vTu2
aaACumIbOaPZ/cSX7fmg55qTgS7o14jbnxccj58fYVu9mwsqwOnzFsyJnBI6P8D5+sOb/YUt5PD+
xp6zAvL9yx6JURLxE3Fb2TfQqdhV5c0fY4+QVCV+E0Iw0dhiesex+RJzJEcutVHqV4TlpUE8XF1X
KOkxq5XlP6njugmp0Q4N3HEIEIym+lLuPypdEXuryqIj7TX9YQAF2Nh2j0Kf57HylWqyfwliEM3d
R+Nj1GmT+eRA6Xj/clkmbw+/atiA2U8LfQqtDkkNu5v694ftqXlaaVIsl4WucNO6YA5fRVb9VoJw
43kV35nu6/BJuS4as0/KHzHWzRxe1ZbYzyy2aXjllRXu/LsynPa7JGvuxwRfhyHpVUQlCZCMmrwp
PqIPY/CBm0sZNoaCn4LgHmw/REf1XLafD3BqMfGwofNw9KH/dYOrmdQf4BCZ7EnB8M4gaCPptrsc
Uzkimrq6KYO9lt7BTF9xHptY9Jxh9ApxCVbAumGrK8d/onu9r1tDi6joPXguIy1HMxfp+dxKkF1D
npbDYDjTaOogXYWUr8xJZAGU0xjVwtmOARJvZCwgLY0owjpvgYCu9l0lMXlaeQhyU1gtXooDkc2C
a5t6w+eI4EGAQKXyova2EFIolFTQ2Gs83pDAXnX51Iv8FnsTZCETtDYElNU1U8JC8vf0u8saxCPi
F5SrAXk5G1rJsophGmdRZ5GMHNcWhnL7q4GqIDBrgrr0rGye9SOYx0ECdK8DeU+0QnBpgVXuMNpY
chX7cuwBTNkFDmjXwbmtuJ8R0pjt+xuUGtRYi6ifheVbNohZAUJjWDHLgHPtbYcbltfW0uJguqlg
r0Z8jQ6Cc8St5xaJTkkpoP6xoaz2EuKIhB3MvRtY9LDbFh729djPA/2zzcCUwlp73hhwpTkGyStP
5GDU/3cPvSuKkNfT6FWTXkkSpHkW/xHO+P5IJ8lTQ7BsE4BaUNozIPfkWVYMHK9UFNIAZ2JWHOYd
GGEY2aWsMnsNqipma9l7puDbH0b2GubVYRUX/WYnRJ0Zz0lRKDzZYo1ToJfB/SWUhX+3GruhyDsM
g5Clwb7Y9/m6+22JaAnz4tJzii2J42wDKzdIgkD9C4cDISU3mrm8HwEUPaphdiFIfc/i5R3/x28I
mkOLuDrbjBiVrBnf5aNWyzCF9Ab3cRz+iZ5oZj2nG5UJ3/4/CAPnYLeEBeFl/pV+Bc+L7Xq9Qexe
SW//FVrXARBURKcwSPICue+jSPTbLfXfnPV0Vtfk4oZXkvjRxc1F3M460nfPEV6b3kmgUA6GkwBX
ZIYLDqalR5vQw6rssFEf/QSJV8HwQbQeDNvZn/02vEsACdArCUIobjEz6+tN5MDJgswnaM2VmU/7
yUObyYghp8v2ipuWv5vm5xKlGco85+kG01X/IyZmmTo9SrVjnFfESt6I/o8cBYbHByfFd/bPRWWg
BZuFdgp2HtpqXJ02oTJfiDN5rdTTw6gL7q9JoE9pyAZ1nBJiCD33c5Wis1SXJ6PfrdEyErChxP/R
5uZNv33tkDKxrxD7M+wpa+AFs+zERgJHmtL0Sn77hfkb6OnRVZJtT6FOQMJyjHkbztP2zDwXnxj4
0yPvNquSHfxpMp6/8TuGx9rHMARGBRp1jWyXk676G96yOMPJa5qcBzqzXFr5mK/GDNBITSY2OrFL
BhR82r+U5WewZQ1dYqtzggbWFIOG/yQfkxEIdnN36CM00HoO69Q9W0Tft1YHliDUYCH0udw0Q8G5
qbWJs83FpwJzifzNbV5U4CdPQ0rVGa7vOZWlqqC5HsMdOnEQcutkD7KQMs9Ge8//rGXAjw1aD7iD
U6aSJ+1qcIRSyRbC5HIomyclhNuO4prpK5aE9pdtLhFyeJrgP8dRtWECxnAgUAWRiqvpISxGk3BK
30FQdiw6ihmBle/iV7nkMi3VWhAUimuepBpLkQTQGq6W6RcJFA8oDmzxCHE7vnKdwpYMXtjjlfzm
amsG/AGGf0jEm4Pq6CZq8hWBd6TNPK4/k0AMWN9isqD3OUYpTaAAx7q6kPscn3SR2oaXUBtLNGer
qBk7AbENGkL38rD/gSL17Ful8gh2Bkj8dsV5EqCKtsYpZ5kuAJXwe9A/pCgwLDOu2eHv4JsjAfwF
IbG8XfM2nmX5DU9VlmOPq7XcWPtBjU9hJNJlBuFFh84dGw/per5f8bIqQsNmlF0pDYcEj6LUhnrh
Ibbz1/MFOHWo1h/GMtCZrAiVg9FPO6pkViO5Bchg6BwuIHGyuKwdrN/1Uzps85fc9VgaIdMdRSM+
kMEtkKm68lGD/9uKuhBtHhpruKd0jlNaBhttkcVit0eHgdN5MzXavRY76Mkk96hw3pjtjSmL53iT
2nmNAJ8HXnyEX/UYB5+y/FJqizwOAco8A/sOYCLzP57F6LCR3pM5/ucYyr1PWpe7sYok5LNnQYc2
i4w3OQl0CPQOYPiXkpMQ9ty50b5hDzJIZPuUK6zqLmDw3/rQWxVvOX1x3kc3gZnRclo1h3VfHpo0
lapqlDZOvKlV3mAxxaVLurQgFfKEt322ufRcckbNJdQyGlO1EUgFJLXQrdQjqDuxpeVCS7VOUhFz
LGSkgy4cwtezzRI1AmG1gBeHdnVRWVTTsG6QaFeYj51ANrEo0yuxkKr2NZRSMgMKKayB0H9BGKgY
9V5fKcmoYwvBbjCuLbLchUiULH63JuTDkVX+wPlUvy0TJsLThtc4VGWHc+BMGZPr36BHBMiFrSuy
TwJifR/3qu0CbHGSFsOTsGGvkp4KycDdAWObRvgdjtqqe1nCVr7VzL2X2kQgFPB7Ko9DdQYLDngO
AFIdGWA5RwW//cuvqa0ipqyc8QREeAgHFjLI5Byp37UTxdzIIpH6cG6MmqUAy/tdXRPbTPaOYGNA
U3nsMhPXwAdc3zOAIx7x+WJqKHYp/iPZCtUQAQlCOJQ5fGhNYoIf7T/BZQZfBWkQyUhYJMr/UAJA
nYyPS8kHCI+05TAGOf/8tsQ9d2RXu8Zph5suCha3lqDcjNTPDwDovpKCllV8V+Et39N8ysoJb1lY
ojAlpnCNLAOKVkiFCtKEMDdDQQVw2Nc4XT/1BGn7UnnvD5+qtzUgEzZwYsNqShcy959i28TXLj+R
JSHHOesebnBAE+2uE6EFQdN/yq85t9K99AtdFkYJcNTlPxHu9yPVB7JDUc/1/s1kg+1NG4Y8RPcq
YHTLVQGGSNHGz5F/s5e8Rq3SgPbJDPoMjteRYW4ONRkeexXXv3QXxwU7s68Dt5s3MS8VSVJXT15x
74O424VJUlktq7vQ3LuFEw8ElMllsL4rXDGOo0XL1mowE8W0GnnXWLLf5jy1hHs3o684tBT+QkG2
D5RGBa+yCIY3Fwo0fopVOgMK5yosQIL2SRfXAwuNTQQQrZ0tEOUJjeuwHYr36WUW7slRyNm2jTVZ
BEoiqptT40oUjT7HyBsslE0nfKhOksPpwd+YCxi2Zm10dJfsKtpdZ3mUSg6vXglHrHySTLNZZktz
BgxIyjgKQuPtpgh70lDg0tCji5n/YPgZsCj3UGgq1gP30tQrGmG5/TGP4ACv3Q7TWRqCCkFZSRWc
0B9IILQfl5DSgoDqgnTxyTLofa6ESqgOQM3W7DiYHtaMz1GXhND/TTOcM2JJwoGh2QnndtgL52H3
Or7wSVRl3j+cRfnIAeTAKCKSQSAjJTWCfs8m180h50BTZKyrreNAOLIKdKFcCFn+aJ1HWfaZ9kaH
RoqYMNCla8ZuJe+YYq7Cx1fr7W29B/QCl3hVD5pdqW5HEMCkuGEjc0uiQArN+BCMPIEQZn8ldZnS
caevZoYU39L3nDI8nKg7bd0PRNKESm9l/89ZzlFQ9naZB7I026X/EMOcZ2ySNzqyH00HHTGrKdxk
L8zfLyDZf5U4Ac+T6BeglvUAoE5kZJ3HK4/UrMeX09Vf+FHu1N0pYHGoV0O/Simt796alAbY/eJR
L+COei4+sReAqQ1PsfHbHY0dFl6UpHsTPMYOmwaRJDoMn1r4lMVmPaxj7ePvJOk+7aOVVjJFGIPq
b+0TgrCGNdLkcZIPnvtc1ZydlBbLmaXtowxrnBCBYOJvT++5F0EwdNtuA49EdQdnOvm6wZi+kWaK
i5XV4Fb/huKJOJCD0yz9adWd8U5HePwQO6cqP+ZWS7w1KM51YbrlwWhRYEeq96ne8OGJnFra/Ypx
hpYz4XTvuPQVqe9ky6r3Yl112hUn8VHFaXGD7SZm+bGtLhvXE4Znxc7RHhhdOQkd7IaThsZM1AVj
XYeUEHmg0jINyk/aBPTid9RWn71GqgzBb95y5+qIQ/KncuhORUS2oxVp39dJUhyoHiWE7wp9VEmt
HeZmyPpjKwFnqNa2IWwP3Zva0xQ56t2vw6KB+2L61JuerMYNGaH7CR5Ge22RZmQc0yH57Ur2m9pO
1ykqNhY0VLAW0/62vYOymoHL7J32mwgVT5W/YTdXnDH7zEJo4uNw7DzbJo4nL2nWxITJencJR95l
/7ufEduT4Ag3dBOzAymmbKysyhHkKWXYD3N3MCujuDNlSvxKlGuqppgstBIljHmfrnHbRSvte0L/
iM72KOsRFzDt1lfSjcfT1xV4Yy+Vu+EpVylPoLM5SPVe8fo7K3nLJXhLkvl1xHQ2vIsY1rPi5+fG
OTY6h/9lcFOWKqkzKduz5OzyqN/htqpwFJw+zxcifNAfEVqOHAipIwosL2+nIjafaF1d6KkheewU
ABVI3riczjUAG47wpKg9jtXIb7pxMNb4bFdxMTqelbluIyo7/4ZaZRb971KmzlJZObc8XXfZR2qx
2/gly7vQPIN7ibPIOfEPOWO4AQ+wlt7QlFlFEDUpB9d+t7ooLOU5io4bTsPmyaETc5QzKyMtelJu
wDUK5iKOqvMqu0y1lvYEvVcdU1UejFxtjaCpIqzlSFBPRaH5i2zB5DMwiNO+GEtG5n55EnbcFAW9
xsPekbA3DVKV6XQHRzGMuZwKfv6oeiBNNmC4uqBkIayGlMvKQ46YRbel44vjQ+TKfox1Tf8t6Clz
zRZMoN/1YdSz25x3NrDRub5LxxRYVIwn1KV6A6KvEqjr6ctljOzJS6Yl5OPodAq0xsDsRngciLV7
CcNx+B4CBE8sH7QuacuuXII6XRlk0lzs2KY2YoZERiB2BT6gjbvYQVsj8M4TwnV5NGNipbC7rBS1
LLGIo1J5gnhpRF9sb+zeqv3xDYqfRau2KMPdarSGTFcsAeA/2EBpGA52lHYF6kivzexHp2fmf4nw
REUdFZxDfqB1nbXhB7FHrc2HormCeM8NBet93gRCYzJLXlZGXVFpV0e+2H4HnB3uZ/vycMXJbhKt
BFUpuKENCJiaBmZXxT2BmV2WUtEpVVU32DB5VlY2NESUf2d8UwmJhb81oVZOedFIRsH+OdPijV+Q
NV89pf9a3DddDBFD3j6UkAicZk94UrxPZKIo+cZ39I5YpFFyBQkydNRKt5FbsOuuSxxEhsirBZoV
9p9wK+RTAmR25c1gMF5FZoecBa2w+eBc/N5TAaGPrgjE/uIy4ApW+UCfOJu0Jf0dPL5zP7sBIFxS
AqT8dva9nYOswomiarS6EhogY1x9UBoQ4h+bvW74PxYzUOvofldM7eku76huBz/NnvYtvF8vxDWW
FfMVSdmAk+DqHjT1SrJ4X8cN0BHbvc8QHncwp7390ShbgheN9O/XF6uToijG+AyjZUPRPyFEu3Nz
yROB+CcKhrGKutHsW3SKhZiccwydP/bH6B8TeXM6GsO5BoEFV6rmqZI/GZ2USgmFEinNWH1eXebd
Wv4GgwvOSD2c/nnEKxYBs1B+sBJRfUWo8yFTjMsK5T9LixlCneQoM104vc6dg29BYhCS4ArZmyhf
cqv8ljhPj1UohqC2nBb/jP2pD2Os6QsY2HKI+dMf9h9CyuFSp5kohn8NzVnh8OAbvIE0mKHI6Iv7
jJtFl/RZ51qlBTF6q1L/kWeEU8V09O36LCJhIqLRTuVvVK+ooHS3OijlB2LnObGxYlCGGqhKDHxs
iwR0k2V53rn41iZaTUt2TiIjfWeNoHCjxfDe2VshInsBFqtmYyTV2HI09byPk6hN/A0BqqSoMsCs
P4HdlZlXGyLvdmgFNzhgDKPcnyTSaIQKiPy4LiHtgffuWAhGM2Ob7/BH0x+Rboeyc4IghebexVpF
FCMzTtEL/u59lyIdUtUzZ41m47Tuncoio+y59C8yXmfz2qphEFNxeAvWpa5fLNOBvSS6iMUOgDtT
OeB169yurHD+402uu6JSHIYbJzR60iH/thHPcVkOGaQptYr7irwGA+h9PMMkDZQheLqx0x82Yk+D
B40tWYv74sC2VLNL5C1cDl/nzv5yRttPG4bQbEkirD2oh5o/ZmDuga2KpWkpq9VrOcvOnT7lvO+A
GvLu4GHIVedagSaHHlWmrr2nhssW8fPO8z1j+ugMNVx9AeecH5b2Qv77OPusi3NaDmavb+2ogehF
4cdgHnSWaeUz0PqE3Zr4KdSw/VNSAWvG+AHU+pCcTGil0V2cxN9FmAlSkP8adfshotG7uHRjPV+G
PmNjA3M6nsHcnD55qGYsmQEAWkGfChkvLmsxy9viVwcQbuFx9JrMMfJ9KqI2Fm1cu2dD4AtePdcc
7VoJDJVsf9OJNXWcEOg2nlZ87L3TR3OAaWBP+UHciDQcffUYfEOiX8u+ku6XAIICu0oUz3PF4VEn
vZlya9WAus91zVMH30BnFB6FSfIf2A2fHhozYhE2qvROFTC6/mu83v6iLGwC9207kKO/7Qxcm0vb
tWq+OQ/ejX8UA2mKArAdE5Uvf9r7YMUhsBuWBPSTK3+lX0DzwfygK2DIOh2ZOwKzE1TBHumlWR/L
/bzzGfIHiWE1AmoIxVpfOk8vCHv4j/bHYte9q94D2h6Wjsp0i2JbaBqH9qRi3aWOw1hHxu6Wa2ZM
kTbNLdfjG0Mc6jgKbvlSIYheMKTlJ1CXVJKatfgBmAyn4UwhlCfTCd2iIJifHFN2kEcS0n1mbPc+
UgrZGbA6js9sM87dY6KWoQUH0lil/Y19pb4+NXQ38ceJqWtciGHtj4xgze5ZmFO8dT53AlEIGcsd
H+f31xtN/chStkZH9r9WLTHE7MbXyXKyV97WV7so9jRwNu8oSJChp6xNVNqiupTgf+BzaSZhocFM
j5papt4gheBeINUGBUuTqNSEdjrDSILm4sk1YW2FPt30XH8e6tJuU4aIGYL5V08ZtdgzxN4y4wEl
xzNiKEmutp2NlaNwOiyAcdqPUdnwaD/cHERJOkBalmH2u5mg21JCTgTNRMf1MPTKG7vFciPPXG2f
ULzIImmKZu+DlIn9KCY+sfdEgu0lxwedrzFRpXYC8wNAL6F76woOQ6fooHdyhFr/YWcci8eyDMcm
hdBB2fU+UfjN+2PR+b/SzaZbLoJnZbLrNcfV48HFDq/RbgNyczmLjqWn1Kb5BrZgz6QI0Wo8Pn0L
1zNIsAIHC8EogHzTXjh7iuPojq8tYcoqH58LQnO71+yBssTDE087fb+cMR7pbAjmFj/u2Rodw9YC
tBdKhiSOqVpQTA2zNCOvVPYlA8y4lrg4wBnqHmj7B7+BTOY0vmPgBlBq8vPV2dusURltRltLlUe1
lAu00zNVVl66c0ki6UkMBVf2P35UnAf8tlIC+jd5YLRhYjbVJxSvSAXFvx/uVgsbQ5KM+DJ1sVkZ
P8JKdeAUmhV+w4ySgtt0GkCYhUdU/wc7fpDvAYU2HZxE8LX57JJGQErnnhdBbJB85RhemrZGTv46
wR6d1YpoIUWYwB9/6mI4s9viKog1Ntb8LVqOnZhNqitA2G91+nmoMNtof75wQBhTn0Yqu+pbaiSp
TOAhYzfUZck1DzFksc25VwmwPGOaeRmFQMIzhSxRarM2Mk8b012GJ1M5PhsahlhazjoiMkUWeweM
DuQIbR/XVJgrzVLgmE/BS9945aDyIdyoWdCQ8POvXwAyw+RC8XcgqsN97dNnW9Bji2Ea2YqL2hKb
TxjFGhqvX1wdPGXR0dtCJE8Dqlu4aZpuD3ITv0jkn5HP8J5lkHouVJtsUeRvnuplf8RbZX6pqivI
LSeMMT+aokx81ckb7a3Z7NFT49BzvLgrxXFwapYbYqdqq40tRHA1svchDMHh7cPPUe3htJ1ZnyaU
B/kgLb0xbnlJsc9F6ftyajQTCcptxnKfo6XcppjxN3QPDebKkTNzA67yiGN9oKXOF/Dibtd6BDe/
h2HPEKzbeF5yMQ5jMEe3XfmaU2UU2MYr/laiVqk8bcL1HZOFS2f7CC9iIJ07RqGfqIKer4pIjZCO
XPVTorfxhAeumeRIQsYF1BpuZ+Knb169RB/MWzdURCw1uo+fc9LihM48KnMOi68TucD+P+h41coU
bMpsa077osT6R6nhbShNL8tOQNi4tOdhzBjcfv5vbIey/aKzFzl7yiEpHD0gx7cIM2ShB+/6gR5j
1T0Novyik++Bn8obiOlTg6HmuebS1JuvOGb6nTQnDJYo67OSF60n89TXePgwE1JpUsqpJ58GS5EO
gK6qAoa4DE7KMP+LWJBI+HBPck55ih3LdRkWcbOyptfX1gud5bM9Pj41fzY3TC/JCPBjpOI97VKz
kHytGOcktz923jaa7idhoewlANoKYmzl6IyVVuJDivjUo6Ki7ujtr3C/1SlPRSfMixVg6QH6pvst
SjuVKtUOLCWGO8KKT3GuVEtIchDqt7uf/BOxQGskm4bJD4mERDXGQbvny+D3V3rXKBDgbCC4+Nhi
0l/ffNLwIMD63sdEivlS2eKNU4PSxYfhs024TciWr3757EFB9dcyWXZQewEKXeWe9PFCD1hBviQ9
yZBo5mwxt2qv4XWZtTdRSqH77aT4DNL/uMTwZkQvF/tq5igglQXlgKZCkrt6voO1rUjDcL3RUCcE
m6DHuCQcpRhwEVrd3wwYPm3VxoKNz1TvONrpW8lzV5e/nvJM8uGHl5qkVFpKQ7C4JZwVj588Z2mf
pETLFzTn6YnY6Y/6u8nVnMCBRsh3giGnkWr8J6xWJes/UY1uzPE39nL//92OK44VEGeGXg5vJah9
csEjKc00H2M9rf4PxXuiJ4VmJEO+ExjNKMR92uh07XGJVIeaK27XJev4HPFUeIwZLIBcgabUDknV
rQWnsXiSI8nVNlnw/1XHjqlWIA/YPNNAyOeg7Lc6d/RJ2ojmo3Fbfj78mzQTeNVSEzI+Dl4xgin7
xuEmmNwVqbBbsvnf7+XEsYNQ8hmuhOOlbjZZbZJ77Ex9Y6pQ5siRLixrSbI61ZckLqbpPf2406eE
c5GBPS2v/EQUG64coX/rEnCZGJjHs5XxAaaQdJdxec3m/OkaxHGyC3J4rAHSNRRMRVh3FwEliD8U
Wbbf1fv/HYXVK5fsz3mhAnleCSl5ZIbJEs+4Klq0BKuGEE6zeTrUsakI7iJ2wc+V/W+NCoUZ9LAX
NRanAU/AcZedDbeE6MhO6MJgfhCevMD0Z0CBk32GhN1En+yZbz1s1T82mobVeBeWyODEUizc8e42
vaZSqEZ3wiy5Uvj+ksH/WI/v3z4yft3tvyv7OjEryx9t+2LUINJKvQEH9C6ep3EzyeRy7gEr61mD
Ds/PS+69oLedJI/pkb/FFx2ZQog08HaDA0j3KHZEFxXbgZQcrfJMDk6Cqrf2MXs31kElUoA5Vtkh
vAcfNREmaFyfdn35kALhKNqIC8KmW8B11jTCNujLxwyFAE3fz0V4hSeoeamQUXL6MQ/rR1hB8tGl
p0xVgRFQIX6rQU+50B71ioldeeYHhZ3sYsjeKPuwigP+GuBq088ku5kNnNLbVeLTERimaqBCdEo9
pcg2J/tITSGTxR+ji4fOCWsJsh9pOI8BZuNpKNdtIGSK+gOTfjBHIZMNcRHK91s9axJ2AcFKddvF
pO6/dLUUVAuR/d/mmQmLvVSmRt/vqooQW4jjHKWGgQcRsIzoWJsExinOpCT7qaiFWc1mx7/XNOF4
WsC7eswq4tCmEnAGKsHYh8uq8lhzFKztSAfS4akUPjbhtxbm/kQ+65nwKmZC0jdKX7AfIJAyvJml
jbHWjN72OVcPeNDhX9m4A2fvB3Q8zg6pCVGZJliAX+PDJC//1UdH4KqWy0cfnW7lBQrmsu4eXPuz
W7C5P41EAJSGJAOIg73lLmh5ngitHQLhuGDUhq8F0S3Xe6TrqNnZAsF+5OfM++f/018xYX9kMelN
MBAdR97S460iixk3vTTdiwNppkgYBkGi99NilVSw83dn2X6J+ssg6Yoha1AntahzugNdWyH5HKB8
i3gZY6I4jvfbv2QiD97b/Fr/cGVRLiqnDJtQdBPMUDRZDBpYmdO4RmJVNmy1GVLDAGi4vXYscdEo
TJ9tHGLdj0RZ1ZiF3L8uC7dB2QqnOeCx47rPqrI90juFCUdmkxsxfSI+Ilu/tuVr0wt+QAQEn6zX
ynFACIZxgurzYnD8Pn/oG2GsKjKtpYKapyaIDP0l0y0syacEq2wZPOb3RxM5MlLj1Ml0aJPfVpWv
N8gopHbSAv+fj96Jjszv8ngaqBkKXZORVR1s/uNP4dd1I+mX4atEKIyRRrup7KIW1r2Z97dplxp+
adAPUxOgpEqNRNYYxDIDcmocyWPVS0KKwFh5HGW2tvc1vGsxlXM+EtNZiquwhSHlsmTaUv6UegWb
GasNsE/lpzqtPQ9v2U1TFiobwSLdzMhMy1lp8lvFJY6NNgd09O3TZt9Shx9XyARTrp5n5FnwYFyB
3aUuU4WeRMA7Lw8OxqpOOZXIQt2s4vYw8TP5E9ZCOYvUuqUJjLu1CzI4efbmOZ6AQKXo4NAh0Fyb
pVSM2OgMDbfiZeMCEseYVzJcjNbkiO8f5kyFFqg7B1rmu/7rrf5MHvSxn1GBl5lMp7wlG/1WvBCo
Exv+y+WcXXaGetsZR78XOkInt5SoRTtenRZ2Y710RHDDczzLkeTBayeCkjCFKMMFC1I+eiyRLh61
0yy+pg1iF02KTPoXVF5N+N3/AAuYbXqfCfGOghhk0Mgb3RIpP2OEiCF0+VrsOKulfpTziphCN85o
fKdI1Z5+7aerydkiWSUAQQEiCf3bF0rGGV/fg9Y28/BeKlRM1fCnGf1La0z4rhXzHq9d0Q+Y/8m2
ZK+WgIshVp3j1BXh1f37qz9+TEGqtIGRK3M5KcGnd4AP5QkCxQbGHl8Orj+ymci0UhaIToQ02S0H
/qJOfZNvQdCuCnUuOa4q1Gj6o5ghKjF7XQniK7nEHyqqgxV9b0koXKJ24iwCoxPCS3g9a1pEv7mJ
4xmskw1MvNKkncuViEvPGF65HlpQTH4ZPDUvI0IWU5uxmjvX6mzLRrj0U0UEbDPE5PC22IK4Knfh
0YqaH0y8tldhtqnbDhdHJjNdFNLjUDyr3RflnqNqjt929ofFPbHIxJjYsKOxCZtxJSI09soQ+dw9
KKAEjJ9+/k1A8M2HN0VfF+1EGRD2T6yaL94hk36dFaToyfNAV0M9A5JS3naZtmpARlTHoWxm85ez
RGNqZG0GbtTl+W+v8zl05I4Kpzi8A2haPfc0mA7NWdf97ebIaLnqwszo7ys97PGqAtAlTqOd7aE+
Dzeq+i8MDjq1VomLAkdoOS3VP3BdRGzQPK5meAvfCbT/ii/eilbosPPn0V72z/BW8QO2SJBceNyF
zozlUt/T8z0J020FgKOzXKIVpyaGPt0BNklP6Gom8tZbCtYtnhFzBNtU2Vr48p8QOLmH2ZjaXKFY
nYegiRCZR5pKLnAjkjKV18O4lbl4VM89M7SNfCRefMvrYfeMas6tc3h/hu2Y8oWVUu31stdtRh5z
BR2LY9W8pn3aJE2tmAdj+g46wgBa+KttX82Yql8KmDNerMA7GVMUbvjWFCtT/jA/e8Zq2r7Ks3Mi
iHyP7ELMgT7Dr5vjPzfcOF/3+SDA3tfeasStc3v88w9Tes0FuHyPgbJolcQC1jKoLap0xFew9/N2
emonKKT3OA7qDqIQBzcO+sRjG+kcKf9cqPURr/M9u1s+EVSV49NRB26+jQnjsxgZ5hfmfGT/vvqo
S5CLhSD7OsRwXqll6REhTMHSYLqzHV1NurFY1srUNzakN5zwcUlZwHgctc3aYRcDTplrbe1RPv/u
ZxX8PtvTK1zHXDDGA/V8TCbKeOq+slidxJFUMthzZ/LyfmnZnoqz6Iknw0lLRYbxTX93zYHM4q9n
719F68J/JKgQcLX+nykzrRspij3246SZjQ2jdUswT1CR5uD8u1N3ZuvwYeV+5YRx0UVs1NXZ4XQp
VCUjJqCFldrsxY1+StTOPWZ0VbnqQdU5+GXru7cY7RzwWCswrX+0d1pK2u9Ca2aeyWRbDvdtNpSp
X2YBytRpl3xtgDNCq+yT4Rc0jn0ZoC7HjxcXBoXlgx8gwAgI/Z6jfmxxuqHElac7irsmyodQIEAl
Dy0XGcwr+wyNDbv/iDVp98s+mjFzRiSKMzQovjbeEbu0vyphxxJhZo7oMSwYkIfS64trbR0CcVlI
dF5vlpG53eDHajxCrKuAC7zaRqQwusE0+MV+BxaCU+WqHCSoqQaZa2YFGWq0sil49ru6afkG3a2g
jFH8TRODwad1ImAOxZmMXx5fWsckF8zkoCFvlV1dN2VGRs3D5euwjvDV5aYErvmKOqso+L8nSF+s
xTprxE3AC3oZ2BE0XOEwYA+Jw8v3/sKSs8EgPIzC80Q5tSPrJ8mYyLfbLMGJXnAd6BsoieYBYpK4
qmRpmIh1obnAhR4WTK1W4U5//qQZdSSfVJPCEBLsYRKN1WOReGkxvPCPLn9zKE1bkNRxFxwUQpTq
xO8bYMgg4NLkgZZaBKZZzLA37YE/hffMjOwlJQP6khKn/KVMFS55BpQVYsT0xmmNOpObLSXyyNm1
ADL7nvqNlrlehAp5X/Jrgl3adMZn8llGSeyn3CE6K7QFzl+B1Uk4ChT4WPcA/WIY3JBt0Gq2kQW1
Ho+ycsBb5jVV/93YYfkbluB8a+V4fGdx65U8WPs2Uc206fnxzZ5/UtJM/6ZsQ2MeAzBhsQS9b+Ld
YZZqyBHZgRt2/9fRtqJwvL9vI/chGRtAI0iEjS8snpn2RVz5qx3ujUN82IEaVIxYcX6h+AvC4cN8
6RTmRSBTGqMtPBmxL1dxq7//d9x+hI45Tk9h82SyxJxxvT9H4RxaMais2ySqSMK2YHxLCNhIC6Z7
QwF2E+66BNoC688R5AVRjrXlQUj/F9qskKDWWb5vIYEHSan5HR9gT6X99Q+y+CjotuVAxKZ4bVO7
+ibH1yCcOES+0uDn4+y3UI8mRGlQhLjOP9KjW1pnIq9x2xmK4I+icFerOB6NrbjolvdcUZ7Ri+hH
wkwIz082qRjmbaa8nOHEuj6WoRIWochzlfUS54qBvieuT4GAi4DHwsHe0Hewti3nZyn0XlulM2gv
WJya101pIKyg1npMNHv0lP3Z5KoqcUyFM/U/ONXvD4RzecnTGXBVYHNWBYz6Hxq5bIEX8UBtHY4/
mHDS/GU8QBXyjCOB1Xp3WBBY1xbOa67bC3C3kRk7VynNrqjGBSHAPeKChjlx9Xu5D+TvSxzLVkTV
rEjBdJKkLnxg49/3Nm9TCMhsEzlyj7FurIqyihLYf3G5vAaEaQ+DtcoxZHMlMfa9darv4m+ffOvw
7cOFk/F+n3UjiD9uZ5lTiCDZElT9xxUhQkQIdzTxfZ3bn+HQm4b4iBK1ShKffjHKLan1yV7sCf56
zeFUeqJzIGidvEg/AQ6GKukMn1LEusIWSXvh4hhJ8EJ7FcmzFV2kjK7EOgjB8BSGZLa7sJ9yDZu4
/Y2kygeMtA+m4VarwMc0lFnkf5ySFvBF/s3BcAoIQ67FkN7B2wuZOLBhLUeNvzc6qKz3gOBBp6Vc
tJHhUELR7pDzDNbNAOy45TrsKTrO2XTCTsv1Yde/AFkbNaM/H9/F8eYbG2iHwfm3KCrUID3cK9AK
K5soYV9NAKlfOTXFKiHuW6MwHkJFEukUEzffPNTF7HS/a4hMd1I+hkCfz2ZXoXIo2nCi843FKb8v
hXmZfoMvz/cb/yFgOn4E9DDEqm6Dx3j5m9kfdI7BxvF1HH2XBLgMcew/4HyG+N1bINnk50I6wt7/
4xQciwP1qKVRUyVKd3teAiB2yTObw500E75cWBCsloi7KT54VxF1n2o7D/DC9g92UKG4PPQYJp3H
7XJlRsQx1eJ/wueQ9kySvgOd++n0aro61nS1NAdHBRl8I6qr4qNDklabyL98vagHIPeakHJd48yl
8ScMCAfxu0USnOuA2LCemNmngF9D28oYwF0r/l1T3Qk7uq5nFqBEdVzVEXj2I8Y/1iiKjCTNDUbV
hhL3fmExaXGDTkosPuuiZPWC2aGEKXJ5FTH8886GVannwXeNUf66xEQnFsRHXldF2osDVz9RwYLE
esL6cRUpsXgaxklatuD/GltxHwjSW5t59Ouxt7xbZwLfxpQW7oSH8T4Cbx6d6mdpSDsbBTJZRqPG
9KyKmDc=
`protect end_protected


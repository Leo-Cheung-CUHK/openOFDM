

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
lqqBNStVsR3PNN5bziChXF/LcKrLaRf7JxqwYLuUUgGOrNZvwy7lLoEJLnGnCpziSpXPmR7X5HZh
Xf7J5qq7dg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sjTjs/fDSJPsCGHSUS9EktJY54hEhhr5FYRsRaamLL3dAsvK6gN44Meg0wVvlVprxMceIl4leIAC
7cb+AETnsSSaFtKVBSShhsh83FUt7Q6IT7FzoD0+4e1cND2VPTvdlHJl3OIgU+csWJWLso5XhnQM
Km5aXV6+liByXYjxBlw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YjBoA9Yu4nJClK9h6ZMZXAp2BeaTIQGH51jfYjEYajbLR+tQu4dfxo4CikZRJV68hbbXRLqZzfSh
ggVaH9ucrYRw/4cy48EzetUi51++4snJMp8ALqNUsVRg9pRUwesDZEOCdnnt3slJwOytjfZ5yxtf
38pORyxZabth8ZeyswkiaPckgQdMx9MrkGD2S5+VIazy0bwLzu+DLVjTigDjnRIqniD2XaKbCq72
kNEKKAlpiYvRh11MyswR1Xws0I702ALKOqxU/VS00SFZFoydC7QdRae5uYXazvF8mZzOl9CALNBl
vJ2hpTkJ7ghO3/W2Bh6NXfbu8jlJKouFyerhMA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
csg1sAAi9ekVxKNWRnvp4HMb5FavHQFGQHo0dQ/BfpfYnbHijtmTQBuyFcIr6XSLkVcZaekCcTgn
sxt6o8CAQ+dAVat+GU2fdIyF73YkIhJUoGJOg7+bQiook4By1skbI/4w6CYcAJNcE5zFZwDRn+BF
BvWDln4mF1fXpqnemRtnjDgSfxTn/07+juXUrCBe3PHxVpGHoDrqv4cNmZjjgmm5QnLg5Zkv2+nM
jQye0cAkvWo0u730NNVF0BKeAKueY7bTp3PHqwMIJ+KubW9UHwFHCe30ckIZovWkHyMCrnpsbugy
169krHvJl0JFxOSpfqiRyA5Xr4lMyRz+RDtW7A==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IZ+vMR9DGAouuE8DO3BNgzsTDuvZ8EeC2H3I1iPomGu82ccQzOxvZTxH5DxQ3v8XXYqmmmxzxOFM
mav52EPAZJbm/ehY79behAoUBTL34BrDTDutoNzPXLvuIvHv1vUxlSliGCGGAnaOqr0+LmmS3m+3
RMb1kJa4r4ybB175qfn+GMd7jEfLzcFnjAuI/AsIa9psXzUA64KgNDUAQf8214nFk+j/+I5Sq/Xx
Dyok9Hg4fO0JDD6GupvV+ZCpbybXnIdt7Oe5YMaxFsdUKp35jjeqvUE9aUIwV4sP0134naoZgc78
Cq+bCzvUKnqQCbP+X0qImsQB+ClLthU1s2mRZA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DvJd8QWvZf9rXVqd/0WOHtl+sZGJO/U870wsLf8uyf5uESXWJnwRm27XK1Fre2BQVYuNp+iN7GYj
BqtQ+Z2vpdAeyKSBeich45E/CuwFwA+qIu7w26D1yHk7YXxRBt3Ol/EtDpVSTYHrp40vOKKrKFKM
mf/F+UNM7/r3BT2Goyc=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nMMdxBwEbvYKYCMPMAuls4fVVr7ptrakIeQGq254dA4Gspt9kBulf3iTJwLztcHrxlQpYR1q3LI8
iN7zLWBMSW/7Ed12KIxwoab3ymANbWoQDXtNuDrpN9fQzQLzgYxExm7SkBN4dqsSEaGifwDQmvFz
HOwJ3yAnp7dyud7PS/g5a25mjqdE0CW33J7agjdJH8OzbVBubZPL7IH+ZmnUWliWlWp9xDNGPKPH
h2ocZPN6idOBUd+6ueKxcw1/3jAP+Skrt07T8VUToAkv82Pt2hzTrMat2enixpyrN13eflp4gStF
cB1CFIg8jqe0kyUBET+oYOp5b1OpNmItOabfhw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 211312)
`protect data_block
J5Auf2gkJI/ujrQLcxA2sO7QKkI+SPYm8gPGw/dXSrZ6c8AFfFynj2MGvwvn4loBIFH5WwtKOZrk
TQkY3jqAKhMIYdWrPl1fbcoiz873xhiOUUhKDgFKZjo5TQDUw71SoE143/XDF+a25BnyfDLO7tc+
YuQyYH6sX0HE021Emm3E0/RWRdSMnfYGeP6pPBb9amD4YU60RDX4K0Re7/OPUx1hzwG00XwHT//U
ceqb5MmFEZH4KPClpLcNseRHPD7usRi1VpX127Qoqr+uZs0Z1V1m4b6/0mmDo+7tgdo1ayDTJ1po
wuuJv3a25CxSuNh14IfBhwX+l9gQE4Qw42fWkn0s3ncBjpLSVcw9yx4UbJswaggaX4JWC6wXg5Rx
nJgxESblG6Zcv//0qeaKCSnlO6eLq8cFuTjohWZoHSNCrbkZMYD3S2X1EkgK/U8ns92PqGS9gfPm
zZdiNJ0SKVCq3rF49lLPkfZSFAilPG+/LfKl7l03wUxkKW+DqZkY6ni+mqUNq4Xb73bdl9XsG+90
STkpsBGpBC5HopkXlVy0PV9vJT4hSQC71/QYMvEqBWwPV8wUJFIQIFyhEKeo10N3ocLCDJ9u21q3
LCXnaygihkRxcUGVikijDXRWEvSJ6OPmHw1jtV7UqmfLuEIf17m2jKz2sEkUbk/bhEhEWsjI5svV
Ac92ZD0PXbEOcFX5siQA4dOcU5rm0UcSGArOlzalScLbRCsCigVGDeP/CseRv2O3/jDXNGqPE6s3
zStEgenxO3JF4durKQOl4JnmqRTCp9pzdG5tVqO7+ZvT7nKAFTwjuGyhOl6yf7YUCWd2d65JTCOc
W7RdplVV9TDJIRTZETUw25EegVXScZj7z54gqc0NEZgMmcuFo+sLmyNj+LkLJD+MskTmtgxo97D7
rwZRfuI6xrqKC2f1XaoBPxiSNXl1tx94vdp/SCLVKBJwoXaL0SHBYuvN02sxWo7VffCwpGU+Y/Rl
OkL1vbyD1uxNfhJ8xW2dBjRsHmANyBINvahArp2GDZcUP7WFco6A7vXrP0mKRa2GSBTP28f6tpro
Rc7z4eDfTOkdvBLp47JCXqsxICqW8M72XwUzVlmiT/4W0PbLjVFbyBwjN9vYwPl7dk7x5Ow7Ncf6
d8ADe3snDnCOp/W6+QXUZtjnvWF3YgllQjyZ6D4M4W9f+qbf8O+G7vCOjxFifwEMiqWau2N1q0pw
7KibMPTts9nJLqkdrgELlOX816OyxtCLsSer8kL2JgGA1x02k2mrCI3OTSfdoSVxPZwvqM5L73/r
5/zGBm16mx9WSIXDa/giAZ9daAIQpXXe36cqnK4X5AaHq7VAw27qdvwEtBLPscMMLg7jXAZhIMLZ
YCQtSzjQp1VDU7NYunP/74KGr+N1nb1mMmyINHWl3otMqsXdYM1+WrKRRfQj3SSlBxAJdVi8RiHN
a25sFhKnarw0yKTb8WhNleB0aN6+4LFtv7caMh0bDCHWsIXptg9Ue2OuDk01t9ZwHZ1PYewTcvUL
KLYSaITplrs+BUkldZVwAMTDKC6bADO8BbfB0zD5iGuUGBq6AwG+sJB/YYGKrwuEH4ZpQu8uMJjk
2e0G4K0jdXN9HJ33OK0f9lgkafGc1xafYE1BnV6P0fUURLhVZ2O17pZO4vCHKuFd0SmWGFkEG3UD
iByR52JrMRp76Qd5bOHKw9RmLl8bfRPLMaIDJGKVyB3KkbeM46FsZY1ZU48oVllCEDiZjlOnqEUM
TKKVw6Cf+Ff8hxyjRKhdjmoDZpr1oB11wyVPPyId/H8cVONNkLdEbBNac+1Bz3Mur2feHJagunTW
4xyZpYJj4GmmXxhBvKZGKB4MHOuqtTdH/nHsYi1VH8tRtwqmS7g8bSc0SMW23oTD8wrHN9IYABnQ
xizvRQ5nAlge9FP5BnqzMponCOso9E72zyxXC7/MNXSbHzwwDPwLgZDYcBrNlYtNaHRnz5g5t4+x
kEkQxJb2jeyHj/rJB0oht4iOSxOPDMLswRvPlavxLTZ3ilrGU6R1Jydg07Lp6NaIOwkTYcWiBIb5
Ds5JG6Eaf4Cn1JGdPTyXl3GooFcmbpm79vHbkuXKv+UEZx43YWym7dGvUreRgwJJiA5n+ocvvpmv
j2/GBDe3KGizui375oJyabXndAWD7WFr1Bd5Bc6VRR88eYGZIzjvoNxiw7U2iD4Ka8PHO9aaObbR
TfovnAQaGC/HjIX+DziZB5XFgW9+aKVwNmgeH/s5BC0G5lBm/Q/A6d9CdG5k0QfdJ8AMivVagaw8
6FrZ6b3b4l6KulVwlbLMnOoei6kFN3XeBeSQGBJUoCTnaR8L7/kM5VTNz2U3ppaHDeMG23UtOS3C
nPHdPKFBjOhOe5Dmr9bk1X/DKl6EDbUdT4HScJtbRJjLhTAt7aYLJFCChNbnOzu4Sqa4kVIchAhA
5NnKmhgawEoeKhV0/SBoCXnc1dmmuIaP4XMZv9u2kqAZb+sziC8jWWIW62JUU0beXpGl1WixFk3c
dgChU0VAU0rpdeuDfIan4WOrYl5x7Manq9frq1oQiw4wAzQXFgfW7wkSoJyyAaW5eL5EJsl63qng
bbJPsJer+cDJSBaiG72kPfnnlqDuUusVHslzirxLxOgundF/MqpllDrrQPqopDfxjmmZcWLngAA8
/NYUcAB7BdhCcSuJoC/WPG6aGofpIK1Um7i2X6JMN8lW5NjETnMSYv6DDCBWVIcHAtGExd5Shpgg
GMdQcLKZOCUbQQwb1BfTknaLHXr4EM828JB4DM+UrRYi7Jh4G2fWqyK7afFoog6ehTpikTZkSxkX
9QdxL4qxiNMqLiVein6EHmmBHQhpBJhU/FVV5MTKUClOvbKfRCTGJRFclLYOI8HNWZGjcc5vx6KQ
gcpipXfbyItS71Jz0dE3SFlsXpZ6DiQh8kI93akctYuDghJ3ntkCXph4E/q7byK//bl/ZsiFefeU
NWgS1LprbqjBHY6x7pipXCYZDy9v0ISESyVr+qeLz+AKoKLlenCm/B0eg/2nHVi2/OWEwKwjdpmY
R5HktTwB9xL4TqO34jDDTnlysMCMHIbN7USYL/BKHAoDyqeT5Bxc56HglfcYqUDF2MIQo0ubZbYB
V1Kt00t5EyCPBBFFvwrhQynTMYw/XWvdsL2RMZuM2eqKGiZCxO3xx/HHnv1bJ8Ovq951frgPg0IR
w/A9/EfroNI/dFCGXIqgJ/d/a6wqVvmsYUYRlhVeAn1eORGmMDbcPaV22gM56yhzDQ72N1+YedlX
q1zDejR1qD2XmoINydCCE3Xc5Srgi0idjkkbo/2r35Wrx+yVtGoIkMVkJWyC1soBxguKjT5W6TNV
fVYGFooONF6fHOAfPHNBkDhemmjPjNhsB88B6Y9g/RPELdP3HR52px1umj6SI129C3pNb/pKZp2Q
kBiEhdVphmAs7RaZEr1sWnyc6GpuFSsQM4mJcK+2w2c4ax/54Q+5w9k1jCvXB7xyhLUeS36iPkN1
JTl7ffVsMEjVoDMqJ6dpCMxo/qcp1kms6Sjqe9tTH7bp5O8rJ3DIrWKtfZ/hZQWYbo8ckDFhHDmc
sXipZ9Op5cmsgVdMZmChrOBRHD9b2CHtacwJBxNTe8yzbIKHWT0F+VIkQcLp43jE8dpZ/1RenS2H
TaPOL2ojL3jqpNoQqpJ7l7IknMmpIr66s9nT24ZQzc8yCJj32+1bJKdsBIMFNWCOaVCNW8etKJYT
wu4SbnMdTnQEN4qAB6G68XkXTpVfASHyF1zwCfOh8PIbpiZU4RS3vazwtBLpyXYBNPDepKh2ovdJ
5GZFiW4HjCn2cWOJTrsu2MpsCTkRM1yr9T5NZAmN8fnlFGgpJ0tX/BTikJYDwwQ8LvdLZ7EcfApC
DMnTXz296ISy7iSmbwAFxMTPVgrsOqoBGBXi9bXYRCRlq4W6pKfsRpyS+X6NdTMt+bCPm/lDN2dk
12Qnyu1vJIptsRPYyDrW0hX47V6kkftbT3MIMVgXh23zaXDrcNB34YZWZDDShtJkzEIZrnk2VBXB
ZLYDMJmZNVcBYrO2JvECCvVOlXDlm7DDlhLuvzgo9Y2Ek8LSgIdigfuQsNkQCnx6iHoJdICyZqDr
/a5JGHldSJLMbHRk4loM7Zcxjsy79Jxbwk1UIPcpLsntgUhe4ZC5vwZW7IqUypJXNdRTSYPpp/LT
HCU9c4+OgMZiZLwIkgfOABNxIOCch86FzlM5xsdG99eQIf0iqJiQq6R4cwa5SvCtDPAgqmKilb7m
zH1XP3YmQtU5bSmY832Dl4sgvunfM0xCMrYy/zSEziB5u14N12H913vQFAw6bsCqWSrBpxoNh2WW
EXiw/kdz+0TLb8R5DFm4R0A39HW1yIf3zcwlh119+0mf00QDICnbLA2/15HO1/Vj6zG1Tp7DvyLs
EjU+UuALai6QDG6wBfavNbNsBLB9OYDn4omb/cLZAForGZPxLoECipCfstBAFVzcVVmQlSinTxp3
3sNHWhf0ujduX1ZxbTtI1nXl5JA3+l+AmzGTLUcPFHpLxnia3ss+MXxtjoIJk11p/5yUqsM9KeTg
CDwbTXcJaSBah4NM9YX/X1dql5Kctq0OyGv7KDcMARPrp9xy62C7+6aXCD6OwvvUFNh9ZLbHZzRU
OLrTKlZV4sU/JbmTNqgQxsr53TEU0Bf43f6bY4eQjbhTNlPvAdYqL3NcFGTTCgsA3KOY7lnC9fyG
3qYRYeyEo/v7jXbxQ0d5LlBCapL3u1Nrh1Cqk92aY9f55Pj0lVVYgau27BDNrpYr/1/QU2QcS/B+
uo1Az9wjl7HqvKknyZOIUqvqixlrxIbHUzsSnBHmc9PrVnJ4RGM/fWXuceRvTCoVcD9FFwuzOGt9
G63XqC8jVHURQx3nzLcFlf8krLA64hJ7kBgTN1wwd9F5bK8qOnjGpq2BwOE3nR8C5arWf/72TeI/
vk6mty0edauYOzc7OAslbQHYyFcMpXhAtB2Qm/pu7jfhT3BCw4CzKHboMwK+H1wFSG8OHJiJ/qRc
PMxyrN1KDVPoYDAxjEAj+zioPfqpqrwbtXSYKOa1yhNvccmf+Wr5deXgRt2M8/Kgbbq4YDHqWOxP
ey6OxYajtnhl5pWkwSED+/D67h+/I0lMVhmOlxzC/T0lDNAdwUh+oOF5AEPBpvRSMG5sEjgvAlyU
oq1Dz3PYrEMSKvbU0XzV7YothIpdnjvw3E3PHDplIkq4Ok6het+xRIZyWJ7zcCN4BgK7usVivOJh
egrBhPc46eyDSdHmKJfwv1FJN8CVRNHh+edwjXh31zlHMbnK4sdRI1JuWhOv7aR5hXO9P8gt8wB2
EjOwJCDuyCKy1rjHtVBMq4ftOFGQ/48FITSdazjH2XduhlGHM1GwbLF/yDc1ro2+fd5kirIRv/wh
u2SEEKJ2rgSJhPt8vLDVPJBLONKypPFmTk4y6HYIq+6iTjM2fXJ9o5t6kS9eB6pqVq6+rF+LvXf6
pzeuMGpo/e8KWMheuRgk9roEgIL6wy7F1SZ3litMDQC3FQuaCoYU+Yv5wAKKb7/z8OsLNwJbiPOC
LctLJ05IRdiZaLEwr3In97aVaf2mgOiTHtHUvc2wF3V/pKJ27LbX/tOBCLKak6e1oTq2V+ttY+T0
V5WCYPzTGfWfnYpUTm/AdBt6ZYBRY+9gaUaVDQqYF0CXH72cwBDtKU1pfpBMkiIvO9/RyZtu18za
VWwmhPc7M8whx2YwjBI217X3j+E8W0WJCMA5uSndHQRJU0ktEAfR+7dWjVP+B4KO2Bm0xs4G2zNl
FYFKdBNMucrGRPW20YWgSNBPzlPpAr8r4B36eykGpuGsN5a5UtMvWi5fyMxj0Te18dN/j0sFvV1L
1iegHNzCSvbFy8MIUzKJd0mj/voBnhBINr8G3TUOeEQQOYClI4FtCS3V4wveWCtSnzmxih6qleOZ
zOaa/7+Xrj41HvJ56A9Ww5cHBoqYEZmX/DkOSIzW3ku8jWbubpE9YmnNsFZJRANP7N1FajbkIp9R
T1YfHxCx4CASKXWdfGrPltqrW4kdZ6oJWNRSJdPair2BP6rxCQXz1/zfS/jchRwv0Gkb8h/oCS4l
tOSL1qfrnTGkUaO8WC0h6xWBbPXI8NkTUxwQ0WK92YxEiniod5f/LZbzuqWaJFWmKdlzaSMR9Whi
PAu6yJKvaoY6gjci5htoDknktHz35rwFl6OIoRZnB3wSkabQXTk2zwzuiw/7EkZ/xiLrEyTFsh0B
FOTD516EgKYPRiVwpGynxdZMf7Wm1oxUvskavorM5WuXCXoymMDgi7AYlZBnIY+3cPs9rArj0MBM
dzIz4dP/Xn58CgUOJuvilbBnxhhMBk0ZDNWpvFueH+fbxA7i9u8ja/ybiRBrgUbhe0CqcCDgS5na
o50/8SLo4ZO4t2ebtOHOwawMMN/jVcSOBnlIutK2orQqVI1ONO/ww1NDo3oFu7v3QQ8NxMDIkJvs
+/Vd408v/lvnYQ0SGW34MYXppgFQnA89eFiqRWs1uHccLFBYtkcRnbpYG5x9uFQl4ZR60k9iV0jv
VKyFK1OqKFoYjTF+4h56FYRkEtZzx7ARUrlBwpWxuSTar7BGvrGVhRNbgXoom0HfqrmB4plgB45N
KPI1BKhOJb4Lr1bmrbjYYZc0+Yh+QfEYpL8nx9h3LiGDWD6TeNJObbwTIwZfYkL24oqutRtx+CUp
Cnb040Oqr/PuY1RHm/Q/bkfKy6zGbkuQdVcG9O6brCLcN3HvHBqjx/BRH3d9HGL07JDOmpMJarUD
4y2vx3EEqp6OnfSzG2IWZg32C3NAjyAHvJO07zPtJQ+ZHUpdAdUeIlTLKt5YwE0AWqj6BPeGiTam
mG4mtJLZmOYvO7diJ0w2JFZf3c7qk8GMAyTYEBuRErInrQ5z3b5s82BiW1g7gJ/yCi18951RaNVt
70FDshQ+ZkAI51iV7JCwfLZJfqviwOWU7lPWVSbXLqLOWagbN1qtkP5OILCvD1PPlEXMyYTy+7U3
HGiFq78+S4tmjfOOQch81nzhgIjB+NXTcxTrpnWoo1sN7JvWNTy4ozXGIhD6mlsGrYY/a4W9jARL
WUZgxWLVKJdHioYCDab6omxSR8Nui/FpJjokd7Pgjdva/VprraCbFTGXKfOhXCIBK0P8PZwtM2TI
ohe6qkqCwtGy/ao8U1z4Yltp1az0FCXfYvCO6xARmsgRqUiMtUhKpiW7EyCjwtYLRjW73zXSvrCt
XXpfxXl2DBfS4zbyJzAjnl3roGZBDneqU0g/cqRhjyFNW/ey/Qlyr4hn1i1b0xT8BokuvL0nRP1e
I+QoA5XF0jixK1EQv4nd/wP9LTDYHmqPTUGZBLB6B5lmXLTgBkHuPGuf8Zpv1fh1s/usrQzWMxK8
x5nXufRzl1bmNx8R/26TW/Xp5QtA4UMgg9DKHu6UEXH05wXNtKg9LjiOVmzQkx2E3f7Bnae4KH1q
KB1V3KG5dPz3WsRMD7EtYgvoSBp3+TbJ0Y5vr5Iz+sVoW7cYMGIFhJvkfF2dRm06c+q+NyTLZd1o
iwWdNWR9FAdMH14xOjiAUGfTQNdP/esYdIYhBCX4VP1JE2yAECvMTD/rf0BA5Tj64V082x0RyV9y
sNtqMzY8F5wtctLxwcOUtPD+vLDurlJ4/mqOGuBbhA3C7fGBPnnqxWTtJ28Pq5JLuWNySEDP04to
+tbWOLNFc27gKhLxVpBqzOTDwkTVWQbrAj4Q8Dw39uJ/5msx/nhv070U4YezXeMlRKmOLO1R5Coj
qsXKrm9bwfk9WncjINdf5TqRXZLX7genxRMCvThbM38wAh/+sOglvN6QsFrCc4yxPE/92vGR6yvb
RYDhNJ3qFaPRnlziUW/T099D1ydOw3JeObWS8oJoq+E9MsLVWBiX8YjtVXknTjWHahIWIK2t06FH
2V7PVmGztqjvogD3Q87E0hKl62fgsx1up+CuXe4hwpmv97LfV9VXSI38kPZW4b+yUpXVC5oFxmxB
c1Dwiuwg37Hde/eMsuu8yBqr0g/BOpqCwZZDHogRfPIA+zMWjLgz8/x57izbTz7hZg86M2baKSw6
dKdmlZir+kj7M4tdkppAqg8PZtCRMk4qWY6WcGhi4Rz88e7oHLEGrrcn3TxTuu7G+FzydWgfx+/r
rt2ulqtkq/ZieNhESNK+wNLAY3u87K12GIwYOVwLYTFDQ0H1XHCfcfrKW2SApCVyB3bFvr391oP0
F6p5PqBNHV9tdn1NbLaP1BMdb/Wx+OyE0WTg03HwGDHs3SaxCyHrhTRcHF3ckgSHu7Rt8DnEO47V
rkcmFz0WvM34WGPr1Y/r1Uc9qS1lEWIbQgEQcFroanUiVzGIKF5hik08HfPBNBmO/nh3mEWA5L85
DQ5ajtsb7wL5Idim2lKooSW+LiE+49W1Nt4+vsbOLBI/6PryZqTHd5cXlDHEwqLtmsMXqkkxx//9
Do3gjboOEXr3x3a+HPbC0inCuAeJK3zkF3X7IvAR4khsJsXIsKpKZV5oaCMPHvK3WqEc25uFscPa
YAMuRGWPeHYveIfS5gm4A1vyhdVWJgjLhkLzblvsYVuL5B47Xf+ygArA8gy+3ztIfAhZtg5znG5B
TereNIrpg910mfvzPZwtKKT6GrxyWP/FOI4sq3WjE8PfZ3344F0FaxycT1UUtuiSVvxYzv6n7/4d
ethP1UsJq06KsqmnEOCYya6PoVOy2JIlijhALfmZzrN2V/lxhRuQDl3PgixA98t+qMQEYRLoOkO+
ck8SW4sxizQuY7roAyjgcInrhNzpq+RtzZ7/+DSKjBEMXuRHs1MK/EivKtXVNaWcNKNykWcjeWPu
HOVcrvzM2TtqW/0AYN/+EwkF2N915YGt6bSYYxdYjdFWpYeGUG8IpYC/G/j6DM+jSasdtxx7W6DZ
EvTu7Bitl+XzOT7Cp4EL3TAM8JYAMjMklMpO/Jcvt9LaSfLoLU3Qu29dH50smrrhVpIBGIsO3cvS
T/ditX3kbZgEazHZ3+uJwGq6a8/lICVQFFVuZRzy0KsdXnVsRwsfjYV00GRR4f53C6G8OnIv1Yyt
8cN7fjDDvl+G2+7MmEHlYJiuER65ZQLa4i7lD6kcSoCllNK/jv9LcoBWQv9ypJCVDz5g7JNCQcbZ
1eYsvcdK8DjWqy2l1fw8CWxNZ05PWuWajweDdMMuaOZ0SpD07JqJ6SEIn9BC7QU9XOkpPQUCHwXN
ZNKsGjumSoCRuPizMbo+VZ09GWzcdLdiPflVf6Yj/EZwF2EbjJDQLStf/gq4vVELCJMLmU7FOjnO
JDgpSOKKYhnhFT7viulTLvE8Jdhbpo7AOpaPzzF76wJkFRkUymf1CLNvraHz68O9B7FxVmkVW8a1
maSnZem5Gm8Xu3HLjRNnZRavKnpBhUBk8Kfs3pH2j7yfjWL3UUH1eVhT71ALYDhMwnUDZeaQGd8t
trzVBMDkztMg7G+E9bdUfgTDFC729X8a18zkSTMjmd3Gw9v7adzVXnxXUxAArzhNCje8B1MMZKJC
PYHdw3ng7EzeQNZ8odamyF7SEO8ZO5s3rmxpq669JKvDTc1sssKLSDqAefcFiufv93uhqJOfxM14
w/ev+o0um4sxz5QidiFfS12ptmYpqu3GCaj1avrN2Xxu8tr0/fKQxhFoAIUmgnR4F/m945sMX1zo
5QdjaMr7CVCVMFnFCgY9ijm4mOOvPg8qw8B100shKpFobGgp7aY4D3bIwvpFJZBrZfH2DL71HtT+
yXykHxnQWUrvmjr4SMd4quWiFhM1m9YGEGZCVIwUlFOqYrX/M28tgSMr567rjRXRd3zVcTXkGA6J
WkQvKEs6O5vviWycgPH6p3CXYpq5gukbna+kFqKZLeGwp6Xn22FIIBsgLSoCg0vQ7iGrSKcZJmpx
r0u9ZgL6sKOt/MkMeD1dGrGMNMNC3PMzpYmsLNSW8ntOjBkllY3AADtpIPIA5NSwpsh89wq45phY
pEI9EM0xWOBB/+Vxz4OgHr2/c2Tq11GmNPV/r7m1yKrEkhQKiR4zSKYKvFkNuADNudYuyGq4iD3n
h3+0PMpUE/OqTGrmHChTPMJmKSH40Z1GGu6Cz5deYQqATaZXo2Rk9lVT3FCGMkhxt9RWCURbYNM6
NgnIaJw7IRdJTPSsCkBWg4Uf7tpvssDA6iQYnLEv2v2aMUMqCbz66huecnXf3skfkOo711CrnNH2
XgSEeYcPkm974iN717DfKhf7IRHDfZf+7QqkzcmpSVuf2UetzUbu7VXdNM9ro60LqLoM86EMxDi0
XrVIhqpUO0p7r5e2bFs1T77D8xwCQef8D6JC8LLmGnhF1MN/m09OkUdl3gltbrvBeynkTShcMSUy
prjwkuGQU3KV50UuEcCd2n+ybGQ/Fp4562thB1ZAJZ9ZlHsmHIZI4ILw1c1G2WFOpP9nXBsahqRE
pJRiLL80Ia2LVR8rWE7Xkv+bl7qmNy+hqbcIOup4IbGwBZ9QSJgikpooNtKN+d6gdGihA/ZDCMwe
xMnSaX6SeGnTGoTqBS54Z4DeziDsc3cICcQSxaWhjNBD3++gTAuAO2p0OH8HTq6PqPCqmbdaXel7
v8woe5sggeY/XS8nCNDhiPlXp3uWmwppSKN+N3Fmokhwu5MZt1mCK/p3ElCDmcZY72rampqlafkY
Cp5F/Eeq3IXHg+C3sQUP4qGe7adZH9FN7fic8MdBAScDHH9XOvtY2amDuTydIztWrzxZVp7tTs0n
eV2DwxGuisoZuBf9qHf0zG1+X55MFrllRiskWJ3cVNEy/u9wzsKqcDTbzVCV4RDSw4VNQGyKYZH/
3qekLt9T4LyK2v3aGN24h3/IWpzdDvwzPiLF1wOIIckYMUruw/GGnQ0K1R6a4l08Ny3C/MvY80hN
9bnb2Wcs6kf2oZP8zvty/05V/6/ub5hM77Gxb3f+YoEJ+9oIC8sP4KFTBQZCpu5s/auHG1+oDp22
BNUe5FUoogwzqyTy5JRgiyaiIJGApYExrA2nmkC3wcpn81mPXh53Y6C7daeAYMuG6YXC6VxIIZSb
bGNiOv9RbhIea0WhvmecezHzmg64jSfeKA+BLGw5BPGdugAR5Cts2Zxpz7wvBQMGNA2tWcEgP009
kQqhwKh0Eh9OOsvpE5C6yZR+3ZnCswj+i79YRO7XUHTe6RzNT37UgLR0RfLbIySrMLmrc2bzve2U
sODEbM4nf9EMlMucfXxErs5+qYkvw4Ufg8B1tHSwMJjUWItP9ZAmFAYEtcCdv8DMGaztBYIlr58G
qjVvTy6EXuX9JHlyY06j2IX93mr/9mhHi5K4DxEMM0+q3FpQKdi0IyO7/AxF9NlRi9oh4wPQtY3R
zCW4soYe10zLWNkUcJeAXmUOSDfFcn41pxgjdN1y4/A+/nZB/1KkEnyWeb7P6sbE3LpGz+o30bk9
0Fvkt/Uz0/wXEUGlG7wT47BR//fLZNbtD68h9KZOkoZyCNexsAC22HY+lS8h8hK82fuDl7USfMjy
owLKhxlnq6xaYAokI2VtPHl8vxEtoxLwN1yIviKU0T8c1k0OLl+hzsZSpAUIeZowavf3v1ViNs2T
f2295evhTOCjH+y7h27/rPjPJKUdpPxoMxIEZtqPPfWZs7vGQsjlM0x3xcCf+IBCIEzcuuXe7fLD
0N6PYjZeU3meSi21HiGuwg97y+iw/7jNXSVu+PCT6L4sOFPPQcbygGR///43mYMBtJAaIBHkcJA2
9RcHDZ0YYZ4OAPBQ8sdCe2uSWG5XXGiq4LW/CalwzfwB7OvtcWmZftiLfa11ZHKxCjz/9Lkst2z+
w2xaa1fkb0/dIVokvmY36KhL2TWkJM9aa+KEiWEmcuRTvJGLZ0ogYPG8X/y24soPg538ON+EZKnw
tOlRKBKR5/1iY+/jSrVDzctEXiQiD0tuY9945OuDRZYYAq2kseSx3z0vkIQIvxA1peY0xI1SurUU
rR7WSOydNebJOPfEwJr0gBJYJNNDrz7AfaRANenw/hxBCAAzEWK0922STz7zoVYJBRKb2qaIqjBv
cvpTqD6AKqY9tBmtT/9ZL921Arb/TjvpXobu5iJmkELc9EsxeRNEVRTehYsTUdk4KGQ97u0izb0a
a3QylWF4Umf72Aar7J/VhMoxJSr7EUOOaMKghkZvqCdvnLlvsBLze3Dj9GAUYlzotFQWA0fX+fge
Z1BrHkmChSkpypw183nSmT17R4hkAVAnnV0hEtxjVVA9o6iGJPkEM0IQRphhhSOa48CJ0KfxYtwu
3QQy4Ak+869nE/8CNoX1URXOeFzDSoHeTqdynTvJeImr6XK97svN732gENu346yNKplObqLiNdZT
OxnsHmgNK3NQTV0mCygti403uEFQnqm2OX7MXAVFqxgMhBkpOC0kdo1d96PtkatWZjVi7StMo58P
FCl4TtIhbt+wFMsmEbCu56npT1inNVCvxorSSbhCFmKKT0XTf3QSpk6bHCY2eEsiP+fyVsqTJ1Xw
ZUBecEzAVlFWsZ5zgfhh3MUWZIi1ZG1/GvQd/bY/SOQagq6n6KRtVRAQtqIn8tJ4fwhavDouqBbi
oThDlYVqVsUu+FguXiIx5pDNTgGhFu+A4PjHoherE9v8R2MxVOXEb/lWJ6Jn/2bXEqhEjL5tB28R
zRZoPhBLONBJLqF2AcGWJGLPplAGtZUKp8Dvo5i++vrjVDsyf67tRBuP1mGKve+mUkYyvwqxuiJl
vT6egn2XDmPCJU2WK+4OYxf3HlVKB0bA6saP1hL/dOlNH+oXBQbebU167r+QwkuwkBTsJP2NDyh1
9MALmxplg6GJU6XPLQhTtVy9X8slIzcjHKmPneZakyidJSZVKeRVE5prLNSWgXa1xtV9Z5mgGkSF
NGvmmymEDFci5qrBXO9r+9m/SCpuNh7CrJjHWwc9uQKpO4qU9ejoDWdZr34+8uBa7M6IRQDvTdCF
qEtONI1TrGzsIG7e8Z2x9untbXOMfR78rXtYEuSWGHUd09jtJij9GDssForkAqJqQhXaVtmPBIdY
W4UpIIXVSGNy99lqzjSuXzB4kegup740FHzmUvBuJDShglF50pc3d64/GtYJpoQQMXIBGtLg1w6h
WTkQXyWLQZoo8s4DzNoszE4+J10ojnAVojA+kVykVd3BkXJB8nzJi/2POUTLRZ9pb9Gl+8gs17pZ
WitlZDiU50JufeYGW8YsLjM4XLkme/JJcR6JsQrIjfUoR/XNMDLvIGccEWEduG1rA+8PtVwgcc0i
VGhfwEbrXU9ZW+HM2PGY2/39h415rTa0Zlk0d9WgYGTj2artDcDBxUo0enSPMWtgfdJ4txmRBMR5
SHN6dsmL7pjVWYKOVZ/s9w/tvO7tC8aZa/DBZiyuEAPdhjebeQZfNMEKLvfP9l13YXwDYEL3BZMo
+u/io+c1RU4Cs7YwWemG5UQz+iW40RPYefPHwZSEWF5d2T6jBhCjwaFCOeaj4EUx0Uz+ewhbiz/3
9eI3mFls39SVJ/d91dEsm6IL7JlFJN0UZHUl1vMkjfdgWdC4+d6VnvBMnOmK+Zw7bLsSarX0aNU5
Bmo6lMnzR1ynt2wdfpRd3DaoB6DaEtf+mBz9H4V7DfMymkpj9ZfO+jVifAyGXOA8hYLbTfDugkgz
FjQJt2Yr7dwwjjSmKENnSskR9P+MCRGsYHYgc7yMzDhtEXkmzRfjFS5Y54KJSRbON4xwmC+vw+KW
TMn9MOI+KlL3+iynTBRlVQxR2tNnLFwd3KMvHPSRGZ4fLbyUEPWL9b5G+jravnxJadoAPzh5CWi+
wlAQE8qaYQ+uPyHP/Mz5s78Vuoce3wwWGt8FvYBD4U/uS/LkTGR7LwtMtcbDKL/6I3woJJq1CvYV
e09BlaXqjcZO484/P/Vap3OtCM0ZCldlH43rDIN/fI1GfzKwbdZb6K2Wy9j132ES8n2YdJZ68KKG
tKT6IRdmcieMq03mMnIaliNcKFP6K9ChZ3HF60OSgYfWpTUG6+ezc9v/a8NX9cFRtmQmdrU7zPzn
aZ3Lbb4a1hUQ6gU3oWJHECJ2mCIHPVxBJsYLwdAgL/aGU3SwxGhGsefLtcIV/VZgJNN0FAtgL3VH
4cX8m+rSa8clGIvRotJfZJLeBjbAA1h7yY8C7iAl8Iy0VC6NrsPKsdWJyB7YuLad9CscKBBlwonk
fny9wD2IrcUxyAzeHmP4aCAXK4i1PO1tILqMnoNarNqun4u/k9Qv93xbUxIleGHhUD9Hk0GGWvkV
G0ySFmC47QWJj6ufayR0o72y23V2MKCsNcEYpghxFE52P+KOnzyuB6UWgevQmfxrhKO9yakqVb+l
OwhgPIQ4cV7DEOITV6cip3VOAJtC+/Fd6KfEzocdXXQ9JqQQDHWcvaEdbgzWRfUyJO9Qq0SunnUD
DyMY0DZDhnlJM3dcCygTWdS5socuxrGP0NiSmK74nznkuGinLaubaZ8TAeSp4nNg0r8IJR/V5Evv
ZdW2z/shS6puvo7LtaZK3Z0Sn4paBoEoB6yHgMNMTjK+4mD7JONk2Y3BeybhIqIof8vF9A1VBpVm
SRj/AsoDVdbQSwovZdxiKFzndlXKx/NbSkcLSdGDQ2yrQzQPiIZZDIJgyFYP5NBwETm1sY9wAY62
1LXpEwePTGgjF10DBH6XsQz4+P508MjhT2KVID0hfOPcDfXFYDGQbeIa8DjOAFexr3nLUH3kBTmo
ZZsFuXYK67O8u4GNiAtmDoz5l73lfJIVafszW5hbkWGsChwdSmoA3ElxO3cbGKlEqdj7iFOgafPX
aaBDWn/DlBcQnXoc95yCCi3hlrkE3x9omyyUtnBXJbHkSJkIXKuyIKREOUDs+rY2fD3fvkszStAa
/2rpJMjHshqJaAzL5w/x4xbC8de9C9xw6kJWqiYthJs5XB5USPGuh0eRmMzbLres7Qsac8DxMcQc
bZewvTxZO7MQWyNAQRQv8V+COa4it7iiI3O8m05cObEtvYiSm5Q9WNu5lUgeC/muIda6GqvcXSS6
RHuSlO2j2V1Nqh+t3bqMuhGgk2gEKmAIWmrVWVCeJCe+WSSS4HEQkLMY479vZAQt7aKSORIpyCs9
9DYssW/LV+Pz9VkU8mEAi7dYwTRw340lQ76/JL3XDeUXegsmR6PiSB7jppf/5fp6Q3WFcX1YZEKK
XpcejmNpqwjTg1kEI47jkQtJ4XHCJ7Zcv2Vz0jFEqeGxAfVP4Qc+EvCwIsxJDvdHsaD3l7+GYTrQ
3qV/bLtgstHcxZaDtgPPytINK6pA6Eq2yKSBUWrY0cluYjsxptSz2+hn+ul6qX0aT7Q3l7eJtyoB
lxncs+IQoGEd+XSemnkJu3x1q2jXcXn9by3RW4rOI6NY9erxpdhRfyfSpEHLo3tzy5F3fGlJWmWy
jPTSUieUgal9apoy/yeUPabyp6uVwvBgGgoSYTvz4WikGRyalKb8jEpgQQS/naAd7SOn0YBcS2LL
if1E02H83d/GA7TudVgLvfxf7+aIu2jxzq47snEFIADl8Uux3KM91VPsmC87ibi8WHS4FosRDBsp
Nu//T3ZHnfMjlFxZJFLHxGnUn3b+cdy+UdXHLtfIoLq0EBxcDyXVZEfSn75yqsxB+XHdZejbrlWx
3sXXpcekx/xx5CHa9LNgpJo7FrXeFNdBcBhdaaT3IqoZyMt3YFrw4vUF2R7rmwbnL/qEn279azpL
GGh2poO6CWVxrpSZqMhWwJBeUklSwfonhFzjOVaq82qVqj4f+QH8pUV/7tgERIyz24tFavvNqFWG
70mNmTDsVqmGNq59znxVmFqlBbkc19ffXqbF33vMGv6lQFhUlmoqbvCLVEv1aBEtwg4KsgKCGHDt
8JdKHCpldcwzriWFJXH7BvEbJC7ycUfaEi60dup1EIpwN+WQwQOuGKbANOaOcnGlV12LTZl2BmRs
RLLQ5Hm42lL0m4uQwjTidyZDpK1mNyyFlG6cYrrCdaR+ao5a2rXW5pXTzxgac36zNb1UnTJyakjm
kuVWN2XqcQ/kM6Vakd2u0PwPmAhcpTECFuREpGyGKcXHlnOTXvUhvX9IVUe1JdzrlvJaJr083VnU
F7np1eG2V5eVZQDuj/MF8Y4pGG9oDWEp7AuC1v7/a1mj9EwV0FrNl70PqpR885RIPK5qk5nWH3Av
QEFsY5FJlAQaPC5LLQO/0TX//RvcKUEnjs/dsLnbnooA0tD+pSjLSADdJI/RxhrC56Ls0VDKZQHS
yTLJRVTcQ5vyqEq0ZM+oOa2S812O/9217ygj5GlBlyklTSFtpXiT1hVFjjpvCssjnV/jppjm70nM
+atVuNa5H+cXP4sLxEcsyyw4Bc4bQfQtDrZT1thnB46k4o10Mr5XqpaQo7XSSV12F9IUxjW43fK2
vZoiRIZGxI0wqbysIIAFIk911c6KPTTtOrxnRcVWIvKnVzuCkgJEyi+ttK0g+BSKiE8FB8+Bb0UT
RP0yMb9bN6NfCNxpU3cQp6jMse0nGvfkgJzKkp4CYdPF3xUOc2VLcptvv415XEC5JeC6yc/zsq9X
OiY5C/dkffnsWUNvi575VTsybj6GMlBcu5XiGeEAQBoAQ9JF0WF/ztqxb968E5hBPBX1EXowWNDO
jDmVZmPtP7FXmbucNPG8hkTc60uZ5P14xL6HCk+35D7cJ3Z7GK9rtw8OSaltyYONGBhGEGs0/CXa
2tvz2yBqbEj9+rVfQQ5C7DMSy/hY/z8kQif5Kqh9KzXbzXTFLYQwBG+r57u9Wxw3HRlq+OywUw8O
0T7T0AHNQfOSCsYlwhlIKY+HgJIY/qMhpSl358r1FQTrbjlzw2ddILa5v1bX2qscwh/JRFudJE3h
vkdsRapvyPXpRZlYnRLZ+NpHDW4zRPOUJSujV1B9WbL1cAGBmkdCtsOf9fH/pwBRAi+G4nCkgaIS
AIQmxGE9dYL/MZMLP8uzFpGzgXRi+56hxwWf56e1iHs415IsZ6aVXIpVS5PKNxSWMfV/636eRp1l
zUF5V4bmozpqUL4aTZo6W/YZ+TfzQBaRXzpJH+FQ3tGsNF8qSjANaWLwxQr9lIKN+gBDiV0exmTC
gwhvXOnh13R5Gd+e+589SFXFgu44skY4NNSiDytCXD/gPKnv+e4TdjC5slpG8rypSHea+SD0LjN8
O1QchtEZvAIUVSUyBZTRkWkqD1MBJE1um6O+Ltp8XSChuychFFu7tXT5ijoASFdMq2Md6TQcIxzh
ayaxdvWueIRfiCxE/EXagwKJB5H+Ck+h2+KBTtM2ovHQQotNh12HIU0Zu0aKOSK+6xThSIHO6tos
sOhqPGS+M6nRnhOOljebrdccW7D25TbEESKiDeumWGAVeINisYnDSxNNK6lQ8GuMwzVOqVx+nBFc
y3XvEXE1ff+4Fa9Zn+/MJA0lyQW7URsypTrOSHhTCUxjAM27QmdbMLLqZb2TA1y54h17n1OPaQSB
99kdpa9WLvYWxLMYG+TaibXyyl2g2DlhSV1RnXR6vP5WmUoY2drLEE7czTc1Zi+zTgV7v1nKF0P2
IFs8UDLWzATmzbExhDQrhHqiby19qnLMmYwhnRVE7MF4f0hj4HotDb2+pWw5E3tdzOr62m8wIqdA
RGja/dE9e0WBkMZ9jqS4pORcP5x/PDHlRttO9SrSYEu4ULN8jBO1dnKBxEXrxx0zxA7jA6SF8lAG
FoCQU845D2oiXcj9xhUk5OHllEus8KjyWLZqCyBd5NXUE0BAMZi7Bl4KVQC1+B6JQp1pzAeqx9v7
fRTMehOpVv25DwH9wDYU8zjMDEYq/jD2/KBKYQoRbr4+kr8uh+PVpBY5oJGYdEZ3fiLzHrOKhekA
kUFzkaXLFxkLzcsKt+ZA8W9LxGmdXFQYvUibPk4zsRPJjsDfOlCrf46G3zaJaCIks/sGBsCA8dW9
gCKZgr2UIlmY3GtmTalL7uE50koNLaWeZ6hVAExnYqjfgrLIE7GKckMqtNJ4mG9cEoyaenE2+bqi
ZPEH//Ok/JMz0sG2M9lSun8y2lCJgHhaBaGpFpD0YJPZ3t3gU/l2q+tWIoMeo/WArhqP6K9mnjZq
L+wBUUvBs98AQ7NZqBkhYpaauPnou6yKf8OXYbAGV9UUPaQ7GMZD9fuBJESB6UoWI9XIc8dWnfcX
XEHH1FdXcv48YwlnLw69U8ef9Bmzs5pRs6sd/Ya8aO3AXxoa6Zq+D52giQTLSafPkrBhD6WQGzVU
nOpzYqEqGoSdaGWGSKqtau4r1m24WqAS9MKb7T3cxl5BlzZrtPJZQyv1IZHCZGoSSFycy6euiSpP
6u6B0okGoS2aRf+TnOL7qWenXYg7oWbIOjauNQDwqk+PWo9VuG1BwLkm9s/ArKDUEp+qeUbmznNY
EgGnQmcLKKcWOcae1qhG5PrC9uSScHJuXSxHkLFD3v5zWkG4s1B14T6GB4NNhrNxP2DT6b4uTmWt
/z1jfcb6iza7VZUHwAZzEbONPecGSRrZHyWkMG2pfp5RyqU16bfx/V0q9WClqn8JKdIBRPatPt52
zEG0rqvNLz+9lpLjZrowBLnsBH6K3+wbnL9wwsSs9NsWldHQ0oMWndVMJY/U3nTkGxsSUqM9um3n
R+ioz/5xXHIvJuzj0MgJDeC5uIIzRIfyLo5xMjA9ibvCOCBjM9RbPzUlNZlHuPVL2tZXbFmlSZ0J
AuZY4qOXLaV7hOXt+pjqmWjXUhpw/JStapEAYzQ7h/FhfzOyOQz73768PGxA8Kz74F84Qcii+Dy9
1ysnqIx8Ca8mCD5kQUe3aN99nUoQg66dpbSMhbu2aIC6zwJzJyVlSX1c7IAotJLSiMjCMvGbf6/0
rwvMTXdgGUiyV/msastIkObO8bEEpMpQXrUcsvHbb1mOhF14PZVVmgL6rxII6dNpod56c2BwZgUk
Q7Qk5lFWyWUPAY8RraXhk59Kz0U/cH0xmOzMCGaqbTMjoiVHTn52SFL3/0DIhvQRVOalmLSsFPo/
pTRim5NjjP6aB7rfifS0YN8/zOTx967Ilc0A4OhwWb3Y7Yu0CKwodhmxmQG1KHMYLEA6tLI987rt
GmAIirGJ1qei1XeaQ+JeLf6djCe1FSznE26wMYnUNpgDraBXXJ2WJuyyPYwp7QFjqWPWRSI4UQFx
p8hFsIAW+khd3erVgVTzxtMsiqiHkGbwoVRjCNFbLfXhc07EdEtDHThVP10ntt1v192VLUzyLQ30
rwFr1VzYXTP837vdPcjDcFc8OxhSUv/tz7xYu6yM/iaFj6PIGqn4aK5XoPx0QJYQLxBWMxF+wP4k
qTYo4yjn60ZwtKclz3giARXzDHbLWvh2uR1HgFAWQXVeAkASdYGA2/F3IFQFoR/LxFgSXMQCyyDB
XvKf4oc98WPnY1F8XHSd12g7srDgPZyBU8HfY5VwhguAZxa7uSd9nTp/mPXztDw0MuAHqXbZsTfJ
62GavTykZLfCRz7zgiO3Vl8p6GHOrKsak/pgciK11gqnE0VE3AqLCdmTh2S5xjPkSDUbb1y1Vp/X
dfkgvIN9x/R7naSeuRpvhwrkIXnEUWsnpuRHbwYWHd27DyiIAlZ3V7YnNBKl76dMWtMosnfZnVYY
H4xp9vi2VF9qiDn6mZESWz0BUmgWvpQ7NXJEm+4veGPifWE+4p6rhA0TV1cO1zCLIklFXGv+Wq7Y
/FBHjh/VLWr5lXsRGGbCX8P/XHVMeC7920BJU8QgHsLIIuOoq363XFeYPd1IQzb3Vkgy0Vz0G+JX
tnpB5FNPyxVoef7ogK8iKzWfmFV+XGu1+EJXNpHG5I1gH7ailR00S6zjL+gyp18t/Y4x9Y+unfJr
scPljJ3ichmLty+JN5OBE2yppqelu3Nw2svqcqp0lXWy3J2mBtQ7KBYePY2/SjCoxNKwMZtB63aS
p10zcU2/jEDbvPA3wF6HmocvHqEcdptpVZkuo/+FMx6wCLFwskspJ0alnz24A6vz5YG6Ut3Oi+ly
hMwneE4AfYSE0lQ8kBNYejqEMqdmPveaMpu3K0IBYlMUiy7fPbo/aTe7xWVxFNKurSVO2KkEVXDU
ZuRIypH9PEvb+ndc00cZaZbNWepC+tiJ79KfzAXbqHd/TCumcZFu3Or2Zd/x6OvBWbe49Ka3OiXK
5ldLHs+X3rXpvGOcDFYDWl94THNR1mVgTwt3nqsYhlJ24IoxC036ZaaUq6XnwYig4whIi85vZJwh
6TrlAjhROlVoQcxmxm29gL1ADk97RATfNZ1uz6TW2fhVM6+F3sQ3zEEydgtT0g8LGIGdJlDzDm6v
BjMG1w2i/paVnuUtK81ZcjR6KOzCzNC6kxqdjgkEtvKlVDrp4nnaz40xAcHtY2xWrj82zHudeR1q
IWWH2gHy9iOr1ymLBcL6q0rEhIC58jC+aqBBtAgqvhS9IZXrey41iw3Nr8pJPPrZnt1/3kMPfoLR
eHgKJKvCC9KlQ6Cp5U5bZemYX53LvTEohJ4bQEDiqTBxHjSBFVLKkxAAvunWYu/gp6f+DOJfJA94
A1hBuDs1aV0E58sB8mSWZYNb0L0+NvIXANMNBkxL2uQiaLVr4z0noOAjoxhdj3K3JDCdn5ZkkLGh
cA0eexvD9MyWoUE8cvCEZHTcfu6Z/NhRMUdH2waIFfQEr4YlyiNPvWgI15YpNK9BVKAZf+wcuLai
LaxU8fvkYwOMg8YXhpJeY+E8k0MY/6AvtZKpohXxZlt4JwEKMvl9YNARDMyW1A8rcuKp/kcJRqQn
CjGEc1rXqU+G091z6zJt/v83jakxc5NpMwIUzD1VnDwshoRmwwK+Axfb++sm/H1W/v+bUHs5gSLz
3TQQiHx/1ZNy1sPzjLZakpqCjgMQhO8kcEt2kX79MwbWZycE8uWOT/DBGG5emHvmxr7ePziWxbDU
ULg5/SN71PM8LwSq3ZQ7NlHmtwmIuMzC4A5Bfnv+juI9MnZki7lmf3oCx2tLHG/M1C1aTeBHQyhp
c/dxO090JPscV0sfFHBRtavTuUr32+lxcEX+mmCEN4N1WJvSuPZNpquYzRoquuCJTQWypjNHvf1S
BC1ldgyyh3GclwR4YhS6zTpNHSTAa3d7E2Y9OM7mb3fELHxirQeL1vRiy7s0iRJ3fO9C7sGWzWAM
FfGhEPcqtHJsinnPGr9XMPjfRqwUjJ3uYyv1yTZOke7TJeUMQCnpBZFoumorLX/eRd3mJ2A6Ip8Z
qT6/WAjcnNFlItz4i2apq4l5q4frwTeUhPZS0wojZdo95xgtNRHSCNZG7V/jtehQoPEs4+uNdLeA
jbqJaFCd+RnnrRld/a7iX2ztagQpkxfmvlkAO9aHFEayGV5kIN1UYFktEfPqo5flRVZvNzAsPtDt
JS2X3nQcJA6NdtNcmQfed1LUYFj+tU77OkFKS47bECPvxuQ0XElW4n7+AaIZQ8cTCEL5snCluJSP
I8ph3apVl+fUY7dVn6bHceTGNeomjNiE8AUL+is0Q0ZpmZsrXVBzSwKfd214GlpscSjxOK8+xZwY
6MZZdaOqcckTKZTsM4F9X62599LmAwM3kdIeulCPoBsjm+Hi6ocQgxxwRXO7LfBwBODbGxqOzEh2
MIuqIfIm+W8fXf4lxVI1eb1QY9mXEo4N4oKOM9rhQOpsODkUAOnJIFZ5erIOR3El/I4EppiwEBMs
tx3mDy7MOURHrWRAldn1D/mMTqEmZoHgJ9ANnp3iU8Bn7WaaWQZIM7PRS+Q/QVYm32R2YU5XrtMI
+sf67PAFS3pAODNBavfdTuxTYTFYda0TcRERTjhNxVj3jGZlHaWEP0LQQ6DOrZAdaeDeY2nVVsaM
oq70KDSGXuSb+p+TMKAx4cZW6Jrcb9bmX6q0gwa+zJrw5R/AwP44cFAzoK+532PkKoMhjQxZSLSK
vk4zlMaWzRmy2+PRXmVJxOLw0Cjqy2UaTF9GNbNBvZCyXEkpVawnH+SaoERwJaxjv2d8jLT9+k/F
CuKTnCG2m3SS0bk146VEZLxIZVix2ijq1mZsXdvi1nrocSd/NRkq7FhoQvL30yxFE+qOhzAwe6DT
GuO8gn/HJ9nL83roJ4DNHrvdYxSyodbumDitaPd6OtjwzmFvEePz4TnhPyQ8VOdjPjO/pH3i9haL
XLo4+0oQtv1ZAHFJ841LqI/NzrlY3ypocxMaJB806GL27qymQWNGusAqrjGxWDkMy8BaS/UBV8j3
gyv5gFWolWD2LqSYs+waI4YbYoeNL5mTqkdVM5KDoQFQt3tNEC2ExCnhns4qIHE9q9kMCAm5i1SX
O4Qot9W4KTnLUBodwzrhDzm2mxHdImGp3XbXxJ6inPUGCkIGn1sh6/67YqqTfs/qljHM0QLrB8wA
9JZno+26CyhgSOMPWTNTEqobIGxzdgskL+G0OFmahchhf+gWyg44caTZ2Uc9P4XUDdxZmfNR0PhW
naXptNEWZr+8X1YBJtXtqHK8uNc0nDrv7fr8EVMFQPOwuZeGhwDBGizjpyrxaNrAZcyxuWE6Qmlh
Oj29ybu+HrCh9ilI/IbtEq8pnhYHw1xn5P+wmuuPC6Qs+dzDoal7XzjfwxCzd8+DfhZYkgr249te
CdGnYm0zx21h2jco6r27VweA06/Vj9JrmuPu0dwaG/rVqSNwUgKcYVRPDDGyeFQTU0Gtbr2arm6V
6qid8XD0AzXrBTxBJqtH3o1/rxDJpjUUYr+p2omuCCXpFXgGMtpRSoQ0yoduE1J+fJnJaaskdE2F
9mbRfnAp2gtWq3I3lIKOWqHjH40aoFrUXnrX8OlvN3NfsbFvnLhl/mZLHUPJ9Gs7/TzOljvT7LbO
36FV2hSELPtH1nHZVNUl09NUsy9ESqSyhfc2ce6qXNP7EyUkryp8qpEUZvKoIK3uOsl8SzCHAct2
J3SNjoLaF039kj+dh9XduP9LJd+hjynzluEtBY8W60Q72DEMrsF/Akll3rnLqSzjwnBX9kYN9BxS
nAiAp0sr1lGyLl8+mv3TGZoihUnZjzNvhKYEXUY5q6bV5/g+H0SNdTGG54Ij0df2BND+VPDtu0NC
wzhblKE0SXIIV8swfoIoIZ3VKyLnuIbapaK8cEHpJme1A4Y88YrqcGCieEBKN/2YRbtY3Lv77MZV
klNbFgMH9HfhBZct4fvJaDRUB1OWWghG7owx+8/m2bPmSlmEhcCJzCpQcXSGThSJAVSZbKQFayCq
fm+NQyNirg71ZbMVfLuuKbiRF5R5P802PlmcgWflu+ljFU74R7irElnwsOmX6O4vOEYmE3wVJhtt
A4yL74fDUwDNdIryZlG3YFqWa2/48Hrv6rtJBAUDp2AJN5xzPHUxeqXOyzkZ52cjLu9sEJW4uQ5z
64wC6+HISrJEgMBgLVcElhau6BG4wfnXOgG2QF3oJVPeNE33ANJnkp7dQudgAbIWO5Ia3tZYgkOY
4sZeEFFK/8l5P/XmaG7eV4xaDPFgdKbOFVQ66ZR7Y/EM6CHGFV2MDaw1ipIcM1Cqke95SjyJXD2S
STwp0qsQlYh43V5/7vxeLsk4mp+rQ6inPmyybUNnak67ERp8ElqPrDCGm6L+BODISBzNRz+f3L7c
B9FI/thGdQEbe3zG2qGvYSZKkwfSX5/srncRih+gndrD4LF6MBYQfo4hikxkctBenI9mSLUIZwhh
/Uu69DOUgrILUr+8PIiWFUIQDrgDHL/Gc3JvkHFqsBz4REwBh8wyOaMkrCdOYwVVSt3/d0ka3GX4
YohH5yEOPHxq5VqcwlSkLzY6Suo6sHGDNHoI0W0310QWOXYK5mZJ73cLcMDMiZ9dN9XNO8vHaW31
E/0GixltaXuyahi3agRrfX5lEiubeL69WetFax7xle1PBKP3n3Pi8QSG+HVWUFn5hpw5akgBycFr
4+7VtqbaaijCJf3of3C0HFItNwln1nkNU2d1x1I+PDMbWnDU9ozi2wT/ShE2eHoPNk0NwjqPHJkL
9XQX/6B5Rl1Qb3b4voTbAfCBbO+S5dVDyAH0JNJSn3ssxZqrVyzlzhZgmS+tt/BWa7Y70tc5SsRw
SuT1iEv9PRTvDrh+H9rADp+XZORyfygY6IeUk+rCVuFNmAOeYFuv2ANXdQ2twPYwLcjQlLf3mL0k
lpMURKW9LAFZ1sZHBf3CDCGoabed3S6oR3HshHHS8iqmBfSCMjawAm1OrW5tizeGhO6C5kf/TJ9F
jh1+dte1honPt8iGQMr305jPvEhEM75mgM+NoIXGrdJInrV87i5XL/s/M9rZZ8O6BsQOh6yWuAYq
LTkioqVoa4JLeLDXgeX74fd1bieIY66ONFsKdege1rImEbgQM3feTAMJnhmVj5IYEP1+x26Zy1A4
efokYafB0xZqKWpNiR528EAvRPCdB7pPTQXpWeeTmSZTluIxCvAqh6GXnAh+mN2iKvS5SAA48cZ8
zEVvQnFHQ72dMiEjYBg6+SygVWokD27vs3ABlleaE0V1nEXYRLwFJ+G100GRwzGGr01DcZ531QJz
0/MO/Y5nA7P76BlnVBlj8/IoF0nLwe6BOyeD51vQOYD3QuDhNl9oUWH7sXOpfy74yFm1QirGHDE6
A4Xkzffmpw+qjExgK10aNXt/lrLlXOfiRqxh/C3MwUfEL9s1S1+wH97F0Gt5wYViLqJxeAI6iIWv
DvYNeb89vb08x62EJaZ2LtFwAZbMF118hVJ3+YVgiZ4l4LbA3eHKRlxb85Nwtk9/v5d6Vw47lkTA
zxAnleDFev1wEDq8a31P72ZAl+DosIx3tYbvmRqBVe7doHPuWxaIGWOiYPQ/K1qJJYZYD5XN5u6N
kVz2nV3bPvYQE0rKjF7s3hP2PevLye7gzk9XGsLy9dBZmOxCNFRFWLr7zN+M19UhAKvBFgF57zB7
Oatj0AJaZC6R3IbWsFtI9oafGmBkHXljD6/2q8+8MGrmTXIChMGUDjuYEEA9gl75jaVu3qaB1YZh
DwQ1KdXcphQqxANn4TtIt6QIjCEnVAAurh8OmcVkJpLpVe+hGrBwIBELjvqLASPUnrcZ755kh129
7n7f9Sg1disu3WBTUWY2qvUl+MgYMTGNSrGjwQDQZqnH4ARRkGA0YkLHlqDNTmPEBiTCUgnmzzYK
xV3VMxwmxC0hX2ywlWekn4S/Q+IO+GjyvfiaRN0ZUDQttCddp8l5mTYYQYNFVE6D3EON7Y/oOD+m
7NkqdNG8AVvwX/ziH9G1mivWhMTlQT01CZC055lvrNa7AJu+dSyEFGolyTS9uxxiurtSrPMCauKn
yIPb+BuvHay4IyenN1NHdWhzRfp4gYxmCCl1LJinfmkFTSIHXzzsaGKKafKN+G0eFAhhrcDOtgQ2
eYYuTvoV1BxMrx0Zqcik7ofIHwkpSBKgV/XTmij3uAxf1bGBWmMPDVtE41LLaWjRkojwlN0FHQMS
ullt9FShZCNAThnF8zqLFYtQhWSlMo+qXa4J/qOiVeTmtIMDswcrSOIXEwC8Ps/Oj31dknxL7v49
Y3oByjPHaIxOhuj422eX6Na9aPMLSFqEj5xFhtRHrTgKgK/4AZ5LJsXnHq+q4nSV/MSeAdczVp07
C1mRLKbqYCFKiygn/zSnSb2Cve27Rq5bSh+/bsnrBiVu87k/iBsuerr3OYgvGd/93RCT/hv1gRa/
1gncwvlB2BBdflXDKIJPLTRt1IEjmgycNjC3Kg4lk6dIio9/ie3YE53F4LJS5WsT2gbKFBWDuxjh
IXM644k2jGyjWWSVTQfNQDnvEWFwOBBTk2fuVpoZusEFfwR2XTQjeuKBqVTKE8Y/zR9TY9Yu8yAN
kOw0Cls9JeCP4GnfD3dP7jgN62MBROh+DZ2NMcdSTQ8exhj7RlrNrCqaeSGAgeTwvj+A1i+jzHXB
anU/CtZZqv6nWVmkAJIK8dWlV/11jUH11pL5HCIFqx7Dtinjfy5tPAf5knepmuloMczbG9uFP8Bb
UEZjsZsVU8dUnqUWlg2w6ZeefV3Il+/Bda2b/AP1uKWaKPBqgrTHZoM/dWxhrzLz9S2RQCrbS5Rh
BbzyGbn/A7/KTxBWGoB0dGG8OmuMCarGHYrnxS/MmKaJfAzfnkC1NrWru/piMKJ8l/C7uW9MjCao
6VSgpiYn2gLWM46wiqnCay+9yDWBRdXLKXTnWaPuevILImqZ/8S2G0oC7BOQMaQSsL44Xl+s/y65
DcKjEbGsG2/UBnGOWT2vGllmUbAp+xvKPyNdgf3QbL0GKftdiYgfeKhQyq81gsWk6mjBTa60TIRw
9t3jDOSMsDqq8nw1PHhlfQ0W5GYmJmf01GFX9xFPpIFGBh5eV7BIe2Plcq6wuYTyY2Tks9Rg77Kx
V0tNe6iArAUdJ9NHS9qEpaqWV1F/gi0q5wK6cqatg0RMfa/Sajim/kgsJ2SrjP/wQxnGyNKF0qAi
0PJBX9QoxpUCVdBd+RF79oZc9rvsX+ORGldLW5xNInPSNIk3Wecl2icjyCB0erRUpoWfbLnlRtOp
pfV5uNv7Pr9n0l6AcxefONPUNjRW87ng+uot6cka8tjm/uFH6XP2kgMkgZJWwQ66UJRSESjSfB3P
C3Q4NOzrfMlLbO6TFsYjpbk5Meuz7cZUlnKxu9Qk030YaoXHRSNeKxnSVPq9svm5ecNjfA2d6TuW
+EwLO+U4nnmFt2hSygX6MLU3SUWiPnGxe5LS3FM+VmKRCYixFYWgnJB7sqAWzgLPASnvEwedUOwe
JGBZzmWeUAhZkEnUB/QorO5KwHImNleJr4f0lSp32X+LJ+98zwzi/fA6BJtv92HPD7Esyxeobwbk
WIW1msaGTPsBIH72irDq/B3eMa7V364YXIm2oNxHT85rDSyq3S4468AayBnQ7+9LZhn1q5F7ys+0
rWd9o34odqPrSuLu8VLKJmscN1brSUAVVpIOwAQCezdOHL8N9kGxW/C20tAr2eaYmkwdMjkBMksj
6c1/TldVbvk5Dv6ub+fsSIkJPGv2R2LSG29Q5MUS0iB8whhQIcmK3pkt60cZwAbKQDPhci69TRuS
Ib+l8Mpmlu0ey3bYDS+6q3QWR6huZDFeDKzZjWH4eBHUeXzsqpk4iZ1/SU+NmHqWpZZ0NUrPqlPU
O9qGyZX1229ufytK0uZ7TTflXseLVZ3qgdHXAu8G2Bx+Ln93YrLpa998D5ln/WFv07aZi6irqc9B
HHMjtOUgkFyLwKbyXxJcLtRQDmcC/mMJQA0lFoBz2Db72xO1iC2xV/f8tJaiZyOMwjriWU0JtZSv
KObR5oWYlWSLdWs+2fhhEIBvwPOPbjUUca1WR3SniEsLtuG4hIqHeda5M3OWvxSjF4oULPrkT50H
GNE/NJxEAKhXh9TrmhidTQ7tue62Dk2NWGT/AzfeumFFsp7DeYQuQfxGLQ6zYCry6SJ8TarkxVNC
B1o/rDDUOZdxhEq1+/TCWYwLM9HrGXOzxcqHijS0ZZw07bYBUyjIKvwvPTyZuHxkDL7BUNSqnxl5
oj5eLpUERWvmUkcbLYVV7iB8bHEcb3RqWgtk08wzZk7JxSQnEJtZPgR1V3jYJpfVY0Y8xu7D2XWI
bcukpWoHdsV8+RA4X2J6bV4e7A9cmYCvsLJ1xhntoQ+11MO+VPgVi8MKRJqmneCkigV3zMJH6jqc
dQm+w/oC3ffrXKE3MwBZ4Ovtnf32qB261Ij2NAHK1Dxf/P4bVgK3Vr49mNeT9MldsOC4E0MAeUB1
5mhvbM3+/0ZJFhz3f1KuRrTADGxW+oajSyiiHVlx9ElHVnh+YnBv0FrGl+rvJLW0Jcu9aGSrjsFl
0NFT1S9uTtnjXc4ayxX0gnRxr+GIEbQ752mWnLTpegzyMAdgMVq9AMMqN9PKid+WY24a5+8tAEEV
k93z/fex8Yui6rcP7QSkFj4Y0FOh8w87f9r0MQvYxUmkZ1owiE0rJ3YEPXF3CJnCvrJ5tE/nwepO
sTk9GPLwG0Jb1CO7OCR310dBEcvxz/dlEiZuZM56bFdbJdbj9hznjL7km/zSYCRlLQZOi3w3E8rv
n+kTLYSRTd7c9C1yq8umsZqT85hrNENAiohi5PDviUbIAlJxjh4yCFR5cbiIYeujM/85ZOD5agH7
GHP4/tPIbs4AWiaw5ZTNH5cdybZgyiv4qpyL/SFl0j8h48yy9AKedf6Wn1xrjUtQWTQgaWYezLn3
n8DB1xXWCXO3tltRLMCzvAMznI5GD0fNUK8U4229Z1p3HTmVZ+bcoKPiik1hu/rldpdmt0AmqOc3
Zgq6tvGp+0Hfw1BxEIWGlzEPhHhZTjJRw5jxCv7k9SEnR6rxqopYTfQgyeIEExsRkZs6d8wJvunH
UmajqvhE8XkNI76jQJSdCj3bJ72P9f+nbDRFGq4wNFNbWgA+z3Iez08DACy9H3RpqY1qVVZBhSCr
bYP6yed+9ZA6YoPLiii2x6ktFsEUPRg0yLf1E7in2GByZRVhxVaplsf8RvacLCFOnnsXuRRR7M4s
XWWHlKSa5fLsY130AgH7Stg2TqTQpGUKEaxJiUTrXlidiOFI5KkwvwZRI4k4LDjgQ9nj5huIT4xG
xLU6qkoJ7IZZWM1/+qb1C54aJAsY9pvFi7ZiO1Mq4ysneHmjQ2BUoXSXbdcjDnV0e9wgkEwB4HCI
PHoQWDVp5RFsE8N/jGh9YXHu05SLZG1SKtHZTKkkuhibV0XCkHtBuHLB6QWq/H2w1G7Fv6Pv7LHK
YppC7FU9YrQXtBaNjmM6WyHqt9pOZqXUAgRgJYjwOZMIOG2HGxXvD65RE71ghBGVKQJ8LRhDp9np
VLPnWLViqrOcgZWa5ouELtw3g/lnFW0bR2NSny/cRu+5ln7hiW+jc0X7KtXOynzku20Xh83XSeSk
c7QAB7h8LF1Aa+2v9BqDmeTrNJY+fSlz7sy28pNRwKAMEzga9VVVQU4KRG0fbCnqLdvZ5ngKhU5N
IebgM4g4RIVeRkI7hK7BqoxSNKywtwik6MOYLMKio98/TA+cp3EvqXPuppXrX/7BxoNw1dboDWbK
sq4Jo9q/Eo1kemZN6elRvGffDVyTlS+MQDEnL4mKD7TmjW2ORFtYR3UPfhb4u25kijWTQbyYgpnM
rgDtecDYq2rncKtfMU/lnomDGWlmHarffenGDmIvRV/NXxxp4Xaj7QQx8T93m0seKge6xi4nt29N
c+v55qPnG/CvfqZjPfGedrKUiRtOM7K4EvriYwTdwdXLClcfUFUo+g9haKalOjdXmcH5CnWVZZrs
yEloWMYb5yzgmKg9lgl1ofsjFLDFJFGw1fRLTlIRirYVi6I0qEBPf8POP9YZf1XAB/5g/r1AgxWz
nKp2GoSYGFJOpWkSb7p9aoHlzoqGAnGxJFLvOU+/Kz8z33Btjddk0/bC4g5hnWSEOfzJ/ShAnMJf
pY872icp6VJyzKueT0dULDe3TK30+Y2ONzkw6BcGGOSiHxzPuHA2XcsThIV79EMTyt0LFOw2VKPs
2UPUiESLg6duOnQ5KMZyMvcBhpCjCqbXGD4toANc7WqK8jFt8yGKrrESRe0gPMrB/fug1pAGRg5Y
CX+nn5bHk44eyC5M47Q/E+sJT17yKSa28phodGv2n+isWxcDDkw606zfsjhNj54Odj6MhTVJ3HLS
xOWGdeei4IG/GDGgyVYEpKGYe+1IhSHjbhymIS5l774cL59Tz2vzFPKSybg57+V1hpLpUFE/mjlF
jA9QMi9HPoV9y1dOpPCqEkcBD4hsDnBJwNr8ZmQSJ9P5rfoBb43gJpLBGR4o14UHB58t5rNWXID3
UsqvzaSfxIP2jg21cF6/NoH0eUyHj8xhV3L/4gnZnwGyqa71wNRxCXsrNZBw6bn79q62V3/kbGZl
F6E8OILUHaAlmxoSP57V3kpztUN/79nTMKmytXPlJB8DeuH2tAQs88R9AAT6rj0db1MUMuWO0Rkw
vnYWskyvZhB2k4vC7eb5Qjc7gBG6VKfL8+lTnLFYrPywuATb1QFmI7p7h8T4505mRX4ZcYKvg0ua
WhBCJ1/6F0Y/SV2/qnwwVbn9EJLePWyOUhSc/49Mb/yC5TmCAFTohAKtPpl6rbW2VSRg+9rwfhw+
8zejXK2F3bdEqUSgorsEysO0j9GEODtyYI5UeDx13C39byRjQebws56Q7DmbtWUFRo+QDulQQUMi
oqloBqiZUlRiYy7jbq45RmWOBo9rBBT8Ej6Pv0XbzgE8cxqGorJLekAGDhjCnVKgD6y9w2a1y5R1
yuzrG1Xy/EVu6pE7Fw5RpfOwC2Ocu9qMW8LSDIDI00tjdkzCxOVOr1svur/ybLl3v3LlwiG+cW79
aPeOOq6agypzerDEYfPJ5uUvWUoVILr+ndo4VQJBPDSHopJ+wpCw0qVNzmdi6FgGLJKoRK4fplZX
uagjHjgp0zPQLn7ht1eFV6ijn/C4OsHxgwOf5RDSZvvqPWr/OnjbuHgsUqJQe0LWbHWJzBVAGKcA
RHnyrEVaHIkX7HqV38uYD6dS0Vq3FmvI9r5AtkW2jr5a737d83+OWvtNK6pluQGoekzGi7GXDxpv
VETw86JAOG6L7GZ64l18OV26ulFaDgj/HTTsy0OFKUM2UA2FJko4+j0ll9WoKL2RWWTur7BwEILv
8bqJ5oMUbJ86mBZj2dKIFOR6thmj43ugaNzs9IAzlo07piruprFEMthAA+pVoByvI6oLX3w4itnw
LwZfOm4RcdSR3i3AIgPZo5NfGQDqHas05+ehQYGcA/RnbX8OhVAYJDvnmEvk1bw0LtSLUu8wNTKk
fFU6+6aZ3nMGYptDcC90uUQjsmytjFhbshgQKm7PlvGqNg30b+iuZqyTUTLTS/Zok5OrUj1weg1H
UpdNFZmzVNPKlwi0KiGchvprZeiKPXUw23/rVXTufdidxzWQ4u1E6O1OlL0utGKiXsYyvpaffQSw
CvbSZ4CS0yyOm9krTebbg2obwAQtzwOLHWR/kCQpUO/MkSkv9OyEPq+uXg3JWJ4KGd3TXRP9531A
uF3P4QvNB2JHtVuOsg2vMlGIg4H1DYNYI4JxcsQ8q2e37LfjD1OwPW3QloHvAEfTdmXRspHTU5ot
EP2q77sjy68hOq8VxM9GatxxURICM3QWDtypvIepMdghjzwJu3C/+tHt4Mvc6RCypJ0hBJsuV4LZ
6nH3yLLm+jdOeOvOqB6i39BAu8lGypOPzcyJhVFWTML9oup9etNNZGG7s6aGWkmf00cc42Aa7yqN
ffpCnOPd80pV0PHsUw0EbL5QsLYCdtCw4zT+L01g6nsEm0qwiR4cDhVdyCg/8CmsRDv1MGwo5D9U
Z2eoVzh1+anaEPoX5JjrpjWjaE0ep1jPSQgSoo56IjpsVMUXMzXUyXmB/04lF5VvN/HNCbDvhDuD
Cv8WUs2P3rvApL50FTuu9IAkJHiKwc1K6Cp9FfgU0xC0Mf7v7JSAid9Ltqvzv1hPT6vh3uCDG0rI
wJLmNHPpbBaFaXjG7ylZzJPLu/XOh+4utJRN6tMroOAkeF/Iim3bjB1/6h7eA96OwwYgGWi1WlMq
gD0OWaKi0sXDe/ABfe70VAvU354iZahO/ZBThg5A8nLOu3ZMZWfJtPpI1xAvB+wzGI5yuHQxTzfU
KaApcAGOt43zLCUbkRmW5IjlswdJh5qx88/MZwfROk5AYVb/nyVsby3rA7iiouai1QnE9JSyo9gW
tif7JqgcSiXdYQCuFnpronU813JPtOdW+QSnz7Das5ZLowGmg3cKQaR9PTCNfQ+L+whni8p6zTt8
zVf1GyuC0ZIVTEqoeyuRh0lIXVWXW2OvDxae+SpwxFvJn2vbqRJqRSBhXVT+SxBSxl9D3WsGCOlY
S0UZQlfTvT2jbFy0j2YddVwJaptiAApqJC9FPRuqa1I6kF9ySfrMy6s4briON+j3ydezbhhYVyHT
QlzwnPgmvMRDQArdzej44+46viVB+TPtrZBVUTdqIbZbbVfOsGYUh2mvCr4mzYbs6kPnE1+v5AeY
gMXKfwz3oRPEmsn5FbDi1IVgP64HJZgrkDXoARcGe5YAM9EtwpQ6ny0P165Y8UiuXhZg707SUD3G
sU17LpaxKBdaegBBY5w4V9ztzOs5Lf4RnX4yBD2pOhVDTcmxfL+EZziEeZZmRfnB3ZmwgZrPUtcF
f4wDjJaiUPLewt2VM450h9jlFjagqxc35FHN/1YJpCqWembkcjxloBtKmKP+XEC4dcdbPi/v2o1K
RIScfEce51Ne8Hl+QN0vmkhuMPMhRJ339mrkGswLSUmLlmXrakL253gnu9qZppje9+2LyuAQThmk
qWZZtcW9UW7D8uNnf+pgzm8RsRhLShgtcyDaSKwo65zek+wlvB3J9pWvWkxa2zvsW1sFqVLvpZMG
qz+GlDqexhWWfkq/5YnWvXjOX/zTvtXmnWg1yLqo2FQKeuL+lzt6okjdWhHAM//qVyFlVDYJQAc8
8rO/w6IpHeXga8EyidBlofLIEQ8yc1dh5VHhH+pYWeJXxnlHq9OMgmICWeuSqgmmRl822kYnw+mQ
VIsNMOXsNb7PZ1AGyFhoo0T8negpCfJqxNwapSk+ZLmo3pvg3fDmziD/57h7Yy7wsjxampnnxsqH
J7aNBJjiQHO/pjn1e1Nm3xjXTGsQjZw85jF03jVYrP4ARjCTzMoZYqMdeCIbdfM6x0OmGePnWDSw
rIQY459mNgyWGTPep+NRN5bu+9R5hLkekD7vbU4eWTgoCQ8ufXj11NM6a+0QDJvczje2fxAGNYS1
q3ffpuYcbBI33XHbZctaNOU7QHr1bsSm+Y1jvaeB3Hv77lfDPWI0MnrH98gc/hdsNqBE3gh5QJR2
lcwfDPibrhI4OTYv7JJwIFG23LJjXP/hIPbuNY7GF2+Xi4nRLmBYTx62xSgwagNWf0Xg8duoVT3j
BoZpTCXd8CPSCUxtiIVIdzjXYpTkbzVSSBPVdFi75MGCQEIJlpoAYtMRo2MgVfAEpfAo+10XC6bd
mLtJl9Zrr1EQlHWjIRhkIt4swcq1xwQHyYxKmnZnfTMk5qI9p74cp0h5FUJBo+QBZ5ofyzsVkz0s
GeUT5GLoZ+CsGAMrY/uNGNKi99C8HHgFsLSIP02bxxWi6igrkHOfbfMjh8ugjD8CgtkB0w7ecXnM
2u8MwEgrWDFxnelpMfAPgMAezyJt8WKS7bJCXF4AEaXUgNMpwVx+5ghvClbDqxDPL9tiDAjaSO1T
kMEwHvncWEGc+mdtIhwr6utv53L19gdEI36KDMvv6zHsN5dygEpkWetP7thRU263pTmXSysX3gQ+
6FswIhnMvN6zWQuoefbg2JliifzIuahT0wbsiL4lbtPSGbJXq1Mazzq3/2EKijAN7DYCCcSAF8iD
MEGE8Rc0VeOxQIc2vTGsouQ5IcuBVfaIm8TVF4CfjU/hmXNMtieWMyfp2N/9nDNnmiyF2pXCQOzx
rnz6IUn7dvnKFBCB4Fp6H4l9AmlLxcRaTsswDWKvzRaf/Bh+JrbrhtGkV4ofHeXxL810VxUecZMF
5MK5A0PWqDC7G/ZsOmxYIRYdAqTlrw2oQwUoCMPhivJy4mr1o1O2XUeCPohjqZwZG5FDSjYYf+th
rf3OyV8I7aix2Pf9HAvrCJN3O22J0T9E5ed4U8e9zKH0McS2kzBG7Q8jNqitpcPABKNLwIi82hoJ
hDuQFxtLqvWqOq6ra0gDi0jf9dyHHss/A5CwUsQkoY0iRw22+zLIYE0PkAuuP6Ks8Aholx6Ymg/Z
8dLo64rtn25xau1p+1PFUWCVobifU6Y59owmR3rLosxzSYGKvqlJOa4vh7fCWDqiNf/EW4llTAWt
zxO37u/vFtLfFjw/NLsmO9s+jOvcLSHfYoJX1M/Kkhc9O8L6JIoDmVC9iAMMpwBZclArIRGNKpjK
k+eCiFggRavUC4a36kVDJqHj7APwzUUNyzDPM6kUq5zgQ7UG8WcRvq7EtiJxzpBui6sXOmlYeLXn
WDPjkD6HNdq4pc8DIuhIlISt3UmXeu+xxfUR0pIVE59b1VrCG9JBR9E4o5Itzr66ME0Zda2B7tlt
D+NCJ2w1G9Z9qYaHzf5RRRP0wTqRi08wvE0iPm4RkULmxtaMwdcSrY+PcH1nczjA80Z9OfNKiVrp
NOBuaH/XTCHGBKvnGXWmFwMqE5nfApicIi8TjPX1Ago5boRw9P5sy9IpmG2D0VrczlujSAZU7dMp
BbuL/ekKTyrgeO9rFcVow10nKcpPD1DLFsBlc6UzY/vsHTW6tLvQKuXT13SHiMQ2ZPk9z9KjYUJv
fhYa7g72/62sormBFMsytViPLw5kypn3GrRQaVBHWbqNi0ejJlX404EIBLG6Dp1Lnp9TV83WLTaR
GPnxahA4+sI5kr/vm2/S0U/Hax+6S5wjpFlYECyNCJLVHDB5cMVqhkJabRi0Zry/0xqjuOY60aGQ
vw7aRrDoC1d0oMeqCLfESdK1Wg7RnvnRY4zH8fH6Uoiky90QXf76I4DZPKzlfhgAXVF6DhpszYC6
sJabhAI5DP6cFH6+PCNgDxiwBduwvDENs6cMOVFtvaOCpvXVZw4BiV4AOE7kaTQzmQ4KweDQAE6u
PxvM5/fcGk3FH9L8X8QpliLJnsYsL94hyyc+yhyneJFznYZj3swDdw3QQaAd6nSxr+zFksQgMswS
qpizeA6kbmjZKZlqfga8x9eUbBkHePKztfVqty/VQrVNRaIabF9U+vSZz/XJo4rU/wa0we10Fch3
O0bCvLDrrPaTnj8/icqb5GO2pTzeTGf/BkQfN5nXpB/Y7QUP0K3FXxGcOHVWnOsysOlCqmw2qzeg
ML4klgGaXnCkXaX/UfkWy90KV6pgYQBsJ6LEHX4dAs/WmF/Ws4StRMXk8kEpjZrn02HDIi6TOQWe
ZjAsxHUcTJmZsRpPDEJsH1igC+hnfIsJmI+E77iNDOk3lhx39rkukx/gimHKBsx1U32jewOGLcq7
jETy0MMIf16exd3YXtQAmq+2rQkQ4o5VqdF6rkxJ78BvY8EtkCLL/JvmouUywZ+7LQnHCak+8Nyi
xZ1JG4Vi2e8FWTPbyP3WDRdOPNLqtoG707oqUcI8NBQVzUOX3xTj51UJcw2u6bIVCKRy9PU0k8ub
fN7B7M/UJ9P9FAKt887GH1dtGrxdjmyr10XEceOj/jkT4ZaP94PiHSts5ZLFqX7kT87nUGr+f9pT
G5MrCZu1er+Ww+LNy/62QOZzP5cvv42rbhfOuJXg+PEfPdhKcQ3EPDozEzHZ9axWyCfILhUncqlq
0BJ3qrIiKqqmzrkuGy+PX9DSVh6h67QV8tLQR/ZfHnYXIAtjwd6iM2pqPJVqBvHL8HpPDQp2MUOA
f+mtCFI6nX8s6zYGNTycpSivyo+o0cz1Cq1kflt8iMS9JzlNsTnW8KLkyd3p2YHBsKCK4hH2WPai
YCU38QSeMEcGyT4fU0jFg6yOvev9iJLHs1GTlMr+dFNe1jrA4rSxFjYmnYitxmGcWvV3nX+2l04S
TG2kWng4pMxtdCm3np+pI2FerHC45i8voLK7yq4eA/AYQ7PXBy+0Mhvcfpkx/NxQf6nVLFfGWzME
SLNDvqXWlk+JVJ6t1lE72/HeBFwSg/SYS4Q1cpWhWP5WK8z4gJZkk8Omu30yQtOyU1rnsbf5oKF6
mmsZ2aHLPnJPqCyICwJy6ex/fOdCEZqhpxRGZY1o8XA+aPyXrk6P57+bG8940f3C+wiPXIh/Lowl
RZ39wIFM8SvBfqlnligoznpXYlXoR2v/ASPzXvHDURnDgVuGX4MTFMQ24NTRSZoxOIeKnLTsaXr2
Mf2Hs2Qyq+DQP+nAMHgOS3o1DtDK7zrdlEAx9wDXoZ8hmEGYcybG5Nshp1H3ozqDkx029/3NKZ05
YExSKVnvjzQvODm3Vf9E4nIYRiGRj8tLOcO3hQ9vgG4aZuoqT8dQHkIO88j/I4A3xdqqRec3RdoT
bY90RJsX+gQ2+LcBpIpkJNV+rUwWAPJAl5bGRctWqylkrKVdnONvwV79Id+vy+ow8YCxDQtp/DBw
BtxrQDFm9xEybLJGco+BFr6aqptqg0O08EvexBjtUF/JliGqhP0KdbklLWnlK8XSOEjQkq0j549l
ZuLmqml4l4ga4/zlVIjM8qjtIECYPZs80iw6wWFljDk6A/7JKUOx+z0JwBQniwbHHoYHxRuKg1Wp
cQJpxGV5kkjuRxbu5fGsmf+c3e1nOPhadE4D4vyaR1RmtFUlfsDjalpnfrI2d4F7T0WgkpzpJdxC
OY81NkwB14pFVpqfdMtE7ylmJN5OtRy3RTfaFlkUth1DASbY4xEnsCSrHqENW/ROu/LRAoAt7bzT
9GA2/mVs6kuZX1fNW2mClNYhjXQ/TmHauD6QBG4Ud5c0sa2J9VPoODzpDKbFvCH7u+ceTZd9dBks
pFQ2HX4dCI2cjqqKOSfDx5GLlqWXtgd7KgGk8MmcRxinTH7q34LfiA89NH1CoZUyiGGooZ4+HRib
0jpetnZIT5oqEDf/QaF5RYUBuH90oRuDE5EYmOaCTeXGj9jADlip2qMeyMPCwbDMo0WF+lR04wjM
LifbwZLmCJviR8qfCs2XxKvI4gPK3/tU8VFyWJDwDURhMT2d8Ce1nCQ94BmlGc6ooWLH32I2fYnK
45dUYjYDgj+0kKjNl0IMiVDLOTa5NadD/Rv5+D4VPwwxL21GvVKhUTvd4vua/Brv7uyxKxS8BoGa
1xG7jf05a7LkYZJXaZhOpN3Pq9KuiCCeYpb2RnGd16jUQydNl0apoqOmceit6+kFY1EdVHUWR1LD
7oiBx3y6AlS823wU9Kzi3dEr/iixIkgIZuhZlgZELGj8MQAaBq7MMr/kdF7qAnEl7Tbv2aNJsYM8
uc4o1a2ww3WhaMYXp6S1qWUX02rSJnif8dNWXKh00vuQ8W322HSCR9RCb/8XFQjr2Y3VolUms7Un
rOurnP5zxQwZiiIwKBmMUclKB3ni4Jh3M+VUo8EsybhLqbUqKhltpuHb/mNsMGa066FDC5b2DUwQ
+Dv+qw5Z3Hu5OlgdxC7SKDDt84XrfPs9elDdu8vZwZWt/ZUGAnoYBizz6mZxfpsGlmVHUQEoYIeB
XA+3KZSLhey7LKWi6qYM8j5A4mG9rX4QKdlT+ojoWno3G8uxuOSFT/0uggcUUfptPqK5+75ciIp3
OFuD4KYbzt/9sEOSvzmXucI7D7ltszZAzaaJVwzW1TcDwOxtYw4EpfN+XOpQE+Is4g4AgOmk7KCM
/HcDXQE/x2jSgX1Rdb2XMuZ7oQokXotba5irfY7bmLWVWq6GKbzJJTT8kBkkq8tSidDiN2F4H/VL
BBfgsuxarJuVBeYNFq7CLYq8uHr5JM3+Ls57CBhYgybAv6XmyAt24DivtkSZfvmme44V+F63nhIH
H/3bsMX/2KaP1ypUzFiBJX/W5x0pC4W8KtXAWOyCdcfyrLCNr23W2XyAheB4rchPHUOBU9g8maHk
smbNRjr54Jy8JXcF3DSNW0wlPr3Gqht7ktoyjRL7g+IrDG8HT3PbEcG7IsghMRbKUGyt4Xjmw8Bf
GTtZg0R80+7C8vUgS3sWp2CmcIqSrhqeD5wg/RxWKglo2Cz6xbgNeT3/uf/hkbM4zED7LnygHd7D
h5ilIpkNl2hUQ2dXIT0PQmaceren+DaiG5GD1/FaDFr6/bFXD8cv2B7CXjS78sUSOjr7DI0/rgoo
f7UJcS0sivqUa5Pkg8C0ejzBDf/x/XLM5yD1chQcJr8EiJ3JVlVWb3dBPoyv4552E5SEFPW/grwU
+mSXAgFf43E02nf8CYXrcMA0p03StB6T/LTfaXNYuCe03ymC9+kCeiN3q+BlmfMAxAwtF0XsvfpG
W4wCDVRWc5mI442/KBMOwoBuxK4NZfIOVjHDGt0FmympixyJhC2FMDYxX8TIiQLWxr3E1U369K2e
zE0UjTnt6Gtbuj7j1XPvM2JrIj3GEPfS3HjceirJ1006IrKYFkPCC61eebssOx18Eg8Xh898nG9j
B9iAD4camXxtFFIs1o2KVNypwGgbIDg7S4Iyq4HOrymm3cJ/Gg7IqL4qMfyw6CDAFBbpomzqxCh4
bTmwVf8T/NiVKWGi/N047IhsD7YxfmluhH52CFNbr229ZMisRSP1xg765fNfForDC7Cz5xc07CC9
hZDoyEubX4kq25GKrvqJRXHmGirjKS3jMird9ar/5b34oEVn3PoVQXTyTyQEYn93/aT3TJOO2KIj
3wqiV0FcuA/rDbBeUcvoz9mlVjdeukgEzgRnnkossSdBnR7WfLlMplWaLkljWinNfQooQbTW1W8x
iwJOGRp+bJPO8lZ0iH/iH006/Q5WgbgGtw6KjEhJzUSsyvU9r63jdYzzABCz6e6syUJc+Vr0+wEZ
z+KtZdGNQWy/UXvXaSQc/kfGqFKt0YlJSastKKW9bgDJBThR/xl4nMk5NuWraAxRuRfhvrlaMqdX
a5yGZoDUMj2SJDk7LSmC0nhgRcCogfkGNE+kQ0Dgt+6Bcj0G9hCeiP6hXt1ArbzLsrNIquKmK6dx
/udHSkxhCBHlSo2AJrpEZpo8I3QX7ptUptcVZv30UzsTtoJv5uEUqM4OPrnl3dy4N2jJJoqJW/sL
+DFXW9V0n+j1j+NJpo0w3zJXDzCp1GmIcPmmBUFa7i5u/qw5elFFkXY0J9cPP2cGJuu56U+/OEqR
mNW8db+FGTap2mQZbWx3cJHcPHJr9PdUCtFsLVPLZD+5xP3CiPildh9XsLHPuNAk+fl3kkfbMZPO
WnONErM5dnW/7CSCKJs0kVjZ2fO1E7LQq68sXwGCCExcQ7s7R2NeYEq2L++FL3hRSbKWY+dRA+Od
y1RBf4UqfWwxxlmngrVp9dI6QJxJz6ULXpdoBhliysN4iGGuww6BZV9izFvNEw0d/+RE/uRQhcl7
DqiKpXJ9nM9WdPewT9ZnDeWb5t0pc99ezKphdYw2m4PqiTfxmgNq6+OX8ZAzRr91CZbBPbglaJSL
P9Aj8nUEveeLD4EHsiF8iiV/z6O3PwEtyAE8ggPHEShv5aJVNP3VsewIi7EE+SR27YoqexogdwoH
RziBG8hMPurMPDsBZMf7SjoRMku/pkL36qOKsM/at5myWNRUEPsmPLiBj3ZnBvVfFb77ZncoNxaR
D5DDJ6L1kjwtZjEEwlTyLH0WiaaRfdKoh2Y+cwqjyIIavZNmq9m+qMym7YSY1LY9lqkTz2zKzqs/
XUZbmcqECVYzpnG9fu1Y6Hyn+Yimzc2lwC3zkRE9O7RzRdYlrzB1uW7CHZL/FzGuiru7H/lAo4TC
39fKhopPe6dMKWPrjdnbYO5x853v+MIycUAsF7tmNQNh1sq7agSA+4xPNztnQRcvzN6Vyf3Xdpea
M2/6UTRQ9ObowHubeKvM7ZsnV5g0pGZBZ19vGL0PO2DGbTcdhxlYf4iNarHZinlu7QnYZDWcLTYh
I2Bc0XWEyiYqhTkaHCRO8U/XP1CQkR6FWleKyZ/ixBerJa+mtZuRAmEN2kTNr59pMrWlZQxUhlAa
rambgynAoJFTA/WQABZlSqFw40BNL+awLrzVY2YFjDjU/Q1dDZ4FIbODv0o3CYlayKnqGJII2YJj
RfqOm/7b0N7oEky4gpmv76poCaemhVIRT3CsjyIEUqTsLrSOTyQ77RGOMH/FdlNEgUOXP2F7LuV7
mjeDPpQLQViFCwGWO18szIq07HASCtvYzYx3AzhJ55ttMVVn2c3EnCVnlGrM/neKgl7PihEpj6uC
hnwbbOmvZ4w1hI1heJ29iBNMWWXmBT/odYjuDye6eWEpASDycjMhUFaNfaUKp5z9Dt5mI3zQVLn3
pl2sUyAogNuYmit7Uk2sM7XJ35gpbPgu0OXqWQmhDKeTLBJ/t2K4/gI7JYNtF2Jx3yu7zGO2xkLv
ZdKeah1BtvGIQKUgd+DNnAoZ8JcPJaxKVX1kaWMD9Coz1KMl8MRBdAzo/y31WZG6Nv+ZYPbXGzMj
kTgCcKS2ySmb0KRPvnRuQEmJUSxi1rA4UmmnWN2gtRg0UwkuuliXSyeDd/ZTt0gTIzEsLPCJAgzO
kIB9D0NmrHeA7REHGJdfryc7CV3PZFvPz5Ui25XIpEP6pPE0svBPgZIXtbakkcDkQf2Q61WvxNui
IJMke6uQGZmcvu8uZaiGbN0vmoZitCPE2Xc4kBzHL7eho+M2MTz0R7IXxgX5OjcUx2x5tKjZGqKX
tIJEZTjY+vQtkrA+pfu/3tEBdrwo/+ekyDJwF05kk9fgHnOWXzwX3goei9SurUtYD43d6q7MvyoO
OgFKCI6EAxh8JGIlTIU5OVwKaEZgyeBEa0LfLt49wKuUJqpIDjW1MOHCoJ4mFa093WR/fPGyBha3
vS3sAvAUpwUUouI6zVxwsdOuP7SWJmJ/pgKgvn6F1ZXjb/rbN8fHU6ZFLCQEz7l1MkeAvebPVa2V
uR/9FTIHHTDDvouqDvFosxrNA+v9C0lmxf77TzgUC3OZ+VaZaQv69ktJS19G5OsERCOfZWbKTNWb
Yv5dIwmKpTXvt+EdnJaXx3hHNJFpdZEgwDyLq9I2GRZdRHBhBnUBbEnRtJViuYMcYHPJzMjbnX9i
pbMkqx29TE4dI6/in9lCEb1zJFdyWB1Vx5UNdB3p4I4yYsJaONDTs3AcVKLEOE60bbwvJTUtjOL4
oPXcaAAVGAr/P7UPiHpK6V4A445xkA+Mt8qTskIvXa3lbMW+e0FdS8kNNmnvIFhHS1cbKkY64vyg
2IxfHEzQWFBfz1v/iewE2eIlnIO0sFFLXjpbAeasG2AeKa5O36XTFLdKpvSBIpy2Qkg1Sf/aF777
IRw8X5tNMjiwaHHCBpcNFzjm7lKrZkD9JaV8/2B9ERR9dwtGn/1nxg91nzNGiAP0i7INje+/oys7
y144OwmA/hZsBhuikpKgJogmzSkWl9y32zsIBXNGFRTAZn2vwmlitkeukS9+6y0JMWY4rVSXFnJX
8olgSNf/0Z9KHKtxG0bCmd5iqn+J2KolgqZdDArcucCtKdIgWeHSgSWISBXp615BVrfNMLpGkTfj
Arjb8pNLdX5gq3ETQaC3cv6o8X4etbwIBM3+Q76vLCJDJnB8iJAy7o6xzDoxUvXj7bKES82Cs8sA
V/kxaLV3eGx0pIwhtWMuA3yUoFIldvaSux+Osy9T3OwopNeQ1LnWjPcjRi27qBU4LT2ZZsx/RjZ7
WspiEx2N4TZ/Uno6qfI5LYH/mRsiJdEQOTH8AE45WpGy2OvPGOiVBwouvQnAmVT0E/vt2aevisir
QAFADJtl91FVOdXR+HYMuOf++3w9LSBWogVuOEcDzIjZkAPjThLaEyHcuANtHKQmL9AHyyDLlpSd
6TmoCZzRq4uhfagY/oKEQyox01h3JxmNvO7WHzgrskIpFmKxh+AV1p7B8+PIgl8tW9t8FRKECymF
JUkEIGoumOOImiQ4hY/aWNU0g5sRz9wYLSfpgeOZ9GCtQ9Hoo4eax+i7zIIfiflSb/xeOxoihllK
omEaobTwXO51EJ4/Sdd/shR8WkjtKXCq3aHXxs+lFsUmVvDACrwi/O17yyUcPSOzUizb02g2jH0C
JUfyvqqzkEp3KYpRxC+bkBLp9N0tJMxnYTfyv5dR16WYCQmBFbTJwTrnrQ88iuVk5Mt3VVxOby0F
7E4UBBuyFBFHI+w61HVD0g12YyvxfHgEnQoGHRSAviJV/BWWck8L+xwjrvxMJnQNCxUmnyJVhHVb
BF+P84fKNB05/uOQIJDHg3WyvOKZIgKZmCcTbXRHcDqWwCQ1ifxFqw1STbGw1gfirBnoz93yF74K
eL82eqrd6h4Sqgc7dALenVuejDARAmsEPBRQDxWVpuApiFfBe9PpIlpi15lzqheO1K/oKpsXcL3Y
xHzDtH8WZjfn2357IwJj7y4GSsvO30cv2LYmvTEz1M+O2pXGasd+4mbwNhDN+DiadrZtm24gojn1
MqFx19aG5AKVzmK0fTOuIpHqt4gKOvV9OFk/PZqKdKh4r3hVer7QZMyCI2EfTcbib4UmeIm80EZ3
uKq0jWOxlNjGfBIqPhO1SWPJJVy2u/KZu1sz682rjuRe2j9HBBWgdqbPeJdrh1kXxqtSJkqrJ0DH
6STIzlDRUztD4n3H2nESJH+RG68zQ1ICmXHHTwU8hhy2/xD7v0uCsg7kGa1M934iTDuDjiKo01yI
sYHoqoWKH05K7eOQm1UZ6VHUItKr/tnBjMkDWMfOOnvK1YFCTPPNk2kdkzG8/e8bNg/y5HuceAXZ
ISnbL+I0IAwa3n1VFKVByk5SNNrKe+XSgDheEcOiEK2frWbegJ3epux3WEEhPhA7QEEZwqMXBbwH
DoEePU4ulTfsMBgXjJJPfIBCXmHykx6OB4FelBZm6LeR5IGzJxGuaKKGsarwewLRYrUUJIsRkGQM
6SurhwUxSTTbReoWFxL0oWzPMvWHPNsUrPeL3TBKV1BA5JuMrnks3WUkMiQjik0Qin6AYIXQD+UC
qHHGtwDWgxYiRbF4yt78jmFgzzoNgjIMxxyy7DroDt0l4z3jasOO/Ir1XO0EZFxtR1goc1Oi9Ode
FTFUEH/3kYQlz2fP8PDMRmp/HJhvQp2PPpamd1xWUhts/Y4HWJeWRJAy5jGTGpp94bb4fz2foVuv
LtX2F9vhnOdlsmA20N04EztbtxeA50qw4guuj3+poKNKXfxxbN70Y8bG2rR+Srn06Hbloq+aZwSk
77T5+8izpK5uLpIPM/YZoweFLjX5XFQFjT9HnFDTAmbFIPPN5pntYqv+r8tuy8b1Z3iXScyCp+Gz
3rVvC4WadIdV2CU6jBzQHsggrrPSWlFq98zBYSBGi53iZRvMXi36JZ49ZU+zhYOqcn3fKusthfDk
oqIIz6mWSuaPeVtc7zX23DOk+qA6JLAnXXDS0JwZwcGVv7NwpEdwdISyu8AB5gitv0pRngP3FL5U
LiffMwOGLuQL+qSnkKv1Kb9ZXNPvgTwbyG5goFWMW9Ia6m6JSIBFRQRR27ZbLnxCtPGYlJl58ZUe
DgtEftEsuQeAT1OqRvUBjV/ePIAS0IHsLwcI4M6TsGAnSPXj3hcOJgVOOWCQ0FL31k+dxPpLGjxr
E8Iuu7CoB1jeoGhi+dEw/KTlMhGrYaet7bQ++rDOrjXvZFxtE41unxuUPZMeqfUpTwGd9xJMXHb0
P4xmDhQQ/8VMGZVdauIDl3RNsHjk7o9+zUmtoXCLK9XF3kqjjRpMZeh2P2KFR9qia5R3K85hlEu4
M4PWA2grRriUEOsHykEpVW/uxiFpKgF9l6qwTJp1UJkkGPLl2oLc4K2I0jgo1Sg/t7wBllwM66tB
IFpQInMIhfgQRtJW2zktzVd4vo0tULu0eNVFv2WMzUNO3OLvZyGRDYbvewiMvej2iuTq4vdvIAha
dXVQ2nZyi5lmMSEXsSFN80iySbsPdKABU6zJjlNTK50PIIUN1d3G3pUkXuWxpOSAPFabPHEBLTpG
5+kUkzhSemLJ9O9jaMTlAEzvFln5wofAxYZ2u370BT5D+633bXV6GwDMkfKLITBDqYgC0gF/rGjL
WnVdxRi4C/YW/AOQ2R9PV5eP29BU5tyM+cdFkG6zYazed5wAsWi3DjpNEfRyy2a2JvEFLTsfPmFR
utjBQ+kP7x1uvgit1yPHBBell3dlSsSOQhN/0cziuCjrcJwCG/WA2nm1PMt+0pAjcRwEvCG21U7E
2tu8QIyYZs44JiYP1C4G/FVlGTfxWb0LKsoWhsbFg9brN6uJXHGwg6h3Zc1kpo87MWpssoD8lwVh
H4OdqYa10C5MuDXvaaQbK58po7CAMehqWi1uypJgXLzRvIDqQ+ngr8F34iLE0kUuvztEElGhY6GE
4cuAfqQAzAtUlhLGEU0TMgUSSk2RM6L6sde0Q+yHD2BMP0bf2h/94jponpen0QRW2Cpx0SEhqCAo
DVtK4P2Bob6Jnnn1JNg5cHPNMd1xcq+jt3leyVv7WOIc/aszWuyX11HAczgv4B+OC+urnDI/7UCZ
Q8jELbc3kVe/95txgYXJv2QSO+h4j7VusABrmSXif3UFf4xgtvshO54/clPIXwji1cjygxGKxSEQ
CGnrHhQfpz8JqW31PgKy8pcBoFjC/fL98J83Z1YIqBjBoRVcVG18FdvM+mHtQ3mypiVrGd2VWJLH
SkhqtI0tt6x1zEKYqcEKuqmrVdZVleCcdzSQRQdbQFjlBA179Xa/xoH9gMQqI+PlsGHFMJYWd9xZ
jz0cBTwVt+fu1nrNNirupjz7g5cR81Poj1sZz3wtQEH1pBSM1on9I7XIrBRxh2fswa03G3KDCJt6
QjCJ6BWlFLer6rvPNb69TaTB3ol6xsSX7Epf4sdIoW32c5YQXLBFWm+ik4pirrpOcmbotxAHFwvO
aEIEyLUN5RUNnFoRYOe58YKtDN2YkIJroP/eh/4c2F6DBAaoWYe7HyibD/DwUNmn/gqgaP3hwefr
y/0Uhp7Ep4SQOXu/Bo9SDvcN5H6Qpjj080cdeujKzRF1sErZwgJUSQ3EL7MRKLHWL+tzEewAhWI1
qOpGb/lgInXqwg2xz7IwJ7BqFdcjt+0vfbnkxwuTD/sfQNID9o3vmB1jDLyDI3bH6lWrVHJZ0Oep
Te/XmRZPb0V48nxo6ar8aJ77pmqDTEUMg00Q0h1NqzBtHO3p4ouOhUFEiNQapRwPMTk9ErbyYdDs
rH88QuTK45HJ2ydV5RWz0rZw+QTt7gaAsE3cDXltYdRdpuyIuEMRLboYFd7jQB+X3BvBLJqzjjHV
2QEzadimoD5O4G3HZFzaiiy8e0a3s+Bed5gurmfNU84xRyTeuXHmtSTo1eNIspdLP5Hkte5wmdcB
C8eFOXlGVgXubmD9iubcYwBdqeAq1S4NcD27Xf5PQvDVzVPFJLKrgE8q/+bTaRUAgtFTIWMiOVR6
eYwFUj5cPyZxaUYLi0w84OD2Y1cY5QS7ycuq20l8Cmt8FiiK5QuSXOJ5wzUHZS4WPJ9PUnRdxsog
nikN2k//OITbYMKgF8uWAKGi6vfrDwE1Y4OO1DdV6MWLKGqq3EVCXzeDNoAug7b1klDjD/uIMVAs
IqeHfcOI3WmZXdxq1QsmCWInuGEQhOMDAseNl85LWqEM1nPDcrbUGyQFMp+FuFGVnGYXCHX1l0RW
/8VSj1G730JnnKy9zPKDG6i0HqpG0C6q94nBkMc4cmn555JUawaCBBNf+bYBsMMt5LTeo/hdoGGJ
faXeDL/282TBOht2CQ/N1w5QKgPxsICyB3HZrHwdYR2zw6UYWDT4X8UsSWHEF3KstQj93TrG7gc7
BtUUOw2lwmRH6FmYAas8L3T2O9IbvqjwowRVoDGwr9+vd8NK68/LdgUInlA9xQNw5/0EpULuhgUR
1glXA+UBuLTpeajWVjrgtC0v0ZeJUhu1L3zygk9pJgpnPNHk0ew6Yopj8ObGVh9RNttr1XVAst0b
qR296QOKRJacoUvSNl+cey5XOpgvgj9hnZAZ1oDx9JzSg3+yE4sSJh0vvQGeLzIE7NeRvS5WExwX
+MEO0IaRsEnAYU4QTCxtHOgiz++xBSCt5haHXxMPsU4wfcUd2mCjX6EpZS6pDdFSuTiM1nn37nUX
76jXhIJJrO7ivGQDvtkmxg2jeH2nUNfGkm3e6J8pgOpxcatkw7rO9fBC4FEf96f2FBKiWCPiDH93
efRu4HMqPmi/+Cy7tBj2XA7OqXsE3jmfTtFaInsZm3cNfG8EAYm5g+Vbw3wN/MrrUZbuqOV9tJJ+
As1GAcRnfHb8MOEo8/3LpACwR0yV+eu+yE2UaTxlgfzuwy7Ac64J8ziodmuMoec1zuk9HSxCxMOv
oLLD02wPD14OoS3tTkQq9uKfxf6+jgbS+e1MXzKfd657ESzHh7vnF/dba3117U+OCBankfe3xO0e
dzu9hOwSR8MWCdprwIqjCh9ZmlLyGuhTzXzr8JEzq0zx4Rf0FT4kFazoKnQm01S8Ynp3NA+cKj0o
GbKb4tVTYf0Gxg7NJYUG03UlvjV8R3sQxx1kYuYs9IcgX5+78FhWuaqi03yvApW7uU3y371DfFl9
VT84k/uRE8BaaNCNeO4QIHM2739nQ0SVKm+C7pv9Xbp1QPM7Ld/MSOfiNi0N3kWLRJbQ4y2Skq6p
+X0avPjTX14BNgG5tZQBxXhMMdKf/MaXB/Z+SM0N3eHArXfIJP81kgc3IxTa3m5S0a7YQ9AaeFPY
KIH/X7HqKGU53pBEVC5LOYrfOsFoJczOmSJ34cHPCZJ0HGZuVgGPLPhrfjE6fvZR1TsuTXJI4he6
371UYtnSZCLDcKwhZJjILZEjbE4Wohl3UO9Ue7sKFJopkZh6psiziyjaIhh3pDOqbKJjpeOPb0sZ
LXnqjE7RI8SDNFe0688BIGWl4pUmqrnop5qTqP7cDzsPq0sBCSGm6FC6BicRPi3jOZdbG8p9vv2k
xbfllYveuxMMmcnw3VQVwFkLMevl+AEa1tw8IYOXVE4o9O1CelDQFRzFxbcdiwvxeHF81DrFvs1Z
rmGflC+vk/JK0OehzTXpMwjxkGkc3D+Cqcd/M52BmU8x82u5/PFsPI5DKAluNgKS+R1qXUbNNG+b
06YY8csqkf3I9BpeswhdhsXyJX2DlcUdjUneQEZjaRYILkTayAJJO5BmeseOyGdU0F7UoI1wtSYD
kIrX7zfWjF/8lqp38sCvyxBzFBrlS7LWzW+l1tVopr6lU7he5pYb04T1VwM2LxxKMR2ErQLcoXsW
otFkkfhhC6r4eGizz4jSbCzpsqtsLU05/rceaZi1o0aAfDdGG1r28DVvjuHYxmXOz3d95V7+BtvS
tclcHkC73uWg/mYfCoIPTfsPuh0jhtRo2ubBZOmXwSqur6rjv5IHx6dXjKsAoXFiWGhTRImTqNxq
ttPgYJa5oxub0U7nz/naSQogWD0JhGHgU8TgEcnj+kKrW7vKSyWnb6ullAQh/r2eoJt56ODna4rg
V8zQaVZt/ViJP+uqLVqZRt1n6ZfUTEJ1Cgr1NhjMma3zGa9xAHo2y9Dohjng0TuaQn+ruq8o9nvH
iFlNNAgVqYtstkar4Mc//SRw7tS0HInC6Z0/V6C1txHVSjsPmiHjMZoTAYJPRoG1NKDiGUdeihv3
FgLytJ+Z9Cg6HVzj/kQRnpSHxC0L5KGAP+MZZpWYG2Fc3798PEGfH2W29kdZObTLtHHYmYVPMG3d
zIbHeDYgSzcReKKWCPd/8z7bDvo+HNwK50tbvmE3tR2x2XHTLxHh8r8N8Y5QLgU0b5lbT1uCtd6O
iSXDMfNkb8wrNZnD8H9EyES1hgCBlFbiQxztxo5A9WYHM5hUCEvXcUZGOnDuYpb67+Tnf55iYiGc
11o2QaR4BSvOtb6mmSPfZmb8KyEvWfYQX4CchbgXhFZV8zGaexxCcADoeHX4ZT6dkJ53sh24CGIC
gnpfZ6QDnzvNTgSRWQ65Fm2TZrRyej6bHpeTOOYBKucf9lUQUJ74bYYvkEYmdV/487VWiSxZ9mf3
NoIF19Pf1zNyPcJolL+7OpacW6vpyMyVhlOiR3Jxjy8c0H7VIxoBfpndmBSlX85X4AxYP2kZJBSc
OnGPDIcoD9On+UMBssDkHwRl3psiIdVeHtfLnb+s6uaK+B/I3+qwrrHEaSUrccHCHkhFEvXot1D7
vb2pBpcEcCP9c9+Ciq4P70qcUz30SJFG2TlUUcRTu2x2RSMyDalE/cQJyl6hUt8tVZGcaVIgkztL
rpzo+vSFABgKCbuWXRVZwdsUPiX2LiCPsC2nZcuGsKN/iK72sfte0oOZsHdF+GHKUEer69UJK8s9
UeEHgaEhEsyj1AQB5uX2aWzSR0WQ0VwxOmnlSY+diemkZQx6UAe/bJTaWy18bQ0iU7eacVwfRexk
nCfWdhthndsfg2N5ummRQQb3aUPe553fhf6NFpzuWCOth4XsMJPCkBS6U108kXLcOjTc3M4qL7EX
LGeQErbS0ZxLnQV4Oe/PLqdoDFkRzAWrM6N0ieLXyv7/apwAzjsYT0iXHtpGR7WSQ+eWzyfgS/Nn
x0IwTQ6J8nJkZPsuYtUQHKDuKeLxcB97zw8yUvltcFrL754mL7j9klL0UnyikK1qo69X415K+6gP
raV4c0CvmUVyQtL/zf/PmQYwhjG4Jfb9r72ockxdY3NNXxlPVBmzlBDYFPFQ+wytJWpldMcsw+nK
wUQBzI6AY3d5iZm3y8gyPdGoqADGcKAa5XK4vQWPoYax7cRqNt93xEHJxLFLq0kMLjC/pXgh7HpZ
LsRubQ/2bTKX5Y7JzKVn6inT6jM1yDZnzuTUCDmeZo+t20bq3/K8IWLmFyPYN9hj7loD0Ba8NvGr
sJ+htgsj0e0GYEWYhk/3/dYZI9d/IafqI3D1rbwfJj3BrvLsncDiAr0PKIB3AcLiXWRYkdRbtPcG
4k6AUFYORvvafO8K1vSj9W/buTvgOxcFvrJs6c0+q8uEl+avx38xCpgZc77IrXgco0llfPOL9Aty
Fipb08Wd98qpkyeVf+u0LDfuStuTTqPEzRCIv6O2RMH9Q0PSitEDa/tyRuo07BG5teFWtVMr+v6h
H2Eo0iz6L+FZev39GopIbgP9MVQF6gv4Mh2tGa1+Cv6L39CGQ9aYv9slv981KpEiXRHky8/ygQQC
/jIaocoEs5TNFXfnXj00VwaD/4E59u+/aF13ipS/s1i+l2wemTKJNZLGlz6awyjrL9ruSTH+/LZy
nHiOV1TFyOcTU/u7yMbq5U6qhOnTupe4QP9ONLrJvKnXh8WJwqNpmBOPByV/W7+NhJJqgwKTaQrY
0qG4Yy6BaN09mWaJ+EeUSdxOnXWL2WHFpvhyTbXroKfRjvM35sE3x2twSLuukDQcCD/Grbv95G7g
Br7/PvN2txHIWXDiS8QSrBkaDwlQjcWzXJCFxfN37sLK2uPqelCn8vwF/uB/pf9f4DMjocauqTcK
UYdaJ03x1ryLjjotqqhHL5C3j0bffYDoRBOHo0I8JYMAIclMgMPDX+jR6JkQvzBS+wgVeHQ1JPjr
VvETUNSo3FBMDIGvfnJwVzL3mNH8uSByFwWUF0jwSUfI7zX93UuBgxoLMY8wHl8pjot8p3LUSHV0
R+bCUwP8ibsaBJmNsnpUdyn0LX4WPAkEWE6qKJEhYW6SpEsAu1YMYXOpF9UajA0Wz7C55LIB0lAu
2Idl2mlWC05FXGiu2lvdldk0csyvz5F0tbRb8MbibQoi/FhpoKt7k6F/d+k9qckIBRCitRAuui7c
3YvX2ZWGjC3+Ozt9D+QypmZMbIrr6rb/6BDP8ZITpH1Dj1/fmxv/R+XLaQstaQ4X15lPrcRV33/w
RsSa0t4YPk5VvkZBdXiKwzU4jiJZP6eexPBbl1C03KgdTsC3/IIUCY9ebw3Gl0EQWhmkcntUREWY
TKJbZEwM52HZzv5CcOB9yCPV98M9bYBkH15peYH6c1ThXx3S5Jx26pZG06zV6y2hsY6TG2LsrcBH
4dUZjDVxsIp/aWingp8AfeQ07VD5uTzd5oFU3MdIBTwSiK9Pvjc9HsZFuP5o8RWRCR7z3PJ1n+rN
YQsCupwxB7IFj2tzrtoYkHWX+fwc2QNUWaOkfB3ke0UUFHqRKPLzTjnSfkMWVSOeLPbVromY6I2r
ezygwLu/Pzn4e5Qusa986qTxkwEVsoZSkwL61qSoYo4lqk1tnwZD+3pzu2SV7vqoZgqYjjSlqZyj
nI4hPFtTgoV3gHKvK4SU5+QBfMv4mhhfp4SrkbpcxlrST89sqtk1XACRzotqsb1RyDlGcuPHPB51
+reyr1IgzZY0r5mMStIEpcpz2T5pCV0UDFSpNgB8E4Gs/8usxd3tnMn/UHURsZwdQPdzK0yEYIAj
o69xnEDRAafS8fiNF8BuKuoDavAVl484dCtNO/yKxWTFqQrtbNKoESxow9BlMj48S20abWhvYpuK
EyL4hyD2L4uDgDm1AeBrqLFjWQJjaogR+JsJQ4zzw+03DVZSoFsPtxhiqaSRhJO3vz3+J97L4OHT
ZDKdnwnxrYMDhSMil/mZ53EmyssIzNUEVszCNh7a9NaRuFTp5kvI4c7QcdZn+9zHhmB/r2Hlxukz
1lWGuYCuWXSurb2SaM7viyA0qwGMuosW0GTTDgaef8gRZ5V/iRECVb7MDXe/lv936kWP2QKJghW0
yuhIpnoHoSxghOojbMMXeJxFgzPfS5V1FCk0lhX7sZynH0vPjPXBbcB2XVmdiL59N+U/qMCUJrcL
t53SjMHl2HNDrR0fgVzmivp5wYXqnBR9/hhxmbfWPErrTLqbn+jdH0TOUzXFGir2v/qshxSmYGoT
NawE86Xh/+/u/gf1V1AlRUKpWhIReUCpASjtdRAQcmBgysPsBPSSSWeajLL1qO30Lax1uRSsw6AK
+GGozIyU+GTJmzO5VmqQtAmN+ePha0nQhKN/DoIWbPHn3pCxQe/yr0unkaoZaefvP2rwQJuIh8SY
k8g3jM9Bn8QHMdezSl+aY63ymPXWpcuVIE6rgLQDBVTyLkoxqUgIC0xXnyyigUUhtjH9k1V607O6
AKrO4uCTPrnJpx5naoLaewOO2i7hXSfxtJytqL2KLcYmhbnFaqErHphzDmf0GfSd1N0rsvGMPylP
sPdyrSy2aMgSCmROIPgl15LLnTNca++7t8knUpD7t3fYSZ1kh5gh0RjYFXt2Px0kbgMa1AQcB22A
U8ZV0vOKHS+FxcQhxjbsP/QEXg82i785o9aHXQ+rlZFL4GinKtiAZ6tIc6l4ti5PpLEqIaNOM862
edNn7x4MRX7jymuamzeLz+eUfg8F5rIn233S1XaoVu2ZHiIA9i3viaIgZZTLUcIxr4E5P0lzQfWB
cEZ6TW3NNSSJIRHQu8Xb35//3aNAwBPZMAN9c8GSpmdbFc9JW46H1dNXlbjBr0oNtjOHU00lk1EO
KpVVi3IlXlQsgudYnIcTrb7sHW/fDBlQ+cr8E/hm1HzTTjiRKUUTULylwPCGQqFs4dLvG4MDpM5x
VUqDLdwO8kTZxtUzwppsXjAGKrvViuHILka8f9skwtwYLCIVJHJwxMqQgU5pGp78/qTuh6Hrq5eA
ZIBx03sSNF3fh49pyrWs0ICGQHJ4+H0A+C2YR7E0Ixf5RZ1ArWQM2UM+S74mh/t60hHa1F6aRLCO
M79lyqdb8lnxcKgI/l5gNJhIrTGDJKCYocglfA4z+10vacXuWAueuvAxNwEHl1jamubfqP/PaQyo
IgUcE4N6NeOx/CjGcKwAu55rPXxDWSeoP8j2mFJUHoiYNMuDbML+Mg+IVuKexmLESjIB7xIhHv+F
MYHEX5O3DogmG4HPYXEIwMFZOntPI8Do99/98qYV0sYiXTG6Qmg/zxuJej+ibfUR3HY44VRbZX1l
dlLRG3q8+iWtAkKiOFjoY6N6lD9pnqZ8+N0g34d07JdAj6bqPJzG3YvPpdKxKQ52SuxggA/DF5j6
0+m6f8lbTclldt0MZktZIu8GksejAyWegdzD/wBi1QrjyAmTYmv0/uEcu+zIbKQsUkMY4yb1++po
iUJDJXYwxoOkmqiqQGf+Lhsjl3qCir3pUdJD0zs2Y/j1lPKCl2S+uGjqVrt8lZHRU5UhaiioeBvt
TK9fT2CW2zH5ILjLpW0xeGlM7+Koq2WOxys2o8KUC6ubivlagMDSoj5o1v7RlbChqo8vUtSZ4LX1
6kNtYlkuIAuLlR48UAL7x8kLYUXyfUeGihruv5kIU1Zk5pmtby3pFEBbS7uQsgJ1wB+mgIxkTDQy
RNURGhbdLtbsf1bm25OwY5fFXKMlARbXrlWK2UMWx3dhiDev7XxPEYXr5oJuL9DCmu5NLGd/ZF4I
VcWeM7Xxq6dsMU6xH4UUwiT5n5rdTslabz6v3eY1CviTMLPRDMF9VvP2DlZk+IFCvnYX6h6Axkzs
6CTIQvLdL2OSU7wEgZtoH2tfBZ1rKPWtZrIbYMsSkcqSPkoeOdSdB5rAI30g/mMFgYQUlzIYKAey
NQV10JbFsvbxzG3UKWWH33m8yG0hVnc0A9vNxFc4TPPqKKHLyzFUh1A61ndCVv3kz4oPKb+PZxi8
us4PBysTXlPxtqKqRdkAs1FI9P2PMD3Ed7ReHrqIoBqLXOGnSFAgR0ejor8Gi8JV8TBJ/H9M8fcQ
+qNJGMDa9Y9KoP4jrgXQzEDdOCpY/Z54vATECV8Bke08qdydX2WwD9eDFk3AQ93LG1+4toz1wDCk
jAsUeeZi2U21KP2uzjw+n5ZDzCCRPxhnr9+Ov3FjZ24QJEhGh1+jM7nsNMOd2jdj6CJ9m3W6Mvza
76+yHy17e0Wb4rnGvIJ/QWps80hTqwbWDC6NMHuBELubuMFPcEuWd4Cdn1Zw/DpFLm2zVMq1X9oj
ymeSeAjnirsoQCFKepFkCBbVqLurugoDtC0dR4ITog8WRiCiBcHWUzxv+4eDphfty0dPPNnAR8Tv
B10rHHjz5x893sdgF6vMCvm8agoCHII4JTT81bOlnw15KkYNqGyAuznQKSEMZIZJ6qnEM72rBFZ8
PqUFogllT2UkAq5SlYHzr40H+Cp8N48h2DMVKJrH/PazYmWxO1oAEK2cYPyBIH6Fj2TBTJ7Tus3e
f3nAxshIhk76L4LYJlo0Vo2BJSd22wvoN3MBYhVr/yElX8u4YHFaq6chdFW41Y1OYIPsk9ifcNzk
2yiyQ1N8TF46ki0KMPC2kBRzSQ7FuV/xU0MZKEcBJoCvfxkeOukgbsFZloLcU7z+Wjxg5BjUMDI4
aXRw3HzkCi3DUlSABYoHVTshk5AS9j1CvyBF7MFoJtnnqv88OO7CLRVbyQCqx1Oar7p714e34VQt
9XDczOUuU1TmvcsmN3l04M6yDY15PWrqiXzmWy4w5CyQH4IJw7lrnEdE/B7yXXV7AGsIhmabR/zp
jRhbowRHy2OVMi/f9wDhLqIDl863S29cW/cwh7ruWKFnQ2ntBEpYIc7jRW1XhcbDdbly/mmK9/+A
OUHf6vUKCHw/nojBtRhYx2VNe0gge3zXJEXYgaORK8trm38tKGWjmvNdUTl26lTUt0tMwkPCRLCP
SdbN59lJw14EWTZMahwooimlb6PlukGZgEAs0FqnVYiwrn+IXtoVw58qRrwVp7UB7WGEoIPIq64t
QnC2K+IWzFOk5KiuR0fDngF37uJ1tmIE1vLoqojs+vjrKiLV5IwcRXhGy17XYcTrROqI3UZIxCHx
BfjIYj1BAj2rgGgVueZMJv9+TijfPsoDlmLY3tiukdhRtvexdyJqDnuSBCI56ZXWzTGXZZLq44AS
bwBLPHKyA5jWz44vAjmUEF2XUa0FETcJnAeJRiIOPPy989ozZV4WnVGUAcvAWfaJLPoURBq+0UTh
81hFWaCVngb/szIyyCuTCTHVZyeda3xVOGnvrvY8/b3Ysp0UCnCdW1pmlVWu4CTMvUEo+5YkhCiu
odTbhc7p787jGlDrCh9K3QjPfAtHgSXyP2HyJORdQ/aHEhnOrIRRtJWNeyukggM4yxHlhkDq5tbl
2NSTnno8CQ6nJt+BBHJnCv4UxhSP84YuqLIs/i8WyO7JSaBtkvTRTTG1ktNfvDr5iVfF3H4tqaLT
AWgtHI/BTpCQmda+luDQ5OQzK5Jjd9UMzcJH+6S5iJXndtkga4Lue7+Yd1guL7O6cQOaO/vlA/vQ
bssF6h/3HX3hwXDURycLwCKRwlpn6H53RdhHSQXoboMNjaILX3J5/6XW0vf2g+LG0XQhILhIeqTU
+6mtZUnMWl2WCBR4b2mUWhI5t0xG/NQLfmpqbDAFZBBYmEJPcP1ZnPUBxI/nuuAzNJDfCizu9UWV
zwAlEPln/CY936a5wqJeZXt8KMFpjsWxdjwhuTvA4moMrQDt8cE56bV+fldFtnRT1usEmP6AoJjo
VeNh4PHXAFGEu8paSROPXlwLVVBXs2nLB+dqMAKL3IsDeTucXi9nvfsc4VeSHB7ztdr+uClszJth
KjzmvftshR0ixbpVsMqqYTPjKc4hGSnrZwmPXvGke9zq33ekg7oRCN4MMLlENuGyYRQBIbxyY2Un
WvILVbhKWdp5/EJ78uK2B4/q98nY0VjKNS0gIg/wF44LrN7pceUNHB4vIJG3VgE69mDV+sqz1nwD
p0U2d60yNFLCr88r5fISZz3pfsQiVftlsYC7h2CFOpPnxelRRl7vFsGSO+pK0cZApQ4fI78Wy4Z0
/htxSyotaeVedbvYslTgGXUUZ5iD/RfLvZskQEo5Fag9XS/s+VV3jRgnyEikAHA7Kb8zbxLKgms3
BEYQq5AsK9Mw/QwUDcXSiv5pznfXGw+OtQEgO1skWR6g/pHB5z0lQCQH1S9PBLWTuNcxR7BpkZAa
ktzOdc67Vhx0xcEIFKPMGQodUtpLGcfQOg+nyDSRe3VDiHux3h2GegwzIC5Pa9C7m9ksXCXWG0E8
BdqdmmTQIPF649d9vwp2q/Uhbaurv/Lpu+sO1faCis18TAlG86vuIkqDx4Y8AMmeV3ia8Menv6EZ
Z5FuDZIBUBLmRRqR1dHqSgx9NeXjeVM4Jlas8ahukzIWEX0GuC8aY0lCx3MH6xlsw2dSPL7yuzQP
kqY7Vgu+ILxV/ZZNGiUssjfxqPLnuO/UpKDMmq8Eggns4LZL08v1I9WPg8+18S2s0FxLH9S17z9I
SJkvAWu0NhMhiek6M02HrfUcPU2LFtgew6W4Mh+xo74C/OasOgIMTkKmKUifumatyc/JzN53Oza7
Z5cwBumMcBe08qzalqD+XSLG/URCRVXeHJYzUBgMFUF7tziDIvkO5C9OHF3EtjvZK3qQKCjQIk10
dpHdqSyT98glYfXSwG/GuNPg3W0Slxg6nW4yhn35mXJjVd+RaNRL7j1D6CbxfwzfToUudADjO+yN
UcDfmQEAW/YiNcg0yxZvqNsV1SrT8XHpKrvkddkJkceFxJi9jT7CDdgZWJm9EkXuc74cK14RjrS4
75QR58hesONrbADWbCdWJvWYvvGQasR34C0uD9rI4wZKONeXXmVbmdXFVtg09b5mikjLYrpJKnkN
2UNmUPf/zZw65FmPESQdelEqzeELVdvpw8DDjOgPki0lmCN9vw4B7asiBE0zSCe72M/BQQZXFn5M
9jnGZ90Kgb+QAxyS6MobBg1r+VmxdFT2i4nk5c9qGnDp8jqT8+rytyqVv/MjxZ09sV63DSO3W2Tz
BDfO4aEzZQlHBO2Xei2hYcbxJLU0qGn4WL2TuqCkB89IfiDjhvQUKF9sE4BYsD0o/Kot5PF546JL
OUVM4OwR3ffwNRX/3MUxbZsX/ypDt2yBFNGIeqhrhX7eCOmEApoXV22jPnImIJUKfM1Lb5vCLECE
/03LAZqnLq8MM78mllj+3bb1m3Gt3ztn/ink3L+YoWh+lSubc//GeTtlTwm6U0ZEK+Tzw+tZbXuT
2CBsdPM8CgbKGFplhhpLPijK6eLz6NmpeV5dQhQYijx9hy5ASUJ5kd5+I9GK4AK0bq5MxU7GX5Ji
rEdy4zGSpew+XKqqvvYkMsVmlZkmeyQniv/IsBkB6XMyrvsdbB2Nhj7WZ1aXvm2Pk0KKdaQ1Y2SM
MvXE4hT1veDR6KO685J/5Kq6qDn+zD1rg4V8hJmx4dR5CRkosUus4SddpTS+rTDhnJqWn10smKjb
QMaVdJZ1e5VzSX3EvMPhj+2zED8kt1TAcSLK5vmn0dPDlemCB/3hxTRPEe3rslZxygY0a9JfM2vn
R1sLbfC1P8AAK60++ejKgbkV2Lymy9ySEjgkB9H3PrrmqN5D26/Hz0VexlFJHNRyh7Ytju2kim0E
am0Vq9yblBMeZO2kSimF9uPScruslAdUsZ0sjGiy/DgVtkbTOX/PD/hpkFvQtpegBH29GvGaUZWE
2m13O9Mx3robX1KHIn1ATnPm/4xUq7cJWbxdU+Jh3BSxEpdEcXTjW4nAby+MXvGUOv7RFsyApZjX
00LbqWH512wn17aKGPdv/40KdSGHM9VddaLcowWt2OADr1OH2B2dlJ4gpcy1ZN3A2QSHeSfokaDr
VpBrFRgSrZqnaP8ybGawnDYl4SNbFPvFMlSvvuR47SjtY0LyWvG83pFG6ctN24DhG6VmpcXhHrsB
m8m+7Nem/dMXkaV6yz2vCljnmQ6XMFE/a3OYmG7NDe092j1zgZuGw3REZY83ybWS9P5fl6QVLkNX
HP6ortPsLO618J+9HOOftX6WlMxlqoBQRGYYNuOj8cltQW5M0dvVjgR6k4BQKRBfjNfXxDEFUyNw
qNSRdYjA8leOisOnn+LsD2gHx+tdvk1dGdYx/SlAYMNRFo16vcx2CVdXthAfXHBdXTlGjv0PcP+a
NnBnTgU2OkP0EXWc6NgsobcbSqGYKAmasHazpS3u61xY3H4r+a/4oW1cG3QW7x86/pPXE0pmCliw
uMnk0BYk6ibn4gjUwIKwjtd47QsEKJ/G3uHWNSWjYEUsUKYw0Jydwcqs3G9XAsiPRCUFpUDTfTt4
tYsz+up4rR/K4kMhYhkhmWswABK4b+VlYaj1EGtcMv95YrM+ncQ3dVPlAt9SI6Qw4fpYouncvEHT
I4RmEv11WkPVgyi41nmoOfB0bb6r03l0e9QIlI/9khqhLpdPdCXcT1yhMGV4KvfblmX7CXOJ9BGZ
gTJ2OJ6x07zuql1otfqt8193oFbObOTQP8G3s+OJms32jMoWuWtI4FxxkbJinadM0TqaeasYvGMy
vn21EL89w11eVqZUw+N7OYNd5/fV8nXRUiJzHDj03LaoNJ0+FH6rqv1qG5vG9MKUfpztMT4/movq
U6jMlenN1SGQT2O6u5xVHiEruzvNQvwjQAycsjWTmWgahy8QzFBAriFbyG0IqMAAUH+WLThpBeeq
CyV++bC9cwejbe3UMfLUZzIBp2qAkxJYs7KnDIH/o0QNvIdelWrn+7kuOzasJ10jkag6zKXU+xXe
zOta9jF0tjMKnYnPK9WvBdYfwP06juU5WHV1t30KKT01VfSKud+82NokG22k986ZPqumtNjJCvfO
wo8wctinqzKzVnpACtfp8DXCQqs7ygRc+GmzX+vdnYvHZ2VeeHOrE2IsCuAug8vP0cTYxgSnbThp
wTDcA+JOC3MsAeSKMtXbZ5zWv3g6JX13aU8nqVw2frwSXH0hKmx4RT8XTIXxKgwfMgDG4O+a1gIA
/ZYSAsvWnCgEO92As9/pOFRbqFhJFiycqh6Jy+Lkcv8eRZ3JG3V9RJqzXUwsr90fg5Ylmvu8Z5vo
KLCIW+8Zai7zw1bAcnp/a3v6W0P3SOEY0VKid6HnOmFRS0LveHGyKzxtiHGrqyjpJwZWhhAgX+Jx
qhvoXcRW6u3LDO+rwFIUF3tH7QIKxOCvRqgTyyO5AjrHCIB781sg1kVftIn6eIFfpf7ZNaV7ajIq
GoJMAhJyyEc93p3bghLPmgJjiZIXYQqu+nrUIvZJru4HzPD9MgbYvWkLLLZJ0tqVs+KkR6vqktRA
/dlkyYaM971Wye/JrTV+PgVl8LjaOpGGG9h2u7m+MJnASUk2u8gZTK7YIqSRZDltqeLhqp1EL7jM
sRHR5tFvEKeJvYSqjGOPxTO9cQe3LMzKS4jhUhVPXDqjzEbqDe7jhShCpHZRXwvqLovAfB5soc0f
d25rgFq5ujs6qRq5PQ2ErKzTWyxeRa4m1VKTA2ji+QGdxsiTauqahKVSmwJNnxbhKE2U69JlYuj/
BQoIn6rL2NznITHML5O2jK3ntJ4NWviJ73o0AYlnK0Fldc5CVssZ64piMSfBRq3pU0b5Mr5dlCxH
esDvdzzAk2qhCJZIriYT5KFwCuekHB1t8HkuXCNw2rjCGAcZMw97hJ7t2afNJFNCTwfGGSRsqt7j
2inZNjxQf8uzydxV0uR84YXmkszIp7UQ55IHMgpsvyp0bQhs9rNkmGEAdaiSUvyBeCYgX+aiMSsI
TJKpAGxF8EtUjUufRW0eHLbt8TqRJfvrjkgh911BehnH+tSwbH6NqMOyipEHw51mCGZ7NuPZoYA0
68xN/nECTxq4OUE2TeqbjUaqkK5tAiaX50Dxa0ncKCeNNpKInogfmB9U5TxweKwqQb5A5HYbPm0D
NUcD3CCzdBmWrMdez8MD6pROOjz9itguwxp3AIXqhoEuoZzci+My7DEkejaEUQNzsUsAI/MwnQhs
8WjB/q4odyVBx4p9Gw/PrC481V9TLGK3zkuWtdpBhNZc7ihwCH+PWOGMk/H8TpUyZj4zvBp0a/fQ
+ZMFv1tpWwgo2jqnuN3enqwQE9jIDbQgTANLfqKTLpFPbLmFhGpyMVa0E7JRatxC7GXlBFD+aS4u
8pRvh+aD46VqEsHEXRfcQa8U72g1sprT+RfAZhODfgczRlRWW0SfUo9DMBFeKmLPrVmxubTyH47M
8m5pNtW0eElVyDlGPz2EUMqsY2TmEf8AmofI6rkY0OKcyfKvjWd5ugbHPXUgMEvWhcb0sDnThkBG
tB+d2KodH1pCF1QcRnFnqdF6JflA0pMKsRqV1udndbjbsSHlG4yoeAg8TRWMyDWnyyieCaSjb7Du
DEPa+aphh8AXd08vNVBgKnIZNxNQI+c2FGb585cxX/aEzp/lxcfgTEvPBqOGAnVLhkNlmkfKAPQ5
wQG3RJfpGrSxb8osii5o1YZZ2KeMXmx18K5BtlHAk2YurVMPFRM4lymX5O+fhtySx+xqMdcImUm5
0QI1egxQ4rW4CxB/OAUKuWlNvsIBKDEg8hmNanex0m0z/w5tKIZt/16TAOb1lurpvqcu3U14AOgR
ctrJ/0/4lkL3cnVSkwx+Q/sgiXxwJ6btvef7TSLqN56o49SMjGMjzoEauPoyr9bceQx9/Pc79f7B
owBltekvKx9b0dGJ+j4JI1gagaX13mca4UvyVQeVbzQU1zXyO/hLbD5cW3EMgLLqnAtbruEwcYhi
6Dy3OkJA9B2ejSGqbpYrfZlGHJ4JyEobW0Dn+pXgd8VU3/V2yEegyW+NLJ8xAhnxcEKlgBmriKVA
ijE3hszfGuw6mDV69CHe5JSNI50u+IeDu8SD4yViYQe2Kev7DWFxUwJxNQuVTSet111Nn0srbx71
GMsc6Pa3nzooqOOuJzSPq12pV95sgn94vcCSlG5wSBXWcPktnWIgTzXzaH/PvzY3UI0zzgqeLtir
WXRwCv4v+TilAOXig0uWo2gt2s8AdGvjzV3ycW0qHEdzatwrSI0Bk1siaHp2g813A9mmQNd27K5v
cbBVil/2HZDt1UecN/NRNSXRbJUl471OmbLYPRGjhuKIWvTWkU8RGe2ZI4EHJ+FD2cWvEfnh/tte
w20yZBnR3xkc0GWhr0vKO9adFXZd0VfhLUXp1+rHZrwA4Xm1k0SYFebeiOYpbSFCQVGU5q9WJLvg
fV3dZ3zvF0GH7trY79Jl180y0kZTzjMqai+zgSoek1FcbCUnCQstDan1kXeuLsNkeOq3CYABYvDd
TKXLr44HHOjmE7LugjHGkLY+6o9UFObAa/Nz7LLV/BtAkuYPeR0wE4U5yjxkcLr8o/ql3Grl5YxA
ZBk4hxoooSQfVZpSN2Zs1CMOfuq5ysfFL7MAW4B6wCAqDjogAM9ygM4Z7rF9jyCMh+PfbEm+jVwe
DM1Z4w6M/7uEJUQ87gKPKGIS4bKqrkX0LR+nqQWFgrLZtiBz/X7ZPFgpMfBgkZJLppOvkB4v2ilS
gI1w4pkwZWFmDmtGZ3CDcMtVmx3MDfwvL3sJxQqJ0YsdaPhCFK9e5rGRcjRlMhMiqdxjZFQc+g94
8nvrldP/mY8TnD6AueFTeJN9SX21aGvkz8dP9Q5ADaFO5Fac4nt2jBAmT0TnkU+G24etnO7HRLhJ
p7U+rb/22lFpwxTRvDpDr47ZgHSpabFMk1/6rEmC7DHeMcWbthu/4NLwh3S3wsWqgSys9yzsFjHb
aKhmjRIFayT3sfCQSpHtlHiwQiar4W7u1+EMTN+HS6xQOFpaQrAo6EG4PlQzJypz+8JZm0aLZpsI
byBGWSvFkD9OHHF59WHnaeSWet7Z5S3QbO7D1gB5EooQio570pxhprEEF5xFJOlyhPmq5BopiaWu
xZguonlwTPrf1xwVTK9GRdegnRXrC9vVF6rcDBKi0JSdCNTj5nQQXSbCC30+xitIbM8+sl/SEXkh
3oCop3OsOujnjPTb1iI3oTb8M5mDVKHgCvCKf/RtEV9DcdjxKFabM/cfdzXdAH/YR8oNhQccmG10
8v1rbSNBqMjepqhNjOi1S/cOIf1iP/X5TwjeQhoz9oD0nFCQMIq3YXhNN+CwqGha6XmXSffbEbBq
lmatV7rkOju8P30bFeddfKOuxrQ6a8G+GVWFNDpiUKFAg1dRrMXd8Q7/R2iSHLfFKWW61vDh2jgv
Ar52Out1Qe9Gw2foBTGNcPo0q/6LbWTyVQHM2YvEXOSrbxbql/wIBUlF+WIVg1mMWgJjGtcK9tNb
ovi+9KyBszWXmNiv+IM6FVH7u3kJ3/a9z7SwIVSe2EGuHZs8wTrrM4NcS+ZpmYmbjyMIoAeBiKGy
3yiw/6e4oe2eeAck+jONLeB23PeEYpooNhjrWtVkXU6CqHzKUVEu1n9xOwY7fwy9MyPBcNEVLWse
zk6N5uCUwBpX8c+3n7s1vaw2MwYrRimyeMIhX9uWmTzgKHvF6qs+nWVcHPudYAmp9oFl5JOhS5+C
Hrje/jY7zPxql/3E1WQIMBj9IPCk/qtS6yoDhCbE+WSZTLUQ0M04QQaeUWoE+PiJDmHkAxY1twMZ
XyFEimG1DC3DJevkzovsyXaGdtwP1qohe9zLbqjkFG+pOY19kxa+aRUt3GWQI+YGFPCP6EglCb/0
W3N/KDYwJlzLAxRsd9g2Ach3AqyU/6d7xqa/A0HvSuqTrosQaHNeeHqcHaNLRi2jlq9vbGMtwxlK
Bwmr7AbOW0dnuadz/lEarxq8/5gYsw49vfXEE78ggyRnlDmOu6hKfc7MWq2Y7CwbVZp4Rg3wlqd1
GaReLw3BiEs7JrLoUMjq+3xvg2AF7jM4CqUF0bLsw6yw2QiwPwrqz08Xs9SjmHyNwJVAM1WR4FqD
5d0xCxHRs0G8H7Awd0pI9IA1BsgcGv9onFdU8JvCcHhcrQK30+b5/JzA+rjR8A2pVhBuE4WaR7Ky
pLbKhWEWDrSLyEJJnlgbwYIVvv6Q3QRylHCoWUokI8yvZMqEh++cnYnWy8WgO9Ml8Nf2t748NF0j
7jTK/q+v1uFs58kJHI3juGeJ7CUifZzYpinK+KTSETIKiyDto8v3ZsLaQslepxgSsq423Pxg+eCO
pHY+09WEGCnTRIAePk04Lbpj8mRbmm4sg/rdrtzQERB9ayAvr7YZoo+vgjJeYhPa3oGiU0LzSuUw
CBkuY0CpuvfPLVdk5D5DfcxUgIFTT2PvZfeRAVjgFP6U5zbn1EpTGGHxPT78ZtMgah+dx6RG1ucf
MrjX5BTGQmwGcqbs0yXbrL2bYEjidAyKqyYv4IEZ+vXRJBqvThlEc1WRjWzDD/GrwVFHVuLyHY/o
3iC5fMtmO4xBuk557g1YCEzJB2yzkoDN0oKp1SQl5Ng7JVx1KB30kb0gt3GfMIkx4KnOx/1QxzkS
f7z66NT+bwY4lMLASveTDtc4D/dioO7bx4EJq88dpBEOpGgrO1lkWetlQP21ST10gBh0LEPZF81H
865Hn3jWyOAxWF7cIbHxB3xqETsamBwAnpqnKzPgj1DdS9cADdXRMOpo05PrJWyrmyAYwmgSEF2p
++rgpikUit+7gWl0j6Xio0/BT6etTCX77terT/lXC7WSr/XPMOOUzBy98oT5/UYe6W8Sr6zsAgAe
pwC06A5CKmNvg8OyIMOyynNXd+7keJG9sHy5aCGM9z1xXTkq1eyaQs0FBQnjHzMYZ0dFITYIQud0
rbLw1l+AKDyRMkwPgcbzC3CNeXohpOgOzCUfui6QKQZj0z6V7yvZJ9xVsjh8FvD0xltwqJ0iuUT1
LKRNqf8Xs1cqqFAb4sNfVKf9cAiFiXHQwPgatbpnF9UAPI49gfOzO2XcgGkb5Iw7BGFtuSLnlYCp
4nAiUlHI7qfEaZjj1WGfrz+Y/sSTI/MiC2YgomwjimWt+fkMtgJoHY4f0Png8syz2nfLrPf/mUqa
vuR1j4iAof2sbEeHVC3NaGzd/mROQeUsn0RIVOch3SCwhFAgMwOwueUUZulrM58syYBVYG9//nVQ
UOZB8+iEWriogAcs1Up9rjxwYuuO/XoeWvOQBX6hVNMj0oB2Jw4N4TuUrCDAyQIxRT6XXMvtN5xH
xcbCjLThW1Bi2BMy0bCwLUpJ+vNQS6rdH8m0G+/Zye7j3JP5sMUWRklx0u8xqk77ARcOsAntgsWZ
xV0/5eZLFvpsQsQ/B5y89cQzYCx2dwWAdqV201aH/tTOZuDNoWMcuJ6HaZ6xtxVzfej2AYN+Makp
kThyJzdgV2R5O6+KGowszS3m7lvk6pqvHVdtvGqKXS5aPCZd41DMopVdprCQLMObjx7xrLQcVbwQ
xOQaS7KqWxgjZNI9/rjzRPmZaWhMgm3dWWHgtK8Wa8nnT2r8Y/xqlG4CvKuEjm1STpZkdY5fTHuv
XRmZiL1y/XtDOcfmHjaRo1vgRoSTMqA6eQsXU16664qNRllUP8sWA7KNDfDmMF+PV9ZBgpYKSogb
XXK9GCANt5Zj52MlFjQuBYO8fJcocS/VAnyKYTZ4t5fmL5OBRFUDnUz7isswnCh0hQKmxiUUV9zc
iREyiHloWO7/D7QrUrHIoxrk2tGrfobwHNvuHpwzl0RpQ+G1oF3FRbUqhkdtEQNKndMn0XB1bIqy
48tPK3GhK81gnkDxRAa15BqOSiSKLSHc7Q1APbWABiAIwm1t6zJk6SvTG3ennS49HzF2Q6SaXJ0R
UgdROXXeuWDEePd8zK7hfJROlST7kQ341mfWVpRwKfEit8ABeQ+kA2iTNSkb+jq3JgntIqCKJoed
hlRfTkwjg7e0skXYQpnWBAlA+oZgMIvt7ZcQ0wevgHWEQ7qRHaTz2762mSNklWaq0Gt9BxeC5Zpd
yyDSl1g/Hn5tHeJXsBvXH0BIS2pErXXxanU/q/8l0EXxzzz1kIYJZC8gSaPTy/3OX8P+tApAGmZW
EoFjA0cQqKCLz3Av8ISRtZE+fDlma4P8mEwS95IQYTfnbNrhqBghPSi0lWZ9Fm4QspkRXwKbC32F
xziEP2bKrdkXY+ZZYcUQ/VoIUx284DOOhbJ51y9HJDb9XCQclmMtzQfawKpkeOzvFX0cDclD2v76
TtACOnpMbytL5XDEUXrqzM9sLQjml0NiJN5TeMr9hOozFYA2QQxibPOcSOgl2WgqFiwGrPcLxnpp
0lriUwXT/x3d00FSPYmsp6wvnYYEaIoGj3vu70KQgHZOT77rIb34gXKRykFBzvHuIn1wrN1KAzmH
LzMpuL8YXKjIcPEEa8S/7QQSnuzqMFt78TWejcaiqrfxxRGvpZehK2BuWy+ivWXzny1bu1UoHh3p
VZcvGMIoDak52uH7cbPR9bsoysMlONAxK8MaXhys5qIcORMSyJzB3GTqbb1V2Q2KbppZdDAbMssM
LdR5uKsqlXj/Lt/BVQhXLXVDieAWpPN2iknJwCfBfQQytSRfSybHJNeVUxPUOa6mf+Hr3Hg4q5k9
AWJoGSyGDaucN2F/KX80uQwWLPKnyRqvhzW8LmK7ywy3G+p4goCP3TtkVYPv+gFG9DeaAIimdk/j
wrvcF2Z9s5tHts5UTbcnKcscBNEwxzY/4ads+Q8gxK+XZj4QkUXnxN0PQpmSFBnVi9/uUTqDRyKq
SjqerCRqplXsxzvJbUPjRWP9fl+4oj2NtE+A/PUcIGp92+HhFPUxF4jNz2qJ2M3I0tTPSSoThiBB
5sZks36rwrTOZDuehp0g3lB0G6GCQe8nXAIniYI5HtdfCO/I2JkIQv994aPl0Jh03NBVjfjDCsgQ
7rXn+mduZUY4QqUBiMxKmHY4tdgWTPBz4KRg4N75HTB3TFGz+kjdDVqePq/uXy4HAD0xN4kxMXry
/EVURuT5IBnIVex/B5JtybOn2lVmgpBys6a39s8ZklsybuouSLfYEjBFkegpILo4QIWf/qgq6QJu
tPTa/8Br9EBEglGWg0dyL5HHuRV8i08WQL8aQZrfp6X2WlljUA8EOIgfkgzTOv0YQgLNP1fNn43K
2jkIgwInuBtAIKdkZl71fPW7zPF6K0312+JHgaXplGpAIElWpoLeUqHC3RHyoN94VqttAshzKP6y
A4+CRJvcsOEMGFNt1L3eiTIwiWOTJBcBt0NzAM3YA45KoY8xV4fc8EZiIM/EKAmDTQx63m32gxlB
TXNxPnbQkflAg4fV65UTXSefT82jGPyrvOixiZW3JOqpbpoF4QVwIj2egWtyJ2PKUkah6uUocRrQ
ub2Ah8V6RxEjaDE4DvP8zohPtA/AIL6e4+IrnIknknB+vqrgIDKVASCQhUJf3JbgaUa6E+/X0zLx
eXLEK+ECgqbuOQKktWwAeE0g0WgsZA4FZrFeDmQmqZnS3R+x54lhKyygPiiwiF2vYU9qHUq3CeSa
ZA/l9DSKJg+UIEra6BIPDVI4Fm3K5pmS9mSp1XLmxSO/7ziQhdAWs1n4xbE7PofFXg7U++j+zfXr
agzKk14hgjggg9+53fiMnZ0LA+4KmWiE+bWLCoMHvsQN70pikN99Vs8lA4yhMkFWDC4+Q3Kd2bme
EVvqwozqlpR44gqp6gXXdckeYLlwN8pgaLUBlLJn8CbX+I416/erAIS5pqvuAvWxnrkK/eQqq9db
yqUvzZG//WM4Eyl89dQNS0bLFFUJYYZo7FFJ5pG7aXagQ7OHUyIGU3Nfpv88XjVxFe7rhDsl8yoD
u6VoNumd5h5e8nj1BxXV/HoviKcGVIGdncY/qCncw/b35VtAq2fvra9fkCK67m73njU0g/EXYYLX
bukPNmRKXmmatLAGLyzgRcOIh8J97lDyFdI2xWxaxvZRO1CBgOi+pYtqjpoU7RFK09lgnrl8kIDl
9TCj0+fsF2o2zXKXg/XudfKwx2k3qVVo/18TUV2/acIJqc7ulc2FvWirqduMTJu7ckS9R48D/Q3M
/QI/AEBXDCGFv1isQlHe+6ODUirsADxGRYDcbhJ+071g2dUJQT9VuY+6IccE2IeUPDeI7phcecH4
KIxzNrwVpooQVl6OKO9qzm1Krip2I5bdQDwT91K1fzRJ+BNePdTwL8AkI46KGpPw5Ya7TTx9L6Q0
viFJ07V9J6aSPS+X0EtuD0MzqbWehDMIqRub1Wkaa+iSf4D5oCIKHioHnqgmXlK/YUpcboP+DsN8
Vje0VTS4Fnxn3KLCBg+IZObK/9p3mppZiAnzYvFcUF9x3JDNJIkJntauY9bRP1VEKgfOnc/HblXS
2HJ+XmRDUmVg9zxTm5JvcsllQfs4g7tvQQ7AsJWoaQbrTMVv6BcJKTzhia+q/uY4IQx9+sELuvld
yqDzGbL3EIAU4sVqgeRhjvuZwAw7h1KmK4Cxk+Y3/cZzWGBMYjM41vIIbLwUJjPyCvzlsEtPCBgM
T3Fig1dmagvIYnBKp24sIntVUgIoWwj/vW41TlIXI7go8pV2yCrYsrJ/skhRqtaXM25U8rt2YHyf
8+hx29N/h9JCsk+R4Ds0OAC/Dm8cnZ4sFluFn1lXnTd3cjdIpNW8N4Edn2FJLWhC/IEap8nk1JN2
IZJC3JL40S/kxlZjGQqBxN9FiU65DyxiA6CelshM5w8fua1Fm9DKt9BA6rQjDVbnmB+o2WEgj3qR
PFGQjEhYM3ndv2rfn/WvNvXOn6oa0uSRosh3CYsQAaXEsSBCCp1StH38lxpPZW1lkZjaCywKKkPQ
yQQ3wa/5m4A/afSELVDLAw8EMHGvkzzoigEsEybp/H68q/C9Vn8OQulY6uPlXoJezMNXh0rC5CuZ
fbTgk6pn/4HihU0SjchbDNBiyiILvZAokmu+fNOX8Pgzg7O6mC+lKSxRkRy+0HeHuCf4kdWbqzoT
QysI4zz3jDv8xKC10dn3BtwR7Nb9Znh9jmeKQxOXjmh4UMiX47s6s/IMDGk55yC65KsT0ftnKNbI
0IPFZsZo+uUkzgVyCjrcl0RSzfYxuSq2iHAGaK4eNZPcVZBIlOOEmosNz4rCIzhKSI+GkQDtEwBM
Y/U2CxZW+a4hjUmtwK5EtIWU3mtXtsgwco1RLIJtaFWvjlwfCz3yYxR6TjlRzJzJRgvNrIZqgiVx
YcsFVW+vWLgq69tFNftV676GyYOayefTnTQTcVg5X2TPQfGC0PN65Yrek9ILfzKy3PDm+UYN1aQl
FnMs+KD6c8sS60fdfJ3zWbZSynOuXkoBLWCx/doqcDfo8EDzjpLi5rTBGuFs19S7vEqWoI+fW61e
3Z6cAOy0Gu2QdoR29cGov/eYUkgSCdhHpOmOhcF1M6i1bkU5qyfqHLTsahapeIwLvaMhErOWfEaB
TD1kD9HgAO6llTZDW0woGK4wJugJ+lIsLgflY2FuhM9q09GEMf+e8Esq2V3XZtJjatvRAoA00qxv
Revejo6bbELG/eBwL0kaUDyfhDk1m7udcuOqE5MmvyYteqNDD1Xauwqz3WKFN4pwos2MJXD/kJ0f
gepZjCZbDDYk+63MzuEXe9cYIhpo7ycWPPnxYqCXBX4AihWyMxq0tntjRbqDxoK6C2suxZ06KJrm
OPgqRG4e2D8LpMLLg4kjzioP4JzknpQhTT2lLyq7P59OAUoT0jQ/V8zmsPMTXDlM7Oo/svYmjz2m
KRKxdcmx1VifK6nR2x001gSB9ZUIfVZVIovAT78L0K7GbW7IL8c2O1U9c9YHBsz/NiB1/nHn0wDF
0E+R1gvmLnpzkS47zGigUG6Ld/XOsJUnjEWyYMviEH2U7zc0+rgOVRR9WKkTux7dFzpRJn8xMlCT
XflOC3+1qgHUPQSbzsOSHKfbd73iT7Gkmk+7vlSTQQPY/n+j8sGBOIw1LjdsqWIzk2OeopSF+e0E
yRKby0lkcJjPJpnolT74AG9HXQhMkIMx1fj8b8F+DGfOQR5+6GOz8otCi7C5Yzu2o53yhEipVjWi
R+2Qs1MswesOZ0sZcm058GktbE9GwfY221XszfzDwjE8VLgq7kOE7y5pZqnkUKKUlOcBfXn1WEmb
nRZs1roYpbfa/eu4BiNt++EA094tcgcK7J6Zq9B7/1MV6d8FFmfv/wk41xz6mGCkKsot/Pdry9G/
Cui2+m1Jb/WqtOaE9NugBDc0O3GitbZtHbJ74v+k56Z6p1lwkTteL/pVSh4h+hP3ShXqAj4ZPfFZ
6tSYajX2IHE2ic2ghcEXYXXexjWATToD8mnUBU6DNWrs6KjvmpPw7NFCVZRCHc0uvAdTZ8wM2055
nZ/lCy0L72bWsFQgrqwNDhgUjgdPiM+wGEadxlVz8pgH5bIQDMO9X7ZnwEyL2sQ5V8WVjPD3/LB3
cQwwphPwuyTW4c1Bfnei11SSsHRmvLPgD5t/bgWiWWO83+DxfcUA7Udco6tNaZRqoPp5ovISXH/v
lWmTKFdknuadDH13u2hy9T69GC9DwmfZjgP6yNmy3IwBUHBxcCnKFjdcz4Dj04sgNaw/QreXzWlm
1rf+LTY73RH2Ke5FhsW/GlMLQr7jhjws1ejlirA3Z21vJwVStA38GOKEzZglESSdQZxSu9KKzD+z
vhtYvwgh0q1a+PJoc5jFq1EXsUisXxKcGGXQ169HXV0+kq0qMNHtfoPFL46Cyrb20HnvhciqLXnB
MQflWciCqR3GLE8M7Kdbf0ccBo9dXhVGA7E2cO0So7mmiMGASJIKyzGj5mqKgFLjT8gEI8C+XSC9
5i+vMMFGDZMNNPDB2vyLp0x+LTzGUczH+nM0BcA/vnqUV2m06Fhl7YsXOYea5FBFbHXQv2xRixxT
mFyF27wZRrAS9x/0snGwW7ZorRcSUfnO8QwwzUJ6V02IHCJ05LA+ZqNNrcI9GJhJ1kMn/blLHgoB
7cZdEQfG1S7v65lj/iqjGYRA4euOktneOgi8g0bYXNofU+wohGgXZFscmyEuIIYK3Kxjzoj6XC34
ovrgfeiyFrg71oQcB6P0/EpW1bzvISuuipn5pizXPQomlHuZp5fscsaJ+LHkJFJ/2A3ca119rVWw
8TExHN1HDoYWHszaSLvrnjCze7b7ChGS5G5vOwgATZzrK+1xwDHNmjy94FTqWxTaS7900QJKa1SZ
lpVsuw8NYzMgOy+4bA4dVt1RMohzeuWor+L5ErUWb1SO7VEH1f9Wy16yIhuKI9vbOmk4yT8DvaNO
O8xWMR23LKhMBI2N6OKHOcbLPe5turgI2VEHKsNwhenKrIsDcTqg1qnxG/Xd91hgsz7uqhLQwzTB
Y8towFMW2k+hifvBJXohhGtI3jkTcmgTVvt9LGXPaQuooNvdtiH0s7YWWRNeJjqNuMAHZB1ZJt+v
dog2fotKy1vhTZsBW4QvF+R87AXT5rxOw/BDiygZgocBQ1bvcxf5ZigNlXC4BImzmeqR9EnCFoav
bUvAnuz3bSDbIz4TIg7BXW1UU6v5uaxCElfglS9CbSNfF2oO78GXDTTlpKgHaAYfXjcc+1/5Uj6o
jKkU2uEiKzmlQubJ2ht/J/sLIYXjWa12CYswnKp5nzrnmU9LQYEwZoTsBKBpoMsKGfD+Ht2fRdcG
PH4evtBKVvOp82q4S3NqF/DRRQz9d1YvEGOOQ9GpcW7Vty+y+a48yMY6LvM2cdEvda67NnXqROeK
MyemEMyMFmM7WL5Dk4UewTVn20D9eh8cMHh76h5LNErhw74F4hHe9IherYPTEURhXZKkcb2ek57M
9smpVynoMTbvxmwAY1s8mwX/6ef9s+fIahv0oyTgbOImLOsIqyiobOv3U+IL2iAw7+/xVY+5VhPc
InqNwbe0v/NOJe2JQfa40JObTP0J23hd9k2Mx21MJqWllfYSQK259mjGjdG8kjS2YeYt4fu7wq9+
hgLRQYKAnmLIBMksP1IoI20iKMDLtDWqS4oyh3NSbO9skMy10QtDngciA8iTLoiUUdFTeevMnTcK
d8hY7Z2d2ScNi60PYIzuBcJzshSBv5XAuQ0vR5s0/wTH9ZR0HDSLU8zMfC5lhqi1jFxmBPTs4IxR
VklvkOQks8x5myqukj8izuBOjPv3s8QHluPYGQUhG/rTz/ZOeDAJeIUHFV1r/HAkyAcuOEuSDGmw
4RZBFmvhXXp9LLjTZIHxwXUQh5GOXl7m2pEjFMf7ONA5IxpAq6O5mHyHAOUbNv/6Jk1Kyni+In3/
vMp8sH3H+mLdhmhFSrY2cOxOqMAJRqbrUs7YRsjWNBKc5ReXL2UM5TeXKfxnDUnwOYLpmPGhU8BX
smEggk3sv1ccq0dZXKGvaHznXwoJPH0+L0XW8ITOyCN474F7g2oQTIqLxMKjQcj5OXJ+iHCw6Nxl
rzFCHx7Uasp0kjJaRVEWpC5hHmH2SrYfED52b4gUDOOCD9yhSmxpwQzvQiwFzsLynK1RIPRhCi/Z
4KItMcEshXX06BRUhIyjmYuzBXfB3Di7R5/2bI5owFKfrrcv00zErMj27WDpPUy7ZpIV2vVeK8WI
fjoEMeZRLs7097OWHWPmN1JVlGRI2oTbH6RnOpg1ddpUwsDWxPWLTKxgU7OYC4illShqZEAy3dCk
SVpTCBg6Ps0vgSA0EW41TpA+1g4H9kc1v2+KaxaAmzWy7muqTFz14XeJCLUX0gvAOCbsOX/Czpao
AU324QQWF+jVe8t2/X2wrIAi9SJJeDajom/6/M29ByfFH8eLUgDaaRbFOO9fGsZjUANHvtDBspK8
RX+lQM2PyLJVCB1+WwEDnmsEGXXfcWtN4W09ou8i0BU/JchwJ8skTHbTlEQotUl3pUdVRV6Bec1E
sxnVq9Yap0d5DAGQIB9s0wJUii7bqFX0JT10lYqYc38PSoMNdh376lLtwYXWGJZu9K/N3Q/JfP8v
8tXPJlZjhMOm/t/5lwCb/DVK8mgDNnAju/ywYRxoCFnO3g5DaUHtH+ZWimE/gNwd1Mnj5cB7lvrH
/ROHzRhd/otDyA5yY8BpHA8iQ8UcU693FRofAKTMJY0jjzK++HhGdOzhGB1HOS+S2w0hMyt7wVA2
2MP+oTAbePUOJgKIUB7QNidHoPwwpicgln9jOmUfK/5Lg5Y+mVARB+1DSmrEbA5VDw8PLmMVkuhr
BV8hPK6RUJmcNZdUIp+ACgnZxZK7T+gOgYABZ6KSk0/bPvMeI4EbMkNUj5BxZxXNsnF3K569ZdNI
f2D7cFHVqj5Czh+NOUmiWu/dy+t6jC2pNDaeznTuOj1W/TMfNBILW2lTSgokXdBLT9s2TDPz3382
0HIzJi7FSlrOww57N7YDA7eL/ezNUx5AsNri1lSDeLC0yFe+55xX0HElmoe2p4sICREyY05aAzKn
QqFWMxmk6159iP8zHogSrE4CkMRqeDEaD6INoLN/OKXgHJmStUP5EXYAb6QaZOlTWnDHiiFh1xpx
XVma794J8CAxdC24/F30D9Zj2zF0L62jGHqt4FAK3HUsBe40Ziboc6+Ieji910VYfGtPLKKBiLB1
Ab/F2oyprSOHRgNzHJvcJaU/R09tltF/QaLpv1aQYNUiN5TNM0axt3RNUucrcoq+UYq8LDtbvF/n
5ad3MdMN4dycmc8nHw2E/M3RiRKkPG0qQGOuQvLCxHys6fzVifuHnaJXmJ5QtwKtRcBmnRo7EcM1
+1BBNT8rY1sEotyftqC2XrHUKSuN1+SOJEWZA3KrkjN5FRBBYWCNRn+WruWRj4g1+vtFYVeKmMCV
faumUbelXWCzQYuGCPhHEq0njM3TX9G0GiGJI9Ci7fOovN2cnN40OTjDP35gKltSTKV5crGc8G66
iLj9d+4wuBj7oeVl7P8QQTLElLUPNGRX9cdDV399tO7pRaIm0m9scwXk1UpfmjIpWdtGLO01Frp9
Nx8xWFoBBM4tWRDEfRrt54EZ/+nuUFx8wOQqaGFrFX0dfw/krTsz9I21U8+auf+lUtIps2C10jA1
0plZVrGsiCjChKxsQG6FQoW2oIYEKdpepDl+cXlcgOStsGLWHL6fVcnJMM0WNHH8uqkC4muzpod5
clDNrlR03Vu33mz046uku+j9r2Yk2Eg6sj2Sb73jX2qJpD3fK1uvZQzl4H9KkYcXiJysOe0UARgB
Qs7CvYAw5l2UIPPTr3TOzR1PIQYvACc/0ZcP30dqj7WQUHALiIGI6cXyMHL7rw14x0gkBytoXvZz
r3na0ePdwclyIYcxNJxmM1IMQvAdni7w8zjjFyAsS8SKRmTIR8tGXiqYijMtZLEN0pIcm5U5iosA
mJql/Z94eRvVUINvXdpizjkd7aMBVGZuEJWJ+8/NWNOKf9qVByOonkJ0YlSQWw6vESyk1E7LF0AR
UrnaGECmzfNbB39bgi6DqI0EyE3i0W+w5dRNKTehUR7khM3oLCH+Fpr2NFm+CRI1EpQNvZTZayul
bb7UW2mYmi18OiZDinOqsNsRK5aYIH38a6TSLnCB8qqQiAgsFDBu94NuY/KMYyGgZrbvyjjqnWyr
YxenZvB8PeSMY2RHpMO7zXLIdCyXqPh3mCgJdFMVClWT52ce0/ayRLL9pPwBueN86Yc44Jyk6Obx
8I4aQiny0UD+3W93tKfWZ/8BrUfyRTHEHKich++fD0RFQ6FpxN3IAcT13s2f/9B3y5QR0hkG5hgw
LlOKolmaL4lz4fFPl9aPvuB7KZlQD01ywkCN/OVWYFF7tjVkgBgP0vjSp5SYk37sLAzv48YiHDPZ
IB7mWPCvJtyFXONBrPLKnFG/cQFk7hjxCczgXPiQ7VTtHsBY1G4S5O0agh7NMcQrLYQCaA92dQIk
NWd6nyjeAdWMnilWLNcokIT7pOPUTJoszVPqN0+J9hvFI66dv+QM6l/mNj/9gveCOJBKyyqQdJ10
0k4eRBeyS+simXkSBc/PLtJwVtKNjhtoFi6QPOYx6TF9IEGqL8OW83WaQJb6NvfRfYL0a1sK5kyg
An6oThokUGXzs0Nd+dbQPI4LnjhirUH0WFzyfAtUamku720FU31vhDvJ9fc5ZAS20fiB0rGO2I6P
q2CRr5SbgogcL9xeGciW+deQ/GFPfouD224EAa58chgGUSrtMJpLvPx385abe6z/1a9hpafxB/Ug
QiMLnY4X3JHQSWtXzdeLmjQxSG1+tHZfjWJSSkZ+w+2O7MN1jwIHbS/Ij2xbsEkI9FQYxPLRmIYI
5YLiQyXmkNrln8qCeV7rKAkZuM6zNMRG8CiXXqUcNlUlgVPHgmBaHo496MrGMcNEPKtXVYiw7qnj
HQniVR7uoHLm0jIHMYbfnB18Tods2S0mXYNr4AX8+kWSVCGAYe8KyF2/d820zPZ66O/8ve29MAGA
0A6+8Osb8KPXs5eZMYZnViu4oFlB5EndwtH3XJ9BYSObrmHHTJup04JLDsLmX87ZdjX6F403q6Xu
YfqAcJCBZWw7hPRAhJFg+0KB3OyeP7LuvS3Pp+j3oyW1Q8ZSAFaDecOg8wZ+kbQfAK7p6hyUVnhV
AcemvNlk+VtfNhpL9Ybgdew+8BtH4G6lfQ1nMkJU1yCEgavxvTkBT5F3IqeRI7uPNq6rQxx5XIIP
m6UdYZR6F5IzzZP9ON87oqLhuyvfYBFQ+qcWOhn8tmIQ+Z1WCshQPIL/lBXyuBCsTUpf1w5TiYZM
kvj7f+hugT7xY61PFDKWVVLI6q51TM0C1raNn7yerkzUM1jHkGxf3i8cUXQKdK45mTfHqF9ljBes
Kk5DTaA9rpYB94kNRn9Uuztrg8fxZIXrlk2jMozrYKTn1W33vlV+6NWEbnFUGyLHBHCqK5XaS+6i
kKDARptSFBoJGogvlGaRR3TprHA2RCAyEFJwpt6fPPaJXBZKv320cMPD+dg42Dd5Mzhyq7axHIZE
L19YXFepxYeZVLlYlGoGtUZD1UI5WD8s+vLWNQx7gfBbsSapiehL2P8h19RkQjghEdJidUI0n12z
xT7wigPLSbUGJKGeXn64rM+RoOfH3htAXOC1qpdXpWIeMEn2KbhkkBswnTXlLdZ7vFfreT0EegQE
FfrpeIZ13a0Ajnb/mSOk7ax25u74k4+W4uJnncPLAiRcWZKmmC6UMJXxaaNledYxnp/t5TlYxVPl
PkuJLGQvva2wwrtdv3XLlSf8UUCJYFTcfkr4qanaUTNwfmnAvz3LFgNTmhrzdhOAGySWCPdOsj53
AY0DjUwcP+tfPAu5FyW6fbjTXhMnkdD8NcO3RFKuqNG4Xu9J9NXPw43IcwcZrusAURBV4DTJKA92
M25WMgJfNgDgCelDyiUUh6wRTHyWXySOkTv5t4TYq6r1xUCZjKXvbusUJDkUVYGHjjl48/ADySaU
qlOUy9ZcVFN90UDdGnca4M3GXjUqc5D1dFYwzJ2flg9M3FLPDZZ49wjYPH7qg/E1C9CN1a/4tRVg
7ozYmQKpFdkpHNq5EK/jDLEcfb5ZrhyTYZlngywOSOPIRChqFfx50iMM+vLprVHgCuZfeTCVcViR
L73e7NVEm6OpMIQ5bQR5vC/66u8iVTJbWS8ELw/SQBu0uyqneX6dNCt0HdVyvC1J89+mKeYPKXaC
E5uBdqfHeI+zJcvRI/KXa9Vymjm66kUrFjvvxdwb7PKCNgLYl5nutOFi8rr6s8Y70Y5aDryfKBTL
zJY90w27hamc7i4S3A136RbB1doJIxCCq8FMZW7p5A2/RttH1uPa1BQW0e/kGd0KLC/QzJpJJlrT
jkZqz2PlxZDEPUlv1AlaJCkb5bqNsBCgZKN68N2lsOMANjNNzL5j6B4eQIjy4fif+FMy/ASGF8pA
K2yA45hO3HK5r21FJJbBLydYw4p9BU4Q8Et9tmjVZpYGmYkmL63VO+PkVrcqFD5Q8uOsY/gZ0HXp
0nppVmJc4Rb0eoJlAAVPTmVQSXd/koYl+UZjEtSbHeR2Vil+XTKt4z/P+Mw8ppuU0s+thwoWTjZy
mr/E2X1qnJhS6sUjTmV9eOs8wN7KHTwWDbsj8kOMac0CtArGPiJq1FRYetQzFFNEFRyPbMSmAEV3
qYhNeWoMZJp4DmInIizxu24kltWiNkEnPIjv3DTgrFn8wg3LglVrrRrwM4Aa9Zv4nmcrZYoZPUf2
fGcw4mw79fBZTI5xQ+XJFFtBUKifeYPHfczPJ/FsQZH11afMLUqJVT//R6oUoOQ0xJzrUfZhY+Jb
R9gtc7tR2fAlaiKi98AuwYFDGbzCyz11BV1d8g0T0jlt7gl6ldChJld8sQASccUmYn3UBR8c+kCy
JLCm5pu2hA6OiIzR8AzHQ/NaddYjpCxI8H4v4EE9dzWOrBbg1SaOw5vIH8ERxAipVFfWJU+0F3Y2
sW8MbQoAP9Z53s4lUTnalUIxmTBqQpWf5/TJHzmNCPjkGihJ2FZ3QsQu+RlS3l8QoltjlL2MoWfW
njbd6pfebhaO76pyhvWrxNPnBObaVxkm9qMgMjXJD/oJFe0Y0whQLmzo/AxxO9jE+Y1Hn5pW24CM
y4NX+u9SD0zlXX2Ty+Es7JgAGj/guIcO8Z0PsPTV1k6sQCa/CEpXVtG5jaNcSPEX8I48XSClg1kz
eljJqRoWXYWszXuj5pRbMrmudYmsZZdu9dDSxo0JvLQekon0XhgtxCU+0lys1E/FmXJET9VOFbru
qZLSoz3KeKx6GlJw2pFE1sJ4hCMENfjJvv03T70Ur3NHaBs1ZnmBYSmWhG2ri9ozRRaOxzDT2idi
YyvKcWr4TgAIn+tkNsSyeJtf4fpj5uqvV6JuEwR2os0au170pb0PQonEjIqnPlMyR7oev7C8qHT5
arQuJnmGSSlwZRsSg6EpESWTrfllH1R1cYtRGLzj6TmFlgmGeSF7Buh6qjIL3vKvQsKHucD7dMD3
+HZoc9mem7QnKZd5TB1tgvCRr6YWlRTCcW2hsWSfgNL4ImUhkKFCJ1lYdyw3o2HCW9IihjFB5vB7
dpMTl4t2VNkFntY6NrGzsFz5owXq3JrSrfAOGQ8u+N7v4ogtNNVVpYA1qNprAVgQNU7w6zFyna2P
1jE/6LzTuNPsYQXF0vbyEIlZKYG4EFWNd7fuGK1HPS5sSUC7DLYzUYNxLUZuTECIixCn84H5F4Kr
DNMttbvwiMzDAjs9ch4luyJ4BRpJy87R9yRjiIGgIaPAA+mYjjgqiE+7A13LVzE+dc10q2UIsdFj
B3sbW1ezYMp4tYXJtkl7FwLTrR48/rR0JAytmnjieYXMXxJ53LkGQwz9NQRzaaOy+Altod7tRtjJ
HpxyPnewvSObVe3CJm1C03GPAiag/5KWX8tUPaqHuGZxC6GU5IZYLPbBhm3YKOjOeVCZJfTiPu82
gVzdDFRKuQOm0Wn+VkTQXI0Ak1d5GN6xU7J8K6dudmnjUdUDD1GEmsZINaTqj4JUN2g0j1wyQhjN
O6VaXng1IPoXsjiBL9hnagbyWyQKPc6LwvOLZLcCMWGiS5P0hzXpRr445p1AftlyF+X75Bnl7ndt
bF0mv391hxK4UsSakZuOkokAJ2KKunBonLowNsYn52ZDKNpELYIFr7wxHYUWFLs3rKE/CbxzUHMw
3R2nuk+kN0thHSUS7t06OxA/v+1e/wHHYoRIFkSVzdTWGRQfjl13cBgOR8cdzRJeyhMC3/EXyNcQ
OfzAfjqFEkgSAI5JzF5QAHMfFb/wUfi4M/k04GqZljfE11NoSEVTj1UgNcfcRgIZQbE2WNmcrO+1
HJeJ9IuZKaq0xitEwGhV1syHVG3tH3vGymJMQV6zNzTf0JUblAaC3bPKCsUJtEZSNGdKvC1IYS5w
tpIMy7B66rhuPJYnw9UNVxbrID3G4n4GKFrkjeMkCJLZMkOEH9X4ddZaa6x+UG9EWJUmDKs9jAjr
SZCcTDGWd+4GTyCOogoVZ1sBTYR5xq+OCDog93+lDFzOTO8MzEFi0GC8M9sa0yP30BVTGkzEGYMT
KAOGJ5LOL34oBpA7Ewp5Bku52KahIagmHkCYl2uVWg+lIdRyTB6vulc8guH1ss9FQQdhRQJl1p4P
0YguTJy5LrdMRgm8iT9tUaBSwOI82KbtHXpZnNle307NfH8uOCgD/FdJG//COFbdWFCZVEmW3DzZ
FB9vSPF5dfoZyM/FZcX3NfdYi840vP7Zl/JDq2Gx6HR/8irAKLj5R4VV2M2p0on0s0VtoZy5VRas
MKdYzmJP24m9PpulxgHJJZ2IKfIps1nxTZ7in5OZ0dN0fQ/XPdtMlS8qTrYbmGt9hT2l8hJdpt84
CV+r7wqSwjvVqhv2vv3BcQHlMD1QNipxeglHUrt5PmK4MhEdU1ROcrTyIMzk1Oh3j5z7Vfhs+Hui
Tsay08KdrsZO/mzaK7OVzzy72zGHsKwgIcZh7UMN8prKz+8rAIVc88rRaGnthb5Nyz2s2nSkwzKt
O5/IDGlEeGKY9PHRq6+WIpBwXm00G9St8T0DilFJpTIua5q8nOWeJuaEu8SLZqge7PSqf+XUVw5r
BCtuK7z6DPLJ9FIj35LUy27FsLForHWi27nEnn4qlFtX+Xml9V+WPnV6dpqNQrqwMUG1fwNbw/wc
OwbJTGHOd7ZdMKqA5V7wNqB94gX9Oo5YdaVG34fe2R1as2NE7PLbHQa0QW+WwILIUPMHy6kCtzmc
Gzw17KwCrBKdR0ne45Vdn5+S/sSpfI9vlKc1K1q9o+Ha+WaX8+4337yMvsRuFky40XITLNWaqwGK
NZxBOzXbQygiYvTt2JcYTP4E0U6R84xUAuFxXsdcSOJ2IWMLYcBPsXZaXtD6p+FOdc2kukDWM2dS
K3l8DQ6E/LG9TNcK+whjW3vjLD3+HY/V8I7vNpQpOH0Iv4bqkP07oE+YjCBAOUXbhz+8YWN7DWm2
zX7iPAu5eSRIZxSi2PYocHdE+8TnReYoIflnGgs4SthuwoROkY4tOMkvE7yYvybjdlz24Iov3Lxx
RljEeTJhYazFRLCJL0gS2fDh2CBJCpW8x456OWO757lYFrdl+UZW2TL8FgjE8+S09wlSSlt4z5J8
osKtB/1Zlr8qylkeqRqYgxrRSQn91Wnydey4/BhgJi/mnVrjhAdUrhn9QEhxPmSYCLVFMCumr51j
eAipYVDcF79QDIpxSfp6fcpbv4MjW0vL8rP6irF2yCQKpo31ZVzTQop61ZM35J6y2YdnYqX4UAwy
hheSXBDz4NqVbswcooyKY/LCh0pSBuj0XDlolvvM8C6G2wi0dmDXK2UW8Cpf+9wJQ4LgPexn9Ec/
g/y3C0BFtEJqjR0x5aRkkyWIuztpjU0ij5EpO/0QwhR6IJuUxs+tehYklwEk5T7Tlh0Fq/qNQlBj
G0flkMrUjlCqtk9Ego74tidyt++doh32ADemDGxaGkYdy36npSisIdYKAH395265EyiArSmjxU8Z
vAvyYbZWTWzYr0RGBVIOsfCF9VprHKfe1cI1H/AKxxQ1mk4ZHPBHxcZXMfS1DZFl075dlwMMeRoz
GcDGVxbbjcDjQGPb7AU4ort89PNgwS7wJ2wp2EfT6sa7xaAcEhKiYOUqs2/Wc8gCEsZ+x2L4ZxuT
hiAzPlZfzJjkqnGaEjY65FjncA4W0OtW4sxNolYKm1QqwTyMAky0xTqKYKaH3oB89KUilOV2gMRU
I0319xgIwP3CCJrAfjJWGqrp17h6+oa9dPCzUczXzZP4VSnjwHaZeahQO9hq5IQg3ZfIiXr+ri9z
SUz4Nij64FdnacP5489TlXHAEPoQkMihYSzY6FDmL3P761DIRPHPrzsaiM4YA67pZe65OY+2Ffep
h0tlfGZUgcNhRLC066/WBrmyYAtCRTpidS6g7GQvu0J67lpVhEr8gyfmhHEPkGMca2i8CDtYr4Pb
oUQ0O8uttH/qbYpoN5yqhrIG2VZwa6VrKvWPU+UaoUKEHzDVWmvntIYPxw1ov4frKqOmQxvJyZ4N
mCmMb0QXhUuCaVRDUhu/Zpt+vfPqy4PbqSbj4ubfbY+9silJUaZyUW0e7KWFxFOR0MI7oNLPtyfR
Jd/2w3encLoOy0zfmA0ihHu/6PCkVyIBUqjBU9GXpX6P5AXaTm+rdyUbvvYz6AisPOAZrilWBFu4
+Tg6AlFhDVElBa99s3JrQu3Wb1Vzbj89W8613SVM7fq4uVNWdKA7zA9iVvtzeZNiUJZCf/5cSM3+
lqhXGK6LbGcIGi3UB38zYXY4lxBRSaTEcPtBhIhPdnFj6aSkMOUFlQX+PYuEACvwg/DK9+Yhvyjm
nZO14FzPSGU+Tbko+qe87c4kROolOZpLzIeXR1rT4yddaX1+9LXvU/0cDz854vTFWQbvLWUlFTvV
+tXJI23EXUygxHa0E+pC1dQRaHTSavBMsL5LOHeMZTWRNkgIJpZCxXWEQcLt6wAqm2dtapQ/yX94
Ny/B87yeczQELYsWiSV8kIod8E8EmKC+M3FoNjSyP2qDmjWNt9iTrOOlGJp0teFT/MmpQ2bgoNY/
jro4RSkrLOyARrz0ZREALL11qtlbmgYq2Opmg822Xbx3+I4bd3rfK/uMKbVvz5YS6DUmLlYoUMe8
SDuvks8bPxpHbJq8CockRl90pSU6VKU7fim0cluscX7HHG4ZMtSw/bNEGXiGGoZ1QL4o4rcdWWbY
eXrq8ZPJUjiVz4y5s8+tM+9DUw0aK+S+9OCboK4WWP+OJelurk0yVW6fxyHlfjCEiTdvzLuSDzIG
rYdnMZkP0JmP5DkAImJa/4oVWFnBVEvD068Z/ap4FtPv+VYVJQdJj8R4lHfDi4UL6xM1a1R/FgB7
XcPScRhhJ6P0nj1DctupTVKpjfWY0jXueTQfZ4TFqsFPC7HoT2GiOK30MLI3U9EIPalZi8HxazNK
JpNZIjHGPrj4tT0wNZT95ibuhOM2W8zvpofUxFDm2Qp4/yBoTS3D7jKxmR6GofH2TYRFv5NZFBuP
tj9jB+C3VlpaUlcrdK9QIO2hrSmqyjYFggsID6qNDxCCghQp9rjOvStDCWRwjNEbtTlMclRvdm7F
dYfk5ahhWC30aNjFO78LxIzlvuQYLg2lmQInQNJy9Y4cbEHzHjWSZalUpM/4NlXeeVkwGl+fw3km
Ld150ayApt9xx46sDN9gocZ0U3vxkdi6xDSKLLM165tm+A3MAAM2F4IKYehB4Cx4sIQpsGbJ3+db
GbmJr7z7VShRRM0+ixqWZNiurHGoidQbSj0VbC4FsZNCy7/iZORo5X6FhMa5J+f/XKqEp+oYN4T/
c+pLQoJKKOum0PLxNQtmOo/PZpjenfKkpdyPnPfUHJ1I+U5YyR13JD2D2A0mcAnBEDuHMEX50XjQ
KpxejgS7dXuLsXmtUgrn8J8vM2BoBhyPvJ/i+uIkm+CLvZ1Vl5f2H/rn5fpOdQw4tRyuIWpGTKyM
/F+joCa7RiXXCqPfZdoTxlphHQk34KJ1cU/Z6VAyPKr86VlFvFcAVzf2CM3fqgQaD2o2RDBO/ks6
Xkpo80T+5a6+Yi1BIlw/HsTL6o3qr2nyHBwxviUzWrvFs+hTe6b56BCUAFbma13FMZeaWCMFBQJD
1SVS2LSwASQQh+PdMkB6L6YnRIKSmhplWyLLnfOezSOu5FFEs6ch2g7oRfFmdTAMbimsz136wTtU
CbCLzyPfnw/lMGD+zasmWQiul730IGo0RwzZTElA4tlJEZXtKiACL5az/ui/fqCSBMaYo0V9Jhsz
wR2oa8cN8fa2mclwu924ZNf0/9XXCK2OjcUKl4clUkW0nMZ1nW60nLN+VGPztzwbpCets8kkR72Z
EUNv7G/nmReQnJsbzmMwk7SZdScB4kIKBBk9zyVK7zFLYXsqrOovNtCjUp0B3ShIqnwXJ+7TcVM2
/8bAzUWS2Jn959Sayndk+VERBDA6t+N/Adk0hTlOl6yEkjgRVreStPlRNeLgqSWFOtgArbyrdgfy
ITSh7IXXni3CdCzwEZE0Ck7eAnBVzDu9cIjBhX/9OAyWtMjlLwGnTvgt5UJUfOIgwrQ5107WfHM/
N7LSp5xaptKcvh1I46XueXZARJ0jUoRcjDUknjPJB3DlaFLgg+CFf6LMjMh8q7HC4Std2GqlNWaM
tM5UxBNQfOL8r+NNoLN4k4i37623uXVRT5l3eODspRULk8JT4oXHvhqnN6lp/4JXnLNCJsMTgM4m
JeSV5DxPLO28cxRZLgZrQEh5SIaQbNcHvRDXiPUQ0Wch3as6jIRkOit3taA3APx7AU1dFD528G3K
+4tSVWJ+Unpa+rj8l1UDneBQGZGnVh67fSkHs4iLbicrIadrmIySEl5xJRZZDy+6HYANaGkOz7NM
a/BoHpETNIwwNNyBEO/0FJzb6lsokoNc13io+j4Nt/xZpLrGJKtbcXFRgcZL+7hA9LUC4tbe7Kk+
Tc2pu7FNf5WJNMjkcgJUWWR3mdq/dixl5kS/wM7i6brfsHYFEHlAJMxbuFlrfE8tgcnK9DUHZqrL
zMJRzL6JKdCEy4GT9XA502OtrIM6a3AFk2fqkR2E9Unvyn2SvfTk3etwdZWtw0oCmdf3XVB/uW+j
jHG+qJ3Wd8LxZqIjFQjZcD08gkzLpX9GJLBU2fDDKPJcqSQve9BXfgdtfinp5Cvjf5fWT48OUe+8
PFB2OFM8NBqAwPpXBCfK45lvmuxuhn6rva5lf4Bgk00/HAZPGXPeq9C2mSjihzSLO+9CGnbI6Nkp
TPK2GOrago2+O/uR+jzwQXol125peTvJGYjH6SKvmYcKe45q/2ZpqmV1vpppsQ+PWc/OZFF3Pdob
jEJKEzTK936kFq4TA4HSt/TdsoYPf/SqyoqPUEVo3l3BDCvIdGgAr99JAqohmswrDHC3kzHbHBUe
cXJpJa7pSkrjbpoQFTb4iCqHzfgYzSOeVwjgFp33OeKf/UuHzosLrtrYlzU4vJZuV0gOSObTCjw9
uUU4EbTuVCo9mNYUiCx1Ex71da6v4M2cjba7CZOpaIHw+z04ivIHixRG442cZs+B/aiNmPIkYx/C
seH+0rVhHLt76v71faDBZ+6jx/NSb1M//znCug43X3iXyBm1njC2Scbbw1FOGH2D74pZax6mCRtd
W2VxtewevE2aQ7tRkyNU3JJCu/EnTVuyYLgDe0AW7b0HxO8YCwSlOfBe5+6lDIwr/uQOd1JhcBCj
kuH2LuZ5xqHjPIxNUlNKFIrpSQr+OW61DDSCjUattLM6ECoHN20OZq966XqrLnTdjRqpWFaexyNP
LRCpDa3WCxRZpqt4rex9gQUShNgVkKQLC0rmTCzBe5SRM2eIbOAxQgQvZPVjDdZW592OT1N9uIpa
+pJuT4IXTsXWhrrN57iWbT0rqG+vlxRDw4JIUED8QESHKdTRhIrWD8Q7NozLLq8NCrbkVoOYHp0b
GBVTMBTyQ48tZAOWMRR7qTb2bpEKPhV09SZGh/o9BLBkL4ZT16xmK0gB7OlUQjJaFJSNCoH1ICxR
clSQ33MwO9C18zyji+54dx8qKlL4jE3kzV5nF8kLfLcAzcMOt5/UoIc3Ik5J0lF2RZP7+4kCpIQt
9MR0D7l/Jk/GLUq+245wFpXGY1cUn4KAqSMDMn0NAX08kJf9zgz9XDEqroWjBIDULgXAU3XhRHJR
WKq1E42OzYCEhwz9LEVFhk1xFa/BGqnXL2X4O9uC7B/sPiuL6UZAXssd8XYwOZFt6ljEKLmwXGzY
vQjPedMsavUWbPGx5fHhnry1Klva8qBFw2+sox4nnCTsRFBuLHDQkzhTAaWwACuiV7O7+YQDF3gA
3oegt33yuT+xx5NtoTCMDOr/bap9TeQqu5pabDaY5TeeoKgrEHLtujWcJFQg9y/ZkJ8CsCWZIDTK
s1z/Lh23BNbP2+bYAn6ZvwCDWoHheXVfMhbyvHymCC23yeLWAqZpii0/DJFO4zYuoooE0IYOw7ip
b5t0oqrPbQDOyE9yr/8+hGewHWEDER9bCBcwVdp7XSyH8M2FWhYIlV/z8mYBBa+lMnHQZYtsdNOR
q/Rmh+RzwZj2yuP0hwt8H3UvIHw2r97Wa1YdJuBLvWBsU9B2/par1nCLJqH4lrQ3ms16502Snr4x
60Y0PV74+pZ6eOZqCBFK4cpStq1bqHk31rGV+AdheO6a8NkKA8tvFQ7RhYc30GD+0z46V+5hvHGn
sfIT9rnu8Tqz8DR4qwIxdvAqWpuJmkTBvC+7M0zucttvO/i/sPgoc8ZCNrUMq+CbTVV5BkaJCVdi
bMbABFnjdbISVTfb4KrIFw3SlKNOHOUE5xU9pIMRCJ8oJg5xBODoRB+slACeSR84VT+ARfc41xVZ
hfdnzJseFgFBP3xL7elmMoXzSOnNh2byPbyezSdJlyomtd2CknMkmEh9RUOX1CT1oYxeATn/wkRR
Tp3tGPUdSre6nTmTP4KAmClx/Mv9vBYo7ho72z2HoWTVzWB2iwOSW8WTXJ2y/hSlQQVj+E+AW7YY
ETuaWhxQX7yDqmzLZFIMmrT0H+qvGa6oLGTgruwLIN8NRQzg0WWJ1alYlbxnM+n2lQ+RKzaR5I85
jpDvpBNNAHu00Vw6Y9XsKwfJH/Is6RUIQOC0rwXyIhH1TCQMrHfoHDCiJzKpi3/26eRyNmVSOUN8
ZwJs5BdbClZEW2AG6L9lx7L1q9HOINppgHyq5b2IVGScZAZOaJXzNa07e1DVvYmfZ9oH3Vtae2hp
7CTVi/tc/ROVBhvsGcP/ZG8Px/LC8UzUMHAOZLBrS1R25Ft+R4NIOWodj0ch+FvRv4yVrv+YOVhP
yjyrTP/EFcHcvYq6kdyyP9+7lTPLM7khjwBkkGzN18MTzoe8YffKU9svxhumItfnZB8SksqzJR5T
Hz8ayBMa7D78sz3IrR5xVO7SYOvmTicbuEKvW6MTSNKI5k80Ypy2JAhHamnXRbR9TarqMz8Zxr48
K5R0aDLlUC2dNONMF0zL5dHx9uzZkttIPaBLHfK5l2X+ITCgiW4zzrRSVVDIjUpAIvgW/k0r7lj1
fV79xsBmkYyO/TzAKW3yKaQcuOYM4AAaNus+khdQWtD4Is/qO623z7s6LsDnca6lzvvPuWHgDWw6
nu2wWC2Btw8YHk+oI1KfVFaQRDsnQpGZa/2DJCBWvUexSuk8vEpCjxs5Uct2z9PgQTTwucI/O06v
9OAjuvwdTAu2clqgEV76ki5JHLBmbROjcKAB76IpZ8dph514SaeeIEvxTRqkw771NJV+9lJWBs1V
D3b/fRR/YKd/GebV++bHbQl8gmykKjtYzjaK0m1DO0pbbkuuo6A3BBexQ47EhUka9Wij6DNSWUgL
3RITlgsj4ViHSrYfk5M63dFGqZYOwwFHkD+13HEHjIVtyXUL7oDYziwpek1r8s1tJYMltVNM4zjX
pe8XxyRXl6vgYtqPyi0VtamOpvheiU1tn3RERvxOF2opfqCAxgzmvcsMSVOYnfVl455gsAxFb6gu
VZUwt6PRyKFRc+7QSoZDTqqFgTWev+phwENJHAP0Kf7OI5jBBXK3p1zy2KehTm7s5te8QbbyAz9J
Y41Zfbj2YhPSKOIVl4uuiNg/ymJeLU2o4a69iWVpRTecQrjw0ngCyT32RSt8UV8Ir55XeNDxGaC3
ckheUiAW0dhlt9nH4Xf0eM7JLaTRaJIkfYVu2li4+Ww6vCPjZsOwC5xRMGar1WsbYT2Cjl4iAaUP
C1opBR2BP9tffIN9NYqUSBsJxLPWZ9wao+1AO54z5aqBsy91iiFkdCsh3Wc3VwQapWn9GHSwNghL
lZzE4S+OegBUavsmEilMq78AahleP8ZIdTdptug2gKmZlD86mHtCDRcaLlHzRIseyNg1An3RS7SX
mVuhd10uJB6GQS161xyp6H2nJZo3Hf8yQneWrmOxyB5ASotf3OFifZDndI7Gc2N1Dr0ihPbnTZLs
RdticAFaqy8e0T+BsFEffWwoHb8zvuMKZrdDHr+UEtQfRVYcEAp5AeQcgRG1cQ6v+LcK1q2Oca8t
EJiMqyUknTp1dg8VxNsfzjCrMmQ+jNjaNjQVR3tJjJdZa9U8UHnmc82D9ob9WBWYRI1+EpM9SQRD
HFzPQKQUchOafn9DbwDBQEfJD7EtZB6yypkbIi0TdNsjYF+ljjblmIhNWA4rsOkVDkZpvUav5AYt
+lxQH8wjFMIdEbCSmewGC/61gl29yOYFTdcmHAoyjx7AY41qPMYi0hBwOYzqaOOJd/W3hb1EGWMg
hEOXanpCqxdMJ2kjS4b2pB49CmujMhWy3r8/3HG1q32nOiFjG5UozBQNAa5En1s0c7BPXazqAOK0
G6jU3JygwOzvKKtbs68m5qH06EolTaR58lhc8wcufsRvarNanLbTpqMV9KPV/VbBcoiz9bkMCGce
VLjjavlFgkrp5jaD+ZCn/fTpxUGA7CJP9nRMhNJaXQgA7VFq9wdX6C46Kzpnup7n4jo3/lGCEiUk
rGoylg1o8Go4HfcslkViAy9PShzUBfyALx9jD3eombGf2UkqrnjqTL6eV1SL1GgY2XpbvZkgTFmk
OoxC7oQbK/9dkOEC/mQ0TEzQ0Sj3P2MA6mj/JxLZpLm9Ku5rCzH7y4WGIqAIxVs0I/PUlBc0VGTt
rU6NVLa61tpRBiWy/KLAPrF2JQ+PHrFk6Rk79jdl3ZpsHBgkO2Vrkb8WkUbZPQgHQEkuGdwOBw0j
n6CaitVSbA1/51JPFQGbua6/OjXqfGIS7VG1gOqbQBJltwp0KjARZ6DUzYjiXnnDyidwAdIAY+cg
HAWcIstoL4TQGzoMNhClGZOuQORabLnCfJ3TEcK+NyqHqOh5Ezst4npCEjOzA6F+pMegabMfA51o
xwGi6cZEywT47uiKb+L5TXaZnRHZJR0vL94cpsQHo9fidtf8ZQqPd+9H/xJmkvfYorYpH2+JgWkS
1F2VkkGifmQOq8NqB1cX/Y0pn7bEK7w8FOJdRrs6+HMVElVbPppEzxoPlhOUXTQV+N3nesiLa10t
G1S2fDOUOMTJ7zf21Do3Tzc1WjjCnxt/xI95UB2kRaAqg3WudLnxj9Os/skcgmpyquaZSwn42x8e
eKI8FtS7nmjAJ8w5hMbCHLdBsMOMwK2ZKsmJCtnPMTryOmi4G0yxo8CSwigV20XaPr0D7bO5v6X5
FJlQXPMMG8zHSYdq+3HY8V8yPSNCBuDvZI+2QoQLt7e3LIhaOMk0dUoJjKBa6dFAskjeVLfQq6Qg
z5Phn1y7uK8kE3lIptSRBN4quJCqNEVcN6YDLRDKw7DsziCoJZFMpHel8fwqRFucAW9ixhZhgvgn
S2awLn1u47E0eRTzoOgBaOoTE805zsUCalX0IzgxAl9M2JdYlD9CMJx0DC7valZOlLL6vHwK5Fc3
1oQxoGix3tdIIHVi4EGCbVlYADPQjz3qP9z6f384q4mhg/UrLKQNIMIZh3VpsvvJC3Kw2nz2GXTq
x71S8SbxdpGISoASMYb8B1z4Z4CUuez/nK7z4hd4UhjBYs5hrNIRSumAUMonwnMsgEwTGrf8BACd
JKX1qxGbNo+zUqORw9faFr8SkSgqGqlTucrmOjdIf86ez7j6wPGd+RWfAKyzwhKLEyZ26C9BT8YB
JIqKu6qCgecMKdSAJn7nooABTLWq4V+knWahalakMIb1ottTzaGkCA+ruXhUwn7KQlItqubuwkoo
G5aikbl+NhWO9hlqW6niPlnfAgln+VgvvfkLrkqGErZxBBVWF7EmkYTaVKZBwtUqnixJ/hzF5SCg
FEkFRxn8kbrWoQ6J4Vvok35mu7yc66AX0rfK+vb16cMivPQ6k4ut3LCYuKjDtJJ09yMNFybtSJ3g
fWvHFRz2PSTZ77zkHzZscM1oHzG0XB6hnIoRYgfjuI7zJOTUtb8N1iYtuvjlVXZf1bx70m4JJIkz
hi+n+H/GnCuneam/dYKWGiD+AnThf+pWB1CfwlliWzJFdPK/zxOM1AhRL8HXojbivfDX2MBAG4pm
xgV2ArBCKEeRzrV0TXRzGhT1IDiWGINv4GCNjBRk5/d/S76pNwS46ByCvHtgMHPJJALgUPwsfONy
ipPCN9iIVfZlsi5koTO3wcdan96KfDbN863GV3JVCfQ8eGWIXSiCnIVa0oNzYCEvL9W4V9NgdrV6
idXx1AAJ+c25rRJlXI1ziYXQjzgUtHg0+AMKxqJsojNuudcIPkEEB2vVA7xpK5Ek9WXsFtku4pxO
XNanpaeIh+CCBBXDTzzJUNN+5nLlv7WTW8JL465X+ntP0mgJz4o0+2lhRjb9MEU8HD/3crhUSoJI
6xueaEpEG0PTRbhNTXBXKDJrZLHe/hJurXZY3iufr3SjDd512rq4zg0I35rY96ytI743ZqNcozTz
fWCOuI+Z3eYonL3zSqRoB+YvfSx874fbZbKt1l6ITTVpZYX0mA1sWGtUeGfneGpt7FBZzlntHM3Y
sUbe5KVjMNedzLmwsyEx8T4L3Bf+1VAcdzbyBLWmbrXzwFnhKycMS561xKXVHGPqmbVBcAoZOJ+V
XHfJLZ02PmqEflSyhsQm4rl+dCl64zCzRnLoFxl6f18sXbl2rAH2zHJsgRmg0WbnLHwS9+7OQjVv
Zm37OCxNC7fdq7/mFN+1kqYkVB4XGp3O2OcR1LmdXpfharW7HHM3n8C85X9SxFu9seIIgwHewHmS
hWh9D+nmOzAPIDVUzGse7Mz+GdX0MsfdET6VUm56RYeMj5HjySmHL0MrNEHXJgWG8HxEW7KSLLwe
b0r3+pufmCfGjYz2IYsrAaIEAEZHFx8fB8QJ6/SJtrYzo0t4tRpGwWqZver//NlcLVkCR4/wSpHX
wYCkHsipAmavASYdmCDOUEXRuNXXldg9DJBvf1YtzEw1NXJrsXy8YWVige/EdovKlIN314n22BnN
w4uCpaGQsU8yisuL2Mwnt5aCmEhLpdbTFpyvtPoBe3wQOYPMqcToMa1wjf0Ge4+j8aqK6iqBC+XX
VQ9xDp6Q64AHHXFSlx9wx/4gsiVl4NW72JTitoiIdRcPyox06Rr2X0RpWaN1MdQZGW5c8ncJubdp
jXBxl9hnrSWj9BkfbcbHvos6SBFvuz8p4uWu5Lxy2cUrf/hELDDFQybLuiwtgXx/N8Mm+JFqn4AL
Gdjtgy+1I24tMdAm4+Mn/hy1iDbB6id2vKZWMpIKf1e+MPOBTMze6m4GJBAE1gi2grBE4qLZfxYX
3dUCNVdRLA6maeo4/3wxj/Vl59fuZt7qKttYfShdXbdBG4+SL9VdaQOmjOfzQ+UpEfpjlxc+XSlk
ofEvcCNAigZCB4iorvXBCB89KrxQAz2RjhFUBnGfQCp+WpqWhLMymt10LENMgx4zd+t2DRzndUUm
KxMg0N1gLUAhbMBLFDFZmkjvO8wSLHGvc0SkanEj1gRXWpPDH9RmfRl0nMvV1YmsveF6/aiifWzm
79LNxJoMtjNEt+aeqo81mZG9gZbNFhj6HEppRd1hgjHhmoj2XfT2y4fK+DFcwP/+matdEDv5QnY6
Nb4SUJfIafCyF/vYynQxcKFHslYzwZtiBVHUMnWHSCcp1yGpxNTa6R7dXqqVwk+xOQcOjJB9tvoh
ml15wrIun5oYnRQ+xxM23ZFfeBehN+UtrLUE4za1T+cH2EQ/pjerPodf674gY+HT+gdyUYP8x3Dn
pAbz+TO30zLs9Lnfuyo0S/z5VmkFSNoNV+64eNRzwjMdFi1UE14QdpGfsEcEDDnZncmByWoCOM0K
BMMiR6yr8QAtK067nyT4jGl+mqaMcK2K8xWotYoK9y+y03AdP6LCBSF+uA2UD55P/UfWikQR3QCs
s91RWglFweV4gB/7eLa3rjqusU2JxJg55lEoVXNEEG0/97CRpE4VxZ+Tue/SG/S4yqOGTMzf5Hna
QZ0vC2skjly6W50Xo4LKxiTuUHtFa0cxVSajkrkdc9bHoFVpkE8r2BbMPUDagAAnuOTbwTlaThoJ
ppGY0v9FdK1rnXKvG0fihTwQ4aMzzCb+b7Z5wa6rAYNS5KoKDGQGcE4Y+f7aErZITX4iUxqaY5dS
/mG6E6CLaHX+LJKQ69fkX7lJm0kH1KWS/vvyrvu8RLkKE2iUaB+6Vbsq9Z9jPTdQGa5lvF3scSr7
GBCQN1maJclB5ViNCC0ofFBhP3RvKJGjxnthvXrLfF9zoyQhWX8g8ljEOLl7cDflxsb8Gq36QQml
F3KZUHKlrJjGcuw2wJL32MXO/ZaxGrUjPYXj6Gm8Qx6jA9VBF1Kas3FG8noMHtxraT88OEqog2ZP
pIKxWuZqLe79l8RsR9x85TsVReyNhIJbvfukUkLPFylDD85AW4dvRy14p+x34ezJp/RoIjyHAa+7
IVhme32VA5DvNUQ+ezp4evRpt/ZxH2Ond3lsPWysk5NuKDT2QI7fBELOYsv56WazaTZ/ZbTJAJnG
R8hnb+q50foe/b1o1KZjMDD385ceL3V84AYPXPOmVG7/WtIfNkMdPzjJmCiIZkwjKLVNoIj8L0a5
2+7torV3DllYZuLD9eucOD9GEoZd9pizF33dFWEBXyvvT8kQ8gVpTkb3t90Ao94ciFUI0zofapgm
qXTM7G7u6Alf7wvFnDtNouBYnCdv2XVX1Q8Ei9qQTWoxgPgsQtNBF6yphjw4KFeThITmfG/5pjAq
3Ypso3JzUI8JBgalkIQ9jxD47EsJzBacF6lMn1Ee//rHFeBaEmKjqyYNbjojYPKM8QHN//EqsR+N
H/AKJS+PwsYn170bv19K7ZiMgsMOzZGTuMktQGnxrTqJsmbRCz94BCDRnTlFBx1Oc5EcZppT001y
W8r45tYlP1O6yqKbQmeQkJF5eoQ6fTlzMLyJ3rpcFk0yN+fHlOPnKXltPDgZJsrA8SkU593NLmLi
BbvUWXvJ4rEDH7o+02kG8eiUBZo8dZbllebcAiegNcacRrFUQSNyG90b0q8JZ1HLHp70d1dDCbeD
pNoYZN4oJN6dTY3JgGW/YsqRpkaMsg+knZX0gVMgQl70+y+kaY7F7ktbqtl3xxc49BfL65o0ZFPX
gOzGllBuF5NKhv2chBULJ3ce2cPlDWQeMWAFzkMBbjsKOQO8Dtkr5W58C6EoyzSO4NvgsCBVa1g5
mxJR7uB3ejF8SpA8ItUSdopovI5nLUqgf8v7jYY5F512voZfYB/8kvm9a1Grv4Lmhaf2VHGva2M7
km8Y2HLvMxli97+TgZQfCsPmaDOyNsULdSwc6u/D4UF5uhze9XKxchXPvaA3tTms2kUTGs4dtNAa
7g6mitkHeZVgqmM9INS3qLaiKuuuDcOXIBObtPi05Ni5lqfp64WQ/yr5TKoqQ9MBqeQcxY2zv8ht
rsx2d3qSEREb8quKzgEsb97dlLlvcrX3HQNt/MUBddSn+D0hJddMj0eBakBT8raq5Av8+m8aLj5A
xxTd8J5W+3oqweOZrWINhdUXU7D8YdUtS6QWJ62dj1c5Yfddswq6j1PP8nEst1KgLYmQ8HYrkswo
5N6SR9aJ6LJwN7O+AkngKZ/Lk/kEJQwh4dm5Mv3rzQgY7ObuRA/9vHnsnMasvv3KtYsNbr9pqPjA
T6xeLptNre/6ma6X4m2LW8S+PNfdnbiroIj0KZ6WazH7xwdUtAplzBJs/QFcihnXy4nvpS3jo7L9
/qzHR3vU92ihPmTOGueaXeJKhitEUBRMMMwYp4TVUVMc0D/atzaCV3k/k2Lk8LAEmrW52P+7H4Aa
naCdKlnfuLNkg07l3r2qmVwN6t/KyTsq6q0CoG6HGZwqiE5d9sxe9smySL7uKka1YraLuK1KR6Qh
MDw8ezfgPo7CdJyIrpj3tAXSD6SosE76ACFBEy9ehB3K1lZgORDlwf4porpfjNVmcmRqkhPqiJjF
Hmi1g+QcQN04gg28sSSfn0UUVLgro260/Ltw9Icz3HAf7spYQci8hjLNQWx10mCYuawfco5ewqkY
DPawhbeOgZ2dd6OSGGFYywVFI77pIk0vj7ZJwGQnU+W4GW528QoRp9QdyQtNdIhBrVK6kMTMp+m7
34vkl3/chEqje9KdXsu46WMonUcKA6U3kwu3d7/4dIqalHKM70Jf8fyUjOOAOIq3yDyuPaPac3sC
zQscYjLEG2xG1wVglbyzIDmTBNJ1VslPPE3c5czRC1wskZtu0kUgTaygSvAouvjhS1R1Q/1xfNGl
3mMJYLjCIuYnkcFklDGsStB5vTuQIHwAAlggsYPvECELFc4Ln60UxYaux6BWVwl6MzAyYi9T0myK
MwgfZ8yspsj+ICTZE2GrBVeNLEMZpeY2UbXtw2vjcOZCc9qwhIbvccx1JMfurQVY9YuHPaYjMbm2
zLurJhpLMR25D0c5/qk3PE4syLp6wiYIL0CWc+L3tyh1gUrd2cnxXAjp5Yj92iuOlZiiskGvpOmC
NFTWsCIcD2L+dySR9YV3x64194AYmUejnQqYEgB8HdYe7NCJMSK/EAyjIWfDyowqn5D911DQDU86
Ztz2qRijHvqM5l0k/fL8EgQgiUT1R18cUrzdNbtvQjWPUrqXdQ8oIXsIV/+kf7JsD8eH4NAOJNPo
imb1CODHqbSi7SfskWlpnbPY1EL0hhT+P9Z5CZXxUayBHCl1/vU9QBgFRyGYdp+ip10Ls4Q69/Mq
bo90dq7UQ22U6KBgyIPguQ9R35vyGlKc4eTmrbJR0MEZfZ83/OP/Ft5Tf4i4d3nJKFQAVYLEE6fl
YOvz4V3Wyrtkitwpx9DOVTrt8ihY9jOQePIw7A1k46fS/geugc8XjTiQcRqNIaNk7EwQ0dB/zwV2
JkjxhndPOKmS4MJHhNHMaCBXZWJBvvuteqQdpIXdH0T0ZvTPDaC6JzwiPsUKn/yJEsItjwTJKEl2
FgHTudya/xqW1YewqQGc7kGcY/UIHbTg95az6bPINKw4hymj+hTzi1HBXwyXZy8HzCVT3pojv2HB
2c7rFQ8Dg5ed1ZT5u1LgjQP61oux444pxI6oHqbmVV1JJTpgJlxQ9EpyJoZj546Y9NSa+WSm4S2P
Dx1CJfCS10853oaih0BwkFm0Bx2Frx0uda0OT8QSudyCMSm0CUVTs4TvlkIxPACDhzjdi6oUou5X
h6l6zUmzsTXKGVKKcWjgRXeU79MjUG/5/D/+SZo3fJ5W7G0qNZRtjbiM15Eu0k7KRvXCVhxRWYKG
fkeqREGN9m+8Kp/3toOpljROTmUcxG3MLpUITjk2enVRNI1K+Mo6NlG1dNlXnn4i1djGqBMGk1R7
V5yPtpvheJUF2SyPqTgyjL4HeD+p5UbeQs/xJtld2llRPa4XCoQazd9KV5didENgD2UNAfTjO0W3
sPr8gAqNSGlifxgM8X2veDa7lxP8BjgJeSNBoWkic2ODMal4FUY8r+JI+4cuexjc8R0jnIXpFiRo
sIgAPxyQWmY5BCX9JxolQXJu9nwbp+4ORgFjohjV2NPnwZg+b/pI75L4flacNiqYFPiObRZxxjLO
EPyaVkqsOMXHc9rEr73mCJuCjLkBvHX2uMowpoWtoW8+U/6173vCp3VP7r5IyUgWTf5zX7ixrBcH
+7IRnsVH4Guc9hBjYpt5Y9R5xSZI1SpHQuzufO8cKcG17c59QAnxVZBKtqv3VwN6OpKEvx0eRRgT
pB9K7/RHvGR6iOf4QOE/ckjl9GVqZ4NqslvO2ecehENfk1g1/HS9OPn5rX/nRfjJaMiVy1GvFEuT
CvochXMnwxiwpQVWMfv1MkcXI+XRoB0R3FyJvN8/qKk54ZKBUeFCka5dWcfQF0tBx0qPHZ8eEzLH
W5CCqyW4VMvYmr4hggCxSb4tyv3/w9Dcw+Rqe9Y+3VDnWpfogHgmeWaWw1VEjiKLXmL3NIOD/MFa
NsOHWWSGoB3axL1lIm3vvsLZwLNUrmp7XqTcqNT7//FaBSfV/gyDQWlEMRzfRdLpS4Z8schGC2CW
3uGf73J2X41Ujh6Ohn8eAwyWgtUeSQWhelVSdKrz+u2bTC6Q1Qkc52/lpNVsg0xLATAxmCJ2niU6
5dspECAp1CaaWrHTi/xZc4BKtMneyazRPkIGwJac/+R8wSM/o13IxTwZI1hvIz3wYPNK/+PuSOO+
flT2SSbAvznBBrEcapyhkNyoOca4VmKlEjZojUIoMw9tnnReUJBuizNmcTB+NFHw9131klu2kymJ
PY2msJfmVTwTFxbGvp0NOVSBCmpryB8J9Pg/laNG1EEHWcRVWrLcKNdgOrbeZp4jXWwvi2V4DV9V
qi8PJjaUG4FNt1yFHWIlExCRJWxdoktNO3/dIkjCSXxpXAt4M3uKRq3D549tgv1lvlyjYMPCeCaI
gGJfjQ9yLrYugHR+3KZjakEtmB2/y1nZSNXzyJgsodfjg9eG1M/L9muEdK7mL7BMSr3qdAUZEUFK
y3A5cn9toKLd5Clz5PLNMpaEeeoGsMT09yTi8WhLWZMGvoKa77LSzqDtP4RN2ku+A8rktP5yUXw5
QfDri0qPf8XEeZvlmD+9fhYgv33pUbu93qv6jakLtgPF/88GqVlifjJemYZ10rDsTQUCWjaMRfUn
C3CfmFqte9Eh17niCsX6xSn3eVsBcI8LcAzkpgr2nWIgpBJQUZR9nG1mx+xwUjV3piK42/idQwYs
qz+wvYFKFOJh0DmSnNCYu+2eckWRj4lQhEEG7A944hbiEEM4vRJoaTk5Z2MZyh2eZ0rYtEdc7KCC
lo/WYMdDVohGMXdreeo2rUUWfHuF1VKG49EugyyDGz1Z6JW1UWWQCmXpLnxZvBkp7z06MeHhNlOw
Vou2wfGInZRLzq3ZfxIsNeoRioS+/Y5fWSn2n1rVEf6581PkT3mbu3HtU/rNtO7PM1T7omkaiMTr
abtLF/u9/ViMdDq5+VG1P4Oe2JCYwZ0ytBlFVR4dfKqfoIGX3BUfvaIMQKzry1zlJOTqIxceqOoO
ss/98RWah2mbre8MIkGEgqQ8C5n7RVJke4zcsb7Rllan2ZPLGBgAoovVEg/iKBKulaoSM0xvTmZl
YmObSAQoprJji4V029BJisS/M2Oqk9UIq60kCAk/iYcoQiEz2Jh5CcjJvEJXAe5DTcPhyXMGQkXS
Bl3phswnj2nl8IBOdZIZ8c6iSnFRHC9GGo38s5nPOjbd7r31xLH5DcAMwzOFboEx0X9GARn9XWPI
Sr1/Q5Umq1UrAglHC3HejyZoYE5FvB/6DQKRdg0JI6B7D5JjKh5nwc4SupYCKNyGbttZu2jMP8Xc
6MI30q+Rvq05iF0qJbvUeJ/XfrmQxPB75WRvprQ3dz54Fr844tg2uN8n4hYv0yA6IVzk/bVXWuc8
aTFrafsCKgKxcTxJJO9yrw1/KY6F0KDF8uAJfjj0v5gWHs9gF85ElUB8fhBBjdVScqgyEX7QdPAJ
LlwcYxUlY3mAWkFz1yUo6YK5xdApjfUMiqkCk3OY7lYwkhbMA0PVmPDNqvM7T3nAHhVXn4L5cRNd
KMsLKmaQKq0o5x+gYv3+/y/pOBks/4UJkUt2EgeIBNftFRXzyMNOjNuqdh7SEmK8Z6OKyrkbgVxF
lXkuyZt2wZIuUP6Vnef4wUvYCSxrz3bwf5G17C8NR6mz+oEWifhviZIDevDW73NuXu5effWTRuwi
yPmCweZyNXdKPi0Qhorgn8gJFDlDDnVswAqNPLHKcGhvpr6SXpTQEtpiSnslFvtTiWOGLTvlVNWY
/7mg2dhEJccFcPp4fHzfSdNN0fqpvUSr+JhEb/HL99Tckjqkyf5lkBkh2AhBJAQGq7dbhBxioamG
uGtwVyNpBlEPOPkYqYXAvRJwsu2nLcELvmT9EzrcB6k+MR3IYcOva9u6MwGCv3XCh54SXxOfPhfX
S0f6jtdnT6GQ8yLth0CwaIrL4KZm5Q0UifoQSAQksv0yPZZaMUCKyIXz3mo7A3QGae90u55aPDxm
9giZnaENmlxZ7Gp0b/CZmpUI9UHRqDqLWKdI8BnuJ1M/LqYtjAd2laV1w+L683HmTqkP55aXkRFV
E/rGGHEbYMlypJqqNDJxpqjeUpVFLodNO8Orprs4DMYbJjwMqYg6DFcj6+MUuq9Okf4UVfB2mRa3
B1PaUMAX9btUwKtdd6xVerPCaTGdqcPLUCyUJZkRaWV3SeE+F/88y1AUJdKanMGI4LfJPdGOJ0ep
5YYiJp5YQBSoYiWZPl2jJQuTcAFCb3g5Eye7QZcZKLXTw7qQZWEXdx7xfXjLojZEA7dNi2Aif/z/
oniVl+TyasOTIOmqTKkjlpOH2LY9RD9s/a7hK/u/XxXgqzApM+C6JebSgzjJoSshrvSUSpkUhlAj
JwQjRg6MTr52IrfWY4kICeIcG67XUh+JsTkS6Bw2BYtQWBElut+8MZBURs6bY2sQgNv8aw4YZvpq
k9DaA3Ch6y4CaFoQCyGABgr4+PMDOEItcdw7LHxCkISEMkbBjaf6avmzJ62x2NT6TNBJA+Yi+SUG
6eo9K6iqn5iWfJbKBoqXIq2tjUsVDQYJuVAhDgUVhrd5ZNSzbWNc+73N6EdAO2Buih+taJIfTPWm
tqUrfUR4JNLCJm96ZXkl7xhoba8zUvHeFeAZiZQ4hzzsudBurSmJTSTrR01pCB+iZ7/4hwh+4JBo
M7WPEJKqgfJDs2T/e1bFHVMZhjEGhWyIkQ/5Y7KVcl0O8uYi+LHZ3zO17MfvvjQlsYV9o95MqLp0
/0307ZGs/D/qiVvX2V1Wns01OZ9sZuYGlBtK4JBdYsbX58BrjJ+fT4Tu7h9fTwOZfMHOs1WbNThM
mXhMQOopGeqgGTDARR4BrDVjy0QrJCJygxt4VUQULuyK4/83N9+CnSkDSknPtLZV/wpOyxR9E0JJ
Cme5DO8zl7bt9UnegSQw/IYMcfW8B8cKtL6F1534uk4uhQe+nPnRQPW2h2dA8pyvtPJZ5nFvaOx2
ZxDU5lj2ZBLBRfu8a2Cd+SwoCivcpsWQ/+ZrRV3gQ12AtsAwvoQOCsLn3P+3L73L8R17MVJmhKF5
EOpIm25XLb5QHudQvt32eJhGQfit+9M8mCg7R4jgRerMukq9wIPkSkJ6J2kH+2KfrYhzU5AZG9U9
Hp6GITIA7SEWKHvGTeIdhPyn1g4/Pa0kU7uqy1dHKzbix9XpgVXppDgYRqLo7hGuqdZW8dHJBf35
bbQ58FMfNolztUg+4jeuzcFJ+0h1fg6ryvWcJqib0Os84Pw0ccLfrVey0gSO6Bwy+qA+hP4XrKAo
oL2PNBKmHvAz1T6W/Osiq1JgYRUXSxMjPMBVlXWIforY48vPm92NWRjdwwebe4WNraeumtdrg4cN
fxsOQja2kElm+II+6k8jie0BWR/CZ3vFPMFTzZqgrlTcWbWINiaukyzFvFoQzKSqGFoppCmDxwjN
BAOsoBaxLyzlXTJ11QzIc7ix+EkOHS7wbSRgOOX5r3fRqv6MDrNsLoKmCr5CEaBdPCd48yQhZxUc
223Zfj+ZERuSPYspytb+GRhssQuJEQ2QK4ygNOp+Pb4dmNiC4x3iCJ8a2bP/aJIXps64kBmiRmWI
aY8eIhDUHsy0eqRgAsHIIHf+OVWmz+HCPlOAuoW7dgXQ29YqQzK0g7yzSmXWoL1WDAmEN4LIBstC
T4/vaZAD6TIf1fsNdXlkCcVOj7XyWZD5hSGjpfNKnYfopwTyKX0h/0NeEGmXyKgLo2Nt0NXUMade
UzmkR2Tr0P2IXreRRA9i+rjDRBUm0Ya4cRIvzT2zwnWjJ2EO6mj7d2Ey74C/VSe8w56K1E29/0n3
5vql7gNwcJCcJRhVDpWkmibiT5glvTXgHWpBGrXjSGv+fYZYDg6KZDO7ZbFDZC0qvjtJVPL3WonX
SYuebFLLgZOdv6aEGg/+RMxuG/MfON4EKYZ3m2T+IBNsHGLeHfvBxPVDS/FTz2SFoyMWCCGlaO+Z
OxnLyd9qDcl4vAgMI4g+VoYlJcnJwjLtrs1HAe6BtUpu/vizVeB3Rh74ar2bXh9hYeSoVgNbnULX
YdNZLo8/88Jjm3H3s9xPsnlW3CB034eJYTltBIY0Lc3LETRNY/OLod/ciAi2i39kFvLFftdQnes5
RmHzzWlEj9ERkakkUlk+5Lax/XwOJ0B+qurYiPaAtL1jgTXhBlELrbgATFR2aO5+D2Y6sCf2sW+M
txWo4d3TENkYb0+JG5XRw1EORb5A+J6AGli3Aw/6k0AtVAMUFIJoFWvKSomNj0hXHJ+GwTt1THjW
MEBNT65Y1MGylbuZwokJfPAvc3WT6YwLmmRRcGNFG04oPPlZaKdumpxt9xyJ3/1BhR9JFTF1qWJ5
MBG6E4AFqDPha+STCiw8ETT37A5YqJ4Wguwz7Q+PKr9DGuAcwlq593UcOxzFIa11rj1uxvGV3BD0
DwD352VvwqjzJ2HSFg1hoNt2RqwKwsB8UzhY7RvdhmGakCiL4Vm3Wr5KB/2XidNos+FnORErYW1X
AM/OFa7reQgPJrku+mg14ABfqa6jdWi9k2s7gGpIH8wdDL42KLUlzDZAb5lb2NeZKWY096Do9j4h
/cpg34FKS+5NIhI1KRuLPzJt3EbWRYE0vb1FyC1L40JkVo+ejSjTmWlU9oj5z5jNgiKlXnqYTCAh
xbW/CXFREHH1opMzpdN2qWIc4SC+xC6Bz/lQTHh+f0JRsM/CSvpRkmaHprk171yS1JNcHFVkb3CM
14Q0xPcVGvIShrD+Ee5izVirpzXI943+hkXuo/KQ2Bc2TIL6SKCAIA/NsffomZwxRVlYb04PKfqF
dDQ3B3s7lBsei/TGCmCGmbdsCZwQFcUbcndjlKM3G9QQnCokKrajfL/IvavqDwO7nPJyS93I3BfZ
JqcvEb6uTmlQbg8awj5BQL0B0dZTOvdRE+DXlkdvkMW8/4uq3fJ3bwUjUtXH88r3gx1PkLk6ZulP
fKiWWx43ozMSf5+HKaRrmsGDeE2oO8BOoncuUZ50SWD8bP12bRL/PuK2adEWBcGRA9EZJDl1Mjtn
PD+hmz9r5jeJAELkk6vqNPwG6NNnCI6iCzwAeZkXy076Uv7O3qOQctKIMlmxchgP1dLPP7VadPS7
uQLVRUzA3m/W7GHnmyIIi61cFopD+rFqqyzqOkiqG+eT/yzpfsU27Bk17oS0zBjb2kGrALn+/wVA
dftPbpeF68LRHRJoCQWx1IXxqqclz2EWDudafF0qLzE08ppnLSzLkKAhKGsqI02hhtBLjaGqgjm5
49WWvOFBaLI+4wGLQw2t2fdmb4C6/2IjbsviDL5qpBN97HPj6Q8ca7SIX0wTPXXWNKlE4WEYA/Tv
fP4EvG2Wkid/w6MqbPOB33ntFLE6Z6aEJp3Av79FwibmG0oIyjnN/qqIjR70MrqqHXM9mPV1P8sX
xiYB/u5PpdKMvRvdAA+7uR+PlSZLeTmIa78iXZLc59IJuzBJEfoHfMSXDUAR6WW00Ey6mJORq7R+
b9zDRm4Qde3jZDLowF8j/93c+HZwKNH1q0Mrg2uneF+a+YpaYgYOFqH4QE67qaxgUoEx70Ro4Ea6
i3vL/IgrfU198burvHvOkYL/tfod5cavZY4xZ7Cct3DpxVXtpIWvANt4A6Yqs4VBCAP5irtvgQm9
qeoehYpnpDUSp+aCoNK7VhWWcd4DWqL+KACN7Tt33WbPf6as+9lI4PD02jJFovvnOlEwMMSYfEss
mlo0QUOoO6cwKYWQv6PKLHK8jpF+GBerTjOq9cen7AEYwa/rKLQd/WB+NORhLiAFXRsZ+Zm9nGsk
E3akAj0jdGrHWdE8JYg8sRW4suIX0sxaSLwMnOuVYwi+714nVv/lgQgWumZB5t8zp2j+tdFGqB1m
PKtTHKiMoyH1iR+aEma9N3LN7TJsKyGhxzK9SOzVeHldHpnpf4KCs10977Bau74i066vKN6zNWxk
Sc8pKyxQBF+gohPRKV7FPp1uXCmmG98z0FRz5ISqPkjQ1n4a5L6RZN0OGxx73Da+eJK+JX0ikafG
trIOrc73cgzwloz+DiXREsYNiePDg8lOJnArhAGTMmQcu8QqpHHcBqA3/y5STRhiDGQgRDro51Mt
SjFqgaf2Oa7TiAQCJIkMEg2lA6xVARtd/hU9kOCjVn8I1vzb30m7IatkkbDJ8iHgxXp8oTBWLnrN
BBUAzCybgX2p+aJZekPT0TNsgstSZZ+6BeGXK/n2e/t5F7PlLs/l1Uo7s18GEkrSQuqLXKwdFL97
++TfLy4vh1b4b5/NUWSGVTJqHM+8zLkMfQZEnc/4Ok6aDxsefCr+w9u0WlW24axx+vwOXTfGr5tq
sDeh5vN4jNIfu+7SH1NpJH5HpoPe8+dPmXk+foneN3p4jnGKuWTMrSEcTXyHXk3SPhcyTl64m27z
qH2KPasVCnkt9Zndg62kzXj91phy0Qh6E3CVBaxgxDjXAfHh7u0Q6Pfb6WXXfkqJxPSvBXu7XQlx
la7AVnuu+O0JQcPZwrdytZp/Y0yxhBS1J96n3Tk7bKPKyPvvT2sL6LSwiaSmQOslwppAfJfhP5Gv
vxdI2WgYP6z1Tcb7s9Gvo8MxkrTt/IzT7Wbd+VwyKwiomBWyPIXpFJ28JWtvEYuK1qxsA3HrLkh7
7Ftp3mTLqq+3erMWNepodk+MKvPCAB5pP24LeHdlDeRSeblI6OmBs7DAsr8dyjr8sGnNjpSSgnW4
U8uLzqxs2S8ohI3bA8IjPcd5blW9Qn57FfpQbequ5X0ov9HrRtr6fKtObG0+TQxT9cltUprpVKqD
9xWGEgi1Oz6nSuLMFo/KsAN13Hq8Qo5cNJMJLHY2FDARBO6652RIVL+9Qtx9HtC/TokjMXuLgO+Q
LC0P9qznaWEHPWOmcC3G88id6bbGJS4EbkzxI/9zi9VcYtZng6GkK8gn2hTP+GBZuQtoLLItjQDp
NRWYG7u+i0IFrcWBUXxwmDLly3nmHyem6s8HT+90LiornNZ10RizYN7bhhgwPC9jsSW5iFhXNiUL
7Xgr1Xqngc859M0zdxRRq2r6HSQws77HhDr+0z1Mo0+cxh+nC+G915iHPTIHfR16FTKCsYS2uwko
aRqttu/RnwvaHUywaFSPXuqj8TyBJqaHDmf7KM/WX5QFObbZHFayITBY8/+C7kVrXBibONt8hzHP
YKWO7SLeTOQGtEB+I5nZm2MsWtImLJexdX3btMaTxypCtjreP3AqTG0yqpDzZiOhXAOFTVABsWkb
MZ6a5a7/2BgDXG8m55voPQq+sWpkl4qkSCpTIw2SqiLyMoOPEkmX0PmVwmlqos2r91MD/So5xNfG
KwwH12p5jiiQnr3jhr5jwP2wtyAvUbYWssrr+UBpPMCEuLH8zRF5CHEZs1flH1wXz9PNjTPILvZl
1fVQykVUOqRMBXvAEwqqAOryz51mb07z2IcR4B9p9lJVz+2B9NTkCE5vhFkPtgU/atkJrn4gbaZY
LkH78sglHY5/XW+hY0eL64nDditflWIojp2j30cpvHqfpn1LFsq7VFViN5EFUq7Yq51ys/VrdBQg
Yi5FLiGOmsQOP5gpMY7LcDqBIeUYIucSLXFuIYpucj/AkUdake5yIm21UhwgVBfz0HIJxFINEaeB
VUfnFZWIrG5wjr3dF3c/eSBafqjalhX3KTg5RKjkZacWuSHHB8zMbnpOY/tWfHkWSt/D4f8oFKIu
KbmM/XzvlIA0WW7kRD+EdrVbZofrLxLfj5wOMX8zoWtAGj7pfICEMLA8jnr+Wj9d/K9SU/Psx7U+
CtP5aS6kpr5ca41OZ9e47Frwm/tfNZuDZoHR/ts53WMSF61y/7LbGggNYLrQd+vCBYgM4TfP1qFn
aOUbzJRznpNWbfCKhWK6pKCZIcpQqkQkaveC4Omx5OBuCUlJN5TLIfwPR/zEYkqGcDyebZXKkwAo
onIbLxkgi2Ay6Ao1RaJJpIhDIcIDQ6RIUn6CafdYlOeWeeApQRI1cbVknydeG7TnyNts9q5Akc3r
mYUc3TKHdF+N/PvRCMckJzzHNqOkcFuavXK5BjlMrp4N2QJBDKLEDKRE52W9vV3yDyZkMR3C6IFJ
+QR0GZrCG/sMlyXKhXc60RoFdPEe0OKjEm7UHrgqKSgPgiqHV0QYAijlP2oKMf2esUQ3zERGhUfx
EsBhO1xDsNA9zlDwxU4yB2bHyxCwTOJbz6iMxt6vaRWPtT6nmaGXbMRFuJaLigLREKGKKbvgDgOp
0slpT5vd5zBKivMYdxAR/o9pXny0VHWd6K4eaWcBNoG1VhcK7pT13Fjw7m85fvRFdWS62IVMA/lA
Psgu9EJblZNz/pXn+UY+rKvWdvVnbuNYDM2+nA9gkKyMDjFp5AJloL0k1a5rfJ11tlRizLUrGuP4
buflddSeaiZXUCIT61P6z0TvWgD4w42wUVGwhtsJLNXE11AOTGPH9WLUyRUWRR0KDdld88obHAP8
XtYa6qeS6dcAfBcKMa/HeX+EETSc9d7oMPv9UNZVTMO8LuTt6+x2JPgwjD1azT/BEgf0oFo1fsV6
Zuyx/DGlouPmZTTlIMDNOzjZT0+kzBl7jY0837pWJeAggBzCa1lY02VSq1OMs79VCcwix0qg8ymV
CsRiI10jrPMOYd4Xzbr7Gi2JyV65Pe7T58HOQhO8PBER8OQeM44KJK0tSdjS5NT2ZxUXW7NSXn+t
g0Wj1eTTfUvS/ANA4tqCjvF5+zMLxkWLu09pEPLYm0SxzNge0Ck2LUznDJwp7eGA6afEnf/YvEyJ
vHwogQQ+4AVTBG8vYrJEkxKO6ZQfj5kJTv8UBhBGvtWip8hsVyrkKqQ1qqYQITRE1PmlFg+svPRP
jA05lzP0oBkXp6ybB57gglLrcEsFEj8xH8dobXwF12yyqOyQ5VopFHf7ef60D9paKa3xlMfAn4mn
msC0A9KtKE8M2ch1wWgT/7SHZLrRXW8inreYrSvMgJbjWrfT8PtR+i9bBhwJQHw1Wp6PFX2RzvjH
TODNpeeM3ykYBAWbFn0lqk0o3TBJP9FuCR9Rym8K+kY976CCpfCZW/Vxp2v6Ok0CAp01Y/0C7m5D
dKWVJ/dpdwz+aWGXXu2Fo9YrOOtYuQPx4cWV74F5QsRdmJk0ZZiz81HSh+Fs+wOYKdq4t7OEVMxH
wf4sz5KHSA1JUl2GOhNO86H/qd298aexYBGZHdwI8/nH2gq9+vV8KuscKGWCtzbwzcGOkLpLVrbS
xgzFgJALNiLRZhrSK4/kUKEHCrlbaSbiWpAcm9wLvh9YYYRVKJoln71JYCXF/Xc4PlbmiWKywsuq
iAC1O4gad+hmXcSj8PgQBG+jCIhElP8tU5gaYCH/R7ADpBDBMR6f4MlpG0GNd3TtIln6+De9wDv5
8DK8ucfSdEx5dwar6NneYruwP0tdhElwaTjXZti/xAGSSh3f22nqqcYlj/z2IBOOlWggn8WhZ+Zv
x0/kEvtA6xqmLsh+eDt9qNwSGPIrJRYIndkPwnbMJG5Iy6NWa7+R6qw31OyAnbMCWxvMx7Rbh9HQ
clm69oh91aAp8N7Mmyk2aJKvxWyvY/ZUlfWIuzCJbhCIndkiHXGtwRaRD+eBZC87AJxmiJ5GxzAP
CmWYmybDzyjxPfet5DUGhQh+T2ozMfOiWwwnbLN/tGD0Gs/etk39cPsZ1dpo3Wsb741aIdGaUGpm
4TXbTe6ujJBK+Cw2fo1TVG8hB7D6ypFjeAdEYjBEwpW73l/gb+R3IrzEs3wlDDQnDJ0Wkt7tvmx+
kVIq/JWwJg+jMnQiMFm1D2QaY+eZXuIvUCk39v8+BKpcaLajt4kJJ89tCYbTAIjriuo0XZvdvlpB
zRVXdW8b2HKPH+lkNsYJ3z9Rj6p2Zlg4+GPM9f31JIWbxKctRYMlxthr4G9LxWVng6slbCG6Cg6q
GMqVl1RAqVyXoULDFgakuVwU8efSaMb1496l6NXe62cFYIYD2+/jSgKIgI4BMy0dHgNCQh8cZwfR
+NwX75hihVOsViL9qDusj/mBdJK/bvf+MWOPB0L0mbetxWhUmGzgsEG9KXxqxlbWne+27BgsgbfD
wlCDU4Em4EVEZmAraBkRB9Zs0+unofrzGuiQagAWiNbwXMJdpImpeZBZsdf8lCUwXKh/mWM0QCoz
EwShseNPdUgAmhODZOiaehg3eomTDzRLt8f2yOAkw0YKesyosV+O2HiJ/GHy9pEOvAzbOWzPoY9G
ZVtVPEhgvzWM/zSTVzGUpOJwYgATRnpQhodG4d2iD8lGhbbwTRpd5rpOwtCG1sXQnvs4AcYXoudC
NWEGHKOIu1JBDwF2+4Rsxx0O0yq12VLYoA55enE+qJvb1V8e6s8jgnkK4Mdm2fW+5rnyeaOCQw+H
iEI3+84K1oSOjKamXUtMWgJxgxzUZhf8Cu+Qz+rtx+A52r/rxW30GpW2YhmLgyS2KHVgYTNRSdhd
kZpOVBEer07ImDa5THP0wn0azX7pqU8Gg7wS7RikLr5d3MeLaZ+BGlkVrK2asoOcjw7QtcCJVxel
BRpepFP37WyBmJqbuelEwSbfQXz2J1J+t6BqrAZXSK/vq9yfrEquFfkTc7UgZiejWE/l9eEbTKri
J56uuJh100u7x7zyaLE59wCZDIzBKhlP4gOA6IIdDmUNgN0B8c1VAzfGgBXrsxo6tEeSQqVCbju5
/Hrk/QIqX3bz8YaHsYJpv77WVBSh28NPa3c2UWJMFrmZh4DZ/UScXK5WUOSGQ+MWVl9n823dfBVM
xR5il94AVdiGXzv3xfTx5ODS0moPiBKInj8xWpPWv8t8UnuE+6NMeXJEQacxFPBYk5LrC1XShvgk
PgMLtXRyqMXxF4Ce8udUi8n8AkR3u9eRswA103D94VLTFsTFETrenZ5OZkpbPacAQzswodff7BlF
mLe40YFbees7PX4fjz0CZ2+cCu8SXedeqSW6vWplAyAQ3iydLVB1YECZhU5GANwNm+q7V7I0Wn1I
EQgJNZtFhXacGsFqnHewjzmzchhzGVZmGgHHRYctHtkQmM3j3ewBIvgGtXhj8AKR1Jq1VpwZPque
cnj1yK4bA+lhq8vvLLvwbsAE4j7/nSRzMZ9bKZnSECYzDD+9wLt2tlDjFj1XPrUTpnzrkV3sUfWS
LG0pJlgrzxPKUW4xm6YeUb5yh5MhAHfb2pgj5Xmdr+g+JUrqTE8T/gudDdRaKY/k74BSvKI1KGU/
lttX5m1KeK9jNEOT9QCP5N767xSQho75e2D8XHVDCY8XWBnnqJNBiLf1EMDaYdh3AnsAuRwhi46z
mqGeeB6G54U0bsEdxtSHJiVao7monfzW0gsyJlCfAtjXZzk3XxNnmNLSd+9PzBf1ULX4+DW7LcLO
h1ZSD5tl2wmbdTuhgc4JLmbNYuAPega5KccqKWvSF7gcogjgo15q1SP0dfVn7O5iGfMw9Swy8ilC
cMphIzDT2ERf8y3Td+u6Ja6AW6nPC/OUi1v3gc0fAZWk/YgRjIj6KG31lZi8DyPz4coPaIdvgg3S
rPuYCYhCoDuh+Kjoev3W+DiF1dQZk8yNPQCaNXHqwp5/vo6EgDI4ovE2tY6LO1YNM3uIcFWsmoQy
0G4XCdWt4vsD5tLGe3VH/DBOb3SaZcioo9nYs6kMPmyeR+M8lSzvo4VRz35fOFbM1AWECww8bU6g
aeAtc3y8KiiHcWkOvRV/f14UKhW+oLb4F9evfxG97j8BRQMpskhCD36aWiBDp0o+JNk67DHYSGLn
c0fEIp8h9k7AHsNAb+18bVoB2P+kV/XFaWSVNkamuy5z2pM9RgY6O7Atd/7kYsr56JdpCTs+TDqU
RMhtfWld+H1A7ySw9x+6aWKeiAznSi/o1PCP86DG5WuI9nmmfPCvB4bgqjT8DFlG5fRdI1JomJDC
ZTR/1NhhCIUdqg8yhshUzkyTdN4Z8DZy8Sj+9L8pKA2VZqBkkFzG0wpeYb75+0T5VUVw5DzIAKXa
jnU2MgAd0966rlwtjtFqVxrYkWvwHv5mFaaKbzRfrkIvaGAxXtWy69PexqSG7Zj+YA7auJE4icz3
5t55+9QLC7VgZ5YSvcn6xdg/9yNDD9gnXPPaT8PMAvpUJBB10SbkxkV/1BQ4pg7zGq8VeEbhybSK
ECqVPTXHtKmgFSdifSPWOdOuNZEuDsvBoI+/FVznQGtTzAl0VfwRjjWKnhJRxOVTDm3rhWY0SGNH
re2yIH159ngBIPGRJXLakNoFjoIEAaycdVtGJ6SCnknPUKX0KLCc08nP/iCO+b7WTDIE+gMn5r+I
iJv7HLpSDeWpBMuKJ3gML1BWhnk9P3p6t5ssQ4cnY075D1B5Mb72OtPQY8zimBW34xGThTAIgD8P
Sori1CXjVrVjaCML3A3bhVihuRV+UKpaZBtvNUypf+TAZWTGPLjDQOYc0+aQcV1GpzkAjv0usLuO
zYmCyvinKlniEIhNbsRjSkajKYz3Vu2iCt/bEDuVNSZ7R8Vq6wtqDSwAKj4KXxRaAilusGdUI2Va
dWaGFv0AWjC8KYCL0hxCg5Z8JsG4ANA5sb/3RahiZ11BcmsnZItYNCJMn4WITfJIBPBH9OTaC1DW
s0Xw9IGAksVlm09s6RvmhKObfJHn78rV+CxL4PYJ/8rNN5iOox5GkE4PFx4kVj7oBzvpHdvMeTop
S1LVgf1waIvdYgudmE2/lPwAoREPlZxq2xuRGaCw/0/aUrJcwnUHgceq8382qCX5wLQMQZiOoftR
bRw7JvfhkuEJW6PeVfTwDPooMr3SKWCdlbmMptEJB2qPg3AEvV8D6OmKYP1UvLJQ7rBTBPbMzrie
P8mTNFNbigQiNyyLvB+x4GMMABOnd9uVIwkeh1geCKR28LRR3jSB+Z1pPXMrvqJkoh05jtO1A98t
UCE7FUMUXpwu70iABSRSDhAncdzB33w+FZ9ESmzVpQUwhmbDDNQoA1QXNcG27X2GA2jtFTBG1Pjj
ea2Wh0QvwnUFeO4qFY6dFQSoVl8qt6x12M2g1k+4Nzzhz0aj0RjMgTFG+00U4AJhtPiewZwc+chw
4/sfZVtb3g+nGwQrRIlpxIDkO3fAA9upf55jn+Uo7Nw0rVLwoNCFnSq/wjzeJ+KwpnLxL5LaAGwQ
inPZEdSVTnfMLNkF0IJXV1f4zW1Cj1MZS3y1Olus3wcFp9Djlqqag7y7keTjhFrWkPBxQCnV920Z
n4/gZMYS46/Ix8ylG2RSWQf7cjJOasmuUr40INHvjvcyNM9oykQf4ccqJ8dZsoLkyU+JezicVD3Z
ZAf4kqDEhj1EjJUry7wQuPOelLUp2Fehcpi9EvloG8iZExJSJVg7YOtFRc7YrKbvY4Udrz+6tGr9
eh2M/dn+s3hdmiQHM2ARosrhAFpPB50hItA19x3Zd903RfBCWo+yV1+iGloBlowV91ZyfEATW1OV
gqEQk6x4n/pv6ktDKFDHe/1Df5XhtVyejhtuIJUAZBpab1XlO1uwNrmOGSV8V0DkIC7QmHrhwc5A
QQyqUpqD2bgvj98Px1hRlc6CK53U3TBA+ytgyMmdGaLXi7lbNCKbG+I9g/Z68f7pdwydYwmmftl2
hWp9IZkvsEHqIne9hE59Ily2n4MBiwKweFllKd4w6EdyMfRVnd2YeMo75IQbiTlHMeNCysRSb7ce
r+/NfPty1R/ux9PXGyo6CwYbSfTBgPKa8TMqzVXDOf7HTbz682DEoltDNAf1pCDmUNKNE4ya4IX1
8lQv7OQvVtE8W34ThoxWECOatG1Rcu0sw8OIIsfZkDCwzspg4J84oWkdgmk6CnvBBgB1oKaYw6B8
VaFVuTdeuYJIM4LVkME1Sj24BK5t9U+fV3As8bzwp75dInhAZ0e1t5ndimcUp2T6jLBY+qTnBXte
AUfAkR7h2C7sFkUq7G15C8UFDLt0ikLSEFkDP3jxa7FTVQEid2Y4YemQMLML/Pn6ihyX7pPdLkVL
S2wjp0B/kuk5xiacEK/hPvkoib7xv3h3pPy9Hsfs4xfqizEvo0kwLUInlaJTfeSLFavRcWLrA1AH
vdDAq8KcvoYSyP/QHB0OSp0G7e47hwwenM02QiIvQXKxdaFSEYp8FDwiszINbbmNqcDYRviZxO+4
yCJfBOwuKE8ueYecaqLXgDX5CpX5ND85cUaxWuIt3skhukMUkPOl+hOxS0ptechrPbfGwfDiuunq
Ka7IOSAevlu6p5DVZx6Cdtce7LsQoScjAa00Qq4gTRbydatvQv2L/1sYYBphc72Av26vcNLXL8H5
ODUKv8O6MYMfBlpT6XJrerRVSiM12F1Ve5q+J61iqIa1HDH6aHpzzYbBHTFO6JeJr3xk7K3xY4rO
pih7+rtwlDCsANYxqVxjlDV9fx12fGo7RAyyKftpqWfNpQxF70x7fd31ycZWidh9g1vw5uDfYPFa
iUu9dJk7wy4vHi9M9pb8EVuqoASsKtILxqd3GozDEUEOjsYgL/8/92vL6oJM1An40ux9NMNOUMPP
0KiG+EKB6tJFl1KoLMWZAT+oG6XH8qrTirXcbM5Qq+G/2RrX7DzFPYp6juh9y6hHH6wV93cAULNF
1n7vCuc6h91TEmUimDiym1lc/SBruwjKDZEnwb7trqyyTmQOH6fQSisKcH+zk4BF4Gv9Uh59y7ZH
XeLQSpN6XhEisriwYIMx93RPwzt/4hjznfZ2GPCBjelZJADjNyq3SAyGzdg2WmUU2DBmheOJM/4k
+jiF1D5Vq69hSi8Q/lY1ZyhNoBtDDx0MOinlK426hZgGbHDx0JHwcISHP3hZJe88iadnJE8nbJuj
8/18Oqlpp+sj+8qAerIH76zAYtYytSg68kDQt+OXbJqZbx/1tjkbgahkysDLqA4QemfxUBPwApqO
P5Xvb8Kq6BCjfuHNFzcsnSundbXe9lRzO4c12+Yf1xuj6hExyZB8otLL9uUoqjpq3Cnd6yV1ns5w
RVFLQp0rusfCqbKapU2+rjbx/ywbJ3bkcbW+TetgGLDKBd4L9AlOQAgzNJAaS7xRUS8m7tZ25yVK
GxZtNb4qqRP0E/gdzXZ2M7emPhwm15hVRQV9KCrWZmN7Pam2ATP65jUANih4iQAcgSqa1+L+JuMv
9pdZfHeJMYHeB+aAe8i0ASONsJR1ijw0qbeNbmU6yvm3JtLzujv1Nr83mGxm9sdvc/Xhw9HnAXTA
KFybht2aAIc/TOs/cTmd5+QWjO4q2ccT9ANx5mVea0G6kKdA42YypCgkaWHcRKJfk3fDkeZZckTA
Xpku0sNZzx8fhUqQRPHy6Gok+9PPt7UegbdoQTdgpUGHc6K/63Su6v82fVLS60VnVR6k44jEIxhD
25LTG3lJbldSMRpDVDE8tQW8P2p0livaiX5qz2LWiuFXNFCGLuxPxk59Y0QYIMriVJTFqcPKsPKz
ZxGvdQioyE/4xjIiPOuybSTf4gkKkRwe/Wh0fF9rqDQkiCMAFhdzEJdjMjvXLlwUl5PCdGJ7gGG9
8pTY2kGARnH/LEC3jglqgLXDKM6rcbJ6JKjzTHRqA/L2gnCMgKrTjpQ198vQu7DiGaQGRMyJDBc1
XhEnxSRdhbV/OPnRf+X/g+dAnXzO31MFTKT8rbXplQRIj0RUw0DZfPyIIvzCcUil9qc4JQcP7JN7
DnH2nXdIx0Fy6uivwY3mnbjUp3skiChWfI+A2wVIltnEnIFMUjFsQsHAPs/va4EtPE8yvZV4lsZW
DFKQUx545haQ+G+uSWXG6FmzYPLz2116hlxcHdEu349Bdi5vCS0jhr7uMtRUr+C1FivAVLV2L5Fr
7RAeFGl1M7YOf5ICqwPvV9kS1VAd/fzKm9YT1CjSjpOu5qIIDVJqlz18zeNKk7cIlOFq6rTUgkYU
m9s+Dt9aEfnP5r5/U4nGnahnq626LHpaLEKsIano22IKA7Jxpbr+QVPNg6ycDaOgz3ADngGIzxPa
OM/FtnsGzTBB4+XE4jgUgBXkCCjR9pbD/sT29O4XvxuoY54+jIdPXE0uw9NTgnSSVsm9+RsaF4Yr
BDoiajjxAOk9SdlPG7FsZ28J4bn3C1IbXGPXsHwFE5hbiIl/ZAJOySJkk+hbXUWTV/5dEnNRJ7yU
BRd0xNGEivf8kOen1faklua9U1UUhzZVG2ytlzjhI0Ii3UyX1kkb5RyN0zqX6GgxzTCqMXesvQIH
LdaDTxTqZdXvGZ4d96bHRbH0eeB0ogKpyYDeHJWfAJutL48F4eEXls+dQTYf2ahKMJJy2coi1n5R
uxb1P2pqSmzQavvekyilAow2aEeJyn3P3PsNJvfOUaxVKjU77Dz5kvzydWXHfgReOiSjwTjfLXdV
ZfnxNgyi4ZEWoLFDpabDDaFYQCdUHaH11bwi3y+GIgpy/6cbJxzES0c7tTVVXNAUisp58TS5N9Zv
bgamAnb32/aJBwTgSh3g9s/ryNEOHJ9cK5lXE/Tuj8F7lX23QSEdayJGkBLf85Bz2az7SDmPltDM
Vmn+aVkZzzWsE/LY3gcG0+aFLzmMHYORh+Jx6eS37rBUKKRUFyHLrRhkrEhCn1T5Rhp24CAVO3lS
D2nB0CysdbHjumLfjRQvILKdMKsYABuKXJvKN7bj2XFyUdGvuQadvVbxT77Kjic3Ao6If7HZJUkX
vRVYbErG0xe/bw3qPbM6vUTFYN5QC3/u0JnMPe2fOoPbbpPG1n8sA80wK7yaIRxXzaKBUZGpP20B
l0uC00ADlOa/fYg+5EeVF0fqJtcPL+lw5N5PCUiEbvhVbTr5hcaPXfSvEZBY9Q2UzKxnbeh6jJD6
0OFnqiU8jl989V0K5Vu6nt2fJk2ogQ0xwm/ZqxoHE6pMwQh7owytOvULYS+bQ84Y72vb/3dZnB1z
M3o/5HVSkpqzCyx3tVopNdhCpHTHSUcGENy+UZJI76b31HAcmB81aGz9Jrt99FXjD7W3Pt2TlQbz
OEgGGXnf5K8lFr/eWFcd1E8irWyINXwubJVjQHk9ez2PbssaTDLEU6NZlkpLJ3YzEttW0zVh1FVi
YSO8j94/nwiJ4TYj9BaATLF6koJAjUqiquco8FqPEIYB+gBlQCc9RoxsfOzqq4blKJeBcJArVIK7
sE1VfOOhkLhmfXcftmfupjlPrixmqni06wzuP0fdxLf3z0Bcps8ywIykdluRwbmc3odok40H77aK
5GFhxrcpfHHI0rIothpus59rjkfLmwYJzaab0f9bmx0ubCtAbP8z6ZgIvUMAtZCLfpC2oj9u5Nxi
gY2MLT/EovEwHfGIbANLJGmx4XQTCTUSVI1SsRNUsT3Gf6PpYPihyk3T87lAUmgEiYRZ6pFgkVkr
wppWyEfS/Hz335oyF2W7BFmz+fDMxtSt4fy2CYr3tFSSHfonFu1/bngMVS9XRwkGCyO3OB7bASDR
CuVsnBtM4dSuhRvPJwGKtHPnTEzmhyYzJA8qmo/aB/n1hmxe/hCILJgYwkDc7AZ7Fw8NF4Hsn1c5
lvL8Gger3TrQ8BFi6P0yteJRDW8il5hsOzELFbFjZdWHMilXo7tkHCA8PsDxaFrmXb84STv7dLfO
iwTMzNRgbJttaZA9yh/j6YBo2ll+LYO8vFvJuvef3qaqrFRp7SbFTOX+zY9tJlInpHOPZM+0zYB8
rvUc1OfZ7yuQqI2vctvRSDb+9UDLK7JjBdoznYzcZ+hmErgMeIc8SB7aIGi17KBF/MhMqTWUb7cl
StVIyPuvPwdOMhq9iLPOKAzPsqROWR/8xno4WSL+iBsoo5sKPDqei4O4934Boz5dQwsSTWevFmmB
LSQoA/QTCEVxWdRcpmear+GRBjk6TRFDGhTrr7gBZV/M1XigL0O/l8JrWgDDgjrDypZ8OWI7c3Rl
pRoVtTBH339d87YxaqP5l27cQYVjzOA3nB6eT7Rsci6BUuXfW4jvTfF1zLGOARL0883t/gEW04jq
YB1XOdoiIURYiMTvuvbOQfTSDVJ+rUugs7sBgCgOki4pgOEJhvybodVck9RtdI0HYXIrWJ2C5y15
cZrlBwRF7ZoWJR/hejXb86A5yD3KzV2ZNIWNeEg0y16/dLldW3VgOp7UeelieyzrwPvxyQVHxL9H
uAuOUpOhUAXQIHMr4I2BhJISJ7iwDDnyLjTymzmVaehzL6oKl9aiC6a1WwhydJOwjnZdJ3hY4nct
ZEab0ZlDdHgyilp1ZiYfjO+jOFDAtfsj6OwGebH7K2WLVqmp+9beVYX40tefdBkd4l4lMV7OitHn
uo27iD57HfCF3NztdTx5ugOvwl4Ez5MhwC89D5RbYnAghnDDz7ubukAXS8oQGUSTfZBwzmFsBfMF
ligMV5IQq2cPQ9pXiBCXEyR0TBVjaqDr8c1KSCW3qCBbRREY/1M3QCApL1h9YWYrVyvF/sFjj6Nt
tyQU76NspyBaVs3bqNdC0XceagmUOA4XgYol7RB2Ps7VrQ98d9Q/VBUdOxtL1/QaSIDXAg3W/WwN
zlcXBu2vumnYm652/5PYTwSDIkuNC6L1Q23aWkojfiibVCcptNXhlGBu3Fe8pMe0ZZnD5hjXWKZi
Gee+p90OZ385+kJKZr7tRcxw9spvRzr6+cxwuVm/J1kk9fuqeODJLC3Iu3RmU0sHZNXCfGEWVQt7
okrK5d8k8l8dyOLz4XspSDslj52DnCtF3g8vKz/fqIUrHd6thlQdz11E7QDTyoeBOt7QAJd+kUvC
rxLNc0mk3tM/ti60W4VJ50GTvEdaQ0rgqnrc402eJjWrU2WiEv/5SXk6YQgIj9r3YfS++c/e1hSl
WAEsfIJZtF5sh1cNZdQsGZj4VC34z6yx56DWuWOGDgCKVHnHQxRVt3OQBjBrNUy3c4cmp3jxjzzz
fSw4/G/BQFOnVSoaIWeVSVRqlSW6igTreZiS6Wn8QY1CtEnltHOt49z+fxlBtFU3PILXqtcGI8IN
kb+AkYGevLTqj4k1C8W/VXBd9xFaICgKPr8uzCwzqLIHY2Ww/QiTMAj01fHCt2qe8ULj5gtkKCfk
0DLQ3IPCxyi4QyQs4764e7VOkSRDQ47hv1feWMSF7z5ukof0e8bvFwI8Tj1+CPRW64u7+s2hFKNu
gk5cVJC5Wcf8M54sHizKLGXGjILbEzyvKn3x0HmYruAlYIET82OwT9HT/NR9m/Gk0X3/xlLc8Qin
YdElX83lwfqryvg72SjRjV34JDyXa9jBg5iDXGCE8lQ6TSijCegVj68pEQfUUScM1OveisALlVeu
TzVx/DbDLTXmn/0bp87y4aPgsDo2ftm15o01XOtHJDeo/78xBwn8q3AqoxU4A7h8ftWHxcXHPush
nU3RU8/0ZryvUz8gOTeibSjMxf32n+iFtxJ0TOfl7YaJNvPm3yJEEVS9hY/pqq15BSyM0RMhA+MH
w+bEV7U6MQwR1LmFkLVMGbi0+f9ZIwphrurQAFnQARDWK0yaBNz7EnFnxkzSxvSSd8JhfEtZiZ/7
K3YSPkZu2Cx97cxCdb21QrLz9u7/IyPp/8f0usq1lrbGGVlWqwHt9X77ZvstL05e8ThiURgNLD9P
Lp5iV4Knvg0OG/VVHFSEKSdBLl2lSzvqEIRLn6TotQGkWuyhDvLXRMemClkhNmmaVc/wj13xy4pt
7nIkBtIZneeeQ6O+eIfOW4uzb/My5y6UcZpKoABnZ+W7QfvFHUob8Lygp4PPhJi3IWZNo5tenMwP
cQRhMzwZtej9i2eB+2J6Ln119utx1WNCXER2DSu7ga083sDVvNn6zNJOOciG4mgVeNUQa/GAbG1Y
AlGvYC3SV7m4n1/0bpPlWsEgqqNQohRuJQ64Eo9e3CuEp81e501WFcWndnl8oYueD7WI7QFv61GI
NsB2vvyze72JmbABjQ1SPIKtVhE3zaYl2aDiB9guYcu1TmjnYC4OFJCLbYR156sLRfXqM5BVvYfY
wgV3jk9Xlw/HUKzAv8cafUBRWe/+jbRlALh2yYiwgyos455hxU94v51KHf9ygLQpVZw2FkTGqh43
S5cygVv9+E11+xtnO7L2f+mKt+y3hoR5UOWXeJYmtBtp4FXREvf4vnwMV1C16SByt2F4W4E9CjKI
V4Vq/238dvlXHkf8YoZn1WoyELfQT1d43cVxoYhGkxF0WnGrF7BFEcjG9VZStMAsOlqY1ktg0/FY
n8akEo2slO4sEv7ftFw6NScyuxTdNDKutSVskiKgpfiMu01YQ2LJ061w7VnFFJqekR1LEBS3/cLn
t2KuvwKBzz9SCEUe74vo2A+I4rW9GBTDNDc3V4LrGUNCrKd4d9RM3b1UcdVGExulyBDB/AHqyLqb
19eQp5DPs+oUWTCTbDYqbB9DsLMi9FvVyQjuteC+4RptxDTaxgLqzRicCinPjQEZCKVyLYBP7Z63
jbO1yInVZdxvDTedW5fne/JscwMvQjnL/Wjj4DMQWKN1HSxqi+Y4vfGlKuMcgNNN6AGikmxmiWIl
DQU3jDU95D/dhLIRo64dYhPlmAr2yBAA/LcwnJr0obexKCsFWzQVAxFNSRGMlRUjTz9a4SbnhHie
7VZEV4bxZiMFXp8ue6AYlYDOhAYkUF44iM7zbbtIAcfiI1Ho97EK8qnB+2VnpWrvfhwopbwOe3EI
ZiPyd0vNTItVsHGo5dJ2B20Gxnt9Qpzvzcm2GMtwrWvA5yUuQbmvsC52oHKOnP/0/v7+0SMjFd/q
XBgHnhh0N2PTmbcz2U/kfOcyObYcA8X0aRcX+sbrp5YGn6GLUBAfcOVyLc5Li0ceuwwfSgGTwgua
3VYUE5RYM/eEH52hpUL8YsOixVVGPzmP3rfGhw9a1oqirrgEnqtZH7y/DCw+M3Q6YNfrNAgeSzXi
g62Iom2bBcob25GlwnIS9OU2vOU75MQxBnw+JwFf22/I0pRrba39E+juCZduN6/1PCfsWvjuus1c
xKXl15jP5IgxlVT7AKP1wfqaOBYrpcpSJZvyUZ/x16eBwYibui6MVsSIvF0eHxW8RFcfaNjoSGTI
E0SSd3CVYqkHjmc7OZwRsSe96tq6JtcvtLhZkiN+uSHA+2BU+x0+Ncwdpqy8AvVIgHv7axnFZm/T
ADOirNn1N6Bos5BPTjusBxrpZyWgOQYIAN1Uk9s971UusxzbOMJMbo8vJjNvtuY3SU+I/NROzHTX
u3+YMtqpfA7jNrY1k08oReYdRsangU2GD7AOqxBhPo5YqmcOJFfU+eyeHA1iDgEGPVkagwFSBDUv
PvF/miVH2hPUCtpZypST2wbQsUksF432l1fWELtzrd3VpksJjeLXb+X1oSRc/PipygdMw8bKg6q6
7AYB6TccPc+Xk5c5Om+/nC7gmGC8/pjIif6Lz7NP0b1j/O2jPwMMPGUq49Llz17vZSZYT4pibVrV
pqprC31Zci3cWWTjpn3Yzywfjapk0EiIXv4Um5dgmBiQtskQ+4g9la/VrfELGYj9S0NAVzUEt8cl
MK4uSAQ8ZaAOpCawZ90fVOFyoILZh4JigbkYXBKjLWtsW8BOKXLoYJ8SZxVnqf9ST3/IOSpoYJKZ
SZNbqTU7jVen0Nz72U1WDXRVT9xjnfZMn+X710e+fJnjANhD1OhWL+73A6/Vjb0+aVi9RdN/fo9U
k6bvfZGCE+6gj+ZnubEoz6J726A3Z9QaSebNekrCoDV35DtT9qe03fLV2+IzYeyneWXT7ZzyjmJn
ZPzgdMhbzStBuai1ZmDk2HKCTQsk5dP8aQJTpHlo/Y65VxSXLiSFUW6iyCdI7hMOsFkqAkvPF/DS
cThDkBnRavTh1BO6zrm/v3ufX5S+Oxl8ZPJEr2LnpgcSMcHGqC79Uvg6s4uIbkL3J9PUfTjWujFc
pyctXbLrdZGhkUR596/IEqJRscDgu0euSdvSAwxP5wsQG8/fTLu5245ZYL2gAu/onbTGkR1texiu
3tJizjMvr7GkI7fuVPNepa7CpIhnjW2vggLbPXoSqp8skjI5bE7i9MnOh9l21tiVwxDqvO4gdzfL
37F5VbVBZpBxl0eHtBqllT254QFv9sXlSCeeRrRWyTvin1D3w0ymcnj+h0XyzTRtDpjXkjNcCiTc
USbw/r+MwGIezEySObO9LoVSiINuMSCfXCQXcKMxSYeYSiJnusgLwGAcZX/lZoYGGXlg5x3GcmrH
tlMmvPgiF3krZPAgxKTxzMZYB4OZUzNDd2oyXKNlnvuTugTweQ1CYF04XKSx0dEjyp1+0mbpv3tn
hhP7VGsfybbABq4fvePjJyrBWb6pPlNmpYHO87CdldWJP0UDhOmzETlEKYXVQejA34ATUOhX0l97
EjQEurLSsQeiukBtsHYOp5ppxQfxvmVIleyecC8nDksxNASq2bXEP//TujqsxKPZihUzarQgEJgy
1tMPt6i0bZVtg85D03hfNbN4koxLZDhPOsyQbsj30nQXjgLTkF4vSNZDHThiXMGZg0e7eeL49L5A
iNLu3P7+j+bQFkn/0zOlXyC568ZTIvlL/liQBV4SSczzM4Z0CUQC4G+4aURM5VciAj2zhd0LJsok
Rn2UfX9agFYJvCg7kcuIAyPMpGWhQJqgXpW+r/4DQTM+MJT7OxHpedieSOh4C4cQUmZdhfZ6PAd/
YjOt/UdoAxhypI1xuVBE7aATMBHuUlmGVr5PJfSA/TU6qpWv5bvb/pj2NuWgT649SFpcriB+8dtc
cZUSxTtjayJ5TwOkp3lrzVfpOzyQUKI6JfFLBkOdA/3ucGymFqMW8XhR7y2AixPQK6Y72QR3+Qnw
oYbu7xFA+5Tcv5fcmcGFjBRBe+8faiwqE8v+KOYKfxyNPeI8KUSqVeTght0NrNzdArNu+suE4GlS
XQkhDnS3YDKZiZi5PJzIS4ALWzXt+UFP3j4qN/NJU0Qh4SHWM/CiRs7TB95KPvcQHYNknkUkIH5N
jU9kpN461ZcjVnHiVDqrF639rTLlWteHn1GQ1sVs/IQe9QgiE8qkA7Y4WmvaSnyc12EYkciPXLUb
Ebc3YCW2Tgd5o77JeQOJuQIsE6k6dD+q6ziuro4crgbskDnoMaWoAzzGIZNbmIJgDTABfPn81DHC
w/ktT+rlugmWQxhooY1UX/EJPC8om3p9uJl+uHtlW6gcFBeWGBMOPEvH6LczvqNsuOG8LzVucrdq
aMsjRNZ3Jqkxp2K8L4pTh2XCy9Mvfb6FpmdNGIZtijwaIUd0CSfbOGUFZThYBPEeYo32UTWzS3pi
WH5cjtRfjrY9AQzajkdv675dt7b+2Q7sTt1qlftLj/J4OfB0LSBNO6crQSfEDEp3HxpaYGaEKRJS
F+C5ZdA1g04snM5GXPK2J4nW55ijsCISDwV4JpkGKGYK35IqTy9SzUM3sJslA+aWyh9oWfOVOHDW
xK2pbaXdcXeCW3yi6yn/uprxm+kGEWa54ZD9Vgcc9fwPRaEiKGcuEZV9ipzXtNeQ2YtIMwQ6ll4W
q4OmIr4YHeOTpIiiLGnXf+yydGLYgZa74CJgECHPX8TP7CCSQzDZeuayshPcQQLZdbwtWuiumJSk
Ag2bonHZ/Id+2wDC0a3gV3cMbTOL/9kmsCaSALipDpKwHRGpFFhOXjVev+XJSs11shXC38Ba6PKk
fRu7UVd/yf3MiNI7jvIZK0YWPSb2zI1kMF1L6QN2X74J3PavAahBqwBynmK2atb9u6rvRQ9NOxPw
A8HotpykKl5UJ3P5VvWRnnkoakm8jXPhCJzJXVFaEpEMQerCNWOzsOIS0J+Db1qRl6AbR8ItzvdQ
wRIzNqyAIsmgBrumRS5LoSs3Vgw+Zd5a9yn/eHfd5u3V77sF7rFPsAyh5vgbfXhI4CCMimVrHCfT
6AjR+TNNhP5TJdPEiVBrLq1Jtdr8RqrJlHvnxv6fqrw9qVpnjclWEBXxpnXgmbxDjYyAY3bNPJIA
r8Kou2B+5wLpHpmMb4irtBuh7fDTSVsvtXscrKbxJaUHtzTEYGJFZwL0/rOrUy/K1sWCHh6Q6iXP
WwORxeiqtPnuHyBDZ98BVxuMY3u7HefyROAjesv5PsM+yi5v3JPj+U0dx3IsYAQKxsB8h3rjrIAh
w72TIieQYyALQLPL4EYDrhkRSQFdq1Z6J0sNZuGFRRVDdNWb5qsnd6mQe1asSbC/U5Nfj88gYraI
cbsbdl9+JCa8aWxHwkyWGeFYLbOBndvNUyKPzKkZ8bze/SXqEklDxt7mN5nMQg2cp1ncLeoHVqXI
9Aa4M6JkdFfepUnLHLF8j7P3hD4PMkbEB//CPZhxkJNQRsF6uQ2RhiEfDLXoNH8fwqtdwL4kVG5i
bL+UX4WvGfjDTWwxl2Rekpa/qRSMcFVzqIqof/nYIOiVeHd7bJIOw9XFVP3ox9O/vm4KTrD7/99F
l6hhHfwm6DDCMxKiGfRxxiZBvbWd78e3GQYrFseoK+RQTDJB04SpefJ4bt2lmjS1mindYeLvF/m4
aRbx/ewsXSs/HNzzGRfAy4lw2L0UXeP/PXPGSV6GN0FJ/GW/tOlHV8+LlPJakTpKI+nw/zCaFsXI
hxHBgaoF4QI7gbaLjX0e0I2x4PtywHcKtMvSvD9FPn2soeFsBpaIjnVbztWpEasvM7Le/QEHia3I
yMUSZvL+qrVF+NP5iMLv9AYf68z8hIu3V5fI2+cOwxpv4YHIdIJMqfkiwSMncNDul72OZGQqLRDk
84JGku514f8KkhVSK0OWUOwPnsHGmMtk1wzeiiSFL2LNQtrZvGHQwxzPdgVkF0a1GglrPpsqEAg6
T1RKFmH66xycrrHhXCQu5VgtiSf4HakeVtNnQSHqPdfmr4k/2UA3miQAmC2TmHYbtjtDhEKygdOo
U9Jx2ZM4HDfGjwT/r8ZdoT3bMV0qeAE6eEKwDW5Q65a4wJ1irN08WzRkMxb7ec0S8vkE9pKi3EUQ
8gCj5XceBEU0PCGtXK6EJ5yefMcyK08XULkXPFDD5YkkKhcR8rIGBAIO3dB4q/c1y+Uj7fCGx13k
wFEqLAYTChNEmYy/EwZArAembHujn9+KmtEvx2rN2I8zoFijSX792365qEkNE9RCsx6YSkOtwqy5
sJqQ8p7GAVoV2YKNstFna+S5KuHbAeqEXKq0h+2JInEAZ62GcMZ7Q0SiTKPPnJ7D7BwYk1Xcevvs
KUsPNeBOmxlL89rNq+C9ThXGBY6tie5QslpHuZh375u2RBnrz3XBtl32F79Vv3NEVI1+coxbbmbc
j5UGXfH4HsZ4IljPLYiXuHmTQoxg4odSQCCLzcHl+ae9KWSBsfetp+waw1dNp27l4jFXqKwpNKAv
++JT34IJMhiZ8/Xbfg73D9pwR3Zfj6wT6KVnaJ/F9kmQZZpwthVymZ79Aj8Sgn2wsOigV9SJ+kBx
1ggHR/14U8uRVNY6kBlN+Z1Z4WCpM/+4tAjCcJdyZVtO471i5ClkC6NIY+LXlr95D6yejuGIBrLc
96nlO57E/4jqCKwvFzOfxUSxKJus+IYfaV3QVBa/n8jMuQI+jlP/bPeUxgvBZxDu3pyss4+1qEMI
2EptP5j933Kg0z0Q6qqGLxeKzm13/IDmm+vJ8dPPVK8rlsZ5k/Eoz4QnQcjnWk29BPYv8opnegGg
O7VniKWyRHknrxEiOdAzSo8yAUd52zkywLQ+wsRkCbf5Gg3Cyyft25CvxP6SOl/QGp7FvYbQXPl5
Vv3dsOCZDWHpho3jKfrN0uwnXx5oSqXHNlbKXdoXKm0R3dRTmeqSmTfrhDUUZ8fLI0u3aL2i1zZR
I8CrWOuUIodDiVeBZIcOLi2gt2g793WDfoov+/Isrsm4wlW1X4or43JCe2EclSdzQlJD6BvLVto9
KaNBDkocjhc95YppMVGLxou1ZAozHPoKoSmSuKw3O8KlSax0En+Ht0f2wQXX1moiVbpvUW3JxWmG
DbEdBcNWk8TNClkx8X0jR88qLDXf3YR2tyFrjG15u6YInUnstsW8Hzdyzz5dp4m/4JJgXdHUYN98
Nswo2xejpKgLTVQOZmdkBt71tU5zhIMWUR2h9uNpzAIG0+WvaGvGM/RRGvNvkUeZc1TSObt5Zf6p
ttdxNtIT4Mz/oxFblEQnx+Cs+LnucEmaB0hVEC6rj/3LYZckmfD3abV6UXZs3FWKkH4sGZOZ8JKJ
L57waGe2cvVoGirL//oP3SBD66yKcFIC/rpB3OQpBKIJjpiwBnPJb72G4H97NgVCXd5/27m1hmKl
uSz8aLHaw4hM5ckEVSHDm0281/170DscrAHcJHHFvxTA3RMiSO7C/26+Hq2yUIjTfhTaE/V4KLDA
/WZRbW/hI4QnbVAzhb9ikrRHFGKlDpvU526dZmiZuK/z2CgWfQVoGmi2MWwsPEDlmCzdCDjysDxa
FjoF3+nt+WG7wR8FAspyNgUCeHGMQYiulO5XQeHTnlctqPpdyMS8UPwyp9i6VhD98ksf1mpGia6D
w1zZdIMrKXN/xdQ0XAfqoo5KJJGcre8CBlj3BCM+Ky6Krc3jVeVZMAFJRvbNhnyCdlRb2d02SEwZ
vKYZ51Vizy4upMR/y1FXrBDWxV/xk1pLbH5TJTi3H4hVwJFCmLLXEfIfKyswiu5tETYqejrDdORf
eqG2fMJFtProKKKdarHD6xnvwIoesQL0RUife6IM4sPeXWqh1RIHZc18MSydkNsa2ygJQVFLPy+5
umHxhYWOmcNOjPbz5+3bT5aLVk39a77vavvcBAnegByWMTDtij19ylB9QTrZUa6O2CgvaVq+SXk7
Jix8fOSUW1oWHVZfZtrZOYI9Wighf9muIC3sAknyK3Z/sC3WdXZPxPqZINXGrfnUiX+b4Ra55/Ov
2cCz12BksVXqeeQJwhiSWFzEWEWbMDYN9TttVnpTHz/uT7YNWZY+UFmN+5al/P1O+xbqS7DwIfLj
517jgXiE9+yOtzTgqIpBZm9PHgn25ER4EKZRSp0xEsoDk9tLxMC3VtAzo0WLb5CQYNLM7On0iwwK
AaqEyEfzWykvsoHPFkyYWzG1aN/wjLNrhE4HW48uE2Glnc9xmiTfTqIxBpV5jlqKeVI7T0alQ4eh
dT4XI7m2lxwkD1LiJdDbQbbpQ8c6tcixbWOxPC7lyFnhLh5Yher4w1O45WgJEy3jeclA7bdKqfMl
TLZmLJzGvZBvFl8mF8b1qBJUp5REsZ2vbYyniaTC+jt8BJU2IKKhnYvF9GLYg97qz8mg574eH5Yd
PxGPu8ASgVLnCa6nc9YXaZwwpxbcYUyifBUB3pcKNS0BNoKErVdTNa7D+Bjc9I2e0aA4pFHdlZ0r
DQ9E8cOYhwjcgjQjcNIQpIXOyHxa/9cSm909AbOHb0v7Y2D3+cY0RnnaK9Oc0ys3a21JFciMNbDm
Cg6flg/yTGk7Mh7kMMXp4BapOra269VSKnxTABOlri6qIitPujU1oP5FrZunMv1xE4GOKHydDWW1
oymcrSLMxaz8jWftbD/aajn2UJ7LSo/Gm4wQVZMLA0echSMyTu0KjTi1Ksr866eEWVQ64CIqsfJo
ROtT8DxVy/ql/BO+GNs8YOJ+jfxjVGQLYq9vR12JX/sswgtYpxK/ABu/XdvplUcR975p62G8JEAi
V9PBeTH5rTma6X35sJ6qbTbINzTv9faAum7vVhvDv4jJQ9BMEkGwiHRgCdgFqCTO1G2+XRTGGI4i
HI5pclIbXicOacrZRfUMITtT/gv1mZdS5yVw9vvitNhm/80ZLdsXTDWIJUI4DyySH8c0EnzY6qxe
bjiqAu4mRiCnf1Iis3YssCktaDM7cuiBAnNSEA/YvRBdIx0l2pXguNHkURWCXl3RQnozgeFqye0V
nubUspjEu0SrQz3LzjuQ7JLxZvIuaSIX33SOiTLhOxUsRd7h8HCplSsDWM50PFCfkGTz8yloZVVs
mX3TGTmpEUkUNN3dLDBaACDPvjh7X4y8i+ECFj7fxSRiN1gEFG6zMvNkf4NDs/4cW4SD9rXYfGIc
jN/oHzr2MHtdrSfdfAvE+9UDfbgmYsqKFEfwwYr8wT6fWuc0dMh0rE43b/MPh9OxPqCftz7YKn4H
ZqeEsExQ8ZAu/MaxkqviUpRvFnAWmqiZ8uLLV+lba2kYbC9ws59YHtrmErUhwZc3cHCGgWvIShyu
gAjpaTRq+Nql9xomecHCuSU8t2Pxfy8sWEhQtmckcA9YdI+HLUncY0uQ9GmDEvzVVQ0pxwRbqXUo
fvnswxCf8+TFOPviSgBHl1Iqcz+REUuLuZag04O/zhwpY7azsICmQwR6ET0wzqd6iYjmiu9fDGzs
8NigFlUmMX8TqwYQDe8dPnQt0aPkrh7hDfjj5NL9Dk2WuNiJb518UTpJXP+uxhSy38+X09/VaGPo
o1I1balQQ+ubE2pI0FKZsVUqnlMU8ACXMCWMP9Jca/NkE0k4gJTxKouSomEaQ2DWLnccVGK0BFfu
PicxpIaLhX3htS2s5zVHkvzbn4W1nvqicurmCLfJebG8+lwhPUdOyAq0k7OXy466c6vpXWsMI5k4
0a5VebLXMBLCz1/FtFP3BO/mBcPuTJZKVMvM/pXp3lcf52H5RfD3tV6TVTRj2RnfAesW1tEZkbit
KWvoPoJfPjsYP+86GH71ppH3nvHYfoxb2J6GWF+qTxbMQSlDFjE6Sfh4DPQY4LfEQP3Ez75UL5W9
rQoItk/pB0wWaCkinXOKUT1c33z0+dSH6eN1ZN6HqFnbHoF4qUkxErFjfqCP4nAk5em5xG7fOEZf
jMaW23VJZy5cCrBW7sC0M1n9ABzVAAmST50QBJ/+kkfuc/qrYBNmUDz6ZcAQBeZ07EEUOmhI2cjR
UpdCEE6/rPQuR+EoF931G2WtzFwdkTEEEk/IkY6RwzQ8eg312Olv888XdYayBOAdNu1fZc6A6h1v
GJORmWHUMzlVUQ72Aa9UpK7Xrjbv80GrI/L9k3g3AM0eQBNQ/b/QuWbaxDd5qZKBZ5wBF/p1q4gW
wABA8t5qQctvPCp/VmQHJgwCfL9ptaOxH1mm5lBH5ZYIA6kuAW9u6Vi32ro3QzGWnTAuJPjVrQf7
7aUCf2n4rDLcMqadkTzRb8LJKFhMgw6WTW8ZyY38/mElkwpLzFe53lzTsDcnYISEjqo3im3Fv5Cs
KHMl4CwhuBPlvOZM88486IKzOD54yqdxlh5EiBRLsg2go9B1fXsQe55hjTpytJM/CCegT782WB83
lPoZ1J3aL87El/iKqnv9PA/QvWsK9ogW5kxWdgZxllU0gLEKiFeEEGY8ZzAxKfeUhs8eD8ioY74K
7m950PioFyDwikPO57Noc29AFAQIOO6k7M4nmARjHnpzNJ8Sj2//vPRA2+ZAZl2Mh12h4Ig57HqI
pnkeEfZNzQX2QAoBgAWy5QwFUHWUM+3sxoHhhhJoX7x5QcByr+aITdi0JN/MuwBM7y/2P8jUNb8j
w9iW5qOv7IkVbC2MWKO7d3DcrF2bbYpsnIm+bCttfpFa59O23R010LiClaH2gF9W/Eszj/fBExJw
/HFBsH5ZBXO8RwfdIwGhY+QibAQCiGVO63KLj08NanQXOp30ex//2CdERLaDuaKrPHhtqxNS5EYm
LUe/LbAVgr0cxsFRVOOX9V8YAEdJ6Tvq2ATEeW/vzZgtE/85dtvfQUsd6nMQKmmGzW6481Hmnbaa
LeKcGEb2C83Jl1x5Yvoxliap0gZySJMyoRTo4I/VhwmlbW8OU6Lv4h7kQ8SImtfHb1r9SlQ3M4bJ
dheBb3qYQpp5bGhKQXdSKBEzm2Cxya5Js7Shex+YoeUFzzYcojq3ocn7AefGW8gxzxLQO2t1xcX7
yjGRbM41D3GeQi7+KUnGMDp9Tqc0yXjoLrrhF4g/Y4RdAzPWnMxe6MiCV24auoFtK6UgChwbbjxd
OzIyYjj2kJAz/ndshpOnrMzKtuq1S5QZcv+3GqQCZ1IC7Jqog4gLb7/yaqSMwNj2nEdrKTc5e0I1
AoO3hcKfqsQiWzXMMOgakloZbY5GqpvvXEuyjlPdYkNOAk2R+urkTjSb54+xcAO1Qwd/v6lOXvay
eZqhL2Hh+Ar0nCFj0T5KZWhONJ+FryQvW5/0k6bqHKsX4mq2W2RlF/+EWhA/rasqoq/HgH6fpspe
Yor2/R1oWJhvAqAmGFTfZBoi56vcKGrCldEGB9QWf3eKUY4zhL4b3n+V7v9u70ZFBnrpBQS7PjGK
vQDWmGr4+v+q77AXCiKrNRXzegmmzEFtL0/JDEkvTACSFFRcGnWfW7F/DnWk0l0IoxPeTJb6woFy
uwcWfEqVRDfIjq48R+t26XaMkDsF4zLzERf4V2s86x023TvFJ5G16PvUhFyETey3e90Nlcz6FVVB
ckK59Sym3fNUSI71k1t6tY+jr99QsSz+Gb4aPhiFT7zxqkovqT3bAy0B/K1p0MBbdNNBSuZ962Ey
OIg+/X2ucm4d2gkK3fRvdHXIOXopR/xcL2sMPYRa3KHhYFZUUyHV/5UCxEQwRVKuSi0Eewntqdfr
O22bBNY1jUQ2J35Ve+pRHgtY2xqSf5tLIC65ZL8gmOUDQKVsE3oUfhLiQUV9V76oP/4HXo7O5xfu
CYMAAnVR2mG256KwLYYspqmOe/REj5WxU6iaIi4UJn0S4aebNJ4rWsWkwrnaBiu7HCF7ofbNYtbx
iOBhln6PCqS96SYCdAFwZAXJ91ZZvajeV3o2m35Afs10dZeyXTNh1+WKSXCNRud4Xnq6sn4Cm9Hr
ZlUe07oU83JlURImHswRAXy5B5GanOZ3+PpO46FGcWbPnu9RfBwn/PUSlIKYGAV3yjWuiRH4wvyN
D4Nb4JkPm34/RO8B12yYS0w7oOsGJ4A+J/00C3uTm3pcZ+z/7717mRAxtMCY1MvplfIGWhsvxxbo
LO27J0RjRpiRrO+Y6DAQ7vCNHUlFYJWf8s67K5trxPHhkX7RCZAx9eM3NwcX5wVf5Bsvqoqa9fN5
JuxAj6tDSsJyExKG8HfXJnm79nd989D2v5iX4wO5bERMaZw8hWloPbLNCEiG/aRkjhuR1gQ4celX
eMAPRqfApb49p/yMPYtWAvD+MJsgoymhyPg2yb6SDRN8auHhpap8XRBKggiHkQYrdIX3EmKw4e8r
EirqhQDH5h0kdhhgzQasuvvVd2NEyV2+6QboQVtQ+Z2KgmsY22gb0JGB72hjhbu4/ASfyr7h1xmS
V32LOoqWEqgOTb4Mx7ta4c24MXH4ugjWL9VKGJbOjtqKAHTQtIQhtGsnMWLvns7DJ5d7LK4QV25i
L/lsjCGwM/88hUPyDcetvuGDxtSZRU7fCNNHA8ibNCYRwnsiLfidE71JKnTOdQkIC2QuZE7an6eV
T7olbS82VKMX+pazbpNMlrMJnkdMd4DNA5oPVN0jSEEwcx3l1iOCMBwuYoSaj7SIeDFKfxHoLaIH
A0ynp+rLk73acFPTY91TZHfdEx0lJrnPkKfpkgPJVBhd56yLM4L0bOoP/2qJOKS3q3UC7MOCQ7vp
y/cZCyt6YVUH4N3rLOSsRpfI4eInvSVzFwod8EDc30GFpC/Kl2rJ2l2HC+1l64ipUr7BrTkEk9wP
wYKpqilIp1mkGw0bkr2/T3geLrJJ4jYam0uO2AvsgGbc98s1F4rie5TD/Cr/iQB2/SbO7xMlaC6R
9HHzKnuBBQVb/TD9SBIghC20AV+YZ9X2my1S6cJS7CllF438lf7Cq7zG5WXzWkeAqiequ+tHZ/07
nQwfvJ2RmcYyLoMoFr0N3PywO5cCEz6vo1yHnMU8Clw1g4Gm+6Jj/R770M+M9WiPNCt8oA1fhoz+
3hsXVKsLuym+dsNQPLK+wBQDN5puc4Vb6bUA0PLrB5GnwAILbqqzdZjlrxlu0956XXJCCxjgTBfj
ldaggss129J42F6WM9zW0DrIzFyKA1D2iRG8h1EAfdkNf3SdWis2oeHXw6NmxZad6KgSibMKkIJW
nLbIiC/gkHCD40gRs7Vb/sXWrDcrchnq0LIfG8XQFikHGhumSyNJcG+afIP1IvPxjaM9vZUCvah9
hyMazorgefFfMs176TNHi28AKfU41X4dP4LkzNMMfJmja4fSGhzlcYFVxBqPqC1cVNaTtqBa/glj
H9Qrd7Jks4UN/zC8FDAfZAxEeuFmk4JyBdGgWw/semJPta7+lwBz9rYIPAmsNL3BsnwPA5liDwyn
Vv5TZciRtNo79PaSZOifeVeGI0Mds6QWlsW64Cbxm54ui7H3KukKI+KRQXP5HeTmgQQjeda7r8jp
fgh9NlDrBsRGK9eEM2TSUKBypzaAEl3fI2pCMCeKSJ8/w6zrj4gMjLLNSNYFzJo6jeiGRMC46wLu
mmxikVF4DWfWwNzuJD4ldjzgmr1PIrPrN1uMXg4dmmWN+jlEypMeiHc62uVaxZXnbxXpcvPHF3Gm
foXD5Yf3D464xoXLuM3CKu4V/i50nr7sIAtN9kIUZZz8dJxMhSX8MSrBFuN/Va8qmODOpGlNwA6S
UdqHts3DbJIQCKfJOPqdSQ/QtrQ+9E1ix7qjr3qR9a67rzmuLmSFnRwumJlYG11vi6nm03V9vIak
+w9fEH2XimOXLjwwa3syvbUZDgYt2M/AO7whxf8kTZS2dVbobQe4MB0UtVulMyv+2blrU01LepUI
wNIjTc7lS4w1+r4EGaO1sGeGYVVjDdKsZmqA1T4/UacKJAkWXza6odES8Ew3KFFSsaSgrVo11xLE
c+Y8EhXyT7VXIR/xijX5h5WyjV8KUmvxZCB441hNRaZAbB2DO8ioUrdNCg3Ym5lomwK4mSunRwS4
eUJqlu0+YSl3DR9xbOaIDuMHqc2zWUOogLHPfCx9pSNy7mVnvJ/cxqLbzIaHE9+jzWalVdns+Uc2
HRUSPvKY9WKMnO9KqcW/LJUdbvCnXBd4BsTr5w3PT4v3BqKjIEuBkfb1fq+sTKlLyXZYVhKkuUHL
3sDXwNIifatv5FpsL8ZgMt/RrlSdCXc7/5641DxMguTpMT0xQG4MAJp0+JonXxXhHCAZGXiKLwhr
XXoFqM1m2JpBs0YMDkkfGaCOipDO0aiPefpiihdt6r5Gh3NkYfn7rDw3YCemckljhH5gYw1NdY/Y
x8cS/aTJ1jLiJxEjGQZpGfQ8vkj0PhRE4xQgL03pCnFCDaZWylcvdr3Ph1vC9eH/oJdPt5lBUBk5
Ivz8aL9Sr2vgSBSqCImuKUXsEsx7RxG41xGb0J7m1G6jRJ83LdhyXncHKAjYHqhRHKg6ssgoxy5U
Af7UD4xS1BhXDKXcuylqC7MgXIjPUvVunpW28NYET8/ANfV+HllwTTPJQdBqCJNyqB/VcMR8fF8R
zYGjQdtfZfXT2y8rtCrgRbKrSQ3hh9pCCfU271GySg1mpkftvw2lBsCgtGYyGKcGj35HVu+DE5KH
tzKsv8DBLQEDThkQkbJj/Yk4xc/k/DPh8xO0sA/XvnMNeXLLA0LooSCVC4v9Ai+0ercaRC3eHELI
zTEU91X6xPqjg/vvBTad2AVfLpcxNB8bSWNjA7ZsaH/fS4j6gycd+RLEusysnTHDvWXCroRyF3MJ
97tnFduMDfIdQ91kPmzz5Fc188Taw5Q7+0VOMJHKH88c7OlZ4DtktsMU5O/p4ognd8vzrAeZnTAZ
37ZA7zqKTYOt+1BfTp/V9ERvXQfj9OXuqRQSdtLSeJPkhotU4/QYi112QlwA/Jk5AoNyghrpps94
qrUtXiuqZePTp4gfLvDJ6BnVX7ah1DzV8e2/AdoQWxf596vbFSRvM15SO5rpPzSgHdACpGevkPmZ
Au1OBoxqM9C0QxHUzt7NB73onzXRRqzv3kDQVI63T4zIXXKVzdon+g8DxXIzIFAO6Q24VZL5aLWX
AJMP3+XiIoY/uxBVzvahVw/yHbFXa6cu43/vQNNAborZEGx8ttBlgtkgkGKiqr49bvzWC32i8yYv
S7FomRbQFDq0rW9crYyfIOMNJW4luxT+CjIUsdeP/umFMpdPbGuCetOl1UwBD+WaNEU2wyv4/NU7
PKh9WGwF0QkielEc1M2EPlGDI9GQ8qQAHZLGwL2foU/4nqSNczCgScUWW6WmfDvd7gycB9ZmByDk
+K/NI9Rf596DJ6hZnyC8JTAV4igYvrwDJp3Bot+RxAEXfZTgXmVI+gYbUPbCcPb5dy3KkBZha0vw
f/l+mRcgx0iw0qpi56kNCmCiefj9togbXWPC/+ZTUWG7FCSNSKM0jj9TtP96bZbJdGohMXLz9Zhi
d+toW5meS35dl3at8i6xnsrx2KdATq98gVfTsoqp79oiX/aFKI1nW9mSje8H1GNRKm7Rfz+pU5xy
cvRmRMkyQSrWUBqf2i8kN1oDE9ANukAyxyRyUuBgdxnhqc1f7OM9vLnkHbG4IePzK5M/ZF6Q62Cf
pTFAmh6AwDD+ZDy8JhKDXJz3kY4EvLJZRlFbCiuBx6lCJY6M6IZ8eKGrG+or4LzRd2iv9AEXl93A
irRLW6MUPUCIpkaMWPtNME1M/025Vc4brBtOw8RvEXw8NivJZYg17LHX3cRnGlta470ph7sanXMR
83+UEYUgIPNTQYTOQPT88FLm4pt2VTHQCwkWE6LcwemzDluigFBgLy6I0myo/y4K5S0CtfO5yIUO
HNlIxeuL2PJcqWhwsCrANQsqZmwaleMdePawIUj0hs7F7GIf3yJClBQs8izrLrrhdLc99JGB15sA
+XoJmF0FLeQ9kEDesTXD6BwCZwblqheHLMMp3v6hgEIC5lrvLRD0wj3g3QjbJYvBDnOgHlo5y0nL
vtNnwaJVfG+cTiD0FF1ZT56lNy4eKjU+5YohPPxIZSBOvX9Ql8bkpYHNSCNAZQgokimAWeLHfx6S
ar5MjKvSWXvZRF2oCEXGH2yuivL0z3UVTBPGlAGnbt+lVgdxTD45hvcS9iOSSgeSWr8g+J7Le+NT
/Q31o2ryEHvzHRBySX0FoFw6FJWu3D/rEgpYEKlrMtNt6XYiLNQQ76tplzU7BPJpRK8pJZyBnP2M
NFaDnkkWVqkMyjQdWr7fWM/SgdC+aCpr+L0wCzuNhbU/1W57LWqF+MFtb/u9zQzH3aTrtoCVGowM
4SslB/lHABOrht0/zUfRSGOdxRLoyaJHTkhb+KgqJKKe1e4WxL7oHxvwzIW1jPeWvoQUKfl4D1Nk
gZnle43GXF/GpzRrobflJ3YOlcauTM2a0iii++tb7z6rf72ntJbW90GxlC381aYT6+LhEdPdSTMy
eAjG2BpXYSqzmGrIAyRK6N2SO73QeRST3x8k8txXpaStgtCtrbPhFyDbgphZQ9RyzFUUumLRvu4W
2mByz2zLV0iYOBhLcawMfMkG0bVIu3aRns7PBXVqf3euO4ESrjSbATpAptBx2aPcdAY5RMeRSNsk
VpKKBYfm2u94rXKQbIFeaol+LIN5SEc7KoKc3LyU/Cqo0em22Ml1Wwi4bdrM8DEky76PZuBYhsjk
DicWtcCbNJzhhGG4e2GOe0NBj5sAjQf5SUK6uWsw4WmrCYH6daU0CmToTkZPiCrkCLiHIqZxuqBy
/H0XgLydE9MEjAwtmgH5vh2NiOPY6D6ASVaUlsxbrhtWKqmANMigEG8zGqhc/bMqQSVwQTBfzIaI
noMpwbWVWrwYANOagFRwzGOAFjR/RV5VBC2pVVm2WpQwVFp9G9/He3iiaDqAX8ucwuvTH/Kw1bv/
RqPYr04uxeDBohmfjaJtuBrpJGgd+EggGJktYSSAUfJM8HqbQBDtgcrK4stn8erNLv8qQPQmDir9
+9Xsij0hAHEBSA4IEN7ZjFxLerBdCGQSoqjM7dHZreisc/ktcfBHHS8vuMVeWs1bwrLx0nlkpYX1
Cap1N7R0tCQjkSQ2tlta/z1CEZVbX/RuCinv4W0UUWKY62Q+Fy+4zKDhx9nj1GRPAVZXCimhztUi
qnclHb8bqzoo+ng943Bbc3hEGxf9da7CbR0qta0k03v9Up/tfdNCIq/8U5k/TAi8ny/5RWtFnBcp
c7HWBMfKGv4mDS/six6SmxcVyD7DPcdSHFxIvqUcaIjVe0xEJVmp8scF1hpSsxSbVmyKnnlHMp1R
INco6eQrqtv9T8AYcgIO/ez4LdBpbTgaZ5sgK26nPsmHp3RjB3Zi5UszQKFSikEdHK2lE8F2+5+3
dUUJ0a7Irwqby3Vn7orglYP/OH08IQAFn16cD4Mgh/+lUo/p1vE69vjxI9tyyI9WTGNIewnGHCv7
6sI5eDfl6RPAEkOaidFXT1T7VI25ZqIoGqqePlsbpGxCQOq7201h4g54O6lrrC/2urbHXAKb6iyN
qm7/wLIhLR0Uvj2Uq6w3ZcX+qjiENJSUoPUde1ENbcToqgZZU3vk9pORAvnt/ztQYfE/l8ulSGHA
/JdeGt2q3jj3fuWpGnRiLaqFci46Ps1XlmARfEc25VNXsZ7Y9q4QiRsQX5ziX7FEiDZqNpfVuQsI
yXU6H/rgRQOUto3P/dhWI5Zexsx9694bfpHFp2KegyzZpSny05B+8R8z3ovjRaGSx4+u/DdwDOwH
BAZGCD8S4mNz9TmhJoN9c0PppP+8u5R/3AmZItftTGrHgtrqOed9ciFDZEB8N/Cf+1RJHCu8PCKg
nsGXR3Qhsw9alZfYVO7viImB587BiNO5tMpXKvQ8jhLcNLGXdQPjZVpledWAOQ91e71h7bA4jAR9
eqrByhIvmCPFlntqBCHPW1Vc/Reb0ob2ItHZ8Q23QumX19X7AjcAAPnt0qMmDIDuUAJNEwTRoHfr
qR2qNhbxIadw/QjPDkAL6YwEU0wQlhtQaYdxsu8MHhMcScTKS8HVtaJuJBuZni3djTOo+kDCM9Vm
fjm9CGi0WnoTu+oZjPhCTJNMF4EnwnAVCbVfZV7s9DBnYDNhibQk2OEqmps64TPaEYh+Ffh5Ddfs
4EWP/clOOGgf1nHxK9RyGuJxxHGucCxXjm12KEw8s2nkRw2D1Wcx79QnLNXo/8YizHcyaL+eHwez
q20GNKviDSaRfiJGyaggz1PVvnFw3q3qIwASu6kKwdVnrntni/TI69OtEsOenMFlEUFDtYEGeXb9
Hjs/i/NSGrdecDVKm5z4uAniK5mLoo5FeP7pD1mTojRevORMQnLOgKMI5lGeIKcMG/UF1ObXGu7o
LG24Z5nY28fhoH8/6KpcIMDWhI2Lnpe9ZTdQlq1L06x26UoSsgT7FJw50wMTBnxGco20MAwUhf7Q
7J9cZU7v34T3AxeT5ssGjnzN7YkWS4ASa0eaBr/6bEuM+Wa8ftrxjNi/++YCCg5YwCRrRBT6VMUH
Tev3siVMp0kYl6g+hkxEu3uz04qBvMRJosrYFpJeLH3sg5fO032OVON5Ud7ZD5qIR/4goK1+LXem
r8VtpQO6CKFjYyA80NGtCW9diKBwcSc7AByp7d/4pvKTErujnOj2neC/udCKCboRBpjxBuO8deVg
jpFHGnzDOtxl0aTpxb4UAQUm72eZBD8rQ2vgkClSfL8RFpKLF6SCrTS8u79K09C+PmCLuEu5CMz3
2jI3oAskl6Jz5v62tZrqbB2qRSn4h66Za3BZWDLwfWth+yjSP0JoFgThfvQvW8AJFkeYmjln3ADW
quNQvQjji518ApDffvc/ppYaZJHnNxAi0stkiwJFD4Y4GQtsa40Lfzu2DmAk861Tg++LLVR8KmWE
Cg9nMkbVaNgFSET2unbvw9SJEkflFR0Z0F0qOh04NMzOll5C3Ag69yEhehkQupE2JCT+BRu0aXLD
9yuMFzJfkJS+nn9ErFNpO5k/tjDA1V5Y162NFw+ChojqcYNEKT6EYTYev9xFdLt+J5niz4zBo8ga
6ByOfcO9q5iNnoTsnI9qMOHQFJzxOFMaan4CespdAr2+YDiNIyJyhy94taWmsAUJ8edIfGUi8Nro
bN9Sxqz0M5dGnF7sT24SIgF58UYRMKsjNqDMenAxWVPHgmdleUd6y1S+aVqdd5Xz1GvSCs8D6Nq+
nRzZz36SfFKGUYrCXdv52tMS7GDDDC+lZ9MHRfjjtC09jt0KUOilPqrQTkRT/1g2nhfPepf3kYtD
DTt06xziVKqTlJYC10tVnP2W/iwFnhoYhad3tEloQWalwXFO9GhYrDM6qCX0HkkiC/zPiJSTyI3Q
3Kpb3nFfIzqsyVT/lZrO60nmqswjZPb6Q6hqbGK7TlR41THg+N5SMSuRfTz0qrkrz/i69QYMO4E5
TMA1C3D6/QDwFzKrivD5t6avwmlQJF573jkJHxMZjfTIZWTLqaCfb/jaZsUmEahFlJZcuK7BIak0
rH6A+HwALzUBkZP1Xi8wqJ9Li445UrJ47fe4CblfjosKLYMU7Ew/5FIio6Lfl+06mDPyd7dgcMTy
5O+t6s2/w4EtPXNrc3qOUlaW+3Ul1PpYeEpfZxoQ01TaRBbXbk8bBVfULLUwVsGD8Aa08DVRfBs0
ddkR9qKpgLWhTFNkHqJ2yQr0z//UJc6VV8TscAIiF1ZHtjQDMV37tTKGSYTQXUxc4SE2d8X46wZu
fC9NHh423h+j0AR2ZptZVH4yVoxP2ZvwL7QTrDVWkTy0qogXWbBleO5if1Y1ZQ8AC/Bc+8kIOwuK
G4nO/sfOWsVlP6hQP0MlhBz5iDL5BktY83QD/h5dCmXqJ2oLWC7OD6XTktS0eG4k5LVLd9wITmgN
jpGcer1dtOoOihjy4JfZKDHLuomiHPcfsd32uiSxIqkjef64NABFNmzuIxyEuRLurfxtv8wXMpDy
PPGTdvh1Xtr2OHN2AxzEax9BY0DpCEyL/kvB7f6pg+oDuF8BEmwbRWhcOCFE8AhtFuvbTx0bbaIT
q7bKlYW90Zk1yUei1+DycI/KwuBexnOA2DNIfI3UzqG247oXERYRMc7ki/b5Pctq+uFK1Mcd5dDA
WPnNVZbRfFWWES8/D7sY2AjX0uN9S6RPuHOc41ou7TsM8V3hjxXhsmuzr0T9ReSL6U8031Gv7sXJ
bDVWiirb3S1aS46LCLcii2PQKPPzW5NFKRkMaWiBfsiPxAH1GZHuDjQkOzcg/eCZAK0Q0SrKvL2c
gx3UGxQeiXDENNbuPAy+6xk8o9WrkE7UAmjnMJrdtHvv9KEwDBKItcuf7nVLfolJBOfzUFpzyboG
5ERDVLxrcLK5lHjF7fe95sc31yD5Q4LIBrmFMIIVcA6Ur+BlMCaOernZjobkPqRLtab/fa/Bbzfa
X/eQESqvMkLv4JbCZ+waeT66kyK4rkMbdkFTbYJ84+eGhNK5YLuvsalQd2vYP/Kyk7ZQhM2G5wLd
f6LbYjK/KWQqctMrghe7bBPQkHzQFrc8pPERC/n9pCLSI+qZNZOXKXMXQZ7lyfONl4DvZWV8GvRB
OARQfUAp1UxpAnyJ6JpdPG+7GZ+ooNqv92mG1B/Q4XQFIevJ79JaUtoi9ijaJZvXD584x9xkDgRZ
56KA0ji6NqhmIoYkfXruD9iIjAU5ZOJNBHDd5cMsAt+a+Abg2V5Uh4HhsWsd0XoKcNAggs/i7zxC
M0JrY2fwGFoZRsEM5kGgerQdLJDvPJwrum4vqQx24Dh+P5TgwA/CiB+bovojx37jWVdDPjyP2sDH
cmjLb+J/43K5pX9gL/IhD/KGYXT6AFuqpshyCEOEK+YnaDAIYJL+0CwWe8uF0y3/qmYiM5pvWdnQ
8YVTDAhz34prtNAVZAwXn5gBKWJYAD3+6ClCjErM496x6M7p3Pmh2hnoxmNLB4BDz0dsB/GgNIiP
V7kYLuHZKTW2jL1aPk8SQVCeIVRH3LOjfgofWoga1i+bG+2vCmKkx/jSiHf8MssQFF2l1t9dSKNp
6zSsSE3iqJyet5Nyppg70o0j2TnS5zltFlLZc0nSHvExxDL99DxAZL4tsO1gRQpxJ5khdafsHxXG
SYiPt7XaWsQsfns3LzNiCNwHkC0kUb/3EEdKoIk7eSoFn8JrIaGnnqPv/aTQmP4PrXVL/hjfKgKY
J4w0fdU3UgoAp+N933XDxDKtb2uLnwJbw+37qSqrQx4/B/rho9YarujqYU+0/B31tf4kUHknTpXh
yC10/4ue7lrY5Tj5Z6fegq+8gURLMwM8xUE1rcLeRzNYawsmkX15xJUR5nWm5FUuuOQxqyyFTuYA
FhalvjLQxxGM6zSoV+O4U+CsxDt81apgfRi0rYHVgAgZApiCpVV4REo+MAHZU96KpOXeeTUnnXzU
P7s0oavsI3nWMhOjd2M8Q40rYHsHqx6AySJsY0w06Kp7PHLpIm5hMBaOFjHCMoMav9RNJsFaAS7l
ulhmpjeqMj+xh4HCh30Ih+tkbC2S1NsCxnlZQN3eXFyjIUbz5d56+cCY+iNVL/XN3ZUpzLAZfYhY
K2Ngvd1r3tr2fs5kqzKDnPhk4EbIgkExurHJGjMaVoEA45oA87rsLHvLNh0msppuf6s84mJGtDYh
cwe2FlyWMhy0Juqw3V62G7+hAW+PhUmaFWYm4CbQ8TfEoACu4rTd3E7aYolLQZGj+oe2NQ7yxlYT
fAdvxD1yc053KYcRNQdPW1Miwtx7PWkrSfzJLS4IwqO802NuYyKcuYMOHjMcTfAacfIGxc2XI1Nd
QijUCUweNDDmsWqjC2A2DQ1nvicc2/8SzVO214PCEUiSPByosuEPUFX4KNmXEvEddeGdZsereOLp
/kbxj/fXYW+S/dBeP4mubiTl2coKjYsZ/ZNQD1tOJ/KC8FyOA75EMM3QDP3oQNUwNaa5Ku8HJEBZ
CbALCli34wUpSASYkVi29rBLGBJQmZmzBofFEwGO3e65d6YsgAZZtgZ9P5jT9qbnysXgM3a0BBi8
Zn17srAQT6s8j974Iq7EyROFtDqU/nw69jGNBLa+Otjqj2apa8jmq1HcvTV8kCzuhgJc97qvkSzQ
FLuyrTQoD/mrG1tFOSe22mrxHHTT2PoQR3tlwVZ4E4/Fqs5t4EWtcGuRm2lLyFV4LemV6INqupi8
GWhHws24U89+1rG85WFndzKjC1pFDJOl462gYhP3rnkzSQR5bEbvW3zRP/ly6jXHN9n+QJVy1Hyf
8DU4sqGS4N3jNJapGRm+w5B6cTcaveX1+Rc0CPwksAQGnivDeNd8wTaztPrxa17Mmgbj+l3Hq2Hk
2DIXN7wRxC9xuDUPlbYZwdJhoCi+zBqkxn3P7+ozQCuRGDNyFuUegi9pEbNewYm+GOTpMk1PUjgN
S+Sg/fvv7/ibQ3QIUxjyQf24NFFWikAcsOuwZGFZ2UHXzTfo6RXMdgpLzww739dCqSLIy7qjYWos
TvhReGhWaCPDl1yL48c58y9MyviaiMEFxsK/wAZreX3b+gFpecahy9OuRBoo2y7Fe6Zhzs4gQ/73
sdws00Pc1zT/nhIfGfNGwYh2Qx08oB9iyg6h6FjRw0JkKFapb8MsXzgX+vdorB1DNmaR9tjt6LOE
xhLnzsXCLqgngHcwR9Lo310yqZH1EmbZCAiOa/rjsmjr+p5nEGcOWQdY2pP06BgqYgYqrVpAAgdQ
3VbzQSQFB8PrJps/GIVS7AQRM4IO3cNWwrTgp0Vvdn3z3B31rm+adlGRe8WtvoCPFNvQIT6DjFrb
Cjpx5rcVHBpHjIdkSAYVn9ULQ3Vxb+NoONrXmAqApMDDH5vPvEXOx0HK0v/Gubhg306i8fRSZBmr
q5MOHOeOUPHcQOEuMZATdCBJst2oua1oe3u7gCFV9fCOZkorywRiqbQsHsd+sPSg18tCzUdKibB+
aLEX8wqCDletEgRUvQFnClEBnIkKT5Pu6r3FaYsE/mRCccXSbqgxBKbvtyhPO0mMIFRqS3EqffbA
FzR2NRizXOJDaHk93VJicMud0RKUlcRkN3vp3yqNyiL6ijALGzGEXqpxliOvjuom+tdl/PH/WSyh
G9hEDvjbg2k/HfixZlrLi9ahKTqiDB+SkXuvL39wiudLuDQSuJ9KhXFfdr0aipcOtlBsJg2Z7j+8
BsucSvU0wKuAz9Vf5Jx90O0nj/nS2TVEhFw0uk3B0pVTPtWvqiANPiaZyj3fpQ+sIEA58ZtsLXQF
dh9hh/+Ro50HxXP1inbl7rlBUTqrqbVAfPYbk+vib5yz3zk3HvhFM7+QbUjMSTYCtLdA07frfUQM
IMFDrj6LNtD1ixWsxFt0hvOXp2GwTFW8IaPriSGBaa6xqfULtV3od5/Rgnk/iZJ3REAnDL6nJFxi
9xvN5RZ8a4Uwz0ZpFUzJCu97xFA+ySXKDvRFjEfWYA4fEUTOayRyLQrDZfZjXkRcES5AqzCMTQWA
oZzvIBHQUY3nWYdOwER2fCv2nKo6+fOdFP79rahavGpwhlSYA4ekmPNHuE25q3xh3Kphs1q/ZTi8
nUxjKv76GEAmDlpsBvda5g7snkNrm9k/DntRycfhXZGDGRBwW5vW4Eo58lKceK4owC4sy/0k8gZT
OU9z3b9EqhLyVJxGTm+4gZeW96oeP4hDBQCIN0+AmMIXPejYwAD0GxNtghxfV21MxVvBq2OfqSB5
sN0sDUQ1R2FC35+cQOtN2SQ0ROWfpHjQw2pAHqZcRkbqrDUyONtr7AjVM55gGYNE5wYEDLvwbOMo
czU/p5glIPvWlqPp2z7gC9herAbmzruSVveswg2isNMmhj5S634Ng0+lczWcLzH5dPyFhnoRQLln
VYPBgKI0q2gaw72+/b9mKOO7FxFMYslDw/LcVonVyYOR4wrd27Y12gKvcFtfgNSN5xlNtMIbj2rZ
8U5u8Cs4GfknkFMKFeBuZgd6SHWhVWfKsu3fnSFH8hSR9y7o+djItdufianCwBBWmkWRfBRiSTxX
YR+LNlLw4VNWBtkDKiR/pQPzzL2pVnFDzjGIB+c7fJ5W1CzLsYtSi8ctr6JeOEyXOLtfZIcbOkin
DYoo/Eb4ZWSCltamtRJv7mY7Y90zL97iG07zdftvsc3e6MeDHaOpABUdtDYr3QYHYhO9q6qxx9sk
jEGMy6AdIzzV3fPv0dx3SWF/w6mJXerPXmBVBM7XePdnGL/3YdO6looxBXPgSEQa2fkAcL/ONNyC
EygkvEPt6CtSA8/efpHXwkzl1Eh6dFhLBdHLMUrHAEfDbwBBLtODs2g5ow4eCiZ6XuYOaii9Thp4
Bl53ehoggqfFZeZliNlRmjJkQvSEIdI3AzXIrqcfU/kEmQtpZ1kX00AnYqTx1c7epr5D6J+KXErL
zr7NfCyB5I/jFx9Ge96xRcJFqE4/AtB6Nm8lIVjDv4v30u0rYdp+uLEwE001H6f5ne/gNllZFjC0
utGAx84qhp3A/ziZUBDvAtsoS9XF++GhWHqdbQC3miODVwTR78KH/2lsfNd9JGSrHISJz7dAYlUD
HwDOkrH7Gs9A3h44t6jhxU0iaa2OJVXmzkwG0RrysNOTR/VEYFEl7JFpaDBsufthw1P0lxrRrmTd
Xk+T/E+ecQt5i/z/3z+0kVdpayZtxh2wRvsln1hR4m9N9xCcgpcGccKl3WIs9PUcDWvsZ2qjmu5u
U2fga8SnKOlh5GhwLe80N0jfKh8/qs3CGg95Pavix/DmQvDhlalbhyrxZXfMXO34jaTuVN1R6cw3
nJ6PM3joTubvWWj2Sh5DK5gMKVfqCuDcLjheVo3dN+dcyOk3MBZBo3BSvG+Hxw+2Tov22RNqJp9U
HLm21EZBw3gwGKwFAYvm57xWSGzzgGfeWrimKl/2TWzeKDyI/d0XdFJvHAU7ZTSDqcsawN2VT4D8
pgZDYFdxF0R6iYVkJum9L8a8JzacXA8r5paO8WysVz4IbWfarB4IoHlLV4lcq9ovE0keS5FELwx9
lwmq0j9cR9vXAsJdbZKKgJtWpjGnP1dP1ZXHx/+iCdhPAVTtxdSdJosjpvoiiQ6GJorvVZ5Sb2mv
GdIRtOHziSxeX065mqdVMXwcZFXG0EsKEVo4/aDHrU5qMifgOYjaJD1yfkcNfBKHdm28qECHtLTr
QmNZOOm96ykCrK7q/OK+xNrhn5YwIYcgJNTwQn7pUMOxCPfoSXuPaEQTUY4dHIvugTaY8elqWtF3
4lD81DOu9hVwoVqu+0S2E5w78umD4/zEOxco419yPOZOE0jmeBLOKs0di17yIS4AB4ixs7Tf2JGj
pTVpcLIhXPu5k925aL+2T1vp8oM7ombzw80IgRYxXjlK/BjgEJoRO99/vzk5CJjz1goRvMKnAvUX
4gCsKPvLyF1nfjRBuilwYvhGsaWiZMfFDQQMeedmZ5lWF1WS1GsrqgubQGXyBbMtFMPXKyrXj0uM
pqrzN2xUPbvLggxqrmGQkc7EZn1kWXYiKWCZNvmBMmA0MP9WpW61V6ax3sZXN93Cgv/0ZPXWaoR6
9TGcBFsF77duURzdf1/AGnyBqjos/r+CMZvyQsnHb8GlAS8x8tifhsfL8VdByPGVajFp+b2IbFoD
WxRR/wJB5Rqi9nHpOQr3Nx8EeO/B/E9/pOzltNivQABb7223SasBFQjjR+Fgz/RHXwMHN3o0OXPv
vU4TuacgxddLmVZJR0KnvvK5TtGtjZJOhiwbGwf8L0ZL4j822YwS5/u8Oss4vOir2/4vUWpbScbY
ZexxGoY8h4nZpXC3FajrRBzBkzFOiGSFRHnYEuSn6wOCel4wzEsK3KlpPpHkQhyp6ZDsYZ79FeLG
qk1ockRVeKu9I9KYnjnPQ7vtJGMdkYgdYOC6d9eOtQ8jWg7AkKNzFJp49tfXXygjsGS95Obex7EL
ZMKjiWXwUZF1TnUdw8cMLZRlDgW2YM6eLxC6DuuwhJ2xMQY2dpNSLajlgigOPLEX1t3qX2/rdNbd
VuMQiTK+7X/btPqs+JDmITV7J7E16tCHRvNWY2Z6t89dqBwxMUkcFwGW3gqtfs2v4u9WYLglV8YW
feRMGqLiyYh2jgZ81PswkdJNLw+Ra4ZJKl0FW/jR0D5h6DDqDpv/U/UeyLjGxB2vbCJr6aXYnkb8
GHd1U93okxITiIaaC1M6+5KhCpHe/OKxVjU3IXOfxrNPDu+1iUNxRIO28pb7BoOdLicZVSc2MN0W
byVd1C3WQkHEDkwQ0bRK7Q9bqWFe98yADErfVYXUID3rfdvrahb5vyyuJ3V8nddvnwCgIXg+In0y
BexJO4LH2nV8GwKlLQh7K/QW3/bbh9GVwgw5FGu4nXq54j9/tLNSUosBYuiH08R60iIZw2dXTcSz
g0Ago6YBeOjqN+lXHMv2vaxvTXj2RL8zPgn5LQzOGwh0l+b3VUeQzMk5K00HM4UMNLdQ6fGEUG+Q
U7Om181nrrgp3jvSmcsIXEN6+MC9CormHui/XKm+0sJRifaTIcLJBLKByKiZz/f7bwruBeaS3qpo
tC8DqbeN9GT32V8kJqm3lf1KUR47bQTLyCIE202ZFVh4AB5285b5hlbXYU0wJ/46N7b7J8p0ahiP
i+LJ6poQHspHWxfWoq9vCmkD3f4AnFNFPHVCLXQduoFvoS1TNulAxMtu1mAG5vSlWdi08R0nhjb4
C2N6vraAIRzjO+cdCB0z5hMLWINFJP1elmxxMSSrmtuCM/R6myjWEsWtSQUB5QdhMSMoR7MJjMCQ
aObWEyeJGpLifGtAMAHpxsNWT8GCRvPojWfQrE01pm7XSlDQnantH3Ea2BB1W81YHBaldeZhMm/B
1LSzHfrf+t4QSX4ISxbRuor3W0mZf3TfUPAhKFTSLu0Q4xxqeYcngSZYtlMKST3HJFlzEMB+IzhH
em7HVoS/tb9BuHoST1F6BaXDGp8p22dD8INKhdk6gOZzqyw9qQZv9oNgLdbaIJzFdx5ID/erBkf6
m+4tj5o//QbJfSYHg9LWU6gxftEzNWMFoxa44jjU8BoSVSbm9erRwELOE2SmoQU9lggHSx3aI0RH
++m9GMeuyxtvlwPY6aUkGeE9ecJz8aMQMkCOpGBV9i5t/Y14mgEWc1m6V0/E/f2+WOHNhPrWpyuL
OwZROFJbk3vJMH7nBrRrvuGoFQypSQY4OzJxhMWZDNEg4pVwdGTvzIDJ5oceWO91/OLHUxHQfOoV
yP4XXNiYx3m2X9pdRcsrIGXev1B+azuSfTKYn9eTXfV7R4hBso4LPOg2N5Wxar9LXOSFqrrHxh+A
rjsK7GdgozjNGFcBX27/GR7WsEw4Qrjs5uxThKlaqmQ19IncABaybbUglxSBslqu17EaRc04tJwb
NhM5WmzvjkxsFUi1Wr9ueuREzxXng3VsDvDMp8VD5rP1vx8f+8yv3FWG/Gw8PKhv/3Mx4F2FuQA8
lIvwthvv6a/MPxCkliEN/m5aZLWmLU7ezFc67Sa3VtbFXDVnXaFZ353X6879oJ4QJDNKHvPrWh90
J2KqqSqb4h9IvcgHXDP9FvAZATbxZ1eleKNnUFi6ylOzew96rgLdVbIpeFj5Y/bcX9FDdQKE3KdH
aZwX8ZbrcLom9KkASuzmkNLLd4jtf1AtJ6Vt6v1E+93ZlzNwh/bQaD4E2w3RW+eGLkWWuoKIYXgz
P+Gb5Q0addaiDmyQ/TqqUY0PMw1HpJ/2oqj/WLQ6iHiUVXrF8mLg+J9CXRKK3dyMtPQKPII8/Wpo
5B9wE0QNQVZhH2zdfr7frpDFbofjY1Weg4qp6q+7i4/Cx20g7cKH3j8U+rpPNOCy6v4S6j+BD++F
FX49pHnq8STIvp05hrXI+y8/s1AED5Dko+gkKBbZVwuZsPwDKRZsG1wrk0ZJMKEB+ORjolIoIpDh
FBNIe1R1VN7zkmEH0Ck8dttr95KnKmkAOsAZDVj7AlTo7KoksfFMu9bs1HMXo1rizt9mhTCOuDns
XRaL5jBftHU6BM+qce9CTUPryyl3i6ri8IyZNwj/ngaadR8bEO9QGbHYKkCPAi+vI5yG9Njr1EwA
+tTW4TJTfZ9EsIU1tXnfJ5vLxQReembbWEmiR2ZUBqff9vG/CdsxX9lwIN86T4V2n4+svH9FuyA0
BhWdQ3pC2PiTwx6BrGGAlLc4ns1JsTmiiCDfkd76gc45ocFsor0V8oUmsV8eGqoWOeLLe7wHqEak
CnF1fUpvC//czmgnTlRS9LoUeFap2MMJ8W0+Y728t1wMtih4uVwMvinunvWRUltKE4KmVIPAkMjO
XU++4uDHrIZtdpYHUloE2JzyG07r80DSK/H8RijN1POArhP5gMTSNgm9riJU2H+Gyx4wgNt1SCSu
R63Sld8TIAMy+6tsS1g2tFB6SRgNz97+ccZYHVJ3TAkkEGgz0dCSw2UMrDiJorHjLc+cqCajXsog
/n4W47BuyKXtyC8n9LuXLw7VmDO55Kh8qFsmDd4dAvl/SbImfl3l7lWMRvsxbV8moyn/DPIQgVdT
+6k8aQ0nYmdwe1IQ/mdFmRjbUNr5Fj1A0sz6ku6EMWtIlEHtL1ZOfJhJ1cuHes5V99mVtM10TJd7
oZNYyIOgMg8JmKaViuNJzkxdFkrFV8hPQ8gFcDjqOCHwOrR5yJPdJ+GBSm/ckpe/GAD/Kzmv4gW6
kX0zzHEYs5nDEn6TxiiYl2SOiifgycrw5v163UWoSKZrUNOaGAlokzegsqq4QWzT3NH3sYfaJVxG
quyQfcQHs6VC03/KtwySFU62YS2iHAKJSpeM4GCdMFCoY5qF/TzP/eozPwi7/fZWhVYc7g6flfcp
jJbwI6ezyFNyo04QQjyVZ5rFNGBJjoiAsW2MYpdAVGKi+IiAeo7JXIHacJlp7sg19Hc8sn5lCcGO
pvdKBZhwY9D5BvK3sgtHYZZ+3/Fyt/vTNRbMM2zNZcCioScOaEu9UGMYpzVfK1ShHVzEpadZUyAq
NlqpankYZE7tB4qYr1ilGvKLJPOEW6syuT3yzNACNiTTioxGpTaQyqMY+qBMWBocZq06dFMAWHmc
uMXORpjHCgRgMeFOgu18hHE/hBvnXDsN/XNc9RGP/tQ8epV5NytH5K/ifXcuoRXmD3S+Sw+zwuHJ
BCnqC6sUz/inEaprZmMR6wAOQqXGGT6CdVWWB33xQ+3UV9tggYpIdRNcE7Z55YpqEjBo/RpPFFlA
zoDYWsh/I1LZEBX4JLgm6HVxUQhg3vn0XMUaikBoMHU2PjL0tC5JaA216+LFYtBfMgZoJTxYDV03
PdHyOW/ZzrT+ptCPp9o5L9bVCQd+snF5bRHvwWXh/DU+xtX3B39gy1+0kb7KRIun1AHXqOt8eWC5
HY+XVfj9KYL2U01xxLlHXlNGZiru7sEHfJFpDzSJHIPuG2zBJLm4P+FMIb6QYgSIi88f8lAwgK1x
5UubTLX4BQwuG8PCN563FkOpbA/VGWin/Eeh+UhrmOdzt46YnXaO8ybZ59w1EvXXezUB9dG9/0+O
xZu9jzfJL/ltwQGvnmOFxXrgIIRrgl95TZGfcuSPhFuDXKVJZl9VCOmUO07aWDtHXo85aj6NBF3j
/zFXtz6DsZRPNjajbs5EJivdDqCT9TfKoV2HDds7dqds4A9L+Xw+NfT685Lern3J3Uky4NND4vrK
cdXPA2OHHD79UjzKAXjgsiJelKbl+5C4c2bnm3knQ+BYJ55jQDUQA4yPUtIVytDDIrHvUavyXT4S
G7mm8SRN7Sqr5X59hdZJGrsU9zmgMCeRUwbGsvnJpxhZ6endmG7/iQ3ZxK+AJz7stX/O8KgDgZox
Q9RwaYtsekmZTa7Px2RerdfEdrXuUlcSFaZyIoLeIjpoHOnIenbssEXlAQ6Hxl4LeS+oW2gHsjeF
K1iNXMHWWiviGrsHD62uVoJKOvNZhpofis/vLoP7GhT2CkdqOFnc/wjCiS1aoY7OxXCuRCeRlzT/
Gz0PoT64zJIwaHQmVPDFDs6iBblQcFQEa5YUyQvjXyzjYjWHd3d8ZWU8qA/gVp85dAFeD3L8GlQx
PB1mtSgFn3/kG2u7ToiuP4fULN7O6qJr4Ve28LElqC9oBmPUt6uto2p8MISSKXwWJLgN/3v8aT1y
EOsmeK4G91Nu6Ulx01pxYKJjCyFuihbL9U5rT6q0HiMOTiBlZo9alVIlxtjDAiTJmAWS9Ulu3d0r
jR0rWZBNQAVsgA/UW6H50HdgA331AUZN2JOps37GW75C8qtkCGSTfQIxqYvbupDbW/W+VWyon0GK
j5e2e/yxUUw4kLvzvRZIkavWKoxj+vpJGyPgUDvQtTt5jnoKAi8AgMsfq+Bl1Uekf7UK2SlHjrZd
4pN0+OA6FObVP03K8n5pNRD2AYP+KeqMvBjzatq+PDlwOKF/+U7wgu3mRwenVdu+Gv71iYzF+xNC
XasSu9HX/P7ZV0rzPWJPqT4oNqEoF12Vccu+n044NpSkJEo8JWZpToJcCzTRjGw2a01gJBxN9Hzp
/IRPAKxqYiRna+95E8c0s9RXrw58f4yf+eZsPqQ0mqcyQAobMZMGNYCkpP9DRRjpVor3MVH+B+cr
vPScgnw+IVBbNTnrtYDa7NolPs6bVnekG0BsKV1XjVyLCSW1D1fNJ2CfkWqeXU4Ga1ppKDHMbLxT
l+Mv1RysjXebknUo4BlHDcb29PzRR0g1j95vP+yJqRmUHorg7OH9ztgsIjtCV0Gd7/ipseU6KbSG
nTy0+JjiArtymsYnLGf1R9M9XDObJBg/VQlM3iMuYR4Qw3NRE0A/XidJh1wYeLyeU1DVP9Qq7LS2
ah9sN25uyuYMHMkQhEQ5xFleExXRVgCw6QA+4VReR3JIqo/s1QdqzUVCvvr6ka366ycGlhqGTlOY
perjUL0NqogIQUim4+7q4K2zJHs6O+XS5lIJBrOExIFrmVIBgsXlJSt1zxtH1+Ifd+aiJJ+RdCrO
1/qEssyUtBIQSKDb38o0DdMGNdpCVAkQob4WOvxVsJuo9+r3U/yfAT7SBW/OkUyQVf0jXRt6pFWl
4xn5b3ERop3LCkoW32yG37jW/xV4U2x49MkQlgqHUye+nJtTh5A6f5EE5lBRjAyfc8bccY5cE2i4
w1SvE4aeScJoIm/rHk//IIpdONSaTPOGBsMu81Lfuc4VcDrCzSxq1tqFGRivbJPZhSn/WRznfDZc
fFKCj/19vMX/wLTVHvEicZpmDJ8S3Z2j86dYMqQh31E8XOnfosUYfgj2M930WEvDvy76u3mNFo/L
MutaHCSQvxJJi/5xJAuRE8vCgaunkaYhsUiyjPGhYmdqAoMmu1PkhwtkxlM/n6wmMXnu1lHUj+rk
fVbtXMGmjgvgGtqmw/ohuIx3Tql7I6AkhUwKKfclr+2lRX16Qhac3k4BPEk2ELzJdBrMheKzSyAu
4F53+6F8kOKPzAdRmFLspAk/NVRXOpGd3uKnyLyfDa+K/Z/QbHZxbn/ItH7YaNykdxvjIl00ko9c
C6MTr6JqChrInYQW1T+aXqPz41xuEVkqccEXxkm/yiFll0dw6UY6rXWxDXaP2cvjCr/3b/bYAPRo
gPjH+uXxoBdXooQtk/WHHjQQPzjOvvuNq9k4mrmaBNxyyaMJiP+aka1XZNdFs8ulYTI+ymewg/91
QXUpiiOe6+JWBtpPjl8Rs7PDwUF2X+Wcn5OD9R+6jbb0zwak+PpW2ZkOf++b0lc3f09JZqjlDmEB
7jTvYsTehY7TkU4F1RagCjRKLnCWtL9GYEcvFLjcJZbEHYRPaX//3emIJ6M029MCX3RVDpJ932LG
dH5y30cyGQb8YcaUoL5zrytWm2X/tTO9X6u8I/RGLWr0IVmmldxcgJZrTOD6I6kAtV2Fs9ezZI7+
qaARthWQ6Pymhxd+zhMeerFMleeMEPA8ai59LQz+kRiQ2Cmegu6sj/2FcV23LDZzy9EKg/3LIRDF
yOomi8Y1M16nFADhr/AfMWX0Qu/iz3Of1DUjWbJJC1Dj5PX5fVCNxk8dfqlbxbsQMjfRrW+X75Tm
WiXW7gcvKolBRkdDIiZA9LvA+KM2WRdLi3+5BJphP/8sOFm9OBnAWUTqYO3EwVI79D0sL+5RlqW9
gyFlbl/oDtZPJceNLIpJi0mtIngAe2d2wV0Dbhz4i47Z3k+xxzAFRm7hDcxaIxIetsnMeLIPQHnv
R1iDwaYmJQwNpbCHP4DImOl4efLn3u3hRpWLZa1AGNjJo6xspfyFvDf2SOvLbqLODQkAHbZUypmZ
2/kYEZcAcIbnamWEmNtIzdJLMGjDMTKfItU1iEPK1DGTdrc6UD0uMhtaAdfVHP5XFY7Z19A5ReGB
Ss/KZIfdk/UKoTyvpVDPU/Amk78fRM/thcmuTN2vuH8Duo6Oo7aJgMleKdBixeY7XjhcMtBVcikq
aF97yWGiR+YRn/LEJqv3evDS+m/YN9n3jaWXglVkUBysJu/dN/VRacyRvM4XKoG4HEpxpLDAzy6X
ieHfnfbG7W9vFh8ingx6XXLS9bKjnLI/COAib9dTNYsiLrniouxekGBYvdssttcOwXOsDF1aqCjr
63P4YLYTJzLBmwTVr17ziAKDLl9nr6eSjRSwLFNWTOUkeU6DffJ9ATBe6up8wYCbPP1QTAsRzq8O
fJKRDS1qzlmN4p8Sj6D5vv45YOVQTnt3DOU/haeq0adkjBSB7ZD8wWQ764Iy4polYkVPUJWgBKi0
pJxuQdNk4e9c9Dse4n4ljmtF1vx+gS11vBZQOLN6eRASe52l3LmyvskPn4J2tVFYvZ374uIsLitU
lOGdApdNwqEzSOTyeszg86SFJ08B2LpTXbkwMESyBIdciS2Wc1+1q4H9Z7Na6xyY3hmRTtoTOqep
I7WOLYVzHi3SIlXxrJ9FUxtN+az/nxOD9e8TPTmZMRUM4qGXH8ZpJGCSoeGSeIVt1MR1qik3rNgj
xMTObpKR90uebMiYaPboOnAzLydMCT6VEacJX9oOtTGJ2QXA6fZNM9go7knoi+uo/jEqBrni3e9O
GW/sOzuUM+4HDeOSguYUjAzOtBi7exXkfccDFo7bb6J9np9n63DW/qL1GPWg5dFro5Ov0IrNup2w
RePxdlbN1WknM4JfiOrtg7W9J/pgv3otORk6JJOIKWyXeY6pDZF5DbUgbatw3UYO8Xgc4sPB5woG
kOLC0M04SZMLaXsV76H5mqTAZYPNZc+4hu/460iZ2zBiBE2TUsmJFoLj6K6YtihdYYjgHJKP8Vwg
zw7WfuVZCeRxSBK+/muDQFLNqH8xwpIL1NplQH7wiqxiUH3oqrkay385xjupa9077ikExeP33sF8
0x0cS/ik3kU9TZYuYJ4XjXvwrnWTCcl2gp31wA5TDHlMdxGj2JmLKZVaxjqeA95x04c6Fh+p+KKA
Lzzk8Z5b9X+kquqwjFlGVW+dNLxRX6EsCcpRJ56vloFsZIuXO2huARSO6Puyseh+Sq6YaJNzDiv1
AQeowroufwvW+p0MTgi9lQBCnScRk0Hl34YkpKT+/3bP8hiUbY6C9iGrkPg6wR3koNUgw7ZjviK0
B28dZ52+uqm2P6lLCm/vls0LykDM8igm2WNQcjWldVa6rMg2kzh+MSONu6338iCW2zqBnDU1mh4j
oR/vu3vF6QEMI6klstAUneHl+ulEK41QG1lxIiJ5N/rbNBF8IWAi/RDEF1sW/UTsyBvVnFhVwjmR
JJMWnqNNcDrK3HbKNQ4JULuBl1+U/PNJ5kJx2kmsYLB0i/V/7g/fmyR5GM/4zVcjSxICvvx9RzWH
Xx6Uq6Zm/iwT6gI+n3z9nAmyUOWBemFvPZzWyCjWH6g2SXglNflpHLe1GKze8G0EQhKpdF+nB+yS
Ws0wL5eWp3x47B0pgYEp110F118M//2Vt4BTMURl9df4gZoBS6OJq7SmWNI19u3H/RgUsCY929nL
WJbM6aShoQVGSxId+XcKkyzcfLuER5EcQ+SvouDlGVPWy+IMUXIokUPkPOA5Sr9XgWryakG8cJ0G
cRfiZc3Ad8ckcDwmHmaLgvV0DWFNXo4ByHRmQQ8yhx0Ud8e9lOQKZTz9gIxn4uMg/ggmMqvaB7G9
7sKuAAeWLr6ajZqsxwJTAWi0jTWHQZa94xRJ9YnSHjaKC/XNfPvflP5/SvLQMh2a4FgpPvqGTHLg
SS73DxHxDRIMEwvbg6pwXZaPRq/qy0MPV2pkSh7pplySTLHL1BO8JoSXiyhriH+iDlAKb6kp4f/F
/+89JTnm5Vr565UYX/963g210+GiwYKQOZU7VffvhWa5VDIYfj8+N5DwxBLnR1Lys3Q/aZXHqqwH
qVRJf5YJg3hbX0pRYs35qd5ZikOR7xUD23i2vUUOAuqy06TCOnjPBhzLA7dz8/9S3MRypZ0U9uht
qBvFvgad2ilsukCU5PioFEUu9iEYwzrdvcCHnomAV1hO6LBV8Y9jPRIpDl720RJ4o24kmee8aNTv
nEiagMkOZOKLqwWl9r0c8fYhwzR8Lg7p8FgvgEDC5/oP40FVB6M5XLDaqzvagWuGOq9pgqTSrKAn
ZxEiopDZmboT8fr1t/5TJ6WuVRy5tl1ZRG1XtSZl4cP7Zb63J7/UDjqFs5mUUESxBKPI0nm0ZYBj
lSlEOvTfi63upQOevrrxm/jji+DEWOx8q56GHFgJN4+k6bPafl+sIt5MA37cCBL9FMUjOCKqP99f
X6tbItL0Gw9N8tGpovWVlq8wq3DDM47lotsnI/n3JUqS1iJokzTjTAvwCSIhpW5MTn8cM6RJ/LnN
xMjYAW5pZpGln478hQyntItb2xN1h1aW8RqJsdYuN9hluF/SUjopKq59aoNdGoe/e1S0rJIjeU2z
RvUEZ9nB+2ZvT+Co0u71WsL7UsIpzWSGRzLCfTpyg6ezr0wiCvphztGTBsvON59dVhKarBbq4R0q
AqBSviwUk/E5iBwhIafND9GcPKkoeV94gvuKIDm2gnj1l7pVcnF/RzHgI2WuIKs1cYJcn5ogs/6H
8g5Ij+6YZOOctvRTX6yWid0enuDtk6e0fk68M9T9EORHqh+JInCjd7XWoWDgXhbSpNUCf3RUDlsH
92rCvIAjoRH6AdI1ahLsQN3lWi8XKXQ+6R/dmIu2L5Yb1jAJbI/hWGRuvP9oF7VidFjTtWSi9YMq
e0a2QPCM0tnlN+3m/MFg5iDtCuY7i8vfOsXyrJhCkH13c4GJ27+SDQzSderpqEftr3Px980aYG8l
LlA79ZdcQHSlVf4xxIyWF9iyScOT3V+WVMifAeWBd8ezAdAz6+v219vR/O4ur68wdhsG8WSEax+j
0fSMPpB8CLsK9s8SBS5+p2hwIaf12hSl1hKPDsM+oQ2FyCJ+LvSJTCU030TaVsGxpD4DO0PJ4LDa
gsO9Aw4fQ1N6kLxLzYhtZ3amtO8o9xrgn8KecgKJylWdHCPwjZrLA7lpu3fnSD8yeU60bgUbuOOe
KKZv/Q2BT9DnWBWLBne4p4Ptug+2DG1SUO1kGZowaRrCpJaBANPj0Jl1wPjYCw5Qj88b/PkgZWHn
kum+IWkxo9elft30SKEjRcFZNGKtooDLq+jBkHcQZ3tE1DkevrRJluhPiSfb0XqM4hFJdxoqQvJP
LIA5JZtCW3zfrU4aLw6bXBon7qeqA1gYGKUnzjfb+uUYDksCka0w6WsU8l0PDAjDRAxqVbXhsC3S
oTlYstAK3JTIo5SnqqCdJg6DfBnsAdUFMhGaX2wzn4p/Sn3Eco3KnTZsJ+E/t+RudEIvFemkwLtl
/ZgV0Z9aq/nj5VcairClHrqzQlYmqTYdmnWs/EN8Mh/gGftra0BamXt7KYpJjqUr0uf45aDt8Fp2
1SB0ghk8oBm20RJ3Co9b5m0FjBQ3JW2X4bicbDRgpvGUoqn/LUqeTyUkKMdDk3PnXLg0aGRYZ5/x
gef4sLMLB8bnfjhZ3FDGxZLEwqc4x2zVALfXj0NfPLsi6W1Us4WzS4uMk9Gimo4KmiMtceKPN333
+iPKZL5lqcSP3sgE8qUwpOnOBqMAoo9Yb8fSYHu0l6E6d0XDXWrawrY/p/nlCQKtESXR5hED6J+8
SICX7Jp8RPOv721G4qu8DiIHPvjOm3bF4q19p1ZmA7229ahFdYa/hvb/rO7PBpVqISdphQDPLw5a
8zIK2Tidzsej/Rh1P+khfCMlGEnNBSvXZ3nj5lLpPna6tSOJQFsCMgIy/6AFeKpAPFtkP+q26mPQ
wzSIEDNF3gqgXG9Ed2I/vFj8JthfxezjAdaQJKRhmcjlxZ22BzYKuciB1s8yVJNy7KlUvjjFej14
03TApfbu+22QVNafyGIL3v2Ts9X5tgWpskyFca/3Q99oWTJVUfxm6Wgud30USeK6MYuzPRwE1IkY
fgCRIMw30WOolh0D4TLxVnD0JHx0PwoTz7J6VqHbIq/zUnsgdxM03vexgmzkNUjVnWkPqHJvShiV
aIj0yBqEHl1lkw7qA24rjrCGOwcUzgcpPrtBqvofc+/FNC0U6tYXbybDgM1h0cj4GF+GcrPtevhG
bHGcl7tEPco08ekvWwVQyox5Y/baZvbQQT4hTXC5B409xO6K0zHvSnmTXKDW0cIsRURFwfd7o4uN
gJttGs8uaDhweKteNEHUObZo1ZmGAZAMJQ3JOuBDp6+oDfyZpV5M+CJ0uEwE6uodMjbYVrnjNNSc
1Nkz3dUv38ZNHy4zpqc5Q3e/6xq6AJxh8dcWvMbcNNMFvk8Nx1Nin4GOJ4gcvHIvrFa4UdkhtzWi
73ZETN9EVT0DCyv32d7tHXtzDKr8bt1QEjd0zhtYvNEEImR7mb2gHE1g1EQQyz92nnXr5vOhD1Mc
kwHM44FOUo8vZavIBqeoRz+1bix9HJa8F7hG1Fr5u0y5cTNYrur3zX0Icwrp0vgnWIL+87xqLxGB
uqVliTCNPj0syDLVLXeOJWnOMxUZUIwSx4Mok2+XYlWh4iS8pCf4a3+TfbU/GeNPo2EeWUI0o+/W
GyjvKxAhZLSYh5MM3f7TO1YovSOevUxTgVgqV14M3pz1lPq5bxK/Xl7SGgoM8uvP5ZP4/pCO+Gwm
JfNJ/XOlNBzjXq07vrFgnbcqoq/vc2KPVjuf5ZIcbBKUqwU06npKKa8TIszzeofmnk6P5qLl6yug
kGfilM3iusAGiAumO3PyoP8/O7XGCOy2ughOjxQ+0E03zSU2mgHYrNbnTNqHjJBX6Rj5r1KwX/zF
v+7ZBKASp72bAIL4nb6eH/e9fEEcfL2vJKCVkWe+/QurwnzBGTGnjDfBpjNfE53zBGZz9QbrXIjg
WTH00MQAsRRymAN6d8uqg618Uka1W3+0h25ACHmcuVRYb7mKXAYF/jV1sDODZPUeS5cQfAV2OT/6
fDDyxW4EQf0/ZOhjzapNiM1/T8Fjifhhoz3yf/78/KNn8VsBip0plV1QPYr8EfcRzNiyBo89cKN/
HbP5Ho7B0OE3AlD5MKzJ4++5GwKYTr3lk4Am+tOVggPJLkFJIOw7owx02oThdkAiJh5WDivo9nnK
5g1tUGo5WU9HOq6E8FzbTQMznjjNz3/+rjnYgeWs593el2xCul1aUNYNV5e8hsp3DH+g7ni6/hRa
i6VABH/g6GnXg0PN+0+JC+NR5NgR8cuLqkFGElUA2Lb8wvhNFbXHRjHaTUqKU8fzZksZZUP6rhpW
cHTOzXiBtFMOOFcM4VxFYTLBOYTWsCBwmOLECh7RV3/RJ5o4BZhB7eD0vMZ4mzcWCHLy9Pt+rISD
6Snq5HauejBVRT1AizKTjf4/UfKsRxzoTtDc86PXGqbN50SNPvY3Kof3xEOfop+BJEwEUXHV/4Wt
m1OW3MACA6jP/MBnZ1Q3lhiJ6kR7D3zpGEQfugPQHvYeWfvaZojoFh0DC9FXbHYhboiCZYAqzg2/
N0pQaCgfKhX24Hiw7NIv3P6Gd0LLcBzG3BG+EmYGMmbmfT+T/cX0/sbOVmy1JBimKYJe3sw1DbGF
4Q5/MmtD6mYoTUfaG7w5exMmuVj9El20qrd2x/pjRiealsoDebg+zEMfrJLns+q91K4r1WWWzJFi
XiZ6DiWuXrm9PKiNm/x0oyhyd5rpnDqigSZ28+GI9W2fFUUNf5SgqnpvuEGAceUcW9oGSki494/I
6QIKBYReVgMwOS3x+qxqTZURi+1zww7btz/jfLlkRtYmdVdRXD/CaNVszhaw7tZGn70g/CTQ9rHc
QevPPiVB5GCjXhE+GkrsAsMi2Laoxo3OiYRmCGJocCapfljdw1Yh7mz7mpNRwLv/s1N3LRh1Qt84
ezG1ENNHXA+bUwWhHekmkXE0KYe5XeZgc4t6wcYtN9ohhk/XPEJ+BWGGEk91SwSCFgTlGayNHSL/
cuFAwdHNNDoqdD5PUnX1yM+sj8fp9G6nPXBF9l3ilCYkKtR26q1OLviKyyriWffu+snzkLowNxlo
2afUzMQGNnXXcEg3tmHEPZ2GjYveZaOwhua2cEKlMiDviHw22TiNs9LcJqci10zPo2d+Kqn9nUUe
o987LnDIV9QeasW7AXcAuC3hWUW7k/bmjTKrkm+jMuFZQdKTBXOwRIdToByVQqThByIFsvZWgM12
id1tdYMmhn577QcWQPxPsFongqoXfwBFk2/++14W5zqi5/s7ar9dyIEyn3+Fjl/zZONbSP40O5q2
fy0r6SqT/mHutG7wtzftbx8WRSZxLOgoYe7AvQTzi46oglfmVHbRPMpOz9LbOXl3jMMXqtbyCN37
UCZYUxJfBzhOFdttO6dd2yVWaOtG8vEpky86btZaEmM0FgdU8usJVwjuecK5vtd1KxOZxMm29dAN
G7nBdAKHGuI7l40NoHkrp195mE4ymn1hLNU0fHZchz6/E832MzzBY5EK1VzThaCfo6Ie6xg1bUdv
NhsQ1y1aQy3CrsNFtYP8/FFtI7KAS5MYosTIaV3MV3EAW6pJl4eAXQ8dDBlgg3ezt7mhncPeZlWm
3RaL5cbpgcHVbUmF6BhsSrjS5iL7sG4NTv8D5JXNa+uPFdoaXrNXS15eIfdjCR//J53UUM1CUasX
A1rEFh9+DlMBxJiEzslEVNwwALfbiV2xbGD/X3eQ1RRovk5sMBzhRN+7OyQASHWvFk3tWCY9kqWJ
/wdNR8P/F65QxbtU259pFcc1j0hlRTvaisX2JX9n6gzAYqXXmKht9ErHZi7a24PG7WZSxcd4reo7
zbvvBMyT6+KojZFg/OCBfQK5j3r+9PYJtccCvYt8A2tPs9lR562k+cPfQkCtElLBgvE9/0d+VLX3
pThDKD9WUH1oHN7h9ozGnUJSh1gldI13fVp/7EtcfszToO04NTD4wc25PkS1w7gDXcqx1uaBJnFT
McMpE9VHQ25B1LNLuXYkBDKVk4NH5OAKJFgz6TjOa5ZRWTGNyTYioVDXM2YLkmw43BsERfifCrTe
axMY5OA3pTIh7+CXTBa8ReK3bSZcFeorfpY2Bj4Q9fjC4JkISHK9IKF/mpdTQ6jU8b3yx4sfKoIM
c78cJKy5S5BODfXDaKorhVFH93kmt4EzRXs0sAnCMLY77sJXleh4wa7uRVrHlby7RQAGnQssTmbS
zjNrHpkwLC2MuU0NBtBucuh+0mZ1a8JQygxWfa/NGS/R1fAjTcA9wiNmrhjQZ2tOwmKyNJTKRggY
cQXyO0Wj2DCjUrzJe3d1EiKS4sudtV6t9y2uGVzgWNSAoglLmKFoVc7FspxJIGLf81xkdwG4F6Lr
9lOsfySQ0RV+YhhDm7ndptArvCNE8exHYz4ZcpsPKw1kbJKtsA8IXaNSc+o/LTVrzg9QsIKP8G8Q
prIubGbIwLWApS9kyUcSJN0dCKWB/ZPYZeaK+95im5PpjVwI+vfltgTAeufp4rluCp6SsGI2vhzH
Ib4ZQwbspIpUxTdlT1Xtx/UYtSAINI7JaQCmFi1+pzj9HCfLR7qPHdWwbeFoSqjjCZz213IQNbpQ
aY6f+25VDccwBkx5yhWB2emiPn5q2oHWtGvw+s1RSIICvGNdVAkYADNsR8bVB0Ovl7GLJR/aYL5v
ESlhR4i0oE7c705xYDi7+bTMZ/LLva7QjydTaa78HZzpKlfpEu7Zkr8ci0THQ6b+MNrNZHmQscBN
dCHggKNFSRb+MQfaWBeh8Zyptw4a0+vmXrGl7RZKdbJiE8V6/TmGBX2EiC7VKXF4suYiavCIOlae
LJ5v+L0B7zrwecEN3a3f3cH2yzO5C9MhAheX06cR52rxt1yX4wYtvZcSchQYBIouJw7juk0TgvZA
dQUgwz9kwWHrvTo1B5wlNDmwWR3wKYYVvkiycaSDOBnBDZ4xt4giOh/Q/5V68o4dAmDZFcz6GWSH
BQssCpSASrrV1QFr3kuIWg4d+fv6bZ9vDMcH7io1Wyu718IHMjyTYYmBbZW82bBAmQzQhgxHANT5
DPohnQ4DnSeIDinpO/7UDyhydNw6S1wx7ZJKJ5puYbXBAcbN2ksbBpfRKVZDepmDou7LiUGoa2ZI
NB0PgAVDeTnXnF4h1or8YpWvuD8MMRRKf6C5CYZIPodV6UhyxpbffuwOt11z1cLKQ5H+2sMjg4bU
BheCd+30fCDwa0H0p++B+ws/mip7aAF6FZ5xPISFTpTb3zlt5ThVlc7ud3vLW6ms9uMQcMaLcs5B
/uoZ0PFFQSU+YnwWxWx87Mm8/qKVCBCn/mOS2wtFomaF/pRJob2OnZrY3A4kh2emeY9NbUlW5suX
0VOVcs9BiStXQQJh12WoHcQvlebQg4WUZrAPIP6CCnejGCsgEXxQSa1mmt5APL3bg0okYP7JI410
oxQ9Np7u7X8VUQuYIs3NLOjvNlcyep0QXPYQ9ww8K2o0G8FGH8nqy5j9EarLWQYVibzGcIbS4AJt
iAOdhDaiIvTDCr1LRoxZdWgb/HX2cLSMZ7EwqfQ8og06c/D839kHY0nKL1Uod6Sy+vWcClFRwzTC
NcqWbzpQq3lEpJNRBsSHhH+iw3z7kFnTgXnNs0OnmJiwU7fhC/f8c64ajCAr3CEVDE75aIdwnW74
5qrxGJJSfQNLZHCSy0qDnQRfFtwGCRwwPE2WKz4dZ9aEgjMY3ZzeSO4jnUyerdrf0jjfPoPZ2NyL
fNxe9a0QPYcSBT7E61cjineTlZapYxT3HDRp7cNqeH2b7t6cv1uRL6Fwc8KPYqyAYu+C5GJzsFDB
T3znVm3ppbmkqjsv9ToIeFOYQZZd1efj9uJz9bV5tKSzH3UxxgM0AryDnZuofAOBL2KZBfbzI321
ypjNbH2DrwDhi7R1wBQNrKS44EHC0EbJzQhcILO2FKvnExCK1MTOzHCn2LIPZe2unAPr5UYFEBVs
SIzzo4dRA31EpnaZNJdIk4v9uRZRWNu+VjubNkNNDtnOEzSQr319orBq2YXJKbFDd1fWY6TyzFJW
Av0moRKOFnGiObfYV2KRki/3tcZ87ChV8LDcnPJs4k7cGiuSdCJy7s5nU2jyjYDeH5WZxtTZWM8m
MdwGuTn6kVYncQweCYGJdMbPR+oof9jgXGyaYdPSRKaIhBFamzioBneIk0uwf0sQ4FZeZrNWS62e
QlaPkRRYMD9hR78m7p26KgLi6smjo2tU/TL8+NTztUZ25pB/zhW2Lx5YJ+fpyl7afFPJap0063Br
gTqPxhtHIFuxHpU/HmO/L+kaeyzkLzzpLXLgbwo5HQb7W0RnWNwpYtxK+c1+p/tUvo5XuDoJ/OWq
i2Xjgcm9qenKnYpt3037ZAztHVje2KbMCkVlM0DPyKZINa0pZcLQWm583ZEUQhvnbFttH8J/FBIJ
JMaQC3LH4YGgDKLR2osOMPDoQz12QE2T7w/1n3GBKCNZQqvRYhwY8s5Lp9aaZFEwGuBbyJ94xFiy
OPwbrMbcAU+wndJDqBtVq1ihvpeqY/u1SRJACTXWliEi4PaVOZmB5w9/QPTD4AwDaUPOokSIpabJ
zxjsekt+5pVzsq2opXld91ZD9dI/DuIFaIB55MCh81PU4ILDwb/Bm9ikUN2rHkDThDoC8CKvAaAS
4D0OE1QxI8UABaeHD4LDSO7arVP6PISU22ki4NKdp8c9kLCd3j74NKDQjrEsfZunHQaAczRHDIzY
9oQOZsOgdpPlfFv0cPgjYYJ77Co4nYR+pDhcb8MzcgSHSZ1RLZhh2+GQjNfpcfQvVSMoFmeXsF/f
oScs3VlP873G2aFjgHiaG60phFsoiXKb5HEicLachmTlGO3n/k+3aF1Ix0ZyA/NVJuBC0EpBUOpL
O3vMnmNm3WVUh+HhhrXgu5cLOoKQaDHYcC8zYABrlErxWH40oM3bc5PVs4heiQo4MjfVAR7UhwV8
SFDLZwKbROWgoFgskCG1SrktBtVH8AJLDqdULy2u5bvMj9L2V1OzIBLtvzbua4bnPEyMkPjfT/QT
Ddumr8+tPuiwCNtSN1H9Q/yGPHhTiPLayUdVFHZPT4qc1F2cxDGW/7v7cQK/I1gkw55h/TsUVLhU
cNwMli3Pkd1UiEeuFiAwvX1449ukurnsMHbDBRiWLOBdSus6OQMCkCzKdCOMYgqoYCKClOUlRnuq
fDITBVbu3ooPHdjoG4HyIboaRPdMIwQ5t3/aE0qYya2TRzPy69DkuR3NSOmM49uBZAXHjipm6lZo
DaR8KyciaKXid6K3cq36soYKri5AbUgjb3qWPFPB5tg+z1+12Q4DaAA1LZSPK9XsSDXshsUaavU+
e+sHXGQwHkF2IfVwKWwTY9LatpFRAnDOxg3vA1QXgSTqEMj8fqJZ6ER3nRmOVYsn2SkomRv0QKf3
KB9AF94X4xc9GMLmjmmxGxD/wOs06O1xg0eBfwvRiCNlusC5CH+h29Fv49CW3bcmmt/DDhXa4E0v
HeS8QzeuWV7uHV5yJqOEkKuLO7FLfFOMhK4wtvnVrD885aKRozxXKIte/TTUuBEYjlxoUhvlRgGn
Qz/2lCjlD7BmbQimO6yRqtqycEohQT4qxLIzzKcBADZEYAq391E/DsrHqaWDbHbGFGRgEPT18pTh
6R1cN+lFh4/HDF8k3njdOeWUXdVoKs2TrWy98V+1YsSCJbsaFLj/lYRSDyfF3nbu4CGF3Nn9y2oH
5SSNppOGWNZLiTAmvwnfx+3eWW39MJCNC2LCBdikiaHH+IjmnBmKCCoJUqtUMdBt7nqgqK4MfXuo
41kI9UX+FgF3nmk7ELRHG2RjazCqgSXkzOUM7xE4iA083247AeD4KioFpfH2FX1xqhYLyVTkPmLk
jGoBiSmBT62HDX7FoiTl3bpjlnyDmHF+cZkDK6n9shRJKBWp4igoVeG/MstwkWI7E0hbyzNwENei
2Gwsj9we07vz68VfPyAQW44UOYpNobZMC2A7eKvGn682Qtd4eyu++Atbn9tpTmr9pRqC8LKubZ+R
Aly0kTKMz6sZP02Wy68Wwbm1+gbr7nZcePrLft2/hBvKBWo8OquQ1YBmL6Zc1oQOUaIDDsdUVe5+
Zad8ZpnMvdDaeJ2VQ/vYyhC6MYg1tqsXG9M75fEtq86eG0q1P7rqcJdMzF4hqX991/GAY1I/boI2
zLinjnfuDdQME8bq/jerSm160jlN/asbzG3He+gzXMyr78ZZI+ga+2/yosauHw8wppytOARUzh8q
0X8GdG+lV+AMjXNCE3IcdNg6Ls2HGxFQlspgBTRmsDZsSg4tsPOZlRa/9dwZYRPH4g2MAnV7clHM
lQmK3x/WpkA7jZgvxdLMp6hpD6QWOW/5kq5GFcPSWa3vZQ6+qehcp0Asf9hcxm9Dvh/9q+YCS+rP
Zk9BRC772kR7TBJHl71uvOe74lcvP3zR85mi5z1tC0Hv1J0KKKhA53m18InmAo3/ySefay4VyRb7
WaCBbySeZRVbJjqEgc6fT8n8rIzrzQiFNOrKNfTaicGV5lS8RC/o3r0ue1kEXhMJw39bi2q/HidV
M36giOlCdo9yaz0PHxzni/Q0YhpqGNb2Oe2Ded265MMeePI2PzzaAbXfDA1+Fq8T4CxU8MheI14b
XVTKOq+s3REBKbMdS6+f/I/SDabkgVgjCeYdmb79ITQejEw19ZOqKRkevp62vhIFuqGWYL8yV5Ua
yK7saQX2PWMsad5DkaPODV/e6oSGDlX4Ee1mEEo29l7A/+78FHPaefGrN1GgxdukkiS7t4Ql343y
Cp4K5R85CcKKMKbWWx9SbEGC4ipJnNUNZDVVOhZ0bW6SDmBj/wDyDHo96ZFxhWc+MuJN224eAoCu
YVviQ+pB/iofnblBRsFMUFJpbKzRvxWIp5tEm8CmIspxfW44aF/+ppmFYQWjJ9ZAlIQ3db2Ip3CD
m/SnT3GA0w3Z78F3kQQXe9tQOvIK53oIW3cRtw3k0DLTsgIm9VfLSFdYBLqtlAffrSNGbEJAGgcE
CPxSMrQxUHAJcjJG4evO0f6DBdqmXlYskGfOudcEjT/TeqSmr3LFECLSdX8nBSMmbh3yms//eQFD
6XKGmmcA40cs71mVp60dU/WWQpLniCmwc+2d8AVBnlJjZqT+Y0lCtCiUW3JRVwtgFQvzg4mUCjUR
n6oKywpbU26lJyJrBPx7CrYCQObwVFPW8cEvhheJ8ZSSsXBZwJJLY9ciuxaxTJCnGlXvGOLl9NyL
8l2EXVBrJn/mBRLdrc3xXYzo/95iETwsHrw0ZE4fenmsUUBhSVrmrPie0liwqcTI3iuqzesYhGgR
E1XmWjT4lw79W6uQkCkZbY/DJTuuWRBAmD5lE9UUuli80je2jt0rJMO3Z3OD9oXR69dHrItwLq5G
SpCE2M0YLTsVflDjmJvu7EtDW+AKzWRI6I+wqHhhktZ0hBaAZ/RjXXlWBzgw4eR/TaKnT39qZm3t
HOis/kT6V7EgmldxnH9Yd7oqeDG8+MGWKxx4I8TS6q3cqiMpKTohGEzGhxwKr6Ms9Z2sC7NYZihU
cNYEFHP6Mjce8jXSC3RHEyggnbfklSZpmjPxrVoa7WpwSIEiZNQJzw25EN22/L01XZF6UTIkNUMc
TsmAfMC+/t29jwdbDY8OuAo4m7UlXEHbz/zfixQpkwfNLBt5X5YLjHsVSEZlaOHqFYRCkHmNUfQd
BO/HKNy2GrUFnpl23Q6J+VcHjeKVEVER8sxat00snelpgtM4p1IomlZt2L/C+aTt8vXaas4KflTa
E1/tOz9APp3DRTaZp60TuPDiU6hT3EmGDkWGmaCpa228o5efsW3xn2HwdQ8+CsCnrHalWBfddk5P
cWAV/sQdDQRmk1tQLjvXWYP6TC92Fwxo0d9Ewf+NtGe/NHs0KbX8aejBcppFPkFFqkPn/piOlq8c
BcX4xzeAqJA+PArBCZIBeLc3N/LMj2X3WDye34YymcwnRefwpfYfyz4XkHh4FfGv24Wl9XufF+Ue
lVYycun5Im2rvz6+hyUd0PLTXUIUpJ6MZToyENGB+tJvh7LxLxHDQwNGw6pamvQy/u+twR8maJ+C
3KBFbWabIVuZAM9nvXGVH6arwc5FTJx5DC+0nh5obSQEi64dWwcE+EwKXL8+weSIRyflrfAk2+U1
8uA3wenBte+3yQa9nqP9l3zE0jV73X9/1yjm/Bb2Y1fxPqLHA306h+CdoReDv9VbO8aGh8DlFNjw
O4idQ+NGTei5tXtYHnvlngiBCrpbcZKPuT7Kkzv8l+AQuFZz7+VB/FyiLMEeqUa+w4aynFMmt+1N
Y7iZwTk0BAi5vDvq0X78u2xYfvt76ZHSTebydrsZeY8tiOrTm6g7r6fALf+jozdEv/D1OTcHDjsn
LKYWTLBHLq7mKeyye3xQtoac/fEj/X1VxG+6BkpfLdsvRzDa7g+Vq7E8LcBxK2bQcd7wj6/MvARN
N0Q5RWK7zzHIeXRxJ4XFOhlfY2IS6Fwv0UTfyvrlSO73YUUWdYcSbWk0xRk1P1TSjWs+/Rw6rcxE
nbfGp4rgf6mcf/BV53psUKdq5ZpmrGHJ4Zj1+0okpwYB0rtoLpVb6aeRcHeiEXkMS4oEjcpC/mT4
TuahOcaEEM7ESuvuG/CJoCtuKEE0uc6x4//DPVgi34tD9JmhZV0bIbIHoEwv4Nsmoy6KqQefZzSp
UZ+vBb29iTO3P6y5AdNZmegocZ3536FOSIh2KtH43Wf+zLkRDcuj8pb6/y24HVdxYHX2Pg5rlu/D
6vSHraad/aPYPdvArq/mdUYx/O9DVhMp7nTV9M7WYNlGlyN9BJnTNrNeZpeG3A2FmabU+ttbifaV
786B8hz4gby5fmxrnmzZUh9Y7VLLL7fMu4IXbSi6RraPAHwLfAo7eSGRDK85e5S38auoWmXIcWs8
t+g5bc/jVSpCFLyvBXmCMmsbUHAeh1v+b9FscjE/GDC32uwkPRa22oP5eomWnGNXpMvoeP8wpdEk
osiQ3VQpOlJ5wpXHbcrfQ/xWSEPj12gi2PVBAMYgj1Cg6/vzlbbNWwUrX0qJ3TJyh/YRPrgFClwC
R+yyzZlFUeSqj8uojlba3c4XUryz2waCeC+VGTOjWUQsJ+TJXed1KyAoR+l/kC9y2v/QMvBi1JQl
DasbUhkaUGghs0nXAFsIaXUv7V3leoHwXmAkMimLzeb2sBqJVh8OwXsutS5GReYys0+FIQMHR1wt
SmzlAyu7ad58C7A9wJ5ibhr6O4s9Ci6baaNyAuWWIfaYnoePg9jzInXF+KC895ff8ZjiFLqXqvdi
o6VHEqedl/hktERReSZisWGL2dH5cQTA+2w9a7Ohw8Jwhe89Kz+1ScqVbHKSAlpSOi65DsIbm+5S
kvU86yIe/c4AXVWcVMr/k7Rz4dIdAhS4VsmSD4N00r/a2uWuSEZXli3vrMPTPEYiRXOQUq19bfyL
84UKmJYaSlFnp6BlEpaiHwDqOqzfbtf2brsnmia32dG7XJQxD/8yg/yqj3fwlY2RPRQ3hQbk4ykT
NXnopN/3dr0pIBRwiGPTNHnkDk0Sv0NFiCdkdKsLEVB6GTnH5u9Iuz8+VSvPlcw9M98BUlbnuZtz
Q+RzV1fiYbPQ8o38tnQx2LuxZE9rnh8YOHhNHiLgaZRvf+HD3Pl6Nrtq8dKTt9lCVipquX3yCnJB
R+WxvrKktvLleouaDdWsUx3UkixKb+rhs+QEAzKmhugR7KKtnjCFhGxr08XKieF4Mi4IELkOTZ9K
FI21G1nHfipEeIZ/J98kUW+ipNFkBpvHtseITTSJDSBEMfcNDsET4RkePSxvCr8WOTeL0kAdOEIE
h8Qb9J1FHq2TiZDwNPiB0740cXL4MSpFMzmTDOoQ02XjKrt/rXLzFg60KSbUafJVtZ9RqvX6U9lr
JLCOjf3DRl2G9x/ncJ2Kk2XbcNojC4ZivCO2T8DM2L9/JiBAnrcVDO5dui6DUygYDtKF/CttSJnF
oFnnAU1BEmpb0EgbxAcbUNWtfhdwigKYIqxsROtnmwi7FB3Fju5TnfkD/6KiR5ciNY4dqBFBQkKo
ohq9MurnjF01pxnRPCN6miGwFedfek61GeZZrbGu/2cpJ3Pp4biQHQNC3xe15b0q1p2SqYtWP+y2
XGvWBTAcKZ70XB+86qxJrBbkBrLeH3eK9lXhM13RpF7RJW30Ntg2TqWNMzhKypp8LIaqTFB480Ty
CkIYBYQ8zxCLXK3HPM4uuwLAv54CnNLQvr0uOelTpgBngcv7jJahqBq5xvCl863loLvsr0kXGhix
e3eSRea23EQjVZF7DFtyCnZ9cBgHNaCSGl3BC6nj0zYGIB2CSxxdjbys7+O609/4li/Lz3BNEVJt
hC8+t7VBlp5belKVmM78QrktmDgLAE3FNI02VcJfiuuUFmroQIYH2MMKJQZQqlXGfVSZJR93F05I
EJ7klkQRnNYrbsPppRysOpRTXAmOnMas6XuLffZ18oj7Po/EKQE/L2KUTBGEfJ+hTReFZWMn6TDz
yUJkXGifHAIwZyFuaGH7kJ9XCb09cpkXXVNeyZUNK/lqlcNVQo29xYm5UmowY4jZ/rc3rDoCGxxv
njHcxsH9azuiMF3xy5S8AX1Z8JAyRmB75lbkcGMCAjiYW2fhzsW2ED3JJLh/EK6pTkSc2iWtYGCL
j3KeoVo+sXQGak5Hwby+/1014RPrHJ8Kq7o5B/vJ39h0cciDUh2+oBkOjx9ofGq/zO1pmGDJ8kws
1gtgNuS9jtKnAH838j8BkXmiucz/iUHtuRN8ZdBCEcg/qVz7yPVM0PAOUOa90T6rf2bK6Y29SYvJ
x82N7276czrK2urx38lqjQ05Gy6YqfIuSWUFoDLbPkGcHZ7g1yeH2NQFjrlDPBRcn3OiPgzwBTZr
AZJaP9cOilDUdMieuqGJly5e22l8T/+XN9wIgVZ1SFhLPQIwtiJbkQDgGrKwxTasEaey6JsYVGkX
X2/wqlLMt+Jug+pvbArAZzQXOsxcouRpjADiSa8ruCy5R/OXm1tLStQH77Pz4wFbdAbtOLKHLuFV
yI1Rc11wmi/CUeU/w6Id5svpWIdSGciMbSyV8EnW0a8/09CEG52VMo0asGYG6aZ45cbFVI73ForP
1eqhxteomOW5YB4Q56yzv9mwmLGDsZcatKw1m0MoYETRraOGbgoJHat0YCNSoaFwzpl+vP23q0dG
/Y0pK0xyk4AThvGfi0umfsDwL/0cPekuEf/oY8e1Ed4MU50Xaeu4RaqvJinvXLOtjhAW2mRwq3Do
mvaxoIRT23u6FKm0lut+2uYHPb2oYRLZz8t7EMpphVh30caWgYnjSZq7DnMtpICV0CWGQvjb3YW9
FQJjtiR7DvuFwpMViRlP8CD6bKDNqBR2INWo6gLmiFR28tGS0S3LRHVHIIOjY8GS5JOb71g+OsEU
vQUdFaMV4hadsd1xgny7rRo8z36iV79TXtuTRUCjI5CZU7xFosrxr2OYgocx5M2woxA5BINcWd/Y
Xry/pn/ZmXaRyzYchdFER0r/1pKbKqsRT15V6QUAmWjlUdSoHb9RsbTvX8mz9qBOWGdSX8Qaasn9
1P8eVOzaSE0D06xErK/ZKrjsTmXrdw4EdKXnIAMEwKIIPryUhM5C8VLrYrzpmjYOJAQwsSR/DsR9
luhGqCz++CYIRyj75nieHwN487QqP+Gvi8sgtPqxcPOPUr+pgJg79FY3U+bdzTeu0/39DlGV54v9
rDHjk7/vNV1ztqdeCumTsnec31Iy5ddpORmqQ+SBEwuam0AFgKClK+qT4eTMteUFAiyQab70L5H0
wys4XLmrFf+jtZur5nncqgWMJNyyPLQk2F72eo4/fjYyCJMlMTe/XdFQ6bxh8nDRLp8wUSVB0ZeK
BWEf6UKnndGoGPOdhgV+knE3GGuq8LfUd4pNkuyfrYF1OT//ghaksP91sgl6N3u7EwZaR8gAG72H
zaJcs2I+4AWtL1ic8RUQfYrIhwdkm+zTSH7+BKdcs82Bx7EJuBGbt/GArNMAWbjesEm4hj4ebMuK
6/12kvRc0BWktVBZhxcxbZpr7VU63BfLB79GsKodyr6tEXc2BKvRvFqH9ivR1+589y6ilCqfDDDM
z6wwZP5/dUI75JTueppSFaymzA6X9CvIdEtoHYabfgB7y3lvds+EnEiOyWHWITvsCG0YtrIguBeL
H1aMd0lFJQTLTyxFGD5bcQXbodPgWhxrBgtSjucOkUO5YEeRqnrnWcAx9sruFweIbLiFBjKgg3QW
YuPTOrcfxtCfe4YZOHANlouInLas57mTX8iFO8Z1LFVbeljlZWi2Jn68/PEho3UckedDiAspERPk
8GbdKd72wprv4oryC5rmK3XKzoTzk0l3AaSm/xTOPLKqlI05ODggB9GAE/Mq2BAm839T87yywX1j
QiQiQqfm41xSLd3yR/UR6D1/FVoJYzhKgRc3OhMVOOZ6eGUHII4YEMQ+ftDJHIuzUx0FcA3LXkaR
z9yrqmjDsZjYJPih+n97d0qS+W7d2biSesfD0qVMtjbClDhtkEhT1MiI+PsjyOagiWkJhKzaF14I
e9F6ZyAhWJSLmTEtoStWp5aaVAbY+OH0Snemj4H+xzevHedUPQXqrK6JpffSmk+IqfuueCoNy/qS
fxX/m/7GLlFw57j9y+XBZAZw4zFDdpumnOsnDN1sGJbtB5sm0jQ5TQG0zrHNijwwDAy8pB4ogQim
LErRhSDQHUYyA/di9w1Az1r+fqcchhllv6INnxci6lDiKMUSE1QOpz6RR7FbK97RG1+eUI89OpEa
ajxA9JrdHpOeC3nY2r2YJl9g7Grd+MFEXjvWlqNH3mP5PLKXBepUptJlBmeor1SeQKmYsVEVJqrh
ET86cW5ZHQxlJhpi3kdHUuZeNh8ni5lgwNRXC8qTcsd//YHHzMlWjgjKcaGdfyz77uatm5+YPyEA
t8Su0wRly+8b2art0lY/4RKPPc+I/9tklHyjO4xIxOvtvP4OX4MCdItP5tTDFsege4aKmx26007c
zh5W29On3Uexm3MslOKEAKLy1VfsrSnQ4QXrXDLEqXLm4bELJ1jQdpvl8rh0Kh1IPYHJvihCehf4
9BLZCH9WPYayshm5N9iCyT3cuT7AH2YItkFwwvrfTiyygLbnrKYWY3ip255ZZFigJaFNw8tBpz1R
26AJOTfXo2AzDCjaT9ABOguH+3KfTLIfz3VgqxNnMjmo5oFn/C4eo7YIn4YYSeqyarGp1PIRuRM6
3jMHAqAB6gxaGWucMNhlJzssAlxnbuuPfbG1ti8QiPrIzDrRUuwOXe56XKTNo1rMebkxMI5y9J+w
ad92HNcYZ7mWbQ8CFm86AjfiVb5/h/v2s6R+/Y3RRMeco9Me8aceA2euwLpdSQwTE9AukxUZk/h8
UZCTUQKknxnkQk8DPfRg9+RvW5zG0MYB5TbozvJGcHA5jh9GezE0N3uyA9c2c4gMCkUkNDoibRt0
66OaYG7nGuVQXBos5Ogrf0FIVTSPzmUpMG7HJiM5HBRDFjpscUomqTuqr9R6dPdwVmUJnqTeDaCo
ArSUzFAsgtBwBvVCs4e4PJpEpiqT4U3bfxuYE5m2vdpMUkjWIyWS6CvEs1OKqldjAw5diP5SBkhm
nS47sHUAYfQQ75hsDJIjpoNMtenKKFDzCsMyRs2hJyGPUumCzf2grZMKwap2WriOqTYI/0Uv74EO
v5TXooP7ibOv5uWN88e8hiS9ikpl3BmlKF/napVQEcoU2sCF8rbiwuWxM1yJ4tm0w9Z06YPiYhtR
k/Uflv2YC6NykgRcYy9ryKZrtcRmyl0pM4OZJBAR5kYyqLyRuRGvli+GzTWC0Tcb/y5nFvchCD/D
wMiZnKbMxvjpzHCNVf+CF3JkOavq+VX4UdeTfZ8p6qWW94CWMyacoziWPbtNosI0idjutXhFirEg
pjQeWugx6xSpidLPkNEJzITPGwxo9RXxCZimx2Bbv1AfeDXvDjCZeXelKl9gD/DWfk7MRv4KeEoZ
V+mCVYITn9qx/NQmfeztqQvD3IR84r+JvB9yEbhFejOv28AEsEpVNdwchR/O0Hl3h71KbYPbp3d5
4VKmPjHsjm+96rsmPDMUCyVussEN+wDX5cGbk76BVLi/gPHFsJROyw6/BuRj9LWdaDhQxnwqaPLC
/STO1v83FKXXf6SP8rFhbAIYqinat+QNzRp6mN7sy29DwEdOvLdmYny9xxREhWO8xzApxMPP3Hmn
dLS+rqVViskaSJm1jNHLhbJNyHQNIBnkhY50wqjwuyEm4/ShnynqbvyvcS3jQcXW46DzwxUbwqJ1
Z3z4Pea3NdGJPYgocLY3D+asQ5Rpd/pnfunBtbiijz1ngOMSgn3eW1s7E4vgiVtWUYHFxwQDVwNe
05u0uKJ2wbi2kERnK/gh8ODXwoWakg+C+QhTvWgRE6fOo51xs6l0AW6cxpfgZXgtdHs/YL8mNDHL
ClUEs0ZjhrXe9pLZ3uGMj8JiLnM9+9BEiNjVrrL1jvxDPBN2Kl4BgA8riIIQrrgHZjNp9cckyp8p
aFCyZR5a2ifmmFCID9Qq6hb1YZESbkN7JKqJyE0YAyBT7U0msxu0kknhQkcBDgXOt/pEZt6r/dNN
ovl/AxUjPft+DzJXuCZFVSpO/p3NAnYg6SiAdpRegB/xE4G93TO+wktZqSLF1RsjNEF2FzI/jMRr
lnlIv+w37Kh/aRWrT4vht+f4evREfUcH1abqH+fjYPuvTpnRtIKbCmBNT/A45AmDubc5biuRYFyg
yNkN+wp6kb0TsClzxit7/GxoLnTiO5EInLUPV7/6XiTXR39OicxA2vJMwq4/TSaELSU3GnJVSiIU
yVek24pas9lZamfIRCbT/chHWcFiVqFBDqLj4r9W/mFKVex11IHpQKss3Cav6QINLZK87IBo800b
YGvYhRPszDVeOzMkdqGabfsAniEvC0scqVTpX6wmo/YbNhjoueKmAkMTgOuxOrf9TGrLFObcWo1M
NoEKYyPM52i9DmV7NKpvba93ffBC9dLMf9ZTPvhDyDFE0abezecwHmCLEFxD3uiXLu/l33GiPtaj
sLrDHgOhIk7KsQdzA4oQHbLsSPrtijzXM/hTVF2jseaM8mt6oL/401pRd2VqT142GTDcgPU3BaHq
52L0SQTC4bjb+qmUtgkqgj+/4pdLf6rXED7lWZIzUBkmalJVryH+LV67H7S19JCpFpyz526pi5p2
eLqF/l+VTAmxEfAcw9yqd86HYcWnIA7M10ECvK6I43NO5fKArVa/6SDt7mL3igwnGIm8KJN1LNd9
F5WLHjfnbm4BgDsxWIugCFwD2zlWvDEPnWfFtmbJl1fJyV79R4JJqVWQAI4mtD6rLKea4F6qeBwn
uOYPE9iX7yRyWCT9C6rUZqI5v1fEv88hiMCwQ5Pc56DqBgw4bO5gsVmUJrX6896zjlAsiABD9Lsm
z0UwuhnXZByOCJWsdmZQwS5C8ju04N82sQ1+thcoRKvIaOrw/oH0+epUH3uQ58xh5E0SRpHB+XRP
MkRc+F7gViq7lsAHTmOhVepktlX9focanU/L2m/QVY5SvBTYRphSFTFb/RW/eEgU1pegaWltlSAK
2WM2jQ9TSC/LgJJeutrp861nMiYiXPj8pwXurgMSrfa2EM5DfLMYxDh9k20kP8f1UFQNTL0Q3SwB
LJUgjuEYYRTACGb+9qelSH0nuwLUAoRgtmQKquqRhqF8DivnShXd7zHyNA03ii4CHB4582+54sJL
wxLS1YvfRsGgnB/o85NiRtRKNHbpopC1XORyvpWiZlvNB/YWtNLkgmFtlvDieKGmFqG2ecb+x748
sl61LQobkOyTJPy6SLEiTbQDjcYZynypTHuCScHf5abYElV5JtWzv+CQKRbTFeUPFql71PrrSFXF
p6Xc3ePGhoE7uU+vj8Ffv/kkVSY37eusL7jXCrSPPiueKRr969oaGSHn+xa1+DuG8DSwUzDooiAl
6ZDJn7QSeH4rK3Rs9uY2Rhz6B09qsFFKxRL7v2z6Mj39cWX4mF0LhzF0OD/bm+PFNc823gLFK36Q
Yn4G8f0y9Oz3ps+/4DgI6BmDGxielh+2s/mhQj8APE/GSuTkt/iPNrwgJ9IPwczW/SP6WGbjQhsq
k6BmdbFIf7Mj2MG8d/PnWBEZNCQRDiLm1T9RsK49lw8o92qtIOpJdPYT2p4q/hRqXS1FigCKumLj
M9O/eUW29802Jo+jIiKVFoXpjge2hk7ct645UTTi8S5E0Bn2Vt4N+sX8jBovx08/SXN5fIgdbj8w
w87tCo5fvcelXBjb6T2+7XorTanzA4m254tPtxjm0cY7nv3u6ZjqeU4H626Y+gigSFslM5XNp8wX
91NRecHA6bZvLQfGmffMxhbvqRCK0GcQaYVAaUU82sxFPrjtkzX2oQq+YKhL3Kc1oSF5JzofvIzN
s5jrCK9qTG1wyuIW1vCo85Wf5G0oJGnzTrWzQMfQLvGpLbhT1oh09YWdtXh/Mu9376OQurQtUGi8
YasbiTaZ71wn4TEeNSLlCfKxjRj5Ad75TBVN2cqshNVKA+a6Q2nv4rLuojhOL3E1WVWF0PpXp6xP
bZAv3Pz6SBPA0nC7mfGp8b+HUx5xy5ukz2HiPVEYZ2VNUsjhXm2lB6z2brwTDAuogElfwYnJjifO
rz4sF187xkAT4D2SEORNulsNyJcKorVSz78YdbzovZcI/ZPly7CVFicGbma+n/Kf8oF/YwSzstG4
rANkfAKjAMIidyu88IksZT1x18g/0RrGSwB4/r0wET3BoiW/SQ/Nz1RxVjmMJnIHQPOwufXL94ZP
ahdQ6HnsV4MKnaXqaQQOUh84srgmMq0N0bmfIXHejRWR6MJCmo7VAWKDZFDzl8fdiCfkv6lpZx5c
WOxDCciY4xbHvRnjnYNlwxtKZG2zu9qIbuMIbu9c+YQG4h4jSXA1ntxm6x7vi5wCJeMd4O/yHA0G
CupgUObRlD1utQQVbEmscY21SRgQfBKrcyf0K87BSzt/zLZ57ol/zKMJUo38xB4DNDqgLViPb3RL
I7lnI7ju4nG1zXZXa6b5Udpb8uk3+zVLhnahxZj5r3iOO3ca5OC+6a/LmG7M6c5BAF+s8e/Vx8Sy
8a1QdfMZH7p2cWQkZIucoVFo9nZzR3F4m2XwwyPKJfVN4XB4C855LWGcVpUEhDmJI3vl0EqhS4fP
A6CEC68qXr2DEbDZNOIRyGIlb4Nv7wXkWsU33nLLr5vrChfkNbRt5sA9HIp6Q+xM8fpAQuSqvafY
+HVaTGzjjPnJLZgtxZcCFEjvjo4W4LSTbG/UHKNn6UwIIzouFNn+n4GVRkKDOCqEcqNShuEPII/u
LchZoZKkA+Tkkg/8NbTZut4kZDjnP0SHsHSiFvbYbxs1CraO0kS4Kfokg/kUr1qxuqjF/Ut2g0Yi
Xqesh1L6+91pRqKYrxiL/+t1YpV8KtJJQrgJst4UNp/L/lt+SwhqBhk4Em7m8YDF5yys3KcGVETh
cNWUCjMtWfJTJOGEHHZkRgOEyh0KB/KLpHut4p6p/tDBTwsBGOEBnkY2lty5Y7/xbe34Mzl9W9z7
WI6++6dAH/xyjXLuHSiWR3sFCcjA+nCjT7Las2Tgf598C8/g+EI9ylalpJSGq0ZB/10eUSUbLh44
TF0iHr1d8/NshOrrZVrK6vpF8tey28GUWCtJhKsIM5Av/Q3+ZFK8Y1zWjLEl390TfJLiKk3M6H8P
hi+YbQblIlLtxeniw13RZTWao1LNWQjUtenVTOqFqvaz7H3qb5FxtCLwIW5XnCo4zc56zwG0+yVl
LAOEARX9SWfGhsSaS6/cbkximD1jvseraGIIRGN6XPsGW8bep4shEGHWSYgyMeXMaHhhwu5xvNxZ
vvPs598KWvbmPAlLS8LpYEyGgITTl7Vq1XuTLmNDkWOzQXBqUnQtVjzqUOaTa8peyFxrqYoy28Q2
o3269eKNfKoCdnP2NUImFqb6eg8wKLXE4fcGn38B04a4rAEqMzvA18O0HGzMIImdEpeN3OexR9Or
66nddSOgqmdmjVGNE62W0bQXtKkv0PLkUyhoaxKZsqFgJGEcZ8YfsHYbJ27dPP/NIJqXZT8hx6IS
n/uMPgjLO3sSgV/QLeQgR5CGQSxQSsWS8uFgHWb6kH/PMvrhQddJYIDxtfD9cF2BwahQ7S1uDJFp
cgR24BlZG3CWBN4lY8/GiwLSR7ruKWR01YoY/PScXh4Y2GEOGDAvSlbXm+r+owk6fxn2kaowwBz7
AGZ4uApuTzBkkGW5SMirq8uOEaQR64v+dG+VXdwvPe3Mng1CZCrAviAXd7/dQht8cODPTnQGYynI
ff9xndGq+7/pIt/ol3WLtFINP9CU2XGXJzxKwT85QjbNpNq6PUje+7QG7wW+jAEVmmOIVksME6pn
ID4AED6HvBs7aW0KVlckKoDKtl6LyXh9mGd6cAMAb4R+qhwoeeqCSiQKi4NiHMk2u1+MCKg7l9lK
NyBvrZqUDqOeJ7UqdYHmKFQS5cDp830Y5ZPoj/pxoJgjeE1Bpsr8Y3bXY3gizu3QlZm+c0YAxngc
91j15GCSZfCiMjQan39CuyHHIYIjpsGczV3dBxrlyIS+cNqs3XF/rjFXMHD6qF7eXZ7mbWWfFkpX
Z0pJJUNVQ8uRrv2SwM+h3fQ5pBkMOpLa2sXNhvWkTWhAwSQM94bNxW2unKe2FctASHV+s3shMcGp
bojiOzw3EA33ubA9VpS/hrHFapusqh7IvIZi6L6iQuaGrgPfbwSnXGmPy5w5rUHII8tQ5nOFX7cV
Ks/05dAJEJFlHe7LxvCrJX/vipAxUV3omFXMnInyS8Mny50B8LaDdHcNvmDKvk67mg56vXsJb5Ai
GHsiqTfJ4EdqmFtH4yaVhZSwOCHz4zCFZrTzCqL5Z5A5KNrnWKI3VIz6wURVjPojTIIe5oNQxfse
SQnLgsys5JkqouVIhcWM+UfiasGSNsIAx3hKtI0LpB6DEf0C/0uXBS0E17Qo9dKNvewG6MxBbnl2
C++sfpqpIIGYyli2fj75LeH1y2fX7svnbJjg42dVtTpHiVcJ0jV48u4gaFaFEk8T0RrXA8nTy3rL
8SPGscEEyjZ0VIS0nmaVPh61Sll98ggGgKLJmKX7o+FdDw6J6aJv7f4Wk26acbPcHmtlmayQUAap
ei3u8vHu6Q8nzDMdCwMbNo2+OyL0lS/hhn0Kn8DGdGW9LLC3PvbAxBUGbBtvIBByVldcED3Q2dPu
jueuMfHSMGcF+7O63abBmjsI5rduLi9M8KoYOPmlSb3tc14Y6ZYQIMaj7M4RgHiqwqsovreq6Lbf
f1tK21D4o3Pp0ui4/wOjNX51LClQJZMVGL6+H+yU6qcFNwixMTAuqyDs3H1SZXAv8mQcfyMXMFNp
dWe1UxQ09EoYN7LZTeycvY7/1K4QhwsfpqlMjRXSxltazovVs0wv+5x8grHKtDRtF3gTaByuxD4o
GLT5MPB3T6nwjBYwOYOtaFoC1h2OQLYM7VcOkil6hoEZZokkZ2ZBr/wl5WZY09d2aJ4NtOwMZOcc
fanag+5GzkMiRQyp5Rmzo+WWDEl0Ykd2lXzLdg50E7iCeQ+bOFKXv6zSi1xXLk4z4ipvJzLhtjjy
OB02CSyrae+nv4k957so4INxVImf27pcDzbnKlDSiQMZnzjpO7SXZz6ADV6whhM8mcD932DokOpp
lK0AZDTsanqu0HtcUe0l6Gg4O6CkqnmUnWXANSx4C2rvg41Snqlk5pxoBU4I3sRw2IYDKtJZBGvr
iI1EwJfMT+Fw/Q+A1n7mtLE0I5175g2PajAjAi/qkLQdVzqWCe8SpqBAdllwyd4jdcl98ppYaP73
BP3+VaQZe8jbW1rYuBwu/eAaYnLVh8cdmAjC6JJIiOAHyJZaXfcBiJ9+dMZvfYxiK+TueQtNYvwL
cRETed7xfTXWCQkmzGCxBwnhCW0pTQ/nAvTRTbjTzbSkS2BIv4EdpJC5mCDRpLLE7GP1d4mRrbzA
Xcx/UPIkG2d2cDP8XT3B51VLd1tkid+VOrRuCPonqoU+pwje9rD4VGnPNA90RvvC1s/zJN9o99ws
P+mzEFQDV8vyGi6CR43QdyMOSY72mEcVd+hm6JHBbqP/dVK0Lc7UK39kTO55S5Y8WcykM0snIAt8
9+iDbcgcoHy2t6+Cv3a53m7xM7XORMluqnXrRMOn1gPkjANFcElXOiEftiQhOLo0016l2LsUp8eQ
INqGjll95VQfnuGsNCRVAeMfPpkMG0uJndcZ2v0/4LBl0KIEtp8JFPUN8je4YCXGXhmRpD0Ah01g
zucGByJ8mRkW2VfwLHApCVboBWfP3QnkB326u25w/OkEFtFKNwdVHiAjl0hJ4Xy6GCzLV3pWucHA
kQOmD9aM88rUmTT4E8sdAe4sV219n+XOcm6p1wJRfEyKgZY1gdR6kXhqq1gHUKk8DzAcN1LRVuBk
esXurtmO/ilFyKzUFR1oKYu1H3bxiDjELh+Ti9KYXbZS8NkPD1weNB1wnA28YlGtSglVfcHPfStI
k2W1tOaxvGAO8ZofSJxwE9NJ4nJmkJReXC67+O9hDJ1LaxhdJ4pgWuwDnJ5BSVljQ8UAFJvuDD14
nzJIJRjSKqLjzjZDP7eo4hK9pKmWX1IIc2hI5vRgCo7S7gg7RSHcyddKzPVKI3mAZqZUbY6MMafO
twNIFndf3W8lIbJ92y3HVXLuujqGm4wNmYIxgCY8GjOeDkvDs+ThWlX5lgFP04dYisuIHafFCyS0
XbIwRjI+7WU2Qsh9dXYx/7UOXKSkcr1nZyaZJ2vA/BAnDSf5xIWexi4kZTQ2K0W3ZeHx6K4Vh73F
wr5vPKgOcgWi5l5Tk1m5iyuyyhU8W2D5uUmhm5tTAa6IhQ+R2t9Q82n0797oG5BO61KTDWjoIJiN
AGKB2qcbItsdGOnQ6zB+ICSDC0w8cOx+LDlVtc2QI1fKx9U34QPjZh7QiRYA/E5BUfJUDUmUQLyt
TbxbwV7IBz+ehl3v/wVfojPxATTgmvg6fq0aoaeNRhZrV83kvhw2WRFdBJa3hOGbJDy2gz89w2NU
WtRhGyO41D+7Lh6554oWnFVT+1QVeqbRXk6Mcf6YkLZPEpeHqdK8xLfto1lFr0ppgexB0B599o/I
aKGrs1aG/15bR6AL4ahgsmyqmP4yoFiNlWZPYU3tdCA4GcsYbwgth74Vw7/tqBeAbhcS85566Utt
pxu1wSj/iNpiajE1Fn/8j8FyQeKzIKDq8DZMmuBGowSA4kIU0P57uctnoRCKgdeKBBAajTMWmYcv
tuGYRaC8M6KTCw5nY04gG6C1RVMmh2afO87K5d8siH60Ff9kTWS5oqsiyYGfwhHMf0KhGImFYC2k
IT81ozK1O32PL7xuGgd7VeA6SibPZ9NSAtgze4xasTN6NO2Hdt2B7blYzv2/x7RwdXKAEfT4PfRM
TcVCC1KQ4k3eAFQz1TB+gZcrVvehyKi0BMJs6l2pfSfCPL4p+RtXY+9WZNPnpeCJQ91gr0SteEO+
wx+fwnBIoW3xgyFkonLg1PEijdCuVm3yDL6SWzn24pkzamxxejedL2KnACYDyZtbrk061tJx+LI9
9k1GlhEqu8jhVz6B0ilwZFe/VTWGcYw3GXwHZu6aVrNLSYb10EYD9rOLkGVtlrWSc9fhHdPjk4yI
+OmvHYCtinHQJSN9fa/MOn6ph1r7f6z0pSsPrH7DP/pPGh8UFnNn4vhsD/z22POFS0c/SgAteHWF
dnwF+xPnUy/y8KJrDKLM/ape2BQ8941pJjmbBLewwViyLaTeQ6g3NNHZMn8KP+N8fVUhoQAA5Jmc
1FRta0D1pWBfBXvPqKte47HurzWDv94XIsRkeHd2WErL6asCY4RieWJePsryvvygSvwa2KLnYJCi
J588QktLnpUlk/ynBprVLe7H8JXLHBv++MmZNNSwDl5mrv7OVMd2NyjB6sYyrQ+rZlYqcdO9l6kW
QijhJWqYn7MlX/nqJSpPo7sPXl7iD48IjhQ7TuHxQK1heV6rUP9pgeo//Qavc97HzJ04hZcTLvrD
Hjd+OG7ETrnbinis1v0kKesJvuyEh6zG7Tgyin83KdwXwn/ytLWT/T1ME24JTagXPVZyB3y3xaB8
lA+z+NxRAcebD8Hpmt5eTlKzptIpJVeCuPIyQhI79czKF4Kwe/2Geg6FyBScVHSctchCTlqQWZz6
70jHrKb1BLth0+Fowl+hrIEyTHOq0yGE1HvYS9zcVsodaUU8oWj8n9afSxr+g0uwXeWQPXin6SK1
oyy4Ma0dGK5QOwfAyvgQ99ubuXvkIYKLU2NmEL+Qaw/pR4ybTxx/JjbH4Es4Xr8aENeUqOnR9Y2l
LEm+25Ig7drVsD2QnrekjKNkbIV/NZx2MxmrxvD999N+Tvh4ROnPR1NYX5spSTrPiJo0ckAXEy0K
GVPpKOmOkrM3ja2qfLTULYUIQrFKnmjkqhHIir2TGnO4jwFCcsFa3i9JJtEJOV5F1xJ5MciNd/GK
8fijo6qImrMIwJYpJ6mgVv/CuuIGfOzhzACCf7+R8JnYwUtsJYs2aWpmMdCXhOE6zhiLOAlEJphI
KeGopX0iTyYxBgSKWADpuSm3LFZfw3qqICaYmPViwbSQFOtnJ1v8fay59poEKL7Y1ONLKNpYsxlF
+pTCvW29sjGQCFfYQTV/zQZStUJCgJr99ZksS984lUbM3o4ZbwIdNgT6Fl8x0jgvUiL6J2BbLZ1H
vxAbnsHmTlUjiX5pkseU/F+2O5tsKuE+QcNxNLMMavmfbW6dqovX6scp4QswXy0gbsXpGn0e0pi2
CvDTzpMbAGB3rfEYd1DCsqijEnXiBzXysYjMXuVlCcv+whp4JipmykJvNFVjI2K0YQzuK1AHImm+
c0OpBfaq/IUxgN7KX+oCrryZi2fi06r6vuOjtBna7qIHw7QI6E5y3VSwD+D1hSfDQqANk5R7XrBO
PWm/7mT/sJP7Bt//whFy1JlSFJ4dDfnAMTizrkUovxYwbMCcT+CBWOg4qC2kvCYNQqukXDOBRdfH
cQgAsaYvZsLzNO7AHdEdWZmQrcJqJ5XV8scf3Bzne2ADD1/N6C4kULnpPj49vzMxlWDC66iiBeNB
4VeBVixflrmFGbhE+0KTQ+VTrpCrxBf2uMe4nH45pj4sH/Mg/qDkJkUioMUI91mww5TF5hf+siXd
w9oc/SNHY2xMBq+GVRG2iWkVSXfP00RVRfMjaRrMq9gz8mvZKgYYoANYLL7MTug36ykZgIWREhb/
SEvYxGxrtiNKiB49W2pgW2a2q1Dl/LSQG0EBPHMk0WO7ImcJaKNH2H4CzJ7rYDEk+MDYYGtEW+sx
vv4AwlZS5HncD4Z15vkp78vw8fg0v1zB6m0ytBvY49y2RMPORBGLgQw89J0Ns/rhuQnNpMlbKWM8
6YgGsePxhBL/p/pUiskrCiPPm+98fov1UUIlHsdWutct4V0h5Xf0FeJj0KQdBfdXSjkdrkGRtxd3
8Tzwqd+Alq+nNFau2tnQfutYQ+RoT0zJ8YKyHom2aqL0fVICUQCj35uEKEt29zkNAgNH9lXsHhJW
MQXL5cZhL2E7EkMfjiyGLHyNNkM4em38KI8xeXPq/Hx0bT5zHgr844GS5o4+pQDNC73Si60ejkjT
TMRIXWGglOLVx/PMbmDgdSwflZ/vafYgdFHeGYDf9AsozykLD7IbkOZsNBqL6n2BCWhhqq5OwaYb
3WZnkDsUSbRWLeIQldw/Rk/+O0OiF9O5Se8oq3bDmNAGwThWDseOtD8mE7ZqNg/KItxl17AAcNiY
zSlNiF/5NN4jSNJmgogPs5jxN2OapJWKU0svHsFJ1CrZsPLyvUvAUeh76VHCb0JIeMVtljn8KGov
3NjjOmdPczfzTXsW6KbuTXVEgvN2mlr9dAp/xNckSK26PtJZFhXkFZbqzYBw9w3GhRerueQdSWJm
SQCZ1JhIq7/xvn28vLEvwZyQqPEpzbPM/VmWI38hiv+n6dHV6uZdyeRcc2/pLq2dC4rdbnJDYRY5
1PcHNVRC5rEcKpGyQ5xOyUAQOr2xENhow+moSa5lhVoXcmWuI4W2hbLnVVgCSYye0amG2fDb3OzV
0ob5lKhvF+x1qiQoxPZRh8PH1FGfk8RN/L+XZ2kVwcKQGVIkYUdITe0e6ubiFJlelxw9NOBTCx21
vaKF/ziO7yFI86E1Z1tN29t82VhoHZh1Cb+IXZFwhEDmozD0Ocx2bYWnhxKmokhYu79BzfUVu1aT
+cqXFEFCFF77Rl11VnNRWQvTizlahsod/IJqadWkRCeNEwn+XlpCC6p5gQHjJxJJMFp3Ngerq1a5
bkZLhSXGjHcFWnQjf5KvaGHQrdZPjdi+GvQQIVahEaZ9qYK74adCaWqXMxLeVi/Rp6hiB5/+588C
3KbsYmfIv0nV4gkhhMK23uca8PMP+uGLltOq9HkzsR3zcbVVZvAgd6Ud8v2YV5pCy+2sfh5N1qg0
PRmYWsyEJpXthyHtBWvcgTv892M6JyH3+tyBuXZo2ZhuerHldCon9rtizdkZMuAZCNqSJa4iLJFV
YOQyQcv/ijjaVGXvdH/uEhZwaANablh9u1tqqoi8KOkRAQkJvARFfuxQP4s3YOJXf8LoWiMPBuov
p01z6dBNXavo4MnPD6qBPSQV4Kbay9Yuo9XPUui+2VpaszDjhFGxjjdEYAVmTvY1lUpDu4pgi6O5
+VJncNkeiWmbqiZjHE1i4wE9IOytvqcKHVPyCwu3B+8gQqryPjTGTlm8aRt8vkC+PHLbnpyG9v5Z
ZkJOh9yc5Y2jnP8625oKG+q7auOqiMkleIOLAAe5k3gOBd96qkmoZqYxphuGkwNnSJjYMifZ6dOm
K0abvJJCOfeEkF5U7CAhpRv54tjCCzSYsC2X9vG6fpC2fINHJ60A97rK/xchf5Tf9okX1TwYUQDe
VRWcyIbPIKDjT5Q1rWC7TTafqVHdCOgTFL2czv691CQr1U8FOabNPZPw1R0AQoPSUIezO/JFeaqg
MMhsI2c5MziruAy1LCvUx2hP/NfjXNib5lscipnAVmvAMeb2t7xyj7zto7Q7pKWAqTFZTy3N7oIL
ODGL7iirUWTmvol8KcA+GKaogIDTCigWETXIlFMGvKKNkT3dEkGP2UOrrB5mIWZggcBjoThLHjq/
ZJAERvZIwCz0SEU2KU63xD4sSEdiN7ZQASvyw8DzSweEqV+yhvWbW35iWdOk1caNgIrEeoCEowli
cUBgwsvkD17qfJWEcZWlGaEvN3bDuQI5h1xPpf7wZVR5krCvlMa8Bn+KM5ljG3r9n1oiA38kh05G
IajadLYP66T+8YfCPEMDhsHUwfPE72YlYJncTxydzcwwN7I0kkamU4W0dNX5Akd0ELhZMRKW1Ayi
B08GecOAIroYh8Ks5583G0wWE1LCjT8xQkuQzkLVC/2VU3534mwenjPleknAKBrjsUAKW+B1MyAT
1znJZFox2W4sykUvJw7Ubn/eNLw8tqsWLEfrCUVJONVNlXvXajPLRanOkuILXeOcKIrpR89S2FaR
dt2JS2yuX6q8HLghFdEuYmnsm9eWFzOmqqL4q15k+XaWxe5EPbSM9jJDAVgwb28OlPNLJsZAw/53
stcphi0+HQxW38UZN/2YhCdcL27PY8wiwdl9Aq474W14aXjrizkw120ASdRVJimhaW1ZYk00CC3f
9FVE4UgLb0l1p939MbjOk/jvDk7K5dvexjsjI7G+s00SNaOzrw0MZ+88O3lQ171NFoaOgIi5/Q4v
FpMbqtF6gXeLhTrLjEbqQ1zht26RbJ4Ex2BHWST/zwYB/W3EP3UdQs9uVVwWvHpYcjEHkkPEBKtj
o/MI6FbQTs58XhmHUi59tJjmrBZ8MvTUriee63nl/Th8q+MM92lQiSH1UYgaX+zg2EtkEAGXltJv
Bba0UEBATw2xsrfR8Auy8aX8D//uOcdXK+ICRMF7dPUgkLAAMVLhGIyEiiOWxmXY1GMpf/a4hA1z
Qejx3IV4hwnK1ca1vOAvdaJh5qZjqZHm3ZsUxItUX246JntexINaFXXifJSaFJGefgXzSmcnGTgC
yeIeIjxVKDQOaqTkfAJqM4tlLDtdVhBiQmAtYxMTesEDc3kFssLXYODgChpk+Tjs0AX9WH/mD3E6
Dzx5buGOH4f9g5z4lhjAYzMtUYHOABLuS/vQ8mZj+5edszrutDN44ZmCslFlPd1Q213mmYxoBBLj
1BDC8gsVZQWDcFkvsBmxVAqljyVE+oLlMzFpE8JKzTvkLbUn21mrE/yD84mh8to+9hdfqjkRJ7uC
B2TENeMg48ovqvsVmgvsAmX/GGcA/9cLL/twsj7NtdONPKvK3FJS5TOlpt4u5cbvI4IZpyw9jkC5
g2zfP1ethw7NfRLRC3NJljhIjS6pFJlfc60k6hzSzsJuGL/Q2Di4RrfPEf2vDfR4mSLLaFjFvTO0
ilfD6sUdbUQ6D0qqL2PG4r4qQ3HZ0Y3gNANoCU4b+O2MDpC66p7W0b2AQB6hV/t001S2mvXf+dYG
53TfO/51RngUNxJfvYISoW17ouGlX2G/sOSpoBBKfEfJ/gTjByscTqQGUNw6ZpCKmB3Aimy4YvCv
j1O8yEdY2KQgj63sBNq0+NJ7pBMtwX4xmgbladVxB0LngYeS8/S4gdSHzmdHCZTmWHCUThxbl0YT
eYTf7xuP+V9NXA3McPxJLSDpyjF8Zp9rqUBj/YTbGcWDgYTquo5svRoNJw/MqotIZ9czuGiJW40h
Tj8KgMQgdn5OxTwZJDbBunzWfAIxu1nszwND8aPndDFhwLG0PJL39lMmh4zQV0C/1o2IeDwVbHpZ
mtGsi/iVAo8/Vo04haUz7Uilj1KZZU+7ws4C3PnRBpV2vNCptO+35zhhQC9AmZgbgQTZoKYtfnqw
tRpfgzFmSN097iQ3b1kLwRHEmmQ/l6BSORMZb3k/f6Gya0sJgLaR5K7NAZwXBRFVaVNRz5szginT
UNktuO+d+NYPydFtgcn3XofscdBn98c/U++dpgV0gyp/PBoK2l6nHbgUTHq0K/mCbF1X+DuOp5Hw
2v1zYAkwZghGfCDOisr1CunA6LQDRLmuDXXsooTjRTiFN4sQXuDFo9aHwrf7vVUNKqrkkkp1LFgb
Zc5eI1U0t6PcxyPZTTk7oBbVg9+IbiqVA7eCYQJD48onnzsBcWZ5W2gzj5ZJWYzxbsIESmVvPyF2
nkZHRzlgpluhpFcHFE5LO/j4Q/qFqcNGacJrAzo1vO/KAsJStOiNadmFHLFAW7funkx/jRnWQP1j
Q9HyYoK4AOE9csw2Ti76jc9FhM1jiyHCiYTaHSRpXG3WB0iJWNUcdSYNNBJe26y6DoUJzhQTJ19v
6qKyfimwQujfvKlSWDOk861yuj1CSf95Rrlo1qAe+9pOI7nAvlHcIcuw9UY8e/rVG3wY4skUNz0m
MLdyFlxuRsAo37ScAALAOqrxwF8I9kDYBrcY+pNqBVw1N1ovbApPXTJeOurujhWpfJao2gQXkUkR
UkbBPa7hMvJrFm1wNVAYpCuyOdFcV5uJzHkdRAJVreVQs6avHLtWbFN1Utrg3jRrRRCs8fws0n9L
PCF8QR7AqLeUbPRM1Ae7BxIDK+mFCUQ5M0wZ3Vf8tHU1FwiPaGRy9HW09CXbJ4NXYtaF78q1jAEu
gPF8WYQsPr5x65N7AFxlB6i3upgLon58tkQ94LE5lf+M4YT6MgxIZUEecDoGadG/AUxDeqlvSmaQ
L7T3LMEmvB+8SMmfSFiTBIjERIaXcJkwOfnJc5N6VP/Z67Iv43VhcPUwiRRBwUgWJKJK32SJb0YW
Ko0lBZLrI1brEQANv3fg5YRFQu+EcUraAYvUwFg7zYHvUvwpzX6XuvmBXXZYEo8KqEaDSpcxCQCF
/IBNMb7SkAfbqyWMckyEIUTM6+uqB4KspCAgtpx6L6p/2RzGVUOjLSfQH2HSJ5+/XMDQd08w6Naw
5SXlB+jFFiL4arFOUVj4VY+j5gNC2xJaq5S3zUiIA5sAer9SC4zQEeqFo+upmJfiLUIIsGnrGOmx
h5oGRcjrywcUXS/CsGg0fGo8PEcP0RYvpMVrKl0jDDO9p/J2ThtlGU6YR1SC/UHhmMzXOm0hRftp
hFPpsJKGv/rhfTS8XXsBoRofUu84bVTRu+lyi7q5gcdKEPObarJcYFIIXXY3kKIxxGtJxAqlvfQW
aoVKnG+BFluXhyD+QARry2clECpX59wjiwx75o4U5QccJqrrnzO1TiAgfwaEHb43YPlQbUtn84vE
qng2kEesH3WM1j8wfyinpzhVgZCfKT3X41cZnRsCl2HUVjlAVfETEVctd9YPmIunn75PrrDj2k82
9dMpa4/TcjtQb6kJK9yntgnjSLykhtaeKfJOUJxUw4B4bDdj7WJ97qGKJgpPsCOrmeliwlGXoxq/
TTpgw1m7RpQE2UFQ6BICkU5S9KUch02m+ruizm1G6KB+y5Q2KXqEIBgbLVMqc3STdwbWlcgLPhbv
mT+RcPp/z0t0esOrzIY659wTwhjctKw+UJ/VA9ixrZ1NiPxRht85Mg7ye/PTTU89njNL79LrSHs4
QE7vt8tgRWGdj2YhJRvS24kXldUhVlAcSWv10bj/QNZqiy4f82IbuvVJW67+8UHl5RZsmcyQGyAj
CY+JdjI7M+ifV5o8iCqhtEhM3LINUOJMpTgN9xlZnBlBVPRo8yufDAdECNhz3vs05iL4sxZapYiA
IeYy5T3ASki0DuUQkZb6NeGA/NnnxaEBmBG4wnvsOtCthv1JsPyrtHfFbn8UlQJmVpw/jRE7bQId
lRs4gtj082TQAEJnST62npnoeIHxzSKiGabgsls2zhr/L+UFrnFacdTBa1HHT0oRFGYS6qrAHxyF
wzgmqpz0qPuxQQ0H7JrhlJ8C4UmXXd1OwNftQelZqn3R+cKXfb94ZxKmW6Bssu/nmfP/Zhh7NNYl
S0o2gxwicaYYPXs9kdkKCbmejBuOmRT/a56OAAP+/OGkGEs1DpKTS7uFySJQKReDJ2v3ulcUxJnC
na5brPeof3jNuIQLtabwByHoSjN+AEGcFzHIMzZUfczL/O3n9USmdZYsMCTpR2K6n0UQgjzrg+Ls
X9xtbEN7UwgdtR38ZYb3ihENaAqrTdLqwMsebp1/kG1Y0bFjiFU7OTZBFU/fTWu4R427COFsf4b3
Mj6zN0BPAjOyLEzK42Dz55I70ydkdbvY18sNXXDYSMaPIJx0FPE7o1G3Zx3BthYHAlLg65u/SoAQ
jA7YpLYwdAdJiR/qBnHPQjzt503HWJofgvDNfjMvyTnu9vrl/hPvEQtbufebfU3rPkMdWOBPQbXr
PW/7AQzZPEzmXebQA4PMMdfgR9UlHxCSNzBJHgRTGAMaZL/hzOXClPsFj6tPGmib7rg+Y8bRllqK
+DkvYZpfYRTUIRO9z16SijzTui5Iev60XWKjbeI7gKCfzhBnTfQbDUNNlpKaS4GoI/X8sWJy+R3N
QLoHSlHE4uXZASibeAx2nLvc9zTE+xGTJQ8n92nzos7b4RFKrEdug64CbRswvEshHSw/gQskvHC9
W4VRdLmbpll93lIMKgwTDyFMF54BNPQD4dnTpAxLYUivEcE+On9Csvk5pSsKgEXwmAUjxqguijJu
gPDLwaTu82WDJ0IdjtllLTEf3oYf2K94LtmXfLyCEb+Qs+p2WOVlPhiLYbcbpOVReHOpFb4AzwI3
GoKRhw47+V/mHUUSzmA7K/nQd3nkWOjSURliGSZdxQzeKpqgFEFP/OZmfaOszX4YlHqq8SDeNweg
lwEvKSXXapbALncXbhntMGQaHzMp4h6xA9k16sc0btTAIV5BexhdKQQzJn2mhgY8JbHatT8veTGR
LfpdSnyUnJ52FEpabhFiRA/WB6a/CtW5Ccs+9wKtF03UmjCiMLp40uzTXCMHuehu//cKBn+r6BVe
M4womlci1t9uIeK0Bzi7K5BROeKrsh8X9n8NFwWlobfbxi1JmzMRP1BOC3bMBF/OIuqszvvAGGz9
EG3zldNQk9OkcI9zdxZVO4wtTXNjwJDIct33b+0F2y+/PcK5e29MRh0Vbmy3WqYmpQDe0ehAZ1yf
XlNGYCbdB0TJq79mBvPpf1X7mYLnrksSDTdv/y+uGM1F+n4j1ulq6YXcU4TG9bn/8q+zdNtnNao/
EJIglWxSj5vpXdXt8+/H9XBvsXH+YhaGkE9NDlEjHS7bZWIF91dpBnzVhMHQtYczPBalr9goWC4X
1PnXQG5ReiAC2PNgpduSLj4y0/H8azWrVuhdCPov80eN32BX7LETN9pJtqlZDGDJFhnaB4LnSnzx
ANRkUTPnzjhYj5k0gQ6MvqhEb9u+NzmOAv+JvaFhA/ld02cexzkrXZidxuEu3u75NNnlgf2xHsf6
SNXYeaRkjrnPsbyqjei5vdDEsdIGFEStpqNOutua2IVP9Wm3UaHm8AFZSYyy45lxw+yhIR7z+D+b
Xce5VIT/ShImB0fPgnjFCR9NPFQwcrMbPodNGPhNoqNKBAwXl/gcGQAChtqw+vlL94BAAPch9rgY
twHWPBbbyWXXA4KEtiqFuZY0SU6m8cJ6REoRFFv7Qyet0fxLe8h40tIjKW9QBRpLrSLWMFEwputU
+s7soQmjh05JU5tlfwbNHMQk9ZOXDJNFu+7KAGthxnUp9W0KFIrsNOFp+lvwIKn/ztQQ3hfzmfd7
cRZVRyi9E48dlJVAQiBaNmxKbgCKgDr6gPLPYo26Yqvt/aymoyUQhMgS19SmA2ULhhvPKIVKf9jd
rTQdYmGm67EvGVg/7h75tJBfSFiB2SmV1g9ZaWMsqtaODxfDl6MjKI+CQAuICf+05j5eO1GBGEHw
g6CN942xBCVwk5QVb+zCwDzGOZH5OTOgSul3QqBj81EY/onHOl1dhfS/1ZSDWaVVY7ywp5ppT51f
E9uTZWbl9rupLKKHYozOO2Uacu3/pqj5OExTAuCYrIZuI4w2hM2UnV7yo6Mv0gqgIPFUuGqW8yKW
B53crF28rHP9PDmd4qxEFiCP9D+rRLRXwymfMbOHJcOS2Dw/7CpxElDdmt2Kgs/ipyKFt7wGinCE
hU5PUkZ7dbXOI3yqUaQVaV96TslTppPjqpumtMQFi4a7v69ypu9cHwbn1vGltN+6zckFpDhIND0x
4U4fVukHzjbsjsJrKZnB9KIpchKg5gB+Etcvby5WQfTKQDADKsiRe0eTwqlSNeMst/qNTzGUCBxl
pcromF1ZYt6+s7VWY5rP0Bhj/Sr3lqEPWusGZqdt0+qalKgoQWt86chQ5h3JhEntzjwcdd8XmpRE
WXFIUk4kfrqBgND9+fFO9Qq8O3ZyWj+1n0L0qF1LvOyfZ36/QjA90HIbkQxv67kIvoFyDG45nBTI
bdWcaVSEc++88lbDlTPGO0aQUhcFDzXxQRzGAd1fy/npe9Vv5+k8W/fvH9dglMbRvOYjY7v8SxKh
LaCHiHfxb2PcAuaOqk6FGbM85/2ODyiCbdpow81LxBTACuXXn4SyPZRzO6XHnuhfDPCBWHZeduKR
bUGjRFq54OAOji5JluZGKDf2mEaEP5WJFSRf2Xlcndrn0BGM9foV8wDqcHgeu52soRdCHnL9OB2F
/Pha6FebPZkBHO5O4L1oQTmubz95VkK4AuVPYwybkJuEZvfuyysstzUI/k4JclzD9QoHJwksyA5j
wcJdyCw/KhvBuBsgo/Vbz8CYkRajllWArGfkUNpjTxb/pzAUksFMnGmkOLY/B6ELxdX5A0vaQVKo
xhCqlQZZZA8wXUq8E0xCae3O1tqOQfIZ9zwqPpbQxy8jooF3aRievD2q2KCtYdMkJ1bhM3BmLGZU
O+VHqimKHWJYItIitDlIiMusKeQDpenxig/xgcMoB7JvPlkGLFAFdLBer/Y5atyU1x2i0Ho4Dcnw
Rnr0LN2GrqY/t56XVJ6ePma0CV02nCrBqWoTBT8eaVJzHocU+gMwtaGxA2kP52EM5u+s7Zg570vW
wOnXBTGCI1t/PNhk4+hA00T3dn67FiLM0Vycyw6rMJYI4X1CRBo2Rhk/LlGmG/KAZk8vNgbbpgOg
130ubgMB752Zz9jTKDeakCE7wPdzg7bdeNI15H6RYDmnga4Tsxl5bCka+HryW2Uyj9ufv7RcaK1J
ZWOTLLkkEzPEJb4Ffjzt7ddfUIhN55+ArUh7l8OpWdLhHhSlWgn7RPBxc4rUJ/AJBqBCfylttAmr
Ja6P6r0fKWNoTTee50ZPQs4miIt+JxwY8zEeQvxUBvF2/EXCImCYnsgY0tSVXLTR4AAtQJZu5eCl
OcT7ObSRVktKn3YXQlVmvFSi7n9qono+ilmZt2tF/H8q+YnMb7gPiHKOrjroPLw787l1yjqx3Lz4
RXyiOjpdzjbCmr12ndhUkGwIZhwnA4jWF+jCDwOuvW4OAt41ZetMT2j4nIVbvshHYEOqQMMff/pU
5+Nfip11Z67sJgwaQ3HO6X/dz81li8Vu3juQubCDCfliYNEAl/apNFwJMCcXidsuq2X/cn6M1ope
YC5dyUP/zHHp6z42xL5vHFeeo3MrbEFoBigl8iObYDqw05v7h8LsTaOoXSFhTVi7EKZu51aPXPWG
IjxjoJK0f5VYxP0YNg79jrWqZUqy3q/STJuy7cLj1tDxcHU6xF5cKtyb9NVO9JSEK3oKKEokC66P
QEOoiYuB2WMa73urNQWKcLuAr8yIt8LsiWiWO/XW//GUFV3KnpeUFv3CMvbih/XOUHND1KUwi3ha
smonBQTB7SdPkFXzb2qoS5LAem020qiLYAASfHs1RilES3bkfxaDINq5YclIaRJ8FIIeMiv2N98o
IZBrzMAdER3uaZiYA5cXAvaw96VgfscBXAb663sp3+dC3EYCVbhQrHSISRECi73Uq/38Z770K4Io
vmTbN1pFjAFuGqECgdYYLGr4eS8YJHwYsDDd+ODLjoDnNvG+SiwRVS1oSRN2/96oHThbOG5H9Eht
CzI74gOnwYesnHWGdOYvEITrim4JHWuwrl3QY3WCyKn6izMyxPXXDJ2esQuBL7ZHiHoVc285H5iD
nNEoQVdPSBWV3Dw7RPPnjEQqVtkowpYrmfc6aS8VrtjTa8oe2Frtqn+lMCbDsIR/JZih2cbOSbcE
vtbcM1YlIkC0xEz93lyDDb7IN1Mm6q0uGmm78OF2mC+yV9inS0J2Se/BRhguwTOLoINtugVTWC91
YatZQ0EsW9psW2hpl15Y3gnPOaHRUxeVoMLIc/wrRk87YCArDg1yPQhWBpajs5Sh5vWMhz+jUm10
nMRbdq5UvpLgWDsAYkl0NCsqvxaBFz4AtFmc83CdQAWr5vAwFEp+lL9Uo38xkHCAAjgj6aYASQH4
MXM0MU0UI3pmP2e6Qa+clhZBJVDNTqXXG5RPJvUCn3YJltDnsE1OfXaCggwlmmWsVodWRmRfvK9I
z4Bp5akLnqKUr+UNwhfQVcGv7RD9eXhBwVmBjvcbnlFOcWNi1n1oOjScBcOs6LByPnNG1BOkpRqO
mGvLdLXRS2tESfyhwDYRmy5Q3dcm/9UWaF6CWxWDn20BrtwtaBo8Bwz0N+zDPtOTgoWd1WH+/5/w
GNqypQkedLOGuU7dMk8rrA9cBkudGKe7egpfJIMCtojIlG63P6LtZ+VTIAtO4PN0WIdKDc6VS4EE
/XSP6e5+g22js7ScXaOcgLzF13UOgd2XI8YvJNRhYR5TrLnhYYnN6bUf+XmEfgFzZhCG556GHDrn
VgrsZ9qMGdoulvztE5mwS5xxz4dsNMe9KDLIjKmBx7axr3+d3Cl6gPJllRufp4WXST9rb0BVlM0g
9/2IeZBctsCZ/qnNT0xECAxFC/p09kgSWPQQcxXk9+M4wC80hW6AkRcY1HWcXZwcKjzDwwxPjExO
vmLEC6bG9h9sdfSTAaLK+VDGDE/8QLJYpXZhexn6dvOx+tTCaimAIZfB4ZXFlBKgRne2kCkV4txS
mUPo4LsOyra2c6ccw5gPRpDRWv7rudY766POBKfTVVxPINYfLWIKMXy9I7E6mrZGL2XFaG1G8XYg
arPKgIccmH86xmgCIIxAtHgZpH1cpoiWPoqaU85j2rTpRnbBML5DV3Tr1NCEsIslXysUM9m1fDsn
mJ6HCiZJAoygWsYLjys+PDUVY3RNZ6d33KfOaYK41PH/q5vEaml8JIHeRgaed91Blc6/MDidnRrK
TQ7yMThbfXFmo+iN141ITNafWJ0JhxFZWzjY+YK2pP+RjeaDO94tIartaP9ESKcSnfnKefjU/u5n
URfTcTZemTGOlR4l5LkqB9Tx6WBHzCzvn1oj5h+r7xbtcpf8FumXsZpFLrDtkPq4gKXPm5lA71Jz
6ckB7QT+Tl8iSjk7bfEG46m5taiLDWcl0M/Dgki9UhrLhREG026jhvkpcoj7HPi3Fq0E7bt9VWP2
S7NFT7X/oU+o9qnxLAsVbu7TwNjlAAuXIdQk9IZ4EtXiJFQN3ppJd1oOwu3QsSfE77AU6JvQHQKY
UwK0fMcrWL+1AjegKmr6AFGsVvhvmn3SBUof0G9dMwF3Gx+5pCTLNvvtwTWPbVu3ap1dUyIeQuiV
FB2a0VvelyYEfjXoMjd6eM9yrxQ1SwfFxdOzcyn2+BycZimkMmFcEHOc/T/nqfMAEuwADMLHoNae
tQXdoJo6S/TMth8pvGAcu/g0WzHRFS1YFp5RdOd4bvktVRmCf+xMFqdS38yAUNkwvBxUsUnBMZdj
OmdHQLmmTmGk1Z++JPMWx5lJYxZStqgkSZbw2bIyTtx7JNsu174sCofE6SpgdI+UTsMxDi1vZFqv
AJZu+PqQo7qDqJXKvJT4gSxf7u9wq2Q+YSFaNu49ITFiJP+s/SDcUoPJJdSyKD4vc+N4cphYVLJS
dLRZXFwZSs/2KqQcAyZPTqMlSKlyefFmoQFPyHXmBzsF6pCUOHXx9eCpleAk7SxBMa4NGmpJWtXg
ipI3aeyxYw4h+pV/KP19sc+XOBUuSDUIEc1UkxHSBr9XknqvDo0Jj4uXq5BmEZ9meq9TmaisRDMM
MtkNzB+f6CeqrCdvCAmjRD1m/4sMgYjbvg0j+eQTUNgacLbId1vBLoo1r9QWT9Q24I8g0rodfKNp
c1LDbAgJwApohzzZwoMzv59EjKKBFoW9axrSWv9fzkBkz+oc1BX6IjxgkgfDo8TJl8tb8u0oqhoZ
AatfJ7FirWXrNXGyUavOIDgK/mEQUejOlEP1F56BoWxe74cOVsvR+V7L0KDjerx8sQ+C1p0LihY3
3Y5qvAiAPdlFV+Ei32oYzYiJ+cuPAM7gDbQ8m+25Kvuf7QO8cUkI4hPt+YGaw1mQH4PODK0RcdzX
hZa8VJIWjV5IdZbQhTUSGb34hjbypOxXVeiD1YAFYaX9jVEcsKyKkkx9xMMlWcKAY3yTajPiusCx
dupcQXadZWGXJ0HM8Wae/4Soc6lJCHVvS57UQZkshmh58br/gjSGUu/uN5kb/7U9wbUgzNPcwxRB
2+JhuC/pXA6tqyQGh6ZR07JblO7vsPoQWTI9HbAuuDBt5Ik2rcelWMSEUpbDelPClUzLvdGpjxMH
bnnSTs1XYZ4zxsSNukCdZfy+k5nkXg1yazTEHzp6aZzsTjHwT2J7IUNJ7/jGLoeflMaAts8SlzUi
S2Qdn4Iv4+iovCV7A8zOWzkPIkfPhGhkVhBCg2Fdv6uyzjJIPDYO3o99luwpnXna32RdtHKv+111
hnD0q64VGAR+j9yx9m8R6Lr8zjp0jr5c9c+hyyNlBJTmSaorbDxcnL2o/jdA8ppJt9Sxrn0CoV+j
/gnJEdtuzqF0y0lhu0P3E+2gN4B4hviE0OVDrPcG+JeO0IvXn16RO+P1gNEdiAozeqe8G3zgGxSv
6QS9GSB56Ocm1Ch8BgtY9yX9yiLS7huZ7PUcS58cVYttUMgjrTCFt/H/LV3rIuvz3AZYCyo1QXiO
TVMM3iS2uS3O9AmKRq6aAk45TcVWaJ4aet4tlAsaoeR6Vpbg3Xbw7y/v6nEFyBf+exDv+bBLDDQR
HFJQ+dd2WFnXj0x9FhST7i3EFjsEj9ED27yyawHFtjOZ+9vopq6VkzzNse4UHdGRln9Ayq5WKjOf
yJJ58gixMFw4kNBQDBBgCH7lzAnDr8Y/gHfpVskB+slZJi+knkAWKkxaDV7ONiUuco/tZdFZcMj3
bwaGACo+6/IUrCoX3zLBrcOYxpDLveB2Iyq9LIMo5lCH1zreQsV1KPc2DcPng4c2h6yovdoPcLcL
qFGZ54fYL8IsezBBecpkdGT0gupOTJ2r1SIXiWPoPOn3u9LskaaR/3TJMx6wqjDIOxRD8P676Zab
GBGQIi1ziqBnRDYzP01l6QFbo/BV1accNocGURbGQva4VuyhVExF+Nj0e2kTdbgEactLm4VD9vuG
c3RxEvrGS5m9KF19gj8f9PaQtXZEl3fTcWRUO2MfNi52DWiC6p+rH9H5UTWCkzRiHcX7NTmerpQz
AMe4qD0nz2Kegzucb5De35H8+m5BGgPMfsQn5pJrVUs7cD24JrglsV7veOSW+l98G2F6QbXrqN+W
sj1PTAz/1r4V7YV0HyagiIOushPhIfmjYI3h+r9SckWbxFnZL+OFL8IS6FJE5ivO1LNdALPPKhk0
sXVLonNxIy+r0aFiztz01CQlnnQMuAxq355VRuQ1dYEUZWscDqzuh0cuFH/S0O3G+CzI7T5q0cO0
3P1JDiALXWplRM5Tw1cxbZ7QzSwawiu8d8H+WshXDGVU1wfKoPqiUqZI07M5jcNEe5ltJP/c6YqC
2+ql2xYXSbcdEWhN/mXvejJ3I9WwPcOnGX5XGOZFvVk0R4Vj2ELCNyINilrGkFLNfkoVFIS5F6UA
ebf815qeIddRjTTxBeoJ+h/Qtjd0GxW+zWQkgWr4F3aRxMQCywWtVmWG23RkrvMkkwf8ph+ZMdoI
1yQK4axzN1s/AXf/WLJFi36vg2LEiKyQ2tT39UgtrgFCmvQFTfb24Zt0/iTXWV1A9j6Pd0tKLODr
A/dhKhvY5cUC1R06dTa57Whlrsi6/KS643WtzSSQ+mLWvKFwTosfZsNo99XZzf+L3gIm/AioZl3E
X73bhu4Ho3LPWIDKw9xoCIBtvCSltSDRa9EWm3vfr/0KppSvs8uVWBk9UMeU3xPNOuSjpvVw6uoe
edbAQLVO7Hokft07f7J7aW9TqELrVmEhvOFIPLgOeqvjDNAlBEx3SJGV7OKtNl5+pXRuPYZl16Hn
pdMZloxXzbwHGHpfE870RNTMN/0qxKQeBrZfTA1bPWPq2HXSToKiqqxi+/AP4zNPmrJ5Sseec4CR
df1P+8ye8vpHeXZhcuvzJnzKRuuTmp+rOeIAqfTneQkHzTFqtCgOJfawEo1FUu+hJCaCWSgWjZq6
TXeDFbMLe9LUx7tknw5K2xXb1ljxR2mtOfI2dmix92S/VbBGw5TvPagp/fo04GxF7bhDZGN9erEB
kVAqEgjVi3ao5VHCJbJYL5qKAHgYZH+5S+6qGApgKpCREe8knSeo7rMqYxAhW9rIpKs+ez++TbEw
tE+rYtRE68e6Vy5hSn74sZPkn17YiwQtYzpXcNbPB0Vr5ysWTZ7etVoeD0s1nYabMI6teHbHg/Yl
gUifin8P+hXE/QlVLbOKmIZv700nu02+KcHbQ6NHdLOflVsC0TJ3PEmGAmiEPLImyRNZxAvsImDp
LzXRLKplc1ev3tHA8vu7GpqDVlQZ2aiUTlJRJYIwvpWIp1xXUr7cty04LiF0pMOg4f1DrzK00R9F
RfciJSJ1c1Xs38vtQNFvKcergcIAplWF9uW3AiaZzfGlY/hrfMPMic5oReyladbSB1GQ/9hdKahK
t83De+s709nzyI21No2RjvkvY5a6rCsqkGH3p84/CJPC0C7O5ALXdEeJ1O6O0sXI+QOBuOX5HoC7
fqYFwFl14aXwnt6MBAnibROOmv727hRXH6QYzwjjOk3azzN2CMohcynjOFFYCoQiyFvt32GYkN2L
ENTTdM/M22zre0XoDoApVv9HdvyHIVYa2pGQAbnffh5XPexdFFUbkgtS2x6yIlUFOX8uQze4PYmm
823bML3PE1AM7oDBelvYeA5He6akIjAyldIcVjnT6V9dgtwcy7NIFeaTsqBT3Dv0TXhZuMyGmr4d
LTNgufsglkHN8tTkPysBSTu1ZEpvLEjevfqN7YwXHvqsVo0kXJud17f1QtFu2qIz36Yf0QrOM8Qj
uO+Ai+Q5XiElCtmS2p1TpPpacUBjT3yrcLWI8T6rdAxH8SLximwFU8nvVO55qodQHpL2hilbxuNw
lyxG1SNMme6tZ9vqiWgPDuoqJ5nqhEFK86dJzFP9u6U/uJVGIXxRVAXhcWoZMDgLjRT5TlwmPflY
qUnZdS1zTp98mpjQrw4KjKsmchlJBz4udUrpXb0iK5LbfEDC1S26kl13t55buEw4Kh3ZWG71+YkO
K0Taaf10Fv4HUBuz5OxCw6rZhjSczxREloBsj7zwRNPqlTjKMZ22+uUKtwCZjXIEaDM1aVpkjTm5
w6UoVmwKC0Q/7aJezyXaz7skhAN5YRlDOLVeI9Ho4fJTBlI02ZLzBfS2kKBz6LYASal+CQG6YrSZ
XogUiqFDCWejpNBEGOD8CldfQkH34zVfnsVjo/KuZaBuF0xr8ZW1N4duBo/nqAIr/smgUUgCOBtO
Z7piVoi5bqD86VAH9jNXXP+GZGXdP/aexKTqOXsTokQzEv2Kjjl4ymuggd5iJFr6gwwX4Ko7T1JI
HaZ7YsbLIBGsJw1swtJhp6WNAjk/EyFHhaYF4yK3lmJSjcxiDTAlgHgTdDZ86QUPmL3J0R3amOAC
+V4pGTidI79Z7613ftV2c92y805d0EYmeF4eN9lvLfPlF2fpAIVpbFVA5aH4yeieNA7HwNlsg7iX
tOgLTHUu+XEVNPgWTv6l9KrSWaJGuQl+mDTeWzcCbNR1Cdg2UkQ5ZoIKcF4wR/EfpGsuXsxDiL7U
d1vkmIFTvPIzeJ2e1AadjiDH4PPn7sjmn55i2OIXRu8P+eRV+ZF6B3p/q1O/0Ytag43CAQDTmnnu
Slsik3Q4KZ5I6vJR/Usy2UIVzbhRmiUvDSS8mTb1tMWfDVlRYuSJ9nNQummjx3yeMNjWOJoJ+o/4
QkEER4/r36qwqDuPWGN3/HJudFzbwn9VwGn21YbllSnfpE9Isb+hUzlHbO1ypEJI3q6Zto0x6+IS
u2f3+2C7V8rB0EB8vKlGNNQq7AYCsssLkmHynPiSzDM9TnT+DaQUgjaZDLZBWLYowNkz18rHD0SK
RKzSgf+QxXeHZwskkc274b3iCyTwYCcBPaa9UfjOe2Lf0EJcQBC1bYVhfPpiO4PBuXOhvLKRZMOC
kh/gUW+NbNnig5bYEQloTy1MSq3eGErCujdbVcKbz+0kuYTIk3IzlQvkORS2RB0hEK2EQ5UluHp5
4gI5XonEFeB7OFrqQA1drB7QhYXK5GpEsnnlbMjuYMwe672EV6//048E3fJay34lEZkKXIP/xc88
zc9RSGUO6mxQ5h7CKC9rj0HRO3zHraCNPz6pWnJCMZIXoDvU09txaVff6d/Xmsvi25d52mEYINzh
AEgY5wHh1bxkaEihIChkusisR5bfe+wvuGRlbbZ71wbp3wrQRCj/lAXNL2ChMT3yMsqyiNaOweVW
kPxS7VOo+oRxuH2V+CXnlkU83peyDLjufJStCuuPd7q8OPJfNr4gAzc9EOPRxxkLNp1RbK6hOvpi
yG++YQ6snFCEkKp+BEKwtSBx302AOwCb0YE1qhlCAVZ4duvSoJbp9GM+Dum3E7rU5ADvu2ldx++b
WZYl4ra5qDrmdvmPdaMp7DW9kYecuxt30HT+2EKoEX0Gm6D8I6IqWvGuyZB+XZf2ehD4kVopVHwV
GM49DJU3AKoAqR7Nj46eDVHxPp7iLy+ku/O11FIjfvCdztZuoD1FV68ro6QDJM1fJp2WIB4pbKk/
echhh7N8AqCMDHRIobYwXX0ckaRkiQ8237pGHHW6cd7Osu6KERydeLdKpbyasesqS76wXOjvq8M/
wiG14Xxs8hTEnFaPGMI9P9gv4EYzx3iTi+eP27OTMIk+It4+dVCAQ699Fb9wXNxbGxzDpwurXDO6
UQUQ5kjZRtqtq4PP5r6+/OSsz+3syi17iMOn4k6ijj39i09I71A3U4aYRkdlLJaHxvy/T+PyBUg2
ctUnzJm2PDWFZNSGVOyGl6BhVTLkA8yLXy4xOwskb4S9Dfjqci/6M4itl6byBpsTTb0qpPDaaT5t
wOs4Y9Bvqw6Ih+RNxlDG7maS0R+ThWf8/i2LatjI285hsmunHZhMTMTHwYmoyWTYWxSeOulOfMxk
3K3M5uDIvcOx/YKjH+9agRhXWVOnQ0dKxmjz/sOtOdCTIJKBgDKV7ddVyiCjb6GcdmRIjYcCFWik
oPio5rQ8kiRToWBLQqZGdLXSfPSUndi76e0ISSG+7m+9W0N+cbsX5uHIVCyMlCMEp2mAWJ5bOSpA
dI0sYk/wmWEk3D5Zs6IwZJnsEmZLI2kQVmRSPeCPNYAbU63QP+4tlF55gK+it0IDEo+xD7SN/lmr
FB7qns4S4HtMeeZ20xZMAYJw+hNPJXo5HwbEY0N3Xnqby/JMj57NB39JyNYubJPmaXV7L2j+edWs
k9ZKkoHGGKo7aJ66Ywb/cvnw8WWqioibiQGbL7MsymZAnacj0JIXw7TMcBRri9Ae598xOs9++IuS
obVZ2mEu+VgLiLJOv1r2qSMro9wBGsqYVzLn7DDPw0CdiTlAHJOa3d50ShbkyK0doN+tnnkdJ3fk
chWoKc/K5zMxtfrs38QLb1OmZkXNPbFKRkORKr5b5ielOdcNDlKkLGS2aRmhiGPNKsBezwvn/gqI
o7KypQ/ig1f5iEyuIYmDhzZC9/vmAoXf7x1q87bu3NkJv6ZrpA7ozvvb3qzPrb5Nb8ZXxj+51O5e
HaS7JB2ogRBvaK07/SEszVeJYE7Hw+Ls9Bn8Q34SVRz/+HVTJmVR8KTU9DqCW/gyUnTOZ2zHI77S
QuIQd/HOkU02ztHcdpnBcyzYmSRzLWNrt1YmYFBcostPFmZr17ft6tO9OSvtLqJSHpQeCnSA+YVf
FEmozDGOyycP2YPR4RZzCmdJ2DXYrDXKak6i2/MoJ8IVbXeUEbd+rXlgduUHOr3ieUHC6Ud/0kdC
AXDatjSPFyG09420sW7kgbk3zSVN59Mm6OtMyAO7FN6T2P1VDtPMaRVNCIxvvqilzBdAc/Sxlet3
EXpj90zio3sfI5jYEGVXuD3UBZv7auOrnCE3u2ibw2DOic8HMD5JH3GYCPGq2vsvqndQntAHJDmj
nJSZvySU/mImSrA3G9FtgJ8dzbPo8m+eTXkGLX9MqrWGzErIueXRy5vHEUnhZ/WAtfDMZebnS1N2
vkTtyQuFz1ZIilKUnhOUIN32ZvO5EXEJJrC49T/ovOQw8/tfiz+xMKF6qF5Yli3KzkpnDbMGC8GP
IpXneWyQ2aRNgYDApz+9ctc9/NnIpWrpKxCiU8dVSIOOSUNoyKcx1WjKxxXFCReNamGG1hQT9mLz
32s8l06Gls+lG2ma5BKsM1DrpoWsJ+k+u03+GTYEB6xlQFQD4vyWG9eDJNf6coT2ox+6Vwl2Oa0m
SrbbrLYxNvd6abaQZhkeTiEsMLK1IJP4/N93dXYSl8rtz4qneBCYHNZe5CwQvqunkto0RbEwGDme
xNgCLVsMsvVTPDdqZm0sFMTSPikOTdgV8YoqZa26TAimkeOoS/aTqA43jdbSMTD6G1pgMeh268vw
twwcfwBBaPZ/iA6Q++jUFVhrrWUs8r25qqD3a7FNXnr95AofKnU/hWNNkgktXapo0Ukgr9xiuSzY
o61CGYaRNIV7Yc4MQZyVFdURvd423Ax5N8ZWJhYpK8st59swZ9j4SbssMp/duAJzqHkEfuDv91j/
ew8YywmRxF1fSaKJbio3NlrpO1mxl/gG67WSQfaR5CxfizCZfCWb9R1l4gHUSaBc8MogyeeFOruU
rHVdPv9oJT54qPW6SfGiqOP0hnT/erymIq4SYPUXyhmW4kJL8GoqxQKOFjimyWhEvjbGYbY8/MxL
jLan1LCahlQooRB912UyBEY6r21u3rPP4AnD7JkuGQJeupo0DsOs1OiYF9O+ApYt1ViHiFIFBjyr
kAUr1iql6fBPvhhn0woDUDdC5Nexd47mq0SkOYVHV2+ct6uUtxJ/R6FVQOGu8uHd93vU0A0HREQo
phGjI38ikevPZ7L+h8fLYvOrVhHgNmsG4uUXuDPZx4/QvBQM0YTndDXnoUp4flSMIRcziUqwABla
bk4NhhcKFvOHzwai15zx/QEAx+bht0GCzjbFaGl4sIWbOxH+VOT0i6b3Z0HnnGA+/jiEzMc8imgj
4FvJY+wvuhI7bEYRYB2gxh5wOjFlB9cmiE0OuKKKbd1eJLGM/26jMUSN0HuB+hCZ/2sRKrmg149Z
fHYGRRlWM5pnl1txHAi909rapU11IK6vB0fIk35T5wNr02yKMfVq9M8f1nNEkvk1sIb4L1/kBhNz
nENwYi5sqHYFxlsG0pWLynCsC0BU+kz4BqSMQa65IgqzCCVkdNQ2rTzdt2Kh3QcCYvzPGcNDc5bd
MRcO3YiGTO4ndWChg/XRQEMOvwz0QKu6vMfVvaakFWrZ24tDWp/clneJMVnjPttMWwPbOEoO9PbE
kxSuTfqC/qCWGapaneqCol7iBl+3ggHpcktZh8u7HzEMxrdizemhgiWk2BidCMT03AHCtSViKvX5
BHhj5+bYNzaJCV7VowZZjnGFlbx6RcSvHMUxSo9uqsBNqAD/piaquBu+77Z4m4hQcgf81iX68fGK
WVPOHpomrnuO+47KbfSXme/e7cyLWc7NNdV+4UmWI/7FwcDJfrUz11Nh4OvL4aEN2LE0sqdpQGUy
i0PTWs2z+/TKcXjy6LXUNlE8cXg8/nQDaCsbzcBNJRDbWq9ZazG4/YJxuiiKma3guRXXsDEAZqkd
yGfoUxf9DGH3t31O+tlEdy1eJTMpGyRah/1WU9u9Sr86039UFWc3cnDWjZtJ4pnuEXjeXEAsdRqN
D83fYRecMbff3Jfu0yyzgxUkQeeWTfm5JcDyFVSK4m6Id0ueHKvqXvqgyvLbIE7WWpd5Vn+OLuRw
FPpHoGYR6Co2JnOmZgjfC3dTooIcy0nPlByyDAay1fWDHSSE397OVtnDUJGEyfTjwpz7LZtBtfuZ
qIwzwDnOS9evbjWkYiWxc5XQXYIYrFM1reOCwJgrJ5PFFmaMOp4EU/ieIY0fay+1TpOy2mLvq+wx
/qB5LWcWLlwYcaM++ohBny562NzUk8kFv8bRdK5y/ExmQdsDCrxGV40P+tyVfkoXeRFCoJfM07N6
vUzOPuQ8WFrTr+BS83UmpjarTHSolk2iU9nwZcCDFHmr430+7uUxLXdvGCfQm/zEEYxL79YFJZTj
kapNn6xmqFTBv/hZxJClPJH8ADnVLnS1gGOqpzqmnMYEA2L2hVBIz0G7TFxFinNcEi1sfwK/ENip
MSg4yFvcVbwDIMTIojf1VuskNU2P1a3dgKQtzPU8AkC9rFqf5g12hBD3tv1ahjLOBwtbZgClGZOC
xu8peP/WZUclX5L9c1jrMtE4rSiynFKCt8Sl32Gjv89MZGJVO8nLVBwhvpLfdRo72gllT7SeUoyE
hdqf2CyG/o4dmL8u1wZfdwwhDXk/5qsClhZAAmWNxIPjh3e7xmgtJeePTFhFpljnY6TSgv9e1mQm
8Lkihi3NnniDWLydsajrANgfNyHkFOFAxeNWtUKfsMSjOqZQKZmjA2S5AxOcjHZontyiXeRawXZQ
ZyG0HVI+eLNrGO2JiDWeTk66n0m6j+EDKiGGfmglxbeX+G+43rEZuTuQntyl67ItU0Pvs1/rqsyd
7cYveB5C4I6qGm0W5CaKDgTuoSQa0Y73+TsVGRRsA5RrneIuvrrUikPRoxTFOy1dH/imhE0JejgN
G9DN/nTpYOLoQNjIgc+SZowZJZShp7DsIIoAjYTUwm81rJa9Re45M+jtKTQlShxXsAgvq01t2CEa
Sbk2N5HX1fup8PEIvZBc0E8kcj5NqoXQnwkJIeiO9h0AretPujHXPnVtrxoPOaRCv5NpZQPODnRI
EGtuPgbKwFxWVgQeIyR5NFb6ur/YZ86DF1ZOtd40H2dxJSWTS7eHqhUnFNqP8Qlqu1dmsdyhgfrg
PMlcfenYkjP/y0KMTmgZ/O4AB1cvEi/TwRX70zoyo/kTjqxr8KNphq+p1x+IteXz1VNhIPYYHlOi
t/XhnjH0Bc+GRjf/1mlyi2T/FlDUoyuoyFl+bgPLAznLjHsLbK81G+sOy1BjvKiDl+5Oq9DMSJnP
vxgXeiJHAmL+ZqBtJla4WpEZGWCkEb4E366Jb/ZrnubRxPIdkQZYnP35tdbCuExGCFYP1ZzhXnQL
hyOuUhHw7XZLtbw1IKms+VEHEa8Ot77Rk0eJXJfGktD5dPOdBHwgUtq80rXQXTHUnm1os9038xIi
vcnf/bpLbjhNZw0SusNrlwKKJORwcUOsLtd7MSfi31itZj5zCHhJVnCveJy8y1LqkS9hxLWfpo+x
IQHVvMLyQQpXBnknE6GHve5GzxeqPvfIj3Vy2gEMaggRWSQx1QRO0iFvZD9p9AJjJiOXp9krTPmh
jf1c9HLkh0l+R9CYbAr10LaHPut2xZOPfRVZWodTpzQHgF6JCvnn1O/D5Al07HAq4aNWkpjHGRJW
ADNeLMwtXBK3IrndhuAuPoUsu2XL4rlhzgQGV+Dh3jyT52sSneub5MLcQkUjldHCNxwCuZlAbfhr
23JzRj6r2ufErTdZkVANt9cYyusJ/eG2eYWjEl/1cWRRH4Vb7G3hlTjiFZZ6WIZNbsPGgAelAx1I
ZAg4ro0JXzPGAsAAoyW93C7R1Xar1572AKw29dq7WA6n/K87gGVRCYzMf7PzPsTc1VVgVbAFbpm/
3ktNCQEIhLlaGY54nKo5GfB1iYxNWIa92aJJtrSt+nCxrcQMAFvwaO9EtfmqS9JHtKKRfwWX1F3/
inzh5e6SBsXrKQF73iQDgR+hamFxKs/k+gb635A541DDB7D3+VURNI76CDx20QueTmdKDTlnihfZ
z7DpK4z5vcqr620+gK8YbTfNgKfZH3SAdAO4y+JeacYNh/R4D+LqT09mIvFMb+SRUdC1S0bRbsvD
R07ExLWC5MqdBEVmZs04W9J6eS9AnRLW0azWb3YlQtks/AEVBQpf7g2TZz+ks7I8/EMISGJzPP7I
Ujwem/d1/ZHCOnuOhYg18pB4j+H9udE2z+uPqFC3L3J7o6PrkkHYBbrDCFUk5uwk1sB0fRL5v0BW
p06IK7nES0dAxT8HghLkDIZm5ZIKHkuNB/AZrKm5qAXfFxm4CxNUXfRZEApkc1mdjI9AEnGcsSyE
2bBKR8VxvqyfXoyv23U43J6ROMIaXbYAlp1S09EX/4sTPdkQODdssb6XpEZUu5utvFm3A1JHZGD6
vPT9k6MvOgXGEApUmKsmPkrcXxIjvsrw8NqLc+GATb5I8qvHvtO1+Cs+F/rycwqdZmR/7i9UmJ0U
SKlximH7aFqotpxalng02+ZF0gG2DbrTVnNPpHqknJO+XdO+7sXpNRhKeuYCaiGh1dQW+bkZV//4
odKmBeEhYjawghqy5x0nYTeQKk4ZGU7/c/Df4pPOhIGPvnQ+qoLhwthyE+vj00DTjXh2WmebSXkO
SV+kFbymBnVrjMiQmQpkNbBCwEL7KjWw+CKR6a9tIYuRbqhPr+fOvgZhhoqXbfUeG3eY3n9G9xqN
gBOA9j8i49vKWaNJ9HiVVsdqaI+iiXT36mGmIfdG57aZ/lgDmup/oTIJFz04do6QLMopvBOHVQbg
XdII8re0eceOgIm7A5sKL1YJY7GAKiNEPUzGag35GZ/QgCxrNk3Io9REPUhruDorePdeis82eynn
sRUhof2SJpVlk5eWTCJMujExIPWN8P01kCKVWBpXMWUE7+DOB4DTG7+xqUYAtmjfjSXdMFtL1N3p
dgH+42nO5mDEiuDB2KT5ilxQ2Q0W3eqb5uGbQ1ZnKLtyqJkOFTyevfTFIJZeUgLXTXPuMDgqA1I8
UzQ7TuuJzVyHDu7HI5oH+8mvibzvjwTxPZzKTEKsmSoyR10iKlZnPSzzkkki+9Ae9yYJoTesxABi
oWbVWH9cPcP2IT2jI/gTux+VzT1RyfIbqAne/JEPZ+FIdpqggedcW4JhLq8KxJnujbKx6gNfLYbE
It75grqjBeeWnTNCcf9ZIEc5xbJIZ7ZB7nSuJcOmF/pLLofg3iNAkFlPWkU4vjmb3PJSj5823PU5
9XTsOUHQjCiZKMM15etmTMVNtIPyGVukqR33i5775ZgHnFUHoKNdAZrkWnlTdsX6/Sokd+P9oqux
Y2RH/5Au/Im2Lkjx6FUILBEQEkDVkmG9nzvtVW/8gK5vTUAR46Dy7ZJB5lSNzEcQVoYwy9u4T1Os
15T8R5cV52bJoxft4UJOdHd04ZBgmgUCiF7L6O4S2+xOR1do1jJ27uBn2g41mMofroROR4WL1RSU
dghXLTLgGnqjoQpOeGF+LFMsKfLQSBvRKGJ9IfU+fEgA0elw0QEwPkQDYcRd7WYKfMDBj+UzCLZf
A9qAx6bpTfWRHm3NWvg2JmtD9vVOgwLw02UeNb7cbxNLPaNhplSTkzKzIfWzlGU+cB8qUBWcRKVb
mq3ZUX76859EDnZst92rlILJPHe87khj2aYus9AwOUk9+e7raEGqP+YSz5uwx2t5mz+d8Bh/FXyO
HdboHfsI5/JfyL0P7MpZR2iIocolB/UwxDcEEeK7YvplPeY9ROLNK9ShXz4l6oGwx5MUjlMTZktv
w4nZS4bOC+DoSJUQ7NSs4iiRnkAtqlUsAF49v/r4leyLWh9vW2oQ5WnFtxELDbEKBtHUWT5uPiN9
kiRjtPrw2TXaTL+iPnzoIM+ihhwhQzidP1ZuqL5GBr6et7W8EsXSmP/TGiyiDy9HgOHyzW0jDkjy
PtAdK8uZDhKLTZ5M/cLuZpQyg88fywFCKoFuFqBuq4M0XngTpXXdMT9vqGDQogszOhsWjoQ4QyBB
u7T4K1ZK1fN528zrZgT85nmGItIzbTGbh5W9lpwAuHYz3dH8VgsLtAz0tQx6yEOVMZwTfMRjS0bc
g27hVlvCIDyjoKLAbZru+wDO67kbkxElyXRtpSy+xMdcxubHUbjmANsY/tzo4tJSEo4/PKwxYy4S
3ejE26fSTsStwkUlsaiYuC2TDlVFQcLa0TIoasoO06jpzKGfWCdomn05j+ARz7c9CHBwEH9z/jDh
GOaldQBkpgvYrKaBoouTa6E87/7/Bi2cIQa02yDly5qoIvv7BH0g5ESEy7FQLiINr/OzAxMy87H1
7PPtwOOD5F/Bxbl5kiTv0V6FUx8rHPO0Q7pJG9lYJ1CsobAY/jUr5FG9a+Wgu/UhIlravwSg23CX
l9fdXduJxelz6JiMjNRuyvo1qy+zHiEZrMtWHoST31jiFqZbTYhbwZbgSyMdzoMgH1hv3v9Ld76f
n0sZb7g85sDhq5CQ6Ec4VrQtLf0I8iGMSHxoHz5T/dgtR+B+a4jLn5cXSQKzVACRrigzjF72fD3a
7hdnEYyM86zVGwthe1Ldq5KPlBrf5DS91GfLRvXHOSFmvO2BwMCBnbvl1KYu1D4SscfOhjyS26AI
HQ7qNPtHDgwvvekkWJ4Nz9B166R+hfWFKJk9LA9OtJqFF6XEv7fEq+dYWVJfGBhoHuDu60TZ6sVP
fVdJA0DzXDrzkgta91Zq6tO9wRKcP0k+U0I6gZWnIm68bvGAy0UrWGLj/NcPZEmWgqJFH0n6crU8
cYX4UtgSl2VODVpTNCFQssZa8cVD01nk8pMbwcTwcm2h96/jaw6PgD7EzFoTjn49MJEOoGNBeiiu
QS2+2NXB48rUQI3wSNzHfbg4xPtYqc7phq9b1RbWg+JRd6M1MbhH3D1jAnKdd4zYsxNLb/pKmWaJ
Uzqx4rvWrev3G+DCPegRyUQNPyEuIoVjg1aG9uDrvhwDAypyZrzCb10M2lqGRQuiBAVJsm8ICOuN
fqEgnvdyoeVxnFEvYznPzcrdmnPufACyX8sAu6j9C01Lsy+r7oBKzA4bFHFJxIuerXisWok7UFoW
cseSweLoAmWOKsdZELc96paYDHpn0+/gE7DD4jvr7CgSIjJScfcz8PZ8972yhkc3HyKxBV9/j7Ya
Qdb5vVCBIRyDVqUmKXVmYdYk/rkI4OXYsVbCmvRmpuSW6YrqDnfTSFVswa3G6fCSlthiX46YtQTw
KcI5GCW2eYRCOUEoY10/CuCSQaTHzIbkUcjdCr+Bgn25hWBbZ2iZf8UjX11a6+Lpo9GcuHawR35x
GACmWl5BvEyjyfMAunTFoJWA9C1Idy76C+v8wZONuAw1X8w8/HPxUT/TcTE8+GZV5cLiAG8YHVZM
tiHrZsxenWbqYld8H/wF1O51rgfPIHDIUioQuVc5oTvNAGK4uTZwSjOuDJDscrjBFjcmRK+koxzl
RHVqlt8qTnTyxzSWb8IxnnCEYebIyU+HrUcbRNGdTVYHlKTq1h5Dn4L0rY4SaXgN+/JnVdEZL+qn
p+56ugKKO+w+kDDChaEHM5hCFRmpg8qHVt/gUYfFDoj2XRhHP01YEqFKFvNKD7By4dwiHAL1RkbX
NfkQ3xdSBI3RbywZzrBkVNE/wMJfTQF1qgexphhsvyKUM81s4Ro1qiXJ8yOGZaFDsHsxj6obbgF/
IwtJEd1884g7tSc1eGc+JtfIRSnE8iVHoTqUGlQUOBMKMzcbxkc3Abw6yxUzG0iDqILYxNM379ct
0iPrFfYjU0/Fd+zdFuBe9ghftg2QbmHZVm8J8jObXJyKqVLfN7OKK6gpbK0eWbdF3Evc8r5s6/ve
ofcoED9TJXSDn2B5J3Wt4QgRBYiLoxq676qdPGJr6lhgKMG6hD7nzEsU1PKMbHEpxgMxVtP6VEre
65FC6qHUaXWeadPSH/DeCjx7JXc5kH9oREooOV5XyOSGwCLCdxEPmUGKWvBXQpV5XHiO3qwHZD7O
iF2Xts6T+jSowpL2Q5sqvF5C/ygMzWTFbBawl1ZGDcG+TqlZx/881o+KkrHi3JPSeY74a1XZp2mW
9tfqG8ohkzlQPeHUSgb66qTjlcx88d57LymJ5eCcUuZzzmWLY8oAbtuRN4mMpn8WGq9qUV7T59uX
kSwQtdiQPT6u2X1VX9wmF9gKS+ObaOueHzzDXOrMLD3MOu4gBND6POOFcjku/xAdKY7zGgE3HwfR
l1T82+MD9kt4oIyTKQkXp33S0YhB+RAmHD2i3ywz1mOjMxjdpd0gfsDS3VDQahbP4gaDXJj96jw9
XrtZFw0rSv/AxUD9c9kvNRcX61gfLRKXgXPnjhynv79LkeIjYM8F2nBYH624mLCZI129tc/alRMT
iPlA3Vbb2TNdQn9On23dc8dXScs3p79QdGBDkg7+A/CIKfwuz2rySHfV6YtYsR+3K92eXACACsyZ
MVWfNrgfi5YPPHYSDuZ8+tzoLRheMxB24xdH+TQzTlFZgn3rZmcLNLFexQ1lVqsGvGa+DmceHDGd
o0Zj/tV4JrXl69Pmf3Tc412zgsFbQ7MetcECYlmZqj7ganAxXdPVcVwthojL18uaClteFKrHx06h
5fenFebwd0WFQ7C2HHhIAYbEPoXCvbCZVUTjt+Guy+F7nyOq75OdznKgDi7127fiYckjbhi+O69j
3LqZNwjcXQFg5qAL7W+Du2nqLCSoP9HMrpo/uLncrHnJfD0bGiJvhF5jhgvXrZ+gbMqFY3+/9mxR
8Oi7yVX/izdlXrayXyWLUVOR9BqTtwycmyRrKsYN9gLDTyJAKuMSbtzfQdyB0Y6i/6wsAXqzaW6v
gS4mCpK+EOLiMWwZuqmDkRRjoIsM0Vb6eJo71dBz45jMTSMqLFcMjdGA+gzcm2ZRQKbVGf+dIqVd
cmSf7H3Xj5ZUkEjLLu0cOfoC8/fsm2dHGcV8QDh6KEGYJOPME6FBVpXmVuc08U0v3TbqgfyHjdal
jqjGpwmzy9NNmMzzifL33wU7CFmP8WfgDLUyApA/lLb5nujgaJlRObdyMMPAH047MoP8AIlaArHS
P9S7rvSADz+PHt+yihn+taIlJD6Y2sOgmcowXge4jvOi0d3L0wi7Ino6VSOuwLdaFfCnBMyCjd5y
QWfeWueLiBm1nIqGGtBzv6dCKSFV1Uno4DnAMcdLg+fzbV0SEL86dHO3zxfBOPdMFegRClyeImbh
RX2F691Th/2SqxfA5e1UxnW63FtAPO6TUtxu0mfSGkyNG2GsWBbRBV5ZsFzgfRKCvoTXpNq7IkDN
y6Op8G0jj+TWBMyS3Y6blZnoK12YNAsZ+iiajkRf3+184qewQODN2FhUQl5bIYaluX3z+ew69Lyh
BAKXWfWhPKWWaJI82eXrwpQNzV4G+3pma2p+ZLtx+q2lSVy2cCZGWgaNFMP+pjzxsJOjpHgGSxsG
omTAbiVCyr5e1T1z4WDBAbP0ECGBwX8o5/fqWXjIYOsMO5/sEmKbR0LrSH1kydu8NlXbGfitsZxN
ai9uZ9as0NZ2YNkEyhKlirvxQue9n7QwQiDZsoocnSlFYl2VMZrWYR9/KRIf4JkxEQd8R+tZR/z5
usLg2vgfx6zlchlpquX7JVaQlK6JhOesORPq0wZmy/LkCyqMG1pOcbpm6gklr16haR5EcHEHJtCt
NrrA2RC0ECsnYdAyekcr0WHN52GiWTEW+TOKwS/dokSPAD+D5ItBGNmUT9cXEcDUky/gOBHQENuP
QqlWsIFnUoJI5D0+7V204t1X4Fu9gJEfZ6VLMFg85gJbjHhIM+8Y6YMoziB7/qTKtRv9mByCgNyL
T2504o0EZwyknjf6Q/jxnws0+3X1ulcgOiWXj12Naks8ePccNN30eMWuNiwl8CQKX2ZMQGLPIrWN
sR9fXYCh8N6LzKWc5ZNvPLwGD29SWqIrSDBqro4WaxtQHiYbezyffmdAHYHKWHu+idX9BNw0+KI+
J92mDf0p5DibBFDTyVs/b/BxVZLFen/qb/3Muw6vW6ch08c8QxB4cD0xmabkqbytdPYbK91aNPvT
aAjWgBCZwdFZQTyrfJtQFGCNhKb0xcbbM+pVgexk+ymsJfvZzbAK0xxY+k+aKQE6oA1Yt3019Pt+
huMit16TY5W5RuYIaJBibpFMf+Nps/laHDdXxhn54nV7eMkw1vVEE426jmp2NlKLSBmL+1jpN3+q
3d736M9Gio17kQqaPWxQYQB3wMlJyDRmr2GM0htNO6Ulzbz4v8k5C1v/89WaAcsnn4y9lrUlOpqq
1LRidFz3YaS9JCkhmRuC7HludQQHcjkLPR3luw144uuRg9zFE4Z11j6O8Qfwv8xej1BFjxi8zobT
3qFcxGGz5Xgzt3CufNyS6/gZCTj/LAcu7tgY2SFi6J4Yn6DqHfM8+OYDbTdEPMdfqmcqJ5lMkn9o
UuPHLiVWacvEfI5ViI6SGeFQRjbQZwbhgrebyd+N0ZPceinlgfCjQaYdRRzYiLXo7Y1QQmLk21Gi
x+VTOqHUdstf3+ddzpH5qKPsl8yoA+HB5F1wPbRQysfEudkr8VHO1wr8K1P96bSw9IHpNqredrjj
KEhESQOflxJxRayEKbByHf1IN1MTLEa8HSNSHQvUbtnOdv/ykpWXbjtt2tKk5AoxaWKe1u+2+hMz
xUKFLk6ugvbIVw3/hS7sCMT+anm7bT5Yqt3/tOVhiU7oCbKwVmhjEHFkv4zfS6IlgDuVGqdQrgET
ptxl8WHxZCxa3D385m875ZTA9VGemqpZBahmZHCKO+DAnE4PW/SOMISZyJwTVUEDHyMUSQrKq21j
GoHD9uIbyJVmvFLY5j6SNzZYEeTowjTn+0AX7FJi4EYYqLfK/RTHOudqLaMX3B7hK/wfqlqd0LVE
scDAuqPZyJDFK45Q136DLFJKJaFLgiRj4hyx5JwWxxqq3LtiOdqK9J86JzbHzHPzM1MSsaV8oLYJ
YPAEx4EEJtWdzhzz2zIFwXikENiNkb82oX9x489z9rLtGZiIRQVA/lJ5Upnxt1mEGrEG3p9NtDqA
bhicI2WB19YZDxppYsj/k3kyuUNPhbHDf7aNvpUIrw7vfSuSDJRH9gJCdVsTbVmXgjvZjTkyi8De
y5nXOcTQreFIOXaJv2JWwWOUkPZipQCkwYwGa8p7iEoTAZu5aqIw1vKnMNEUhuIglsjz/EBxGXBj
S0Ms+BClLwASOyJ8GLWsY8pcGSjuoS9uqE9pkjnN1fs87qCimAbxI2Wr0wNTFzkqIlNGn4xR5FBu
eaYaHo/M1rI5c+jHSKBTVzblgKSIzFpujMwohBV3gBSSvFDNPszVKyqnDSGrf3M5x6IyVjllSnSG
1RDotF3HqWIo5HzNVoPlrg0EsDfSRWj8qbdH7VL/plGuERv/wcR94oft1eERaY2GwfXXCzS8DSOg
sOn9SPYcZQMchYhzKfbzT7j/xABgmuGz1vmBfT5dhH9MMGHqLAadRuAJsmhWvVjJtv2kM1+ZfCh1
tX/6OeQcunHj1c9DJC+2ve6B9biRywMii4DL4kDSPRAno7r0z7I1NzjBOS4TSQWVRtW4Eprd+gTV
qfjEMJEt14VifJafcTgJGMppMorOzvSo0xqD35YZraDKOMLXCnvHNxLLZL0ZjdJDa3/E2WI/vaXV
anKQgIUcVZ9xEYN0JJtfFSBhT5BDjiJr6WA6FfvqdB0qPCQtO5r3vCP8RIuHsP8rNlz0hma6IkTQ
aRwBxAXZ09YRi1Ju3NtvCkWnfForsgF76+Jv9zJEH46BKBL0VMH93zliRrTrYNXJot5II2QKQR96
c1AbjJ3Iw2QV24S0mfbV00kKCxKsg2iXe1dB0F7+bowUdLBxKjfFiiXCZN7N+qaPtRJ6wXmygSpA
T1mDo4XkIeWIMiuslNS0Mab89e7ZcnigOyyMJchaNOWIq26LQrXRQjZtiwi1d7BCXIDr6//2GfLf
kDTXOSven+H+LhZo294uebRbKf+oAraI2FMXqrA/1eMbBNTpZwGaBQQSrDHIXuDE1Ye6F0z5EoEj
pyogfikeIC4z5jXqc8JscD/aQMMb8cMCGts9BlXMSJax1rVfMp5YeUjBWl3YfNrexnxZHVhjFiWI
pkxVr7Ki/RpVlIbAp8kXoK0I/GvpSNbhg5OrFTHkppqWf+joOh8qfCmPzcqzL+ouFE/ecFuvZkKj
rj2nVtA5GqioNFD1yIaTrxswUnNjDwYlWyfELC9NyjwdCsTQ8/7eKNoJowdp0IL4iw5CYwXRtIJI
6SpHgDQaBeJLCfdYLvmdO2EiPyNr/TITEnZvLO97rxOFl7IUL8loOUWOYzXjTH6JMRwRDB3Vseo5
Q91X6fCDqBUDUqM3ZRYUi0pG5lFqtzENy6oIawGePVeaO2ymZEoC0vyKXWGzt61csZMTywNIonlL
ZGN6ah7xKRlddWBAEgtCQGa1jdjZzMbKkq8zFXz+m1/nsxgso83w7mgD4/GnIQgGhJhWSbXAd6dS
XC2UXrydoeTkh4jGg+KTqVhZTATz9HqYegKTplzL0wnA1jXcAYu7f1HlwBUOQGeRQj/7FMFUMrZp
gpYpKgtcG/4xlal25m9ztDK3h27p96FmZMQ+i/d6vQiW6fcVPui5njWOZ0naexMQSW9YOTFsqUMT
NACanqjnr3XFUZrldB9X+ba5AhvNTKBY4ts/mB5LeyXMMBTJdKfZxRpgCn8YklhHZVdxXIKIF92s
FpWVbd/VrV9g/+h/aBlya4mS3+06Euwy1A9DIXh+MBRzPOJWP6UIV3xFrhWI00tjQ7D5ol3DW2E7
wjrTpY+IBayEouuDrvoNODWmNueKBRNCWbQ4Md/f8fU1HCqdmeGchfBYHanPiNFE2yKDre50V05/
iuB9yHyaW6SUuSqHppXb5kgCCKfpoqq/pPrqWUkIYcaiJTPcr5q2Tu1h3jAe4mRfT80mI0RyUABV
IzH8upQRpHIiQXrg+8AIiKaTkBSord73YJ4FEsBc9Y7gvUC6HdVsLb1U90wIdN7vSchz3PL9Enwo
VxEw4djryLZTHdbosbrQ8wNKPZ0mz2YvzxILTwdAIpo4qdicCOpM0HEa2D9ALzgyynyM8Df31slS
Ok7OVaLylBgrP/ey14LeUkB33zHvFAJHAignrIgMRWAzl5m6qW30MrKKKvX5buI7IxMmBGK84LQY
PHQALTImvXC2Xaei75pgeYHNJ+qONadGLV3Nl8ZOvJMdTC1FQHn5IhBOGbvRNhcdPIv5brzpT3PM
538QEoWj7gwurkoLtQ6cj2HilE3LSQmbeuxAu10/yf3gJAMuE87jMveu9Ls/qdGg1pEPaQq/idX/
Dilda1flJWfWfjBc5ULWyysGbmW9wnf3XIrdMPDXXFLwhTwIkwR2X6eSGAGm/vjPzcS2oQP4O/kw
BFKZAQWop7Hgr7ER7BQjWt6KAGlI5hPzzoN9X4AdRpyMuQZZmoMdHkepySYj7hE5uNOsUCRSDxwr
jzxfHNA3Ru/Rzih+OwKQ+5Wy8HB9nkj+IutmOhpDvj+q1gV3UR3dI0Zs2IqAt7pxqM0fZl6tqhAp
h0qiQAZC5IXCC2/4vfLQ9MOX43uAooQ93GUr2+eSHl7OjzlGoCZeDVUOnzRcdv1Do+Ggjxy08oDS
2BPFq3Rw15sklcuC/csv+9i5lge+4OVO+3c4rxGFZqiPQTr1RwaN6+/slxbz8IXWHOqq/YG1nWQi
HVqls9hk8dqKTJb8I9CuozGRHh38zq13d1diIfBgq9kWwWw8g+Zgfb0A2GV0T/ltyKbLyOKWnz8l
4wrVlBeiV91hslXFttZ4hWa4qpnnjvWXaxZlFDRWa5MiNy5FYlJhmc0nrv3dlF4SefojSO2xxB3T
UMtAGEZMsZWI0m9TXYY2eZMpxAeKJdljcrzSMQKSt3aFjKOFE+bfcWBKoestVdPY4gSKZ3gllRWc
seeboWJVfiVNurucWLgdpjVgEsIiKnv3GBO+nm7m1XgdWzBQXHqtD7oa1WXdiXC97C5Y1zIsTmTD
Q4aW6mBWTlWy9zGzFhlikIfrf2hWPfGDbTy2tTlj/OnQdFP7Am6IkFFytMUDQNYhGgDU5tw3NVgA
CKvoWHtVu1Emvuk1FPyCSAHE7r98okQVITCedBw+1wRrGDnw4N1fZ2Y9wp3gjUrR8yU4+tUjXAh+
5yPUQpL0zkqZnS4I5jM2sTa2HaOE1/Pf3x0vjRo6LEqX9NvsfOb5nU8uLnY5gk50b88YgQRgzuG1
7Qth8SB4VJinjr738/vpZSaM6xuUDPR2+5TX7FR9FtXPK8/o2W2gbCZlfb0k38g3aTxopDidGvk9
vuaO8klTMGkHiEsWTfRqd9P8kCxn1rUtwuf3JrGjolp+Wu1F2p+mFSGU2+ZbTI8cHiojadXC3Th/
MrazcX0ihWruBC5gF5U8YXDLvsasZ3vNw1ywgoNfUNu8QccxUURRqnR2shuBlxhb9pzp1Jr50ThE
/5XNXvh4emrcEb9VEE+eEBHHkQtyCnXoXqzfKMIUNcDt6X3SpC8dZCiK49rnsvLGUZ1Lg01XHBSy
PlFzkSWHi2b8bpRG4BNrXFrSydryOHphmOEtFXblQGbivNJnr1mKgkzANHdUndMj88pU3A8yGENZ
pG8eG45tcIn9fCvxfceYwzfrW1Y9Mv1jeSZdxS6I59gMu57CNzOV/Y4oRENmCNiuwHf2MUNZaYFZ
zyARdVqiCVPVfD0Jb0gf3Z8YXHYAIo+VwarwjWwlwgC1jcLeUDXM2SMqTyN+e7LiIncntqH1UYJT
Tej1eIhWUUXptPtzMqHLAOMhIPKsl4KjOLEcmKtEDsivS46K1w/TUhEYvokaSAmfVJCkQ4dzfoAR
n5/vP1z6XdY54cANAyKRKFsa18C/P7vWbD/1eo51t8ptt4XHHAVWuQf7SeaOIjfxLXt4PAdGTdff
XFnsgGa/D3IVx+p5jqCm6dNSLsOt6atJe4jdlciEm4NytQwP2fvzVU71fHrKeXQTb3UAM7xC19mz
uMHwhY0nvVYc76d4ER9Es0WQUh5MpmfRsCF4xPFJBK+AbWF+iCc1zEaYP/xObgbwCbeUKpOVlAej
+Q+hnLV4Di9S+Hu/6keNHbInzjh4oT7RsxmJ+emv8rz0MYTJhY7RU5b/FB71m03vroICorMxY8kP
S1Sq4b/qD4K5m34f6ntWrqjUeT2i0kiqVfJICs7w0+05Cf9grUMJ2mJZk39VrwpAs9kN7OPFAXdw
KBJTB6MAxgdrvZ5pwI8xn+fgUJz+Wf2Tgjt088qqXViwDpXn/mltkSH99I1XL82qWnQW7kXsIPXz
kUldDrSVBdqFA0vWLHtQXrNvbsrHWr/Hv3qfjUep7A6k0z7+bcsJO5Paapa8/6uOvcNOUv8yJMxI
KhFP96rR9OiPpScY8Vt7h/Riboqwi57nsM5a1Fu1+bXj2+69krK4rbXAUnEovgKspRdSuCZqqKig
70stvdDY6f1fI2vHTDzQFU5g0wPgSLHmvefgWsb330awHuKs6axqvcKCMXAasR6TrgZ3cXMrzABd
itll2PAnLHnF0+7ztqdrqiOy7OljRrik2goRQbrnBERmkseuJko5bhmIO/eTSyHCAZXcxhsVvMBY
1PTelwozF3Vlhl4a/TK/bGg53BIOj2/BrTBNEST7dm7zShBahaKzIwAJJKeD7f0YlwTdJcwqdZaE
y52tCYofGtS0CSb7GW/NkosvnviWcu8z+VHpnp8+oU5JLLTAPbaHxpHVS2MvqdlkwrE+QEixr9TX
osQgaQnvyT/V1YalufWyetyAgHfJ4y7khtZFC7xbvGkjtdLehNEiQpxXyrFL9kKjh2KX3QOjV9Sm
7Z6SiBf/f8T8jmoTzW+Zn/fsXgBn+/9y4gNmJsIivQe57W4vn5N3C8iu9wIQHcbjNB2zFvQyqHcl
IGZMaqqzpfqcT3BvOTMOjSCFGCpo0ErD2q4YyEYpNdEDzG2sYJXZrr8+0fsCZsZ2TxdiY9x519lw
AHSTahrwyDpbTrWAbRCIN0ZvwMvhhmN7N2zvU2a8DGaPRxlnmK1nthn/HnuHp7A3pAtCfMBRclu/
3hi21ul9nhbBWQzTjpsZlSUIlXwNgviBtwprgyblE1afDCIN9PpwAOdhiBJ3C0sby89j6WUTgqd3
rVZ+2EaxdL68Pza8rZYucJ+UAj4ogZhzeDLOHOCxty+2St4vL9wLFPHHUtimflbDhY6yUYyeKSex
pq11V2TmGm2xgDBcsdsE5clSLhy0AyrRkHkNS01RJXYeDz8xJc4vVcrbIRNTfihCu+gyp45qpO+z
Ekl0WfTN6RYHjEnXKlcmuVhNvv5rs89tX+dxVIDtB0+Piye31hEphpN6mi+dxHQ649TH8+LxTaGA
ckKOWJOQ9K5btTrbAy2hIcS57CuZPjPeWQj7bEUcukavF7RFuuafopoivnA27qj75Tqom/aZsfGT
OrIaeVeX+7gaXchox11iSwIMzm9vM5gwS9Nm5eUz+82qk/rvHfpN+BlCMIGPJYi72zgEgb9t2wvh
SEBoNLK9hBGmUJAV6r+9Sh7cOr3Z70a9OV2FonMT91oYAk6TeTmEL05ze9/Q8Oht6ra6Qmokr9uZ
opqN2We0i3MLuloD11WYjUiPtfQB07T5dEmzuy8bU23fZQvHuggg4s7eq9udcV/+OgcKktSR4Lx2
yaO8Vt/lm+ywVkE8d86HXy4YsudYclWwTA3zv0C3ko0a/6DAkJ+Ua4nIeFZjzzgMv6PI2cCmiHhI
R4LSQN1/iyE5ufrgfUlIz2cXaQb3h3KPwgKdGWhNMd33oUi3UutmwH4sYDBPaphX9No+AzaJZUOh
UEd3TkCTPNpqu6EtFOtAvP14CuuQxvMSxypDM6EJy172iQpA9pzVkSzhuT9K3zQzcN2jKdmmM+lT
7ae80aipognob9Vw4AeUaUEHDcp+Z/5UEd3MVCMBxP+KwR2wZpulwDzymg3LM+oPx6qaC4RJ2x8F
A0RDBzkAgsYHVZmEf7mGi8Olua0SiyD1NejCgVdMjU1vQWsb2ZqF6IQBhFiGy5yWrfBNbKdFBVnu
EvvkbMq2RmzidWHWC6nTnhxowBUTbN3i1zHSIQqG36AOR2C4uixgn0AQA6SHGDSzON7TYdRo5jId
kEY1bZLy56+KWYdHu3yqozmM0CK69ztWvWXqOHCVmaNI+VNSuWi2rzuZuersp+8I7kZf8iNuOK1d
W4LCgAaEdhopYiSZSRa1cT9mdCQbNyMecwc27C3jhSFYgeTk8NjTaUq4DOcToBoeW2R7GVPQC6UR
rVumD+sZ4mvWcBoaWHTQ+Ytqzz0vJZ5mfwnZVNnZRxQe8ywgS8MbGB6KUo0W0nUXLXhzjFakMTev
ndD2ZaJlDAHMCZLzIktNZeWd/9DscJcJIlhIpl+FfRJ4uaMQLPb5z17YqnfCrS3Ae1+oLxq5Nf+Z
Y7TgXO17KxkgfJUCOZX8xGov9QQNtaSxGGWCu4es4lO2Qstcu6vyaXSFTobMfF5v/DqEOFKIJ+ir
MNozcHo0es8NUTWQRMqhMIxFDAPhD6EX12VeY5meICTnVcO7r9G4DadToqnLzl4DgGpJeisZpLbp
AFETRllaaaTYfXiAUYAzM/BbV3oUw9xUXGka6a6MN/ZqYlZnANlxMkjQbr3XQKjXZ/r+zH/SSdQd
7ILpxgiULgDe6Sia+tKBzGR0FSPmrWyGCpNKo+nXNLfuHO0QB8UER2/MoI9ChaZFml3v6n/KQtHj
6H+RATx6irWmgr1SEfdnJfrwj4VtVP/3JDrQSlBwMuyawMX2Pnhp1aVo2WP0Q1oQkkH6UX2GWpHT
KbbGKtb+sPNuwWOBmcVPVNeXpnP4PHSKMzda3Nur0at/L8zyIR+mwAgCYWfIhFlu3j7mFiPFG5sE
EvPYlLWXZQG3B/8ylA4uQjEeY66NMu28ownqzG6bs7eW0kFoWUPOPX4LgTAlfG20M9vjDPsdWqzu
p5hMj1ckU64MsgKik8kZEAo8ylRd+HQLAzEstccn/v7HxTBPilW/QkK+TFaAMwQJ+TxzccGIZxBh
F0HddRWiJd5lmhsrJLmGjH1SQSne+SO8b64KgjPVVVpTbII2u+mfLVrH+C+sN8n/7IkSero/1x7k
3N+HbrSf9NfsnIxOW3N1THpGsm2FNPjs3LYREk3Up5gXPjsqeQXaNaH8i3Yhvaa0sJ0bBA/Pa5qb
cWCIqjeGBNnlIB2tjodO5vLiBdkwJHvuzipABJG/k43YGEEOTsYGFWUaY0By3ihOfjCWWz/3CWtC
H9I75rP6JQtG4ZjsBOgrqVEH8XTn3uZw8REGNLlwLlS3j2traA8fsLtHZDXjnnPnQgjc/OxkBHuo
HBSdjROkaQHbfp3qcQ7ffT++/sMJc0QNeqh67XMYsK/53Z4TwSLlS7rIzeGTocbrJ6zXl3z7tLeQ
d/Fr7EE46VGypuC49Qg/J/SJGAVjEudcPQn6kMwsM39vzFm3nfF1y+GFfomBG+Sut1DkjgHHaT1+
Udct4o0ADH5nttUuxjEM71HxsHFkcyf7M7UiTA5zPSfrF3ylpmTYbEklxGAyMP8Pt9Z83rUTcYzU
AhP7a8vaA1ZnbTa66DNVFjaBP4sVWIwsNLCXbe2HmK37gbX5E/PgI/5UJcvVsq0SImMZkDAZr6sI
wffXb++F6S6B0QZiGJNWxTnp5qRADpMJqe/PB5czvtZzk9i6RRGv+bPUM/Jsu/OhrYEY6n7h3ueP
64yyioAgF0Qv2nZFcPmKw8CZZWokSuG2hgcXE5y/q9PuZELvI/AvfqxnpLzen1Gu75igbm8zulEH
a0W+Se/z4IWmguVgyH1iEvEYHliKWx6kpeyQwE/B9JmXID9ppNn/2TW7rgzs5Js4Pi8xZ2S8udkB
IrX9gLrGIFsb9Wr+2IvpKeiubIHme5CNEO9kK3yA2b5NFLASwb4q1ARweX7w23GSodRTk88oDqnG
YZ9QKXN7F9FCDYLChwmShI7d6bE4dsXIk8dYlsc5/8EaR8dZ7gWtPR5zMKETFQd5V8uw7NKgQYkf
9S3FsdZZqyICb5hM2v8uCFbSzPPnIcMYXIrb9B4jVbWNlG01heOahdPbFCptNGPm4IIdtPmtpiRB
nU92K2i4RcJCYM5pJ4QRBq54MaB4EFGUrjIIVX1Tu470IjobWL3P7BgjBxQVpdwBNp7hPcTpxKLE
MfTVrRaAu3pgkYZDoMsxSiZdCoGaETaf/HsycFJUuPim2BFkG9OyMNXtitaT/DPjyjUj4E1LEsyb
nh/0sl2XTAD+5ReKs1vjNZgd6vbdLXJAAiEVVO34Kj0pGmOBu4aUhFgByUaDlndlNgzeDigDNGIn
uEf9GyFB8h6y9uDvtO+07cmUQ3tKxFYXXD+RoLFhFMP+S7JxZCJnhN2NQ9ErqMYUbyF0kP7DzIqA
WlUPJ3e8Xgti/hkR7XmwYvTaSQjB7nasTiEAZAwtI3zd/+dRDL5NTXSTDyqjDjD3TIICS0r0puxG
u3DaDMCRhUeyrRbThbvNraEsc/VCx1V2XdNnEOn6FIa3mUYOzdUiYLM5R5Jlk1anXcqXwm6Hbcu7
L7RlvLx9tx2xR//j+QT4t+JBEs20U/KFhBF2Mg1mGjF2Ta4T+lCWlGJndW2MHFaY28KbgkH88K4N
do2S2UJDq4E76g2IUIjxi82KO5G0vsYSIPoArl71/w89Z72rGm6zMzlQNc4RaH2Y8P/PDoi5wxW5
hX7B/YS006asAELpnPZejMBGJaMlMWeuxD4LCp6UJ7Khmk/g86FlnGengSmTznSwpMc5CJbfiie2
0/+FKMHSi0cLfIIP41CeI9suURGPSspgFjco4/jSxVO3SMxTrw0W3mWTVrZW++P8DkJwQk944jxt
rOQfMlFOE7As7ZHBOm+Ydp8w1ixb4v5mujVSiw9yrpqY/4FmkyIhtgRfiNO1GFM1ZrJfL8l95wCh
W99len5PrZ49UJXkJu7Dh84owRv+vnmDX1LQSW/Via1n08JQN2+fpokIufnDgEIAZSclgd7uMaEz
Hl7y6EHDb1L9RICY8H1KJtY8v0SYhiYDlmgGK6vN2sc2bUC0MPLnPsEy7qTcY5n5BLaS3qLcvCD6
LrAMylnqcPhWIBw9oHoE+RKTk204hNPJfVsR2l4XgvlSQRFHzaEJ9NEBTVUeSNN/UCc4l1i2pPmN
8KS8uiUXSsHqkmtcgxrfDuSONZqOpIw/ny5J/DBtpiYLKbsQFttEcEzxAkeX+QaZEw3omErj165K
rjjY4iT7GLJ2G9PAHzqM/y5zr0C0nIAguXb+xi+B2VPoq2ioInjN5KXXcPfaaZK4Qv4f5gQ4ttsA
VMm+D2+Lx8WoPK3SR50T24OoSVrTUwSoQ09DLxqNNHcqiUD8C/PqaaeD5FFMxqy1NQUEZbp++B11
mYaLFH6tjscC9GwteF08Lx1f29isGzB2vCRDO+q+qDiB9GhhK/zAsMZlB7o5ZDau3cjE9H2LofJO
Jwo/e+GZ9l4v5Hw0JJ8dpxcIs/ciytJDhU/rDzhPNamYV0SKvIWd0gPQzzfsxqnuiI7XhhsMTxlR
b2QZv7DBf7p5BFYjhcmtB+piG51FXaIJUmNtAbu1iYAVB4v6To482q4iOafuBQMDejt4/hmBWWKS
OTq8AXRamP2Tl8bO0ZB2GhVcr96o8KHvDtA2UVrNOyqy3pqG4+EZDGXB1G0m2nDo4r7ttTrYRYxA
fWDEHxUKnt7+15fGo5YVrGzKk4IVei+XNXvI4hmvYEx9KUOsyKoHaJsVLaEpHwggXlwSsJsvr7Qp
nClZ1n5Dx2pz8MzuhiZMR9qxXAg4I0bEqoN2gGpkG3s/mSMzXoJU6vOTzTPZgqrhQAhAfL1FtSI8
DclB5K+FtB9pb3hiEpOghYkZeHEB3StKxroptqPIAvAA32/LofyS19ykyM/IyyK1KzdQZxup614g
23lZqBCyR1UaPUmLgCogm6TYNdrpqObSQXBk7ESVsBqJJ77Pj4t+PoGletY7uk3wFNJTQjeJmpKU
RyrKGky43korvJrfMMVoG84LlTl5Xqw1YKVvZMCwPD5oloElOAdOzRPauaMFgzVmG82ijRUUCJOM
npBEteUjcJhL2VnRYW2QshUJ3Ep+3rR37w7EFCptBFO3Sy/WthSCeGmw0Ne20QEwNuJ2MjxM7VWy
nX/CDO/e2AnqGjgXhoZkb/EOAilCb5KXEgnvyRq9XHT9RUYUrQ2vEF4dH7MmUdKPTtYBVYzejPEN
3HP21gpUO5AoasrpFv1ZRA2mhCopCwmaad6c5YFvtixbP3aLrTjhfg/nZ7N11p+hqUr0+JXxs8R1
Ftr31maN9HdUwkwJF1UMXhLjm94hFeZnscp41PgGkbj8jusd3Qnlxo5uy0Rt2uj/YeMRrvK7b+rI
PKuGjFdAuHzUzl7Rr9+YlaqFMNP39xGc9qu4lp7zWLcbrddEJK+NKylFAjOcJV3Itrx/EQkhj4wh
HGPEpOLcnhiOmCQhpEt3f9HjNlC0DSs4C1xYYYlqV/Bzi+tAZOCL3h7QhKe+Qi4SGh3bH/kfzE72
jS3dQBiKCi7eXWAa4dJ2O5PnwRG8PhzD9Ikwx2Ok62xeLJevKBFyoY8a5/tFXbG6/ghk2JkYrF1L
mw18Trhw532/8bEaCAsgbAlj9pb7IiodUy2igOsiU7R9uwcM+mMErmSYXvjs2zzsiMDMeJmSLOVr
rghly6m4vErmHwDXgD6lbheafawIH9eNp5kz6TBtId4WoYzB0cg6G4ACorHxOsa7sxVOZhlGhg49
3mLkSmnkHSiXZuwHAQ8CtPCHNVp+P9vxcA0+QLXEtNbvXs7nuawxBlmG7ZH+wf0tsCxMXKiEEHbB
AipDp5DU1iyb0gYp/U/Duc+MsPbmFtpfEq7Bk48zqk3KGt3dKILUhSbURFusGlpivTaTuvFvG/dg
HujSsrACk0lGLwkTjFjKeDYCCd7mbPg/13PkRT+XZwxxURRfjASKT76NK2Q/kOMLiNiD2UtF8fk+
QuA//m4IqANdnal+Krwq/19DHTkSHwmS3dRV0GB6u21HFb7tlls2nu3DURVXZNV2I2KTgfgx0Kd3
8GziPQ/473Fp+bqbtt06Aw9efMzPxt5RQxY7To2PITziy1Rt+T8Sz0+KLc+UaR9wtRLVgk8zoQgB
UlDMU4CovIvmFLJk+n7MtjFHS7wDLDd03XDALo/yihp1OzoNz7e02aSMtVcduWEpIUcH0Si0Utqe
ZNyapu1WY6nyv76EbJsIlPIxRkmtiQZ1nQuEjMzIFqyqmP4dL8hInN8DNowVDjQi7GOTis7TCeFc
89R1YcV0yNWOqr7oGk5ujSOFUPx3f/6BLpoHDf7ZTJqq7WSCGDV46jkYTcGDm3lCuCuNU2yKv3lu
zZVgpYemjJsmaxA0D80JZK2qElvrgDDtVna6fY8qQsn1aHBM+txnStQN0IAXENtmBbEemli2J6yt
rx9KkWr8/c6pHQLWGg9ladFIoPhiHtW2iKJlVV+6I8JrDzcnNxIFIM2HigmfJxNVexZ+esyJZYmO
V13p6EUhA1ahJzuEb07rAIgDNBuuFRcd9Q4M6WaIXbe/Nk1miNWnOml9lAdVk38pssfN1mdVqSVZ
VJuBGRI5heAiCwrZFdRzxU2UMaGCJxiCUx0HJOzWE5U6FuJCjqtF6eKwbQ9KMyi2j0gm1yI9GSAo
hLWSqAjBUi3613u4sV5u9G3W1deqlPVTvRNhCBzi5f/SgwqwK+5oDwofpoasfKN4xVi5eAxVyNBa
Lnz+i98uZcD1Nr01QXCpFy7Ob+MiWRw4ul4Ah8gGfL/uTDWvMb+vTING/EmM/arUq8ogkk2mVdXp
2pTvUtSQfbYu5syszfuUoaMRS+F6Bs3uoOtEgV4qZ0KWX+/z612Z1a4n7q+3DWqvu0tf8aDnjwJ2
t6kA8HGXPmqQi3M9mGMsfgMuf6M1FhT00/R6Qy8D7YqiPqHI4dcIkNsXs2EVsSfAQBU5LvEAlbUq
6wc03XCoAZYeAIZOPWvMP157NnAdvO0EkEZKIpCP49cQxXtDssskvh6Gfc9bw4Yr61TyqxA6wRTX
cGASCwt1ptWu2ybpJ4CH/sZrj2KFe0PBkmAgyGSMuCW7nqBgwAM9GZYcNnz7RecilaBRIkYO0siS
Hx6+2rDBVn+njBIwKefzd3KpQo5Mv6HLTC6B1ooduPzRWvZb1slz+uqq9EqIsLUEafAolKW1uXIs
1da9SBUNXtEnOszKZxvhhtT+seYxQuC0hENXdgSRoCcm1bVDw94Kn6AJOQKdebKsUW5/thBg2iF5
ljgkIja0EPx+twuT1Uxx6o39FdOTwnQEgGX3h1LOttRI+Hgl0TUp9/wukNGXxmiuAzf3sjMs6FX2
TY84kmiRaDUvDgtgbAmymnTcx8sys8jCbdkwN1OGQ3H24rDmY1VZKuc5kGWbYg83jC6AGb0aYGAr
F1wKpYFtAYZs0hL35/HqQn2i3475UWx+C0gjwb5Hi9/zurJtUG6Nd9UNXsNtYI7/aRXILYmKEFX6
WzEklzMJmUx5ricuk6odOYPENCmZUN2BEVeBH2eL6ZzNNVvv2NBjlhbZa1a8nSocmHlXuvhv9BX1
o8lZ9rqqWR1TVwP/teLyg2aJPkwS1irN9UxGlxhXlK8b2wtf+1qIbIyeHABUpa846uKKx0bt4/5p
AVV8HfyLXg2xYRqBM19kvMJvXxXLjqTJIiT/fg+z7398r5C2Qd1i7e4IBVOvzIZ1HCTYvrYzgnR5
Im4tzNZWtGSCubvaNM+boX40t/yjYdXe8HCOZpsa8TH/OEIPafpvUYGz8ii6wuDe4e8OA8cY3ip3
aJtab5W33RrhSpB8OhwS45YBrjMRRgC547epGCi9yF8t9/jLCXL+/+Az31AFsdXWQnfaMmXsekQ9
Ma/DpA9KWeY5eMQhr6TpVoc6w7sqYnL/S0+AjwzT2kTQOMosshaUKYn2EExgCegnlocUuUyLfpmT
PBYRK+2bzcCL/4bWIRBGxHwZlo4AbFPGvKbG/9+WZ/1468h/pGG8rrk5iU/Qu+ClAkprp0RZVhAu
uPjWz8GvpsKA+YEbst3x7wBCo3xORlddT84SSYVTdCFsAW5aQdEU4Ug1BMNGN5mKGM3S47MGVjWV
W5YAQr8+j8nApMYOxlWM0o2OaABxxMtjGjgqbJeSVK5KCjCydG4x/ywq+WW9HGKoFeVY+efbpFfb
2OYnz7BhTMMrrdKk39ow4755XFi65Cx8aGKYqBLsjYO8eKOuYxXYd401YfQLeltitw6wK/taf4so
V3Uoh6V8bpggi9geI4Kkx5GQpvEtTkGxHp2s1ylytRpHEtgIOmtylGgR5O6LQ6hOU5i98Nv275uU
9y+58Hmav1Cdr3KwfUgF7tz7VOWT9peNk26ldtj/1d6dAqhIvogCF4gpuxrxLIhsOHu6jsXTwCF3
A1DbWsNxJqO1r7KiSk8waPHODV11RJNiWFKdWUwblo5ycblTCztPnEzkQfYevBKudpuZnBT6pK3z
vSSXPkcRMXZDugOAD2c8Q927OSyC1WxFyMC0ac9l7VLm/HPmF9J4e3FmBDORlfN2Xs5WZlzNK8KP
UaxcNAQ8KF4uAwZq6Ggb2Jl0HSotB3kErYqiCgOw/FVu3HjZftMebgN5h/cvRU2XiM2qnuPGMYVN
hSoiqSQATlnqR/iZB5nzV9NkatQ1mzVhTYbk+y+F8DLxVOyX5FVJ4aFjADbSzP5PupiSyvy8uS3B
tgpmMzQwZWUazMAe4E3B2OuFFjETikWkHBHPTXGDNObRnLYoouRpmxSvSEQ/VrbO5Lhs/OKHBiDc
vcIzU8ZsDAD8PnH2arzb06DMCJyG9I/z+/hMul5W1gcfLZREdk9ukoz2lIgnZEiTbp/TnYbASpCh
9prQzFHfL/PKru58eWTSE27DaZrHQhnp4OZWzCpH14YTzdZK7L7/zErFsJmKLdh62Ac7PBHpmXb5
gskhaWMBWQl8t3qfrfFZbC0ebK7Qi4JM1XLTZ0nsPOt+IfywNuxrozE5bLAe5gaW8P8SIOBqWRS7
cyndJKmkQHP9+7TwpHlezm00IORTj/C673ITNpflWExrbr5Mu9feDf+DWdBlENvHhrI6zfcPvOWS
FMOg7eLAXNQH5NZY/fHMBO0Z4/9GuKV8y5ivN5qUnfXE/06gj8qX835JbVZOkj4H1cXzZrQzOI21
SyD9ZaPPkwvjoPGLkkQ0OrSu1wBmaPgMF8P8Pk7kreM4hQhkMUDuIlQAPGkUUBTWT5mBrmvn8+dO
2Hu7qpYLvoOMQ8LWV4RMlIknnURcelIgHzfoOBpJdF8qiUnevUJPn1CSRjQgVvMMQi3sK3dh0Wn3
ipK4RpFjcTyLISs93JKMTtD3W4pDnBDAuWe9yFQ8fD5eq/wdPY9TQ9a7a3KgxjHfRF3QhS0tHAST
6hbYJ6/1IIfwNN4yW0+3Hdy7pa15c649LOB2J05qFim7JRYPC+iW4TOLq8bFztBQM6Fy1nWzUJnX
pjrK3m3fNgjJJhv9T3QhBS/0msQjfk0J/La0Fn1FyfzGZfuCupfnRaCdGpYsnVD4f4JNrl3XCJzM
3/YX/cC5sisldy6OTwfP5uJKEGGb1HKeFDAzOoPyzjP7jygL8HmIX0lLSgtBbIPXu2p8Q8WkYakt
OslmIWMf5EAeEBMNZ/PP73F8ZkLJ46qkycijUS6KqpkFxaXLyfhkPGd8TI33VoUBG/PY4aBwG6YM
tS6rkLjUfLQPHlsmS3lKwTvRnKCp91HqetMLxwlVylBVZta6CjqN/Ub6MEvYtkQ7KO1Og27uPLOM
lO8IQDOlusEzu38vmOrSGlejXvBRjhgM0FPWTQYpW4f+7I9WZH/Pxw7bFlgBxQJ+4vtb0pPH2Jjp
dou41GAxGA+Cp/3EGTZBqM/LPI21ViO6I9f6go8wtdfjdukUgXsuO+pu5/rZ4xflXm18MpazIQFp
KMOVlodyjs3E3A/1GjgCDPdYR+YCu5Wv3hJzamZ6FTn56Xpu/E2A57ajfWN5n8192dPxfgNoCBQz
p//vwVcbs2f87/LHyyA016wYoZksyINzEEEgaAJHbnjKJ6TuZZyhaBo9cyDaYn/PzZJeX9rETF1o
Z3o3lAVOpoIQts8Nzm8StAKBuaUB2213qL/jzDAuEm9QruZ8kwdL8XObu4hXvtzAsLkHbGB3KucD
Id5ukvflJXXDO2vNK6P27NdBA5D0e9Afo5QKg1qNQuolIBZQyy8B6YOdxg3NZVMt5HUH6PV4uLve
pp77iNC+O/cKtEx1Bw/sl71iloU1Jkri9ry/6spml/MHKOkTOzqGmcseLx3G3jYWDnGGSySnxJf5
KixELLIbmCrA8jrCvKVEzWGpsnB9jAk2xNANw+a7QpVnIZ1K98YvQsykH6hH8FoMYQdo02BWRTQK
JmzY4+csBySafIcxVCbK3VlrDCGkqZH/GeBDqNjfgpEqY8LnQvDijXwJnqf/vL9WKovbyrHSY01T
dwPlvZYqjAqedevxKJtEJjydm7OMyONRl6Vy2pzgqMGv4TpRHEct6i1aE8ZpJZPE5CUb05nagrBS
HzzKYIhikNmHhB+pcr+82K+are7ZXumCopbHK4I8JoRqTJGJH8Kayxjiht072yCKgwPLBR3LwYUk
6/pzJlPd+F6LyZulFJjXwlDV1eeqRItIHIx6aU9+aHomFTIkd5NVoILlXFo8IGdW0C1k+GrQuuP6
q4ZLUZe3VmbU94v3EuWDczYx0yzZM9qroSlwIhfUla4LsVmusDpuWKiNA15OmiKxoIlYVLRZ36Wf
YXmH+Ye25bTaUEMaKkT4Dfo7SFkbN2cDyHftx/kchzzczI8rufDCjOti/eNUfGU6FqZSe6KHrBv4
uOknVLnzxFBmWfrdO8pbrhePqoa99mxcefYrbDui7IlnaVz1f5IxSthLZsIDB8qY8kxlbpWeCynI
nmCQ+8k7E/8zW7t6aqgtlldNWDSQbaoq4VAgBlJjPY66pxH5Sfb8ZzfwpV7jjiiHpQ/NkZrb/FxA
Hh0FfdOtXRl00dtzi/kXBBBEAv3uot0poeCegCMyLc39W4g0sjhRS7CQV48Ob2YY4t/zUADW8DkU
iCCP2iI+NKdtlba3StTLmQ9NjABFtOA2d5AyjxGs927d0uAv/9VMLS7RiSaBSr1Xw/hjDc/Z2mNN
PtpS2Db6A+GasKctwKJZ+FjWGGndogJ0PmaJ9eZCf5CesRzOeWYSVDu8uatfe3z9qJBtJVU/01Ku
ic0Z1WLstfO2sT2bpCe0ht85NoPAFaRAkNJW92bKvIPZs+Va2iCLgsFxFwgJWZGBWPeK/KIZLcaM
NsM0qpsAG9Aqeu+8gka1TM41bIbIHgg95bK/f2DwzzLsiZcf7sRuvs4aP7f0agIVJC6FZ32yjPQ8
VHgHczds1hI44TuK8ZcO+BMUOp5e0CYy66ksXWqVjZO3X2vX5KtIGhhe/HJ+669LE6Y9xSACKH9T
OE5+xxaWeN5Z7HpzSKdxMbN17XgRFWqPj/e6mVtpXhhxhhhD3DVb0fk5Cstj8+bx8EgkDx9tsNOT
TFzJAx+pztBxovQDYrLdjkrFoOK3yVumPooENBSmJiQ2F5yhq+imvzSrt+DAquw/2Vo/ZtbJ9Fei
STmVN+G2ItqoZ2ts1OJpPX9S5+1Kw2ssSBk9VITkiROt4SZzGBJBMXB5Rm3L9aKrMRy+5aYEyqfR
NL0RDG2pc6nDheYo6F7OqWIotjBRXQgSgFIVNemnxMVkAl5x8RM/nO1ct/ROVLh8oWp4y6C0hGwH
a4vgWeIxYtxbUAYYzjpUkt6p1QyBBjImx7HGdJWDkYlkgMdkrl51HqjWjdGjU4dpBYxHN+WrmX74
gTbVtWZoctmSYV2uDG9mCa2ctdiCqaT/9OnaKfaf9CwJugdJo9v7Tl2WWDh4EFNUi2RQAMQPhIR8
gumVyHhoLRteE3f2PoX6mTvwkAZUgJ65zj5evwpWjZijmAIuq55BB5aKve2EQIEHRfssRX7hB927
Q+ksHGxj48g/zTMHnQ71GEa4tkh/fnri8gQia9DlCYC0OtNu01/f5YumgKYLPPXhBw4ZA2kgmk89
evQZow1gd7xspMCID/giETZSMP8YH8e2rraN7FAErdWZfQJcEQf0JqFEiPZnPS/MmWVTi1A8WxHy
wcz3xIYrU8Wa63ldf9vrsz0BIF9Cge2NX8HAOmN6lYFKLLKciJriXt/+sx4qzSs610UuXtYIaLXB
AZjc4bakJ2NlJdazQ6XsfiDt6Bbm5VEENDoDFiprjXWRD0EB2hDIxe6f/5U75V6R/VfkA6cM4PJV
dXAIEhSHh74o8EowKQg/KqyqncLpvnm6shC+bozkKHNFpF5+zWMclbBSUPbImTBDbbykmEIDTOow
A0qB++NFilNIM2acHeTJWOpwBvVXmECAo67a9SzBLrzkNDpreoQcxcqVC9ZoWRP8DP6YmolR7AkM
AiaLtbVofgoPrSmAV144pC+8IygQUAHA1lkn9vJts1mvR7FWFvIgGt4BVKuswlh8NNxMTlq56+eX
xpkBq4AZ24PqDZwpenXpoXYK83tTUAE8xqyxEMQSY0oED6dTeCoKVpX1tGwwCH547e5dyVahBgAy
WHjY5BTIbX61Bwbtj1JJnrrlt1hRDlLraxrp+pkkf6tXH6A0ZUB6AaogRl+VzU2Nrnf5Mrh72Fsf
+xDwVx1PPWQdxGjFnMese4p4xNjG7RDdQmdqLEM0oHOopKLIL2O7+GQwh8km7lsIN1cR0PkFHDzd
iRiC8hzFJv8MMCZyGTlcwvNEhI//a/q6LKpqcjSiKaKIHfpWjKuie3IAO9kksYYKcIVANcs8bzgH
2C+Erb3RBeo/sRuf0xgU6wWahqP19hwEoZPOs1qQaX6omOtek/Qk48xEJgJdaCx9yfjkNqJfzJD7
xwVVN30SrFUq8WaU1U0WFIFoI80iHPuDAUayX8pAs3fOfKQIKhnawbzUk5Yrf+gMeG71wYjHLMOP
6aetWl3NmkPUHdFoT17l1XdO0S699cqukeK5jcj/iaMuTl7947RWQ0LpKYo7gg8/wmSxFo5ze3Bf
2+xpkHUp0U83CGlyUsdFI2jOZYMnTs50DoRiUaxe4O8AjogsRs09fPmxa7B6F16yB7Qd7hLNk9RU
d+5BTwrkhH6/upSupBXaKmLgnTxw+qtkNjuuRIaAIxKgO9wSx9lwTBaeKbfU6OugeNEgJ0SDNlao
2AmfU0PrB9/FuHKzj3vJaOZahf+BVNusSpIkvIGcxeJstYjQ3GsFynq9AumvK/J4sIVAIoh8l94y
osE/0hao0yRDb+JPFgwjroHt6AxoPriygDvvCziNeiiuy9aKZWCII+hoSAeXTDG3f86DbabsRuYe
8+JdB7unca4AMZmMc24bhNpWcyUbC9fURXQG9AW2MTmG3l0nrZWUA6KB61Klu7skV/uKadVgFN71
UX9s+aXojdxrzMM42LFsYfINZPsqtBFPPaWnNPDcqtqGcOYIgWDGQWov0Ip8x49gY9T0C2u9Vx2B
d/tLo7gzq8IKMr2MB88onopCH88yvMC6a9I/roN9o0mpyXliDpDpzX349S1HXX6ME2qoxNXSqNct
8b4LwestLw4vW/vbtkv6N3ZIZsDeGUGjUdlT/gjtZ1vJsPYBioIznO2iaCYmC0Pq380E6bawCbvR
0Vgdv804ccTK8PCYYVHN4h3cIzpUs+c44jWP9q9+b9DRFJNvjBuvZIcoOnMb2yZyHU2TbdMloJnE
rg8r+KUzD1vG9U7uFyj4G76C4Mkbwk/L844nO6FWlaB6C0EgBXWB3We0Q2IzaSzDZNW+Dep7nXJz
cHQcmqX1Cy7aLtbxx1RLk78c453C6PX/5pLA4IR4XtW3CUyR5K8/sUPvj+L0rDBRqXyp7+7VAmco
3EDI8MZvkzFs+YJ+GZFCLiZMryi60Ca0F004Us/qeNuP9FWS8xAi7i2RpMDkpHzxh6W3iJVRhag4
tJIs1fSsKY8Ccmnwyi1MJ3uZiSkYfEyeqHx/FEBDX9VLmvWB9PWXSslerCA2n5sQ+FcDRJrj0BKM
/UVTLcXgwlqRvcrvXWFqP7pB9Bu3soCxSvOXfVRMm0pQtrgFZolkccsmPpFEyskQCREXDxLRD7iI
KMXljHq8Epcw6H4Y0PMoing+9QR7cANZFo0agx1mnklgPnApeONv0a7pZc+ikDkTY/XKT/KALV2m
VuhFEziY86XZKzAdAvJIEfhDUxZcbOmOjUEB43/uuznmDjoFw5hOlZ2zeONzRc9nJA52Eqg9+CDw
NwRmbyYcXoP9wr6RocaFrjnfBOwoD287EtYrLb/8D30Y1LHOkkNkn4ngIXXDv5QEBB43NXBPVKsC
WKCSmPGcg0oKz5mAPfjUgj3V/1z/K1v8OC4/4ePjljCoNLIO2wgpKJRD9nzpD00aKflFw0InzM6p
bRYu3hQFFJxOLW1EUUsUZJ3CmLB65g9TNGZUz1N9AACndmKfNErkCYcKDiEP1huRU5dQP3O8+K3x
FwWK74qDd39wEr+/KPMcnLF4I4ldv9oDZwnnt2wY4ywEFBPS3AJ+rPWsbFtXc2bUgnohxYbj/nCr
v2TgCiZ+HyW6OvnhftV9sJJKct3fiGsrFLAfmtSfCUz82WdLBpk1o5xD7iU79jjoNTCG8nmKenew
9IKBqbliTpCoUrppm+uscJB0uMoYhm5BfIxtftm6z8oNWkfqU40AlWeyCOEPLQ9OwseYiq1FxKEv
4vaJw2RGOuQ6Uj7Ri0hTeVBgC4n7Pu1VinZjMoPo2KimvQfpOUsJ6foyIJqR0G7Ov44HEzHgDRrW
ttCgVNbg8cbnBJAWT4OetL7sF3+OgC7FcHIQBEsm6MwPSK6R/MMFf8nkWIDQrvHEQqp1bOzBp2YR
ZCVQ9EsJm0qvuoELMkL3CoSB0ZhU0b1ZQKv+UfnB6+uZottaUIQRV1voOnxVlV8mqmsBrykbH98l
OA21noTgwdIyxLyPMkeTDndBnBhs51j0YYvudcDmCkRFM5xUVoKbOEjqG4Y8UBhYRXOfysn58CCG
KjlPllyxXIDXos/CGdO1x9SkaBkyH88RYlwMY41NGaBnsXEC/j21P5HlQATObt7nVj51mREn8hip
jkFYdBWEwJEs1MzmYAaMbVDMjQdOicRIfCNDwqkBtnNNFL+1TR6IPH7pL65OSof4R0owH2J0w31r
gZxerURG5ZJukEiqj7mAAeo9w4bBU1S48Cxm9/zhbVA6uOFb5kkqBejOtj3zJ6+LNUimne/3MNbp
+b5Utenax8qwEO5mRkEyA5rOWPCl2b/Ry07ZZnQVgeipGgtj6m8XJBvDHaeENy5smzfhMpzm2P8T
aM686CZT/gdW+NndwOEPdUvxlZL30xJGUBB75kibwOIlePJMkH6KTmtSJZD6MEQLDTbhYJ8G1AJr
YCQ1/pf+65fyjuiAghuVqLZV0idBj0LOMzekkm549LEModqTmmW/z7ShG9qU78aMd1vLUdkotFih
un3kdFQw4BfUVhr7CudW1UyRDGCCJcC1WsMEMTSdi6NWGfr+RSBjsn4addi1/nsWMXiaa7fiJKHL
Lb9BbS9NqhdCLV822ufr2V5CzFchAQEo6x5XL7LQ3R2hUo//J/woiAs251csneDvoFJl1p2y12zW
Oi+sN8qJF097CWkkWBQd3CYTx6U7YgjvCWQtRMJH53Y7+58vp9A9x/kYPv2KyU5wlD7uLMGxZu8f
lJs7zpzrRQJZFGDsACo4EK0yHq7UVE/rT0QclE+1oh9QNYvaJrHbVC57qtKDjxoLoZAYNTA31QYn
qZD5i//FdljpgJCwiWPCx12t7QhRlTH6e2Vncj+iDZr+F+jbwuet5K/W7CqCDVUJQ4LUctQJcJp6
FrnDtCRHzQG6qiMrkOQbVSY4BVDdqF3I5cRn4XeU3KnIrJeDCaYZ+kidkxpSaSo22TBXINLnfTRw
P0E+PKr6oQ4f2uIXqXpbIsioo/tQBy2+mj6f5o30y5IvpuyuIPru/EVnEgBk4I1muGg+W794TEr9
LH5CZaVJ9gJgmH6KGVmS1Bt72k9AfzaQEvxEKgQqo58gGwdVlKqyuxvFDppWLDmDiOeKLRlXwGmr
fa+AS3/6z+KAfs9b1HyO5lwyGWCrHQWjHExKKygVp67x0c1NJp+lnlSw/DYJe6StFxm9pRr36A6z
XgYhZ6hRe23XwJ7AKYC3tyj4lkX4rFrYuigcJ4rWVYcPP9CshcPpmn1cvPJpGN4ia6Ikl6WICYAu
YsuBMpHyFdWiQ4nirQGvSdMgYq800IsIDN7bm4KNcCHa/WmFe26Wv/rtBw1TubNMxlO58MNryel1
hkU65meBeH2eQX5IbuoYbchhlhEZ1utahW41DCUvFfqBi52JiReakJZ+3+zlHX0fdYnVu6IyNx4f
wiq5PKpuUAOiTBbXWoICyS7q0zDh7KUej55rYamxQwmAlxWiJ3ytYkef22xZQqjxG+btqGTR0A9S
7UXIUKB2m2j6K3KlvuI/QUKOwhAq4DCAGmcxD5fCuOw+9YJ1CXvFP3tjFXl7Ugmbv1Lc69B50RSo
xmll44hs0bxN1zP28/aUc5FBS4ZCNZGV4xC4Au5rFlJx2tPXne5TILBpKfRTBIXagNvLAM+KTAOI
i9d0Jh06UjpMHm1a8lWRMxGoumv48Cwc8kTMJnKEW3L/EElE4SyTZjnzHPDbbbSGkLu/FzJ3ialy
rQUy8XKdJqdoBz7eBw1EuypwAFFzmHE43jHV9Yr1Zf5nE0mnqGzWltvgzJqJ00Cx2vEQtfdRQxnk
5/fevDqhpzIPK/TgYkM2VbV1n+BNlzRYGTJfgSxsUBaUw1wJ5TFEeB2Qtj8Uy92u4rSkpJuHtTCr
zqAcToxJFsYD1YRttB0FA25HSxO6i5tsZnCdnR0ZA30ikKwqZB7ofIHgdJQ7XvyN+cRpqRkBfYqS
wdpi5yWpRbRdanmKBzpVG0+LkaD2yJ6qTMtKZFXRh7dqoDY07aypoSTQiHInybucVbNhTkglq/wg
Zd2hnRSqavaQRIWHbXqwMZdB9X7xam3R8pismXFiggFD2jhks9hmDQIg5Jnor40MUATTPfN+B8ND
0v+JbGuV6Ouwj49VTN0GXPwke8+wDmGzMAs3wClUEms9F1wCbvQPb2kCq+ZrSBJblnomhJm0AJOW
ZiuhG5jaoW0XifEQsi5ZViYFGo/xz8xNpSqY+XoB7IIGWZUe6ko5ejSm3sM9FPKgEoTciNRL1ri/
4xMT9CLKSEU1dmx7tyVZ00Klhh9PozTdC1S/lUyzo7a6wiPeaGnnIEdDNVMx6MYr0agEvCUdygWt
mxTdGZGijthvVfHvtAOGmRiD8pQl1bHRGoOKLB32QJDHccuIS3xnGHivL2BC+FvwWmN3yzPlUXDE
9MFqLWfg0+EIRJC2ZxluM6XNZYREmQXKY7J1Bn61p6JXPKYFpCyJo95elztt7C4o91BXWRxeROik
on4qioNEhQIbY2IABrm+BVlVfduJBkVZcvlF9So2y1Npq5iti4FPiyFEa5eMxo6xbhnNC1o5i8i5
aTHH44ocj1aSDqnuGVV8hG/Q+gudnr8Ux1THeUyAN5YVc/LLqiXRfR3+OMs1dQSOF86J+8juHBbo
uIpyVJ1uydrDog/qr1MNtVYwnr6P+8hffHpuN4TXldJIIFQsQ8YdYItOIIFTJNkvaMLVj9iqCRLJ
WdiYhfHPZRBJhdTzSg2h4Gdk4u/uWI9OL6QGrSiMnmyJDNpCPjoIhxeJfYG8t7ju+u4+5tKgcMZy
107cPMdB0K08u4V33uax5qgPu8vDDLB63s0udGOB4PHLa1CuRa2sEaBhtRPbo6Etx00EOb4r/QEJ
I7GY7KCd3gGug7/7pP0jYhl+NRzWhwGksi0skvgxWc1SiJFGFNOkryyWObizjeiTxT4mACIVNFuN
ARGSVBwc+Lwu+A0/A8v7Txc2aqljlH9vod/NpZPMajkz82Li+4Vgg4q23X6l0RUeTJXmo+0wPn7h
dmIwmtwdExUCcGolKekh8YNTwM+e6K5HcP6OzCpO56u9Lyfr4kE8P8Tc65U/cIJHmDQyE++uoHAJ
v1wCmIqW/RbIErYnX4gne6neWipl0QR1ylK2Crbw543/nLU89jlaHmT4SpuxbuMhIRhrx1dzhN4n
dNp8nREZWJ+JQu/YAw5aamIjJ/N0N86Q0UhFVhHb9ayZW0sWPyDwHymgUqhA8iT/c3j2TKrrmfXu
R3PvLLugoACKmNAYi16fQR4nnsoh5KX3zMmTMGoo04MNj/ecBkUQEKfYQyB/wmwpi76YUCTEFsHn
5Kwd3fbpuj9oSX1skSGha2ChT4z8GeHe2pA3enrkKHPHuJrnQSWruOF4aadsLl7+mna17k/7XsP1
PzGxYvsQtE9miSUx3VyRQiuP1qwvZ1sgb3FsG1j4PJRrMwgPV2K8QU9mu/GIIwVlN2E+155cAnWQ
wp3iITOS+5AOAtRJ73O0XZ1UMYmJ0Trpx+4AglEr8Cc0+pbVKK4WnukPvWloPjqoz7VpqOl2DUls
SdkPdOb7K88HqWYde0X3nVjbbZTthCGEA8tmftrv1xTAfHPjZ67k4kPojS98p86WgLv3IZRO3k/k
Wfb6ZEjI9P1bz5vFNbxmSEDTIXB4BouWlJfQ/NovTqIPeGqkDLtTcuzjjc1ndeOzy+0etHLZBFj0
fnm0ysPb+Lp2LnFBme6ENiCNaVD8NTaul+R1ezgnXIOpmBvzF4URNImmGsoJ/Htxr2bKnv7NLXxB
tcsezfH3sABDkr371lNVqiP+sAV4s4hSslfiUWL4AcB6eNiDW6zMf37oogR0/MdevBVVPz2pDN7I
MormL9+aXH71T9onCpQkYpphICnR0XuNzB+cDboDsqdCKA09Wn6IMpmnfkfoaWneCzWZW5pzoy//
boewRJD4AhSwMHN0qWX4EvR8/9PlKHisQyip4272UUbfA8wN0lOMQpJHYq6JxYkt5H1oKgGEjaw4
sYXbnTUIvDQyjK/TOq9FDUHftxKEgUp2p4b9QCwaeyB988pfPUQFBJYk5v1N4kubH6gcJz/60A53
OZF88qQstfBdMJfQw7fGzV3yXgvH+AWnglP9WGf3EfSJ30eM47FMDPZNYBeZPXrqOXHq5ArKu01o
2IYr3WtpowSj6hx8PuO8UuLDO0f+8Fy/2D3QIhq3lpuSVes/2Z8hUXO7srW3h9DOKf7SOPry8HtD
giCTwJByrAWAt58/8ERI6eF+DNKHfUoFDqoP7a8fZTP4oEb2dT9U3TyzztLh6rhI3dreEC1mLlEY
fA/Lw+aahJzSoCPgMCGRpQBKmXVx82Wu7AIFe6wLSvidYh6G6Dnvrv5EOrnivfnB3yEecXDWGKfh
ROcqtf63HBmp+ZTaGE6W7Mlcf+AuJAd+5DB3BfB/MzTI/JWg0N9fJ0PEMarzRL1hp7Qwc/uDQsAL
4ktwxBGSnhihYM2akhdoIcqGbK/HDwkox9prOTRhmMzwSSUlXKTvgytZe8oNmVcBW5PQhMYm/lDm
t10d6tew4EG3UM3eV0svyH+WSGJMM50mCZ1B+5tcYat+67DfeoU2NGP+EEv2LSepfQH9IWLLRC9L
HVdJkWee3CBpUdhsa69zV3Jh5DV4lPpImQvZdzj0Mvkzj1wXVQE/ePu0yo1rzlAW3KuwKh+kinpI
in0OXqEeguF/lRxCx63fJ3Q5FMBlQ0rQQsYjc3q+dHR/5LDYeo1NOeFxtmNGz8AJkhCRzWogjqtt
RboWi70u2o53fAkO6h84zSvJP5dKJd0diTfbHjFtxxeUuzTCrLOvwaL4gUANEbl3U7MvIqY+bBEA
tlzE4B/sd3FKpSx+eU04Ywxp5L3ib1AHhMTaYhTeIa0iXQZVZYwyB5/xs608Ml6lWdJ1XeQL1Bu6
FPWO5KDSdSv3jd0rEUpDS+7+DVSjMIvefemlsjYtJnRF/r9N1APexvb46FZO9vePAoW27KurjZB7
w+7kZ8AlzpKM/V7hDwtmwcJWWxIE/uwhFv72tByIMPkSnYKuKLsLpstXRo+1bvfoWEklwO4bjqzg
dTyPXCmmTdmuoNjK0RGKEgaB+vM3fHt2CqorSAxtOrONsLh4AZVmdbMRlkogJESi/JwhFdVPflsZ
wcwkmigDK/7AgH87JsT2tfhjv+MGL4nZ269e4jCr6LXYEW00WJUPm+YP0MbeE42iIZ+VLNX7gLk4
zkyr6WoUa4t2N4Ie8ROfKLBqFZ4mTrAZ10GlCxsi0h+9t8r7AsQJmiDvcGaWw+D2t9gPne076RaI
p6x/vVgIImpHdHw1oVyDnf5h9roTgKaUaJ3zo2AKAhYcVU3uosB9a4Ek9VSFjVsSWStASaew06il
VpB6ikt2IJ7Z5q+rs21b/qGzaKLCpGhAHIa7H9RYlur7TZFh0uuzv7HZIpjnq1iAECkcZVURuRu7
frhQqGdSLr1zYK3ltWYk/lpdmqLPAUlw/7hEc8kBu87S50siuC495b8c5NcH2B+jC4wUAK3nFgSu
8T+V7DDi5SHbv9Y65pE9r83c55wUPz86wDxqiv4jEVWpgHfzOf1k3empHYuez06HxG0GaSHVTWW4
zRJiWOEcJ+Cyl2Q7+qr1ZlxMOcU1m5rQCNbJcvzlguAGB4wKNoYUwx7lFUbwCSarLfgh/ffdBFre
oW8qNYr/B1Ij4N9EaTSaNzTJSJTdZzrR07nq3Ol7hJ29H+zTCI3jnubaBfuKCDUOmS/enBdNBpJJ
8qn9sHuk8PzzwJsptydzikTOAYJI9txLAKQsj3dHuwa1bEnPzJtsqmJn+JtBuO0JDoffjagUkIHe
ZeusM3T24zaKfe/3duGrf9uRFp+I8xMtd1olhOQpgOhxeTCOCX3JntRBzO+iRzzZOjjLT6JO8iKy
cEtQFEVaXJ3KCWUAzQ5M+Bs/UUiHqNVm0dXg5W8/i7ov0PN3aGkaBObojrQR0Xx1qSLD+dp/JHZB
3tJkCUToEvB4qxb6eDT7xF2kyZwpAirhIiCW+nF63DXd9HETiMDuv6yTj9pwKzq5UFVzvY2rn1Ud
VzBBZ1yCJfmR1LQ0P3QgyCuCLGGPgaKZoTRgvYanTlww6J+f+gb2Y3qpriK/y31LWeDZH8oUBThB
Xf8gC7lOlVfip9Pwlo/QtfhXIiXcfgA8pGKkaQbLyrgeNhLnDuWg0JpPU6zM40ytYmjiNjcz9/VP
cq0CZl1W8INVn2iRAvnJ9aYayLK3bmtZ9DlA6Eapp+0Dtq+oYxMKHaZS6kW/8UEvHgEBrZIqNSC+
ZHWz84UeY78ABjY5b6ovMi7ursBDWm5a1h0c0tv0D6TMBjlF8DjK0M5ugbcE6kR90r0X7zFi1D3V
vmabZVS1WVOaK2NqeM8NkIhUg9hIywsMCSOs7UjrY2VfSbhKhlZpl4/C9gQFZsN+wwDdg7SojsAt
N+S/nK85dPqPcY5rLZ0hV8dPnJ1v98Ss4GFXSxhpptejWhfeP9CvTfA7wxr2Ih+yCt/NdI+v+n2r
t2KMziP14lGXGbK29KhrB/GDiLRdDrf8J2ZztAfFvVLn4l7AUquLDoGZDAoCOnzupKK5OINt7veg
E+uuHYrVpkWVcoQGSYG0aGUnDM9LXfQqwtNgtkYbUCbe8KU6seuBgxf5ik/kfhVicedwJY5f8R7Q
il/qFekqOqGcNksWyd1xeQu14EiVA1u2AtdNf/DODf1Hhci49M2v/Civmdeb1e9Jfj7ykcgdG+MD
G4ku7MhpmbywkJlFrIRkTS7i2XWVh19p1fXki+saH7frT2VFn4Lsnjei1F0eHWXKkbA9bvKZZCsq
bBo2vpdtkFrtNL74yFl6fuZBKCtgfrQrMZY2NHuchsjCWslOysL6ZP9Nk+KV8rMk4GF3aCO+Roki
F92r3gMldM6RiUmiRD360gpVDxv1+t1B6um+8RQhuHGTFfcEIyDbs3DhZpHrF66cXI2msYwNZMEL
HYjF3ogYy1on89v8AMJL4dC8gQTxymWzUwt3jVOQN5Ht8CZb6DQ4rA/WkUuxW479u4EeIxxxnXbD
Cq9jO644jtQUvs0ahDP8+aGjW3qg8B2B/GzntafNBmAtmfG+CRSE+ATlvuTNLhs4YRtehcLVQqna
pLtIfE4OmeX5LXgpoy5+akOFTR7E1OdhRZdSmmmSKZA9UFBEFGjeCpbj/7uhLCMNGgPbGk8/VN4i
MogbjOiNuJBr3ysWuritWpWvpfhI5e9L8GTg+0JCL6Fd4zSLUqteHaChN4IDFb+p7u+L0vofVnJG
GKOmBjhtcIqzfL5tLSVWRFm4xr1PjUY2jjGaVNO2xgJ2gUPlCc7LLP1u59Kv7RIiJeIowI8Ziw2n
PcaMzlvojMZhO7q2veCB+Z+sjtCIP6twq4ZOs+VxRns1wp/DF4Pulhebzy8IlY0AxPgtLvxb2KhW
yPklIeTeD/pciWQLfJgtM2zcyUksAg1x8sjqDl588ypKC9XJzmcp41mnMKBBX0OytpXOwnDNZ78J
nomadPaZ6guGOJYC4DFjwdBzHjg9Jrpqx3X/UHdFuOkB5V3XwDZ7lC8vsqtVnkplch4dZeBsjx3w
xwE5Ej7DNOkzRvLVoMa7Ptsd/hht7vhf7dxQij0iBRexhhLpEhigwjSU0ZXZQn75lxdCZFcp0Y01
Jau7Ko2MMNYqAXnzo2b2Osw5Y2oIKTK/HjULbsbzM0KyD9fk0yvj+SwQBE70YtrhH12PqUH6niiv
5fEXtn1j0eGkbhFajyQFYUY6NKCebjCqT6nS4h/QC5qTwWzPsm5oZrEAXTU5E6H+n8+/VPzlzlj+
tZrxpP4kD4nyphTC1C5zDYLFwa3e81MRJcdErzbEiF53e3YBW8W7tIiSdng9bb+DAuaAvV6qdthB
gkxjjhoDQl1Lc/QDtfW3B9qyx8iOSS9CrLWQeIPdXgneN98Ig0Vrr5xOoAz0w7csbd1WuFGO1vfZ
KzjE4x+N8FhNT0B1xdelSWvgJHEeHkP+cAbSZOwWHniVV8+oFNeTwe8joTc05nUnoQBE4uiRXptK
HOAPVWw0wP1TW607fG6ROe7TC5XcuaC3R5OqsDVsLFKoU/Qz/e3eR3l3V3zRvF6kgjQe+GRN2Qna
g1FhecdODSJset14Z8kqTGhxxJVsTpv7k7lsOjIsf4qD+Bvk0OSaH/GbekexPGrgzQJmLQ1qZsHC
u9rlHZPVlOdbfgG6rlEE8TBaM4OewoyXz9sUvM1HsplzcUpGsY8XlMUJaD5wQonrI+lNeaOGGjtf
Yx8JW/ODFhVAKSh2fvCyLcJf2znWQL+DEU1Flzt3jIrPwbEoqjcb1H+q0YUnkUdr6XaYD2hfBEX1
ZQR/arWGxEbWPxEvoMOK7buKhE3Hg4Xt8UQCkzZ1g3oiVxkPaVNB0P+rYnIeaoRxRu1ygueMKbe1
JyiS8YxnuoivUZIBsDBg37Yw3hZuUDpmHfCcKw+dCbM99xWFG1lVgrnMktPETvDe8rWjHPlzbn7X
fSyx6D9Bt682TTyHf+2O5SSiOlaEgBbOPYec5M/qOpf8g/CfEPTDq1fmj6IPQrARA9iKPGjD1WJ8
tDurAphw3Su6wPuX3klW1wNUdepC2CUt5bOmXZyUjiGuwtcIb4t1CNMZ+5cn/Y+Gfi1AKIAEDuUG
JoEhXMxBpJYlqOrOrtzcAZPC80MdFhX4k/dL95plSzQ2aIUIEhvhkcQAN03aWdySw/N6LtgEUEF8
SkSv23o1cI3cSS9kxLp69o1i3D/p7NNTBafiyAy+uqfWa1apgJ1eCwh2au/k9YVGxmnwWk935mMi
tU4Sd11Z7G4NmkVs+A9uzHdfHSPWTPMfZgs3ta8PsiZWetnjcH6pgEMvmU/q6kJxYpUafQ5SaM87
bC7Cd/cWb9NA1AYhqJGlDNPmd/9vW315Ni9uRnkpZq4uH/JAkvhtI2jvFzGt0Tdogxw9pkB84yww
LEmbZwhD7DK+BMVh53mfksclbC/OnpXKe613YAkZQXKrnrk8Z8ys8y2wfdqyc3FGfMXKRPs5PWop
ox2LCzcJdTllzPCpSNcFYg3Y40Z6kOIilSfVh2mg+mXw4SUaha+za42XCGdJgA2PdvaJ/RkPQ3Ym
pMr3M+anFaPFi0b49ZjjHDGhWjL91HA5uZyEf6xoFvAb/yhd+64QB3at5Vv1ziVLc4hfnYpSBi5Z
iDww3HqqDGcA/mFWulfSQAONrpo0yV09TXYcKj47DSB92Z9wdUmdEUgUlC+FDYxUfmxI3qw99ToW
gPiDVpxFQk7p6KKgYQ3wGkhp407BnlSIEiIgC7401IFfmezkZHDaL9JaFtSG+C6V37abCKxYY4lD
etclyqAGaUsiodRi7+8bKWIM8Ko6JWu6uMP3HlbB1Zes09xDBTUE/SOb2DFYMjX5N81H+RLzhr6x
A9wURdJPvBOzo34I6fYtFFW1gk5ZrFKSbd5QB0nD0oLyyURW3189bG0/8og/T8HCVQzkhvT36POy
wh7uot81nuVghCLVl7vpsbDRkw+XF1HVCJsr4r0F4J3OStERVBCMojDYt79B0nJ+LKtPkiyamdOC
zm6MuDUrLTxjAykXqsmnpb4Hi+353jZOZ9zZrrtGTGV/2PQe0wig1WuyPEN8AqkN51S5UXgiTN03
v9Ulv/bIdayDf/5PnxpCzVWFXnceeoJ5wzXjZrmlkzmpC5h7Yr9s1eCpUniOJVG+SJoSYpIfibbv
xcJLaGlxBq3eqY4/IRxTbhniGQQbXHIiqfkpJFJ0Ng9rTqotTiUXLc0+Nq8+dBtRGiAdqmlld9Tv
bKFuuzyUQJbMerSX3POCbsjgDpzyU42BgOvInI7vgAetCm4EJRp/xyxmHVFAX+3Dlhxy6cdF22gW
gcDEhF9ojxz7bdNKNvwAtwQlXspUzN60lz4BH1NTpFceQd7xZf4DhcBya2WlcYBB38fktFYYfxH5
wXEtYcVfQ1hEJoukn3W6er//JvcOXGIA9RQIb5FZq9b5r2l+GD9eF5l5mQebS4Bb5yTjQtrsIcOM
wujIt1pWbOpPpcT0Q888WncvZie/1vZkIdBeev0Hik1fZMWiL6bhxbCwUXmHGAJYar34NOq9I3/f
Iw055YVS5TaPbevy2DPmPwOPcW4N8ZzCH6k41J03mu/xvj7kcFmmqZMuFKr6nQ0/tP6uFvR2JQ2t
wjISF8oFgE4H7OkmS4Ur0ZNb900TaiP2xoI4CXlurVEGhhfAPrnoYk35Yre+iislz4CO77tlrA2t
GPgExv4SZXKzTP1HSCkXt1SXbU3Tb14aCMqkKkDABVFfCT8FyOCchpB3gZf9TavtvrAznQw2gDVs
W2Wz/LCNVZ+JjS7FjsswT68+LtAUQtm9uTXj0tSBKgPE3lfb1DPIzKIj8n5FQwqybB6v2qB7WoNe
Me3r5rlXdbYh928VP0gH16bKCLyvuA5DKzU2XGdHcn0W6CpcIrGzbUiQhDlh93/+kWKlAXjC6qws
c909pdsdg+liXmc3i/mIGVeVHC/v2Ihm8W62sqcPu7gksClektQVk9IJcLXoC8EKTURinxjwzccf
kgqL69Y3AL6RQxx8kdoHQwueOSeR+jMDuJ4vPPBZ5jBuEy1To8h4rXS9tycS0bYGexgVD711SSui
O/D/d9E2JZUeeYznGZCPk9dsYH7shqoSD8P6GFoxWqFM2mvnLjfsS8NzQAAPGaRXTdjSqEnVPmgl
WBTD62iTT3sfvosTKjOizsAIYKi5sJUOJf5BuIcuYzTTYRZkmD1ZQkAIeK7cB/hUrgouCqHPM8ey
mGpWfptfxtxcDpseaEFofWYZfrDrW86w2Kbe/eZSnzvsFGfqf+H9TClCroAPjQHEXptTvy7iVPcb
yKn1YbHKvOqkNJckK5LuVJS48yvblbnbdMi9gzpULvOuJDTwhFt00MTnd75nS/ROTKlxkBsisY8q
D/a6jOtLletf8D4WpE60npa2IIpRYDVfvl64OqycvKvrnrRVLj9gEuxP4rhJUAVZ3UHtUgyDFDHm
7jTGI5tCDG5IjjrknhGt+XJEzJ24apy3V29iz9OuN0r8V94iSqZxXmgAOS9dvO22sH88xrFCgAo/
0OagNY3QW6W5SSCUgFSx/WVsj3cc3/M5y2z7g95TXUVXVKphLRWvi0rk70rO6EgPKeba0k0T8TQW
HXKXSpUkcVaHof/j+cZSs1twx+C5IPqGcVTRHSvO8rhpq3vNCZ/40GShz2AI9fAdetXCoV/712or
IdO9L1gkIrVWCiWZxP0KdmNB5jAryqCgRQrPTxMB3eOs6lLAFag0WXKlQgR89EHj9gBCYK/elgZ/
UsZwvw75eL8s9Yg5b6e1j95Obf0O2tiFBngOi9mZs9+5Pu6qiT7WaAIJiAfApezocI1aAqVKrhrf
ZJ6JoLDiVhnqJHlhRbcD33rvnZ0Q96wQIT6KAv4OoakZ1si/DodEL2k8s6EH5Q5Ja5OAZIzN4oDY
2COJ0fq/S88WSWPxzhEPczAyZLrC8EwIOHDg+X+HX5lY/MWKpiOatpwcrnNZPtIvi+oExBZ3n4Jc
0LsKbwifEdJYno8vwZrBLYDBUSK2WltzpRVGiC1pm+zdvQpKWkYJKnjyk+KgEXPMcIvr6svWA+75
IHH4pgT7bJbTaXtl7PNizq9xlALF84Ch8ATYRaIOF8+h8cDvMUPPdw7+/A4aZVT0bAwf1dsOtoz2
m+Xf65WHXaoBBztEDuJNkz9qWeZAmWbBkXUFZ1Qb+LrV3Ic/lZdYhR59gvWI+ZOe8gGTND4I8tJ2
raujZVssBFyPTctcMlmanCStn70OHEvoxjp6cUdZ1gbEfXFiReXSyFAI3SB/u+8W/fCVoA7n7TyD
PvHQQlX90uxZm0QDRcy04uHFsk9sNpBslc+0AWyFm1AzlZOLvztKTUENb/R7obdZgpAqnJP11YOY
8L/pjEEjgaSqfNEt2I4Pq5C4Jejt8R4+O0JYwt968WzgMWa48ZDn6TEIInNOBfammrv5iLOzcpIm
gC+qf4jgSJrIJGap1tS2Bjs4dWa6V3GidVH3MNvUdJigMqZ5aI1GuOM6dVaV2RLDyXwR6UNj6MI8
GutOh5hsnbUmzBl3XOfCkHfwuMMkYahdaAlK/H/8Zdxq4HGctZ0H8U8dA3fmbq9Sk9vgsJoOItyq
FP5pnjZ/3hFynjb8mwKOtwuAieQ11mKGWGdK/m9CS4M5OwBLPZOzoJzPx2uH6/Epl1h9O5z3Gv9V
ejImtzP9gl7K8hjb98lNEjMVxiqXvzPZkqq0o3NSCwZKZqMe0Wc7SXyPFfzVraMiF3CQJG9X88OE
5NHCrAg00177HFMtHWF/8UXGKUpH+zmRiY7ZfXrqa2DM6CriDIvxxSGjx4kyw64TC5TwnkYhBmsQ
qY+LVdVoiubylPynChsDpAfJqZXtziAsuqzOsqkTDfJmCt2DJEMEk3LRRVRnqLHP6XnlOPvn6cPe
+Vvhw/YtpODdE3dZxsqAisxMIyefMCG20WoojHeqkPubtknV0KNbyk0wlVgPIjtOQt0eRZkEIBDh
sxC2tgWJ2Lp6F/LACJFzvSAYOJ6nbRHDgJFHG4MUug5Z8Z8JG2rqXYN8EUPb6bjbfltD5KFy3NeP
mXTvJZUB8e7JlG/lV6djczpd98P/1TiciU2WW+r/SwSilKvAbA4dTmuzzV1mWNxlrpJ7qNijaFWR
Ikbw7rt75yJ1VhhL+2DbOz6f/FznBPcbwyqXPperCGvAmZUjeSN3mP3apmXhBs3b5DmNapQG/v2u
50P7b6hY71t2YT/FQKpc1wQSBb0lG9siKUQVvsejrhXK2vV32F/qc88zrJxNPuXjtT8J88Ir58/9
RHmsFFePhMM4eoIvcJ85P0XkrP+Kb/EavVYdoy/V9lOPy4ZHjAYCNLfQRDrc8uJzXUFqfwM74TmN
EX3GbE41Os58Us69eueZcitS9Zd9/LY5tgtmrB+PqWfyf19JoaLpCXepTBiHuCwT4x/Nlwe1gmWm
2H+2cgTIcmSaviBie9dMgCbIx1d5h24LOhBg49BBUHnb2lHraoVTryd5NKTOvpr/YKVZmHvbl0F0
GWRWchnxXnn4xZWBAXXsWYsin9zgxXV68uNs2tRMdK97ma45PkLruudmYFcoaq1TddqVhcTBDK4z
03LZ1goN+u+T2GVl9kUHp24hOgoXW0aXIQF3/JtY+HZ3AZDDXkaCQ6PE2vdac/HLdya5L26kTlNa
3bouv2mzI9tuoNe4ihHiQSiNUzNmSipoJ9lD5hTwn0fRB0GqFJ3pbv6lUYXiAHI1Z3ATESDL809q
U1aK4ZCOfk2SRphxBR/aw3r7ZxTWrBbZWWJ15LMViFnzLLE+lDgIhXeEhXucYDcCswR3peWEY1h5
zb+ZQJ6vAtP3EAeai/lHSTNGgt4nNXCX5kejRHcdhuUOMFJCIB+rO+6kv+RtYedyF07oXXasnic3
FOwjxHf4+4WYB1AREq7UX+vc8evEByr7SCSiy7NYE/HznoafsWYC0L+e284lO2O81wPOjJ9aUtaa
+rxFOTaLT8qN/QDwH4nAAyhB4dpifxsncJhjnwtyKdW1pmbloUnDsjTpuDh4TU6gwS15YNHhnNIP
fipXRdqL/PHFETQvXemndSn835qQtNMNvmnb7twJ7wjcvhoTfZsawN+1IdbLfCZKwrki+yoBNAwv
5m7m/SscuDo6aZDW3BTziSkADTBFJmCkanDiO79Agc2vzGQMs3eCirxfnYIOyp4Kq+OzG3DXVLfz
JIg0kNo7d0xXkohjZ02KBwiqe5EKarfVLilMJNlwb+7IOd8VYlvzBkWv2Hye27OSbTkKMuB+9GQZ
cZ4kaOHtkirhTuePWJv9aibJZUE56XKVZCJ4hGTbW5QWHXCDySmLx2uBQwYL6BX8CJSvuaPpoEyW
Y4UsQFK0/rN0PueWzao9ZZ+yFzsTh9TJxLbhxJaPNu2jFTc8TOs/Nn5VDy4DvRLiDrDYIP8Be7E5
1a/XIltD/F7pZ12ihlz+yJszgvnATffuq17Cs3mXkgrYcBGKGC9dIFxGWhetcIUynqZOwXb1L/4T
GcEonQuO05s1ADoKpuk3Om0slonv5xM79f6FwfVmCNAiJoZ5bqi8iIOwIixVcHjZF+AuL/j88iYK
CUuxst9S/5vnlV5YT9JaIgvT402Gs+8NKh3LkpSFSnsgLPBQnNvJmcm2OM4tyOt85iz4ENvdHwOg
LF54Gj5GwuPH8qkh4fcXwC8hUseHPzKCHZpPcyin7SAA+UIkQp4m87Vi4UaiowBZ7SNm/EnhmUQW
X7XySQkxBMxeHaxqYiqulB4sELgk62DTqd2B6Kt0+4Ho1jav+cRQxMdnkgHPRf9GtztdbfKe+ugP
7YG/eDAy+FSXQuDE86ib+kyG50PGKYuemgF0rdPb17ACRlYhlzsgr/XdoqLWS7JMJ5IoJeIQlt7y
hIYJyBeKpwWj/tDE0DOFV8VaEItGdt868kcNTUvE76m+AxP2L69gs3vhO8tpeN6bcEeKiUGv0eYF
fh4ycxhmxU4rT4TtZZTuXLwQWap7S9/kfzDFM9lMxygzYvOXmRBcE5ucNxYYLNRdNUGYLm8Fzjcn
PRH7ituo+48huXJecQJLjjKlOhY0w5aGfXQQDGqpwF8DBpt5Xfb27SCpnSGqV4I1X37r0EpOJPc6
JY7WH2iJh9vE5UJHTXrD42xYRmIkCYcjQesVp3wFjjaKYgjmQrkkmAt7u3ZWNenIGFnuYdwOcqDQ
LaAv0/BdV/wQegEEG5Nz4SO21KhLzhZ2WEZQFYEnjIp4s/EU3HDzkscJZlQ8WUyOcZpM2wQCW4WC
V6XLHOdDMdSf1MWNcNxUyXITACj1DVqYW0esQBevoPW0KAdQr3YW5z/+ZHs7lh0U/O7gSGMEc/a6
Ia7qs+Eu5WN+D071X6iEYqd0tX5HtEwj9SEDQ6vr4LYXDNILMv9R49MOZAssERrEcmrH5Midq1OQ
gghlCnGKuWT+odH5XDeIYqKOgSdw4S+18RV6rl5NK1JxnURt0/HVfN0TpnNqat45xAt82IXfXHNl
5p5dAah21gtijUqgNZFzK9oMgo+JBvZogeRuWstv2GTrzmEtEPxgkWKVPWRKbqbnxfRugOwxYG7E
BQc1rpiKFJAgyo3ravU1p2VwvhpC69zY5iFrv47mSaMbcL9Z2TJD3Txi3JeGALcj3RNply43UU8T
QF7h1WNl+HXu8YSHn5Ca2DoAopZ2m+MhelzqHaZANSRfnbx88nGRW5AdY9flOu/1PwQxxKdkR4rS
hQRDoRFHpNFs58Rkvw+uqjKjDqi71CYpxghtuuPcv5wMvSaUZIhXmHnvPqUa46jwfhRb2HrJoQiz
37EA4rD5mYLB5rJgRLQpXlt+r1EWN0WxpRRO1Qa1bRhyAftm7MxeYplAk4/gJf/q3pBpSK5MJmXN
efri7BR1c/aWfmuTn0uaC+BEPLxHUtNpylsR2CKztxZzoR623MxotIDjNEXuzUMcgf44zp9O8Izk
xHtooGe61IDHaQ4JYYIWIMPBay57IGcBZy+YKvAdgLfjXreyFMbMBpqcMvQjMz7Ss2YNI/mhE7xs
lXCXNRqOEVId6eRHi5hxUTh+sdiF1WyZpiQkacpjHaH4ID/JluNHVNBwFhIbnfL1od9gDSdcF2sE
ZSq+HuvSVKORiwkf63lI5FswrZPHOsQwTCzcDP16Vo0QswQRLvbjAeheHdW/SSgVtKE+1D7EOwOZ
i2bzG+flxDgwVeNoTN70Xd5zcsf+coj2snx0UPrVz42Tx/pKWg10dzG5IxLgcEZNRB10KsgIvU6X
PWtAENxSshW6VQhBU1btMLNjL2r82A8yvYGEhWYHhYou7kSy5pH25Wg47ILatiH9zbgGE5YsbYvJ
EstZJog6q7m9LP0fE7dDsr4r7V0DDxOmMhtBOLj8a5uytdaGVW6ifmkfQm5TNFmCV+HLqwA+F1Dc
mmWACmdvwIDEUiDPLqqaWqx66/gAQOnAXB7syLGn0pchGAnJN+36GUKLq4DbBGbAdhPMYb/q9rvh
PvShn088uEVYlkZfu3GPWaqzqrSNkz4h1E4QxIYPA11B3UhQY9ztSKPoYYOPHxnWOw90I2a5KvDC
SvRIHaVFjt+nefBKwbOITRtH6fes411sGXySWaDJe5qlQ0LmUCNdXz7Gi/BhdTw5eUVJVL55LprD
ysDoFa02D4EHI1FwOIIFAXGt5vDhpwA1LdrZLT5nK/CkbzRy/TO6VDcxYWCqtemFVMr+m5ax/R2F
sWcFEH2Gc71cCZ78nISCW8V+zjcbIOhvo120Lia6TROY5+dwMI4rhNbrSYj4TOhpq0YEst7F6ybD
88aNIdPppmuiYPyfNT5flBepdtKVy9vNU17bVS23RWZW7mwTuAC/pfHG/utUmF7EdS8P0h3h6q8m
MKCLSmCF0Hp4YG38al4ZkZQpiK5+beV2Wr1lqprIvirxMtG9Kp6YnhIjPcIQBTiKes1ne8njlvZ/
wXU8Pi6JlHpz5nPduBJhOxxu/ugEOuGSGd719ZrxO7mpEXDys1ryKQ9+2zT0fYlJjoRHPh7rdgki
HS/B/q9kKEGkHv3uIJBejlLH0TGQhcklNCRqo4V+tT8duHYuWh0E2eLBJCq7azt6y2a5BOOzuVvC
S9xArX6UsC4G8rCywEpuv0B52UfEOmdDDvMbjMbp4QwB5YZmzHbMnoheSC8r65bY2jpPUgknjtKD
D2dthlIZUwCtAvcKmaCT6i2df7aBFu/CVuT6hCKdaeJNewHxAWZkAB1mbHNCD3IAj05HtqXP+CfZ
i7O7BNimUGesXNv1CEQWdSIPrZecuk8IpObvRfoDhOitAc2NpGalYm9uv62j64jVe4rmrDHZzQxq
0yMC56uVUyz7FlhPNaWLABe3Q2fKhMWyr69x7YB9/y+28/SzsVmb4fSDORjKfqz/2LEhcFGP9FHn
Jl13j4e5jmg4zDHJ9V5ErfC0mf7p+sJPxNN8yEsnay0lZ6+o9YG6vonGVwSQ7x8fOEPfNUM7f2TB
FYebOUI434x7DmTZtFbiMyOCJJU5lBKr37RjRS0cWiqQRQV0f6zbE4u3zQYqTmhy50ppzj3bx9YQ
DuyoiPM8j4bEsKDoAp4HdetKP3F75riS08WFkhrudxRE2y2Gq3h9sKusyQ3UOuSjx2gQHGCF20wF
oRwKwIlt6eecJBSwBxY4IhJeNw+3w/+6B6goIw+Nkxf0twaVDLzcdOGx6Qg9Mg97pg/J21Mtexa5
w7iYfEHDKaJifW3zI/tabPqvuAvxFTmiRzoDtcq1w3WpgYJgJlTmn/08zv9LoLOy0Cg5ugQBAkE7
92J9jJOiFK+v9FqgQZ3S6gKCdEEkU7mgG/Fxhg/b4hnfPgZUFekxU/sqL4dWvwYMe24aeuOOsVDZ
oC0sCmivrSSEZh94GgF4g04xFQLY8rgQ8cSJeq0zrDtJYi69mpcytQMRdK2iuwX4TSKOUshbcqbX
YQYwyjjgv/HwTld9ocKsEVNVl38hdcEzxT7WDnGQxXY8dfrcxXNNaTbUbTKL4O/bCDC3RID5/ruJ
cUlTpFvXvW8X/zGLJ+eiQJeQ2ZlWxifUHl5HcQaeE/Et0ipmxGjhgBR4qSbwzFkNBTkc2JPhOINE
/t8FNPYolETJoQAKJ66kQvTZ0cf/VkXTdrfcYzftAFgm+BBVyySWHKjAwmYbYLa7C9Zoh6PDsveb
z9CjXfYuMxY3Y3V9kNAugOPXud9QSDVxgf5wDlv1Wg1eJPj7i7zZ+J/M5qq5XGZ9nFjRszK/c/4y
G/FJ094mEQQe3jG+QYUzqdDcYohdrhFZXCfPkOs5E+XNMRfgnwO+M01c7oZZ+6qbcwaLyLC3d5nx
FQbZ4mZ+AdkCcKmBSbj47nzQj9xubarTK4J1jdnXAKEPjpfxTqpsKOmTbpdSZOqugnDZyavcAx5L
qAW/UcEvooC3iQrcYAXJbobvhu7z122p8UTXEx2BYC6URbCQl09WvgG6TdgBrfJ6G/9DFStrPuza
ulnK1fvoh5ztDRppyRmKuJEIHZPIPtf0gPEcwpWSO9JUHyZN9U+Ec0sbF41WPCsvE/6mLkITG/vS
sAWcWO2KsSDWSRaQE281q1ICq3QPfTx+uh4192BRlhDqlQGwTeKvr6yJu0dI8+TY8f2z2umdCvsm
fsF8G/LrKOPN2+/ic8YtjKhaYoP52zPxx6PBO6oNfxO3XeOnfx6V6zQ2HzIOHMZ7mW9zWOq3aUXy
OfEH/rerdvVpvTU1tarWnHUHWK2Chz8Ve7CIdJiR6/KXhjLsMgU6zbYdNSiTbmdbQcDQ/G88+6ei
ZogVHvBVURkP2dgOyjs/0dAyCcGzi5mCfQ39jIwcgOqB4JyvK/m68C23yKnKDfxLLK9uKIj+UyPS
RikmJuFmZ9tsrwvBQY7kFSJ4JPZD/molas9CkDs4yeRc5aoo7FzL/JURBfZSMm1mlUZ93ej9TORM
ouX6mSyQZOLp242mapPzG/CX9GxnKLx7RA5fvs4kscJqNU5gKnDdkvitX/CO3O6B9/5CmyPWIYuY
Zd0fJxu6YhLJxuYSxvlYdERaPEbjTMG91Js2kqvz+T3Nv7YQz4I0ckY5dU2R9Oy9iqBCVXCt/AlO
yPzg2I7Ue1FnvMVOJ9rz1oSqKEUsxALasOqL2AvD8na6Va3fXFyqlutQdw/SFC9OInsDrnISxomt
c/Z6cPuTvGmo3QvXOQNsM7oeGPsbjnmDRvCCr+B8Z0v/pEaznh9OrGiwlEnZfub3j+36Hw9AMbI4
KbKenxZ3rUDD+aW36f6SYNWJU53d1NG2uWjEoee0gfce6ifShuLkvzGrjMK5A8yaNpUkaC8XE1yO
Nd3Pm/bm9kvgkJ02OYiO4T21kk2khb7UiDpXzPB+WMg3qql9IsMTpXHBjnjsD395XakwYAPi1xtf
8mO9gDAyCJ31sfcoiPk6QYcpWYnBDAoo81m515Mog3sMEz/1zXlRQTcrK3CEE08sGKPuSmT9VR/O
WQAB7CsFRQ8N8RWcbXxUkjdXmq/XpFZv8+m8ERPFNA3GVwMtB4LRxmKiuUXx5uI/p9WuseR82KI9
Voqxx7aomlz51DW1YcI+Qb5cjdo5RMFfnKUbktl6md8gXZ453jQwG8W1M9wpXitjD0O/pShTxn1c
i4mjAHFh/X6W9pO5mhLh3pcI7g6CFXyYHyvsileY6Su0wtN4NIQlwWEuW+VVMRYd9jhAP41fbvIH
82JX2wac0NKXExfSDN1DsuC++TZoCm3KjMBWfErh/pItPpyUcnzFsA4QLNptvBLaHClFwOa+liiR
kcgtbRbZADOmQGInRLvL0olqrQk4EycV4VBo7o24xbNkNP45lnZeh4rpZ6ab2DiL4MGgwyJ91QG6
G4CrzPa7VFGMoseATluROFS33DSUS5vyE/1szx+JGhlUe5Z+2SM5bGGDFZ2KDExsV+Fbj6QzqkxO
2MLU8joDR3DhxdaU0eTvBpbINxt/0MhCvxP2zHnRY9fX0+FI/RobGWvUD6Br04ql2yxmfgWwikna
ceUb4E0PYUq2UcppBugPJ0xCulXj1oqBCIXuINGCMii2GN6FRGPe/xXcJakDtIUqVH8lvGld6Ina
/jzlWjBQMvTFEkQZZrQMZGgDhzKjnmVK/T6FZJbXSuJSHk1CNLUO//z+CYqtuJ8glGrhqN1rMAAD
IcIl3G69Qa4OyEqrl/exn1FMJNRlkjryYFV8alxrbQPEEKDpHDdcxcEPrYNyEknJZ6pQ528Ai3SP
iBUaM//UWirPmbMM7a5Sw/bsOIRQ1DC6C0O+39YICg4d/Mc514yNZnd91Nx6FccJy5WOx8G0ronF
FBITCGw5jmOESoncLCsYkbwON9SATSyZvRwQKi6vUmuykB2YZjeezuha4FCwHs7k5HH503g+6r7K
KYDImj5AgIAMUpvKKbX/OZOmUH/aWSJT2ZgBGqPSCTNzEtb4378Em3T0rHm/aFOn4/y0WDB/bszZ
uEAvR3fFW07ipnKgu+bDbkZaKaVcI1K05fyWC0qxPRaSBjZpx085WuugygCv3K67YnaGDRKdM/X+
aeFsArWOBruQ4Y2esnqgp9EbxSowW+wV201Ziirf2/8c2CxkN7b7WT3dI2/DuAm1l9eeypscBpxT
bXRyVs33gx376ef5KDhr6mvXzq9wvQmM3PaxdJmv1k7cvvFFDRITyD9Xrqx/Dwzj8nJA3/7yx6EF
22t23FNgLUdbZx5iuE22IrEtUas+OQO4ZRMl7VtVj3ptjX7T+JkeJhF+UWsrB8eQJpdvUxklLqoj
u15v4bsHiPKNrlBspYvS6wQAUytJ8J31/dulw9ZgMVkQ9luPIHql+FthhR3CjfEa51mnY33HtOnV
GNCOL/kNYR5LKhNgo2PcRKQRjI/SWF9w7WZI4icUTB/8/T8WkzpXquQHrLnqugvUNTCAsUzJ6Gp7
lVoqFuo1EhIfoQU/gR997gF8cORaVMh2Zl99+kTRFwenEIP29hSRXnZCFO8HO/zMGSfqFa15GAWF
4cxZ7BpdhWbQK06HOGmG6pt2G3sNrGErO9IQLJ0tjljE66zONATyccbD5Xv6prpBkt6Sr1RbLnph
NdUzTUrQaT5mxPsh0CZ18K4pJdgwuG5eFymIXMPMn1hbpdFZof8lzEqSXf9/UiIWCyzTgdelBqPf
3gEIdWLpH9wogVqwIjj4UiBtD/m4XfhmeD3FQN8QY4kQml3iap1xr2T7qNmMFAImHdYcxKMPqncE
Rs7/A9PkOW/hJn86ZQQIRqBYGYpQCJVXgWwD781ZRBPoPSAzmUXR8xCoiFTpJh/jJLvYSEd+6nv+
N7b6b8RwduxwfYW3k4Suo4cWRJIuPpU7vayxZlt4jUzlP9bgQRhlZrhsVuV9DXgrqEWS3y1j/WMs
SEZU8mrnu+DgUAYC+psD082nXlvixjyMBBOtEjaVLN5KmyYV7sego1hKoRJ4c3DYD6d9CWhfk4Rw
sVZHoHjl7ChEpT7flIbfwoSFWQ4xTZ8pZuL6RtDvMelHB5INy8mbO9h7ecGX7XRMbYtfCzSea1D4
vjGqYgvySKpE32Rd7Pxfjb2prUtiXCcuwOslBsDOmNsY4ZSq9EzteH0YjY8S5GztUhK8AI4DXJdL
wMEK0nu1J5qJO4XziF/iAA97mNn/7f6nC6iY8I9C922isboUVsyX+tVyl4i/mzZgTpxbw6KEEKPH
MM1sUZtegFBOn0Dz7/Jcgnsm+2J9DbwnfjqL1FWDny6AYrvSPNE+IyclrlbumXHtcP0ozkTYG20u
qb+g3DtE2Q6MLSfV9/khbZXFzKhwPfPDJBMGlRPC6wVYtodIgc95Ep8/kEBF2jugCvNaIviimLoT
EwiiuYxAEwAKq3NqZA6T+bxxBdmuYRQRPKBDXZy0vNpAYFFgMEhKUCbZ17FDMX5Gyd/g6lx2xbjR
un58odMot4LLc86rBHHY5NIlaVXWHV6YE9LGwYQuCx966DAhzCKbozSndBqXGAepyN1/D3nBORoD
WG2MZln4S1Tq1ZPhj/yGpFpgTmXztgX328GozeRDm+3xI3/azj+ER5vv2sFaRa1KUzETPnV4M8X9
FQCJCSYwa/QSfYgvnSEQZ54gxCQs2tkMAnDVdfj2D6OSGTrfx0f9BSkXbi0nt81uDg/VdFoEcnIu
Krbxan1ml+/NQ8IYrVs2OHXUFmvCIcJRPqA9iPqOawU1L68+9QmiJ0Qf7/Rt2IyPvcEk3Q73T0VA
zyGWgJHZjgjEDNPVaEDQ0UnqTk+SsJIELE9lwRm9bB4HSa6JJSAAy35gvtZgb9iEk5uCEtTbgGCC
Zrqyrx3M/xRvp9rkvABr7bAPKPFIwqnRWqWnL53Lb8cQFN7QAUuemZjZViIwcaIjol1aa6wWx04U
6St4E0Ba12e7czMg6RgI39XBhwpRqIM57UkFs3otFdenJ53yr+lEMgd1HlpuBYhXEgPVMKzgkh3k
8mjbpP7ttmQD9kkQCcd1Jxu/NN/ZCk1OhfCDm3K97fueJN0zBU0zqnf6KFHxkw8/iGqPUgur4nT4
Er6FXKqPMcrszm0aDi4Smk+egU8toF3E2j4LnmwxhDJB9QZFZOqrmXUegErOryQz4jHVJb2lwpbe
rVr9IpAMO/HIH147AhyWe3yC/HoedT+RXpnCaNaW1fZchf4nWB8Okn0n9R3gBQsk5hxYyv4SKsPm
L9Tb755JP+Rg19FHOj0wbMJ0A5aKHUqq8XrMvYPknezgHUzZKy+9KQj6++Qt6618d9HDXMsucCL0
lCMKPF2k9uMAjkajhw49jFickuTeAHtNhdk2jZiSL8yw84AJQujXJeJNoOK/Bb2fRvlbstwM+uaz
KFufRQvPBBY/hYwfSkHE25D4bZcOrUXxKfMGlY4HDecmRpBur/mAjKeak2dOqswjwvbz2JUwbaCR
OcEFl+O2aEsB9tPR7l76HysPXpUBJfWXbKX7dMpZLDDxjumbiUMGpcGrbqJE4FlitWQe/kdwg2Cs
5+/QFW5NoczGlw/otWSv170rx4+/MFrUCrlbIt/lRjolbSx7rEYGl4wUhk1tQKw3YiSB7tQ3IHMs
d/l8qamuJgw1CeWMgPNAQtk/idK5eA9SAugA/qapEujnJfRQaalAloc1zB0iIvoPHw364wLAVtqk
q7GwaSsiUWhuceKNxPySM7I/Vv33fwjKB4XN9WAGGoUs/tyDMXV+jzSllO+xz3tgqtV/jLXzhQnq
rGTJaa423DgLj/mHGh031V04bIoOLQW8ZeJEn9/LHjd+7FbJpZCuM2EWNmgvPzDNGm4Muzqq/7gh
tC5HuH1aAnYL8gRcpLa3v0ZbC2sROr/oESH+z5q9WxUv4p6yfh/SW9eOcBKbjXY2RBGPbXZHjZtK
w0l+ckvJJLWG+2e8TWWCfb/8mIqCdI/h8hep6HjTZI0FLpcnPHSgXaUmw0D48CWdw8hxYqWCZQp3
P3wWOe9ijmTvfFTyPfrftlcCswHG421HgbvAs5KnW3fkx2cC9+aIG0CaHD35x6E43oHebWEQR98x
orQPyT6QrfjKKSQxjH4QSXYbIbl3pyFLNFCKuRv1fDulh+WbCmQtdMXtXC/lpjpkGttJlD+OUutx
a/0HXaOeh3VJ4WhYiFnfVH3GkgBqubyslFsx6+iP1kfq3Q1lbIe/ELvm85KlPwJ+VvkAQNTCKYpG
1ZKjXU12tLseqZkbkLREDZOw+Mna5mFMopbLt53ehnwJgnGDKez3cSi0WOqzjzqJlQXOqHB3O0c2
vAnygLKLe25q3X37pwc3J7LZ/H82Y071fV9uy7NLs3O7qZM+/W1PPOTWRXS2GwR/CikLO/uhRHai
fOLchINuzQgjA0/N8IcHd9qI3iqPZX9f5+lp9Ih3GYsuisvavUUQLZ9F45lp0GT0XfEE4G/ZJALC
1Mf4cf33nlRo4PnjVjGcK8UGFM3e+bdkjNR96N4pQDUXLQrfs/QxEnGmUUCtot52BH29h3/9rSTH
BmF2cB3J5DGF5ptLDxJ3MDeQmoO2RlOGH6EKI5yDuroL3mUmgbDTqDHTSLc1XD3tpeDha08XzKYz
2SQLhhnt01MjT7nD+ps6uQlf4KZ1hvq4V0maxDcKkpLBYSyYWp0pcs9fLU9bO6ZHECt73uS2xdJg
qvmqmQShW3oIhq3iC4XmhIdyI2duPj0DXgoKLu141f0U1kQkAXk5m9Q8ZeY+IHL0QPvx1CCBpEf8
qlbyQ5RZCA1vtzswjoH+lKDmDjOmW8BMIig1dbjbmfGw07sV18S2Wk9+GwrxiQT8KVWomzOA0bOW
m46+Phv3GFQL8nd+2mxdDNP2q/6LJ78wCaqyJgJ9t5LR2OncWUW9mtKiYRWAWln8ucYgqLGdcf1P
At/k7tWMUZax64rJ7hG0Gg4Va+uY7t9NpvU66+JOvlVgY2fcod+HFPwOb09VsVSK6J7UbVTiNtoF
LQMh96Q9Yh6I2ME7jdLzODa9iJNT0sGOHNRXiR0aZE2TgLhUuPn+aSxaFBUX7aYAST3XnEcViM3o
trJE8NPALjzoMhH6yg91OfzzZph6LHWa7XZKdutCD/LvjuJbizfo556OYsoPWlOQbGGEMxv0r60O
2GVSdTUUBCbxgkHzSlgC3KECajJZvmFF3MylX+sKxgiqceVZuvlEB5ozfn1nQBJ67sY3B1lx0PTu
n0uKcJjMie95RJSuVsICfxjemm4n2JHcgoKwJFkimSXOzTTKZy1L0NX7HuPqMPq1XkaeJnX82Azo
uhuV4p5EcHSPxCMqQYDq/xihSDlktqsik86E644mXPmkHaQBV+ZfaAB6x4QU+9dbgiySTa6tVHZe
BWpNtLCRSphf7k/RaIRUk4TeDtuNvLTqzyLoJlIqZ7whg4ukV0751kDD4TX0FkNx/Tkgr0oSszKZ
fEPg3oPepXeEEawrL/zkaHWvMy6gpd7VF3cVBA5Y7YJnN2b6qAmJMqCJMyvnBlnRL3slGuTVeSYD
GPzKPBxw397i0dE+z9dR6qrghTk2ceB1mLVNCfBU407oC8/GLnB7KZme+xrYEf5vbp2ooAO/jQ37
Zl8LhrtSN4IU3qibFUODfPWwU/ASaLCf/zhx4vhNjOluX+kgS7UaysyqXunnQjvgAin6u5xaZ5dI
iuOn9jbiJ0BXseIBGliePVclORbAorNS4ynZLySaTPlj2DF0FKRGCTtzyuy28wJZowNvGyhMRiY8
gZzYHhwYbGB9YJO7r8HVtZ72utJGwBj00XGKt+ubufkdJA7C8V/ijjoQlYr6KuITRm53DNLSdl66
jp5e4yJshsDbWC3fw7f0U30pxMVMtTJSdrP2HmRwkUuN1NQYL5gan5tiXii7hTKhvwj/wk9Jlyf3
IrIlFSGpUP9RiYe5VKihpVu9CtMrHtj12S0Fqmxsh8ElILz/Rvvsv+M7Y9z9LcT7oPSxMLeDshH4
fQ8ehwKqTbZtc30zCzuhvmekwIXFvBRtJtV12mzz3rbMLX82IvNno3rcH5iHFl1y7McX/s4JG1A6
kMq/uOKEh/Bv1GEA9IyBhJIkyDSbuaGPkXZJDMOuuQ4gNk0MFFEQ7L8s482Nj2+f1QT8nr5bC/AQ
R/LNzNk8HEGnNOfTDQ317rp77YzszVbc8g3mBWSqWOYvcKajE7/ITeOhZxhbRJKcJp41Gw38V413
hMpmCWjTklKQI6KXr/Fw63tP4qPOWu13+J0KP5r51ifvcxT10K9DvrOM6YQJ7Df1Va4zZI4d9nsO
bxNKMh+FW6fZIhtx9kViIpomdWFdj/F3voZ56jRbdN9e0ZgMCahhsHFpkRcScDS1TQ8WyaQHXUXB
HNJWkbILoD7LRafIexlQRh3dNDLcC/zaelBeRozJs/7QMHzM6LxRXwERPq2awAZN8JfFR1mHrgZL
STIw0BtVJzq1PGt4xyPX3zSzrBHGKJhrUrZLeMUH7P/CvZUomBIukkInVMNk/0+kJOH8n62NodXx
PsMsNDUDyRstUATn/x5TRE6IhD6hzDWo7BWR+ic7PM2H8Dpl/4HpKAd36LcSIGpsK+3xYiPSWhMS
TBAJV1XqipURkBYJQR03qQd1gxAc7f8p0XL4/aebwXEDp6LzCSSl1R5JtGkfBQgWgKdL8GHBKItH
fzmaEGiS/yQ0J9rnxeKHQQa0jrcyWl45xo5TcV0+i0/t24kWVysxAN1i7t4Xwx+cbsErwhqncZrw
WRB1W7yIFqHVjveHWuaDVQwFbQQ++Zx1v2xZqMO/boLHnw4cUn/lQ0G/w6zcXw8itRcMkunf+Ivn
lYA6wVl2J8g9DfR7kE/CBOMmXMDyUU3oYpOPz/edYHX38mNLp1F3k3aFKa1Sn0pJQRMlEtxs2MO5
6BR/LD2Gto44v1BCPZOlGp46prZoo01sxVz/5Sllq6xoxR3mUJuw9Hk7MEMVcbdTB96FmFBJQBzw
dsWjbRMqpoIbTD+B4lo9+N/Hi50L14+DnrfuhisqeoaYIJFcvpYGMBOzPIShMfz33GlO7Hv0lQvd
OLY9x+zknBKde+DsuTQmjpO6TuYuWNbfmEhRM7KznKYrBoYS2R/dBzHgpazp8MaITSuxMBjNvd6E
ETZq27XaCOEKYFQiy6qi9oCcig9CmZDKrPdVQbOAwh7Em0OxZuUiKevuIz1jEmhmGOZnzDDoQx7C
vJRMz2e3TXFAY2v/cS8+LAhu8h4mYJ7Iv0Yksh+uj48DT3k0nLmJmG7s2qdfL6NE9NgMs0NQx4+J
JcZN4stGLBeCC51Tyb8xA6SaN9MHJkGZS5SVwdDOjgTXQpAc33OTC0C4DpEivp33pX14sGJ7BPh+
dS7Wahq6xOvM8DsyGDzkfDN3Is6I/7adGXsHgInYLAH36Gf31dvaxZq+/rWDABUPnLZyldUzsyFP
o+Hr30vnrFOhAzBXQB7Knr8rR5LHYAQJPEh90+xtPv73gMuPQOtDWxCzzbFp9hCKp3taMAxVv6uz
5RJFl4CUQh+q3nd8CYKPnRT0VstlX8decqR554oBD4V0TznYTC8lPa9thZZPKMjQSJxJNF+TG2e/
iAZZILiSa0lYzZp7GR6mj0kph6btNHMZpONxw7UglE16lHfhm9ab5r4tqFBsms+x08EMdaVG2F6K
9YM2KthcvEM5PXrhv96Fx2lkgEL+yt/T/4FJDREIvL0qUyI6VOwK+s4NaQQJ/izgbdteU8IHOUk6
D3RauJG7FluClJfWj0/iMxomtRA4uZw6Rvgi14hJY4lM+MDKPKYFH9i9hUre+FklRSZn2KzMEpmw
NadF+XxTByPYPyH16GdqmVq29EDZs46eKjH4V17i+z5sCAlbKcRcIjkbEoSC3Mn/3XX/CyR5DAct
KzcAsH1/BEjDmjtW7vv/FWciLd7qCG3xraOEgzqN0QC1Mp2BfQnQ/jgZVMvpmHPlG0VgQow7HuZy
M0azoZFYQ1K7zxv/Hh+Xpg+cSiTc8ckCDO7wjrxvUjeHSn2CpX7HunlM3NADuV6fRhLR7kHkO1GS
TFj10Y73pZ6k3crKd4SoqctLLZieZpLMZ1C08AOi8Gc0A4F4Rif0Hk3oCU2h9YeyMBrz2Bpv43/x
EedUEALBmOzcGWTDc/E4KLdMvKKdwSHwwagt7OoPi6+aaCJR9jnAHXZfnv+umWDOGiL33vq56iW8
LMIiGQZEOGb5a8O0alRqR6wFMxwrM69PZArvN4WMZaOSURl6x7p1JDfurI/hGFuUr+GT8p96QYbJ
A5A5HDvZYHgvA0pVPFXx5HcWD9tJOxCP3rjZJIhmSe0xNMVZZMPkNMncOUVJD8pDTpdMi7RJFcdS
NzAaxjfwDdPN34P3ib3cDUefJ6iH9lxCRJ1zUfYXj817T17BNvoMsTLMUEXHWlAIBMMrTo2vXanM
/L3sIoS+rNfPEnvAJ9k5AtaYzxS33nqRsWxCGzOS72irKo8eE8aNVGMVyUTyrnIZX6vLkDXeMPwo
f/GtpVeeEeQkybQKboPRkqpxXAwV1DE+PdHSyyeC0eb8BcKrpmlAR8EkzmaLopOvYLLv6uxE2JBq
vK3G2dKng+YZWjaV+lQIlTUsvp4rwr1s1lQuNWV/npGkdyFn9EAq3PP55wM1uFsUHnnKegiVDx0E
UEcmr7CxVVrV8z9kAziIPIApm2nlu6hltRo3wcNcLu4+n+5dh3rZlXLddqQWafoyB1ALVTqba/Om
D4uDVyUSXj45NtGfyQi5noNO8HCOKv1Gpdf8SWGjsdiBRP7MSMc4QMl5Y5keMidOw/6mcun0qgQB
iuwO7+5jWy/gVS4jrZO5bPIIkt8t6NQ5A39s4sIcifL960nLQkhpC2OrvbOMw82c2jUhVKyWTMXQ
rN/QN25csyrhQb8ZdkY36fQJxb1LeXO86nJkfTQIe1YKQwV92jZhhqfJKnUJcjdtW6fuczD8F2Yo
LQmBHx9uQuwg4J6871/l8bmLdaVM1X8DMjG4uUEmCqpZg2lyM6e4PDbQgaH0m0q2UiTtB75syxOP
8GeIpsDjwgihnnBrvZkoFUq4HtLyC93bWCQi72JGZ7FtOICishl0Mq7afyQp5S9PMuRJu7Z8SyFJ
NvtltgmwGvKP3d5y4z3ANd4SaAOQKyYmbInm4+8+IYxpDhY3YCJ6HwPwTl1HssemcLfxTMsur6/X
mVx8417U69wWooTjvCwuJdhGi0rqrIdx/wKUwRPUSio5f/FjFX5vqw/K+fP9XmV99OMvpithbjM8
5Sxd5OrVjA1XiQrb2Sg/tBQBOVO8d1pQ2wOAB5PJFxs1PxuucoCA+HN7+7gI/QVMxmx3UH/gvKaf
EsQLw2Ew0WtW2Krc5DPv3Eia7UTyDrP02ib/IIqc8csjiWz+jcEAuBXSQ22steCIKiduv3PYcUrZ
7GYk1Q6wLP4oiWn4+nIdq6AImMTCd/JURD0iK5qREBkYf4g2jACefnjdurkZAq3Bc6uGG7/bkaQJ
h6m0zHwAoK1N+5inNXuNH62H6eHPi3xS2tS3qMPZqA/p6f+vmsCIFgT9M4UYTyFtbY5654qg97+K
CA2EOY79cuxfCDn1hp2vaKv1KR6/HFD8IS9hD9QDzTjV45tzJF98G4GDGQywyx8Wt6S+2RqZEUcd
AUXlPno08fL5DvbqcLWilF+5N3cEaN8JIiF+KdapkQTAbiBrvbypvvH79ca3eMAhASPhS8jDHkkj
NvJNYsE4cHGXgNg+Dd590S4wUiGqTqjYQyrW0zuL00DEEibJfNcg74KcUisz6icT+5VnFoHg+nN1
Su7M+M712ohT5OYGEujHRymQqnaEQdLlOXILK0Hxb5TbXL5ofsiLuvHaVkSjtsZ/YJLU9bz45FcK
vBYHualBq24ujRISX/0I2p13Xtp+IPqXlAsDXnJ9rHd/EkR6Wpd0WOVppgg/5XVsJaKFoUxpO+9j
R1VtumOPq0oNkMXGa1Y8yQ5L3y1bQwsgMTLhBFsZvaNFW0P+ou0HdaMLX3aQpqTTj3u3vOtCBGNW
U/Bjw7iTg8L8rBq60elLJWljZl99nLDUJEq9Jw4BnFU4zMt0FvPaHp9nkC5N95JSGxgbC396d7dT
fNFRX3vP5E/wMrydU5ZGDxgk7hKrv7oPuxZjNYP9cGGZ7yVXlMysxaiacPTfgtnhUIIsyhk1zpVB
pHGn9kSPg+LLbBV/jQE0KDIpX7G+aHPY5HIzjrQGZ9tjc1CnKpbBY6Y8YkaYHKXb26I9TNg0Asnr
zdDQDN0NqSPxMFdtUd8vF6USjeJhnjz2Lf1dZNPJ9w1yumn2wPbPggGIpk0628LXuRq/imEZbtyR
Rm0nzVyJMrGox0aWOsHEGrLSWSKQBwcMGqEVOz+FBVAEU63qdGYfFBuENn4lv1T+3zAVMykTwcej
nAwRotwMDMV5sg+8BhFCxPYN65vwbT00JzNSZdWUSIwY81JjgfR+m36KL1r1nqYSE75qAPof9NuW
B3UGipXeFq5lW0R4Baksc6wTfTlM9eu/Yzmv2PDQaCzlzZcEYN94gRei9HXRop6kNIpKPhpFXcOj
hJT06HvNjjh2tiCl6dMEW0s5/IDJT/oSn4AY9o5nJB+Pl2dKGSJL2JAUaGqsnFjph7GlEHNWMDkg
1QfcS+g1JEY04SgKYlcofhHzqaT9tD3h1r6NlxXlXRgNqG+NUJx8/S686sPpjRi8DH/dDd/7qxjg
fORJ9KmyewAHU5fcYaXZwhg2xlC09CXxwZqdQOHsc8/a0ijFGMl7gRZHVKDbplzZtg/bemMZPHgh
eGCAqHDf3ef9ObxPZQZ/TczEiWJiho+mdieQh7Xed8WL90ybPeOeGoi/csC3WHwWmKBOacWnWduV
wBZClYO1/6V2RAUjy3zBkACppihxRRWdBM1EyZ1i8oWf0YxvoBdi3nTl1uOfWS/1/YwBLHh1SGZv
S9Tc84o3R9L5bgzxmPgs/ewx2vd0CEWRHFHquZ4snEg5RgDaPGvXzPAlL0X6O/GIKxcdiCLIhyye
hA3GYjSjJRqGieEaUaOmhr1dfFDCvbt3dcg9D92SCl3839f3w3ZE3UXqpD4kmxIEIG71zBwP5RvV
/EItMYCmTWirB9gajDOXpO/YjhpmeYbwAKLmHoFlXd74Q8+bJ18gkYWsjHBNgA/Takx95INxsRmY
aGbJ29kD1nc9ao4Zy9ecQY1yZMc5uw6xbQIgPRWob2hNjjDSyJ78TbO93IeJsu9UL1KTYMMU8yf+
GywuxRud0Kcmiid0HiqB+q5jDiZ4nxOXRvUHD5BSk2FImD6UTW2ob4IF6u+5zepSa6OpP6ny/HHX
LQwodG6LMTBiJPKqBpDFfES/zeodSpA8tJ2dT5GmwurZKluyeYRq1Wsgbrg+Ck1Vr4jPVrMMhijK
RVa8uWhyMm6Q0OtX/D9Sp8F3PNWSLS56PzYRxotDdTH7CvYPJMe5WNZIajOlKoERhHCgG7bh0ZGs
icCGw1ecmuYtfa64yo2YZxami9iOWWN4Iv9EgB03YUELBWWrwEm+MLuCh9LPz58ZiilIjQ+8JeYu
N43er6uDy8GXd571uqV2ej2Sr+mkCihAiJmWziQksu3U39VQzTMUGpPl24GclgUiSC/P/AYeI/1n
hDxkcey82mh2+e+AgW0Gel5n7UABZ2uTi79M7CZsMZ06n/ydB+2bFmpvBz84wbecx2vLUpxb6vJO
0haJy15k49ed3xWHR004fA8iuyTRGinvYekjNrjRadAd98fZeacgo0qfhApQsDWhExXz0paOv0I2
/6XrhMxwKFvLQcLjSAeqyoVsxgp6ctxWs36bJhNbQjQy4/Ku4WXzXAlOK1bz0wD5+zdPhkUyHEIX
al/YX8zCi5kGrJCYOsB+QCu7aPZ4MKoveipmon0G0IB6Io73T39LTHrbWSmLH87+F17nQ+Vrt/q3
/Ca25ZcFlN4G/KRS4zRcv1lyT7H/e9K5vh6KsY9JpPihgWd6oM2cbj5cXp8V7EbeaUQhZNputzuK
mYOZ7lA5MSqWsuhL4B0S0Fn7mokrYzNm9T8yGmq13+GMzndxIXmguUsvnpk03G89vzZ2zBfW1Ipl
CbV3q//ZXuU5JVhk4TV6BXkTZx+B10ZknqJjJifkEZ5WaCqEQaIRT0cXb3P7yggNiK+P0DO+u/qj
kj2U6dv+ackVNg3fy1f1QvnEOJ0BYyagBPpOo7imlFG7bsnH6/1AhENO4sCvV+qAWBMKc+vqTY+a
xrAaAmaKqWWFLccpBvB/5yk3GsQb5aNOgLH28PB1q5prIG7Q0EzGWcdn8mB4r8YwZGn58dS6Qgc6
GJqTYtnhN+rqz9QktJMMjM6tR0w6Uydrn0dAiAydeHLLxRCMYx6x9SKpw87QRg0D0QO3Znd+AvEa
X+uFsS+eFfCTLd/YkwkvuWlY8zApTQFMlFh5QID8dnYjf7jr9pPSaJxy8+3EPGjy9nf/ur4MdOtl
j2Dk0ZDVdXvlkaDyxOHXv0g8lEy6Lf+8gF2vejVCJH8ocDhQB8Ha9OPcB7OeMmyHpYhOpk6QMoVG
5TK+10PeCsMWkBoBJ/AB70JUkCHYeOYeMy32m55W/eGmT0zYHV2tfo2vSibZUqW0KiMjPRg0FUZW
EPzSuh45UkeIcZQ9ylqDR1tuKVdSowxUq57NbG07mdrKpmAtFGWbArIOQ2JNyo3hxlWeK+EQBsCV
yMWeDSLQRunOOartSBw3PS+4H3iH4XA6I4LICe27XqLGLKOJW14oFrLTa+yXHm5cMXiXk+kAq6pb
YW+X8du1ytOYjjbTIfnDT8Fjnle/fx5KifMgiiEy/1TUJOxmiMi4CAsK7bk8XmQ3O5HKDYSvgpYe
90E64gJ3I+s8E3nYNiQd2YLVMHnJ4IDVGKUTgJ+KDiDzutp54OAsObBbrKrFsVJ+Cgoui1KQXBcN
uVYwEA6fXKSn5zdC7WxtVOgHhKHAaMOv3FtzHD6si1erxo/qslsiA3men3cMhrXzbbj7Nu92P8YZ
g89Q32US3OZfXp5AtDQFy5qWFDVY2U/R4iYT1lDIPgy7jV6WB4OkSuWtUpT7vnD6wIZTYXU/p7i9
lAtU+QEwJMKmmhfU/NDQ1mfgPu1sGb7HP/1FgEv0evmgKm3t8AOZdJhN+X5SvMm5jApI60DHtHTp
T3TYZUeXBzdP8IZSyYbPWDA5e/P3UjKaAujI84SLfgebJZs7eJMN/4IMt/et6Q9XnIaxve1NgwFH
q93UMX7nzqP359GjD45wieA8AObkoVt0JiWE26DMiFT1e5ABIRDl7xuaJ2tEQyxApC20TGOxyC9x
EUBuI79Zpt8tUHX7Y20U6bLzzXw5ad1pi5SCDru/CfGnKS13gpYUKd5MyjYIsTV/mkSWwSLkEoFd
uSkxwJYMSjD4GdeUOsRF+8rF22B8P87Ib/QhjHlOCTmJL7sWHuaAV2iobTUqcPfkG0fDEwETDh6i
DoYtwc7KHM7biaMxNBMMIajRdxI3lJ+OYW7zP5LEidf6qwdtYYYtnyrJJn6/G/CiAHejQrzG2Yzw
tvHJl4XRr5AxKl9w6LLqbBk7soAPgAntV+TUSVo/7TLkcjQxta/6ya2En81bA9ivu9YErn1a2GB+
phY/TBLrfyP1kgn8VOmfCAfGYCNDUoZ1ONoSjF3hXObLe82YjXShTa+lnaG6cFPd09rkle3mc+fz
K0SgWo/UGGh98dGqc6vt4XZQUnYH+QdRZcY/+0aCpzeStF8ARcN+DVL1fmNQuzv/JBRGc7xq08Hk
ZLyGWMVDFvkxhKw7AGkDmSWpfcMpyNsYbTyG+Arhg6xMYDQVEvFGGnKnXpfv3bqW4c3ZM9Sl0m5i
8hTLvjbKfZ0ITh3RtOBp70X0FAV0TbMLXiTGO5o9GXst63dHRvPIgRzaqp96yLg8p6Jpe6KCB82W
kASJm7e6gilbJDv3gdyB+H7kOa5IAqiGyKQmGfdoq8WTughmuLGWMmsJ3jutJsxv4UCLi2LF7/A0
3nXlrMk2hHwl6VOrJUpBi0RCzehTQH+ujJbdFqP4CwUYsB4QAjkthfQ9InB9EnM58YXQFPno7xBI
40itSTABiJntE1ZtBHFM96T8zfmA6VH866oUpeFIRkNxIQ4HzvuLa+fAMxfcMY63VgLkW2tciiar
b49jHaS17RjL+oss872iWcfrAIG6X2LnRrW4uBYLrecZtSTh3ivKuU0ccTQRY7r7dW2SSV24/KN2
eZ0y4W0T6urnfYSRhRaTquN0BWjVdoOTzuzgu6MOxxsa7AGSTnFlMxvProDyIYIx141GYRQgja6w
Zl2qC443lCj1Gg0Vl0GJyCStvxzj2c89uDmMHHy5k6QQC+/scN4A6s7hwtZlCVcAzIvvfmaCQ/GT
i49NiuPy+YRf2/fZh1awDhvih9efAIjUvz9ivKhAJIBPJyy3rLqRnUq5BO6qJjbYNFLMJw6N/uiT
ZzNCCL9WJ5sZ996k/IYz0X+DuUx5rh3gu+YffekI63G5kQhL/0XCTeFb9FDO53h2QyJdMzvXHy/K
Rjvj2ofMaFEETpQJhBye7dM0Gs9CaONZvqTosTPrTCESVwcLfW3o7Le+JOjyCH7TXOyizBeEKJgg
vmeyjmk/e454wZAptY4UNr2R6DNVXooQarzZGo5SMUfrUXFYpQXdjMQeUwtevOupfIDK9w/nGeCg
FQiUuQmCprBhxAmkeDz6uKjwDIGsQQw/VmSOZAQnrbR/nOyzKLamTpXqKE0MKF44HNzsEviCuJ1R
EfJCsZwuh816MVlYHYqvj6CjvAo9vXtJf0K7//xTNhVL/YF2ejGHI2RNHvL5hz29YpbuWMQ5mExu
uyMHMBJM/SGllgTevSboyF7IqMX+stmgcoH7igHGgYaovB9XgMHThjL50qng/gLQo0llZiV7LkMU
FOZNGFT7lhsYpEDI9JhvRZPU37TD5uIhxfVOKMsF0MPTR7GroqOBwNGi/D/fWFPPILhuZ5zG6zd2
T4cXJSwViBH0i2RbKHSK/hST+R9gzfo3xGBE22hVIqksIgQlNTYElc3hUlZ/WTTr13w39eyr518X
XabFEsQOcrFQTHXBqcWA2zW0SLeGvIRd91wpyLw44SfGo7ashi5k3PCH3i409mL8FKvMTgy6L82+
rxIw6WHJPvUyJp/QNqz+GHEFa8Y/+Y2rswvWKneHeI+ndgRIFUhK1vglOO5nANu5824yQcr2IpXP
AtZTFRv3/iY6+Vs6+lEPylZryhLWXrSq2P+X07Cu2OeWV3Ikos41IDLKatYR7bUr+oCtY5ASBuPW
8bNkxUrjz/JNcWXG9cHRQe6xJ4FEjAQgNZ5cy7aV4Cdogrm4soKkZY6gAAFxrbqndlRH9qJvnoMS
h8lCM8xOoHGuO40gL43IPxw2TMmSn8+8aWdoyfqAaDoeggip8qIv7DkiCYK9QD8PJvel85lcI4PY
6zGtoMAnfSpL1NfNr7d1syPWIKoTW086NI/iHDgQvaWlQExF18Rxlw6YgWkXtSDL8S35x5am381s
UgaXadoGP8fEzlFyGDDaxlBO5WcdPOepEOoWx6xR9g/iTFhsPs4MET++vDVLtHWGUQbs94pwWk5w
Ml9X0Onw4n5zvaf218oaVQPV9YhiIXbtiJcONXgGl9YKBgV8+fiCYqEhD1LUNmRZHy88CQFLVAjC
7vcJGhkcGt+rnOau+xu/zRzBI4RC18Wb8EjU8d8lNezTd4y6FGPU1rz7zYTwaydRKXqO7t6mhBGX
1Io8V15XC0Pg6jWgilM71ZTPqNB0BAK3V6+5mJBtNEFt2H00sOynXlNmm97/gL/OHcuN7KF2xyQC
wh8EcMApK1LaWwPVYLkyMy3F0u7xvUfyuLsR5Yyes1cqCE03dkdRPzCanvQypqXQAkSXRxJZk8t6
QFViCnE/vZ9BBHuLv3mamAQ/SeJkSOWnkd7P1+DVmmaSMvcwXclooYYz6JWQxTtAZMb5JGbG9FZP
ahtlv2jFafNDddpkZlmIanLo5nAiBbWHyXHS1ZLKy9uah174CfMw0zXezzSbdYgbmt185kJRy4AF
Z7P/ZJmPXmp8CKd/ZuPOtuaCmCUxgp1VLfKs3IJcpLFhvXLzW1BOXrawnOaJi1okcX6ClQws+heK
lZG9FWaRQwL+L4D4Lx0UgmApWRXr1AgcSaYVyRshdMABy3GBeGF2Pgm1V2qx7JaXgt9ol2mx08AB
QWpmiXCsaLo+ZmNKZj/iNGiJkqG63YCfF5im+iRSRyJJaekBThonUM4ojXQd7Uqsw96otEu7PMXs
cuCKHwGkWLZuMJydVi465HxobyeFywCX0NVKilug5z27cuIxVKrHkT0+tHlwYizSB3MVz4kj3WEQ
uHgA3cVJa2na0zMPq6bH6jufjv4pv8il9GnHPLHkInFRvXcEIJTPtXUODV6GdWLktsV+EBPzTEqt
3Af6PCWL5PaCd6wdMLcZeXs0pazQXBN5j3ic9QqhDnLRe7YkG3+/hOtOP8YNDc7z+HeZ9+rcUVuL
2I4W/E3MxdtDRmhmVplL54Mgc/sV6OR2pnDFen1JQ+yGcS40t3aZU8R5L666EZyZJlwf41Ni9w/n
6y+8IBwkxy/BaPflR09+sNoVksA3aXDWIVpEYaxNNsFYqC+2zkqn7+8qUXz3dStrUl+oYZH/xTgN
5nCzQSJlhTPC5ZdoB7dxMQfOHAb6ZMWR03vbmZnAqWjbUSAIfivF8vP70N4uC3TC7rHw9cDerNre
gYcuu54uw/is+mULQ38I1rkWT6I+3P5lh+GVrxfNBnutgGTiQqoD/06/bfyXZ7IfSe8BACD6Jfpc
5KedxXyo14YXcZVAj32BoK6raEQDH1x7R2UnSbNfLImONTOwPY7lT2v2S7lsnp+1L8B1FSddmoJ/
fR3qfi+yTXhf1hj63BCiIruPqme+Ugkwr5oGwfdkTJL2Yku5oX2wJ7VjeCCsvkHd6hbLH4jjX+3e
aotomk7WWbByCgLRygtTiUSQLPsL3x3H9nbd8bT6Uf6i+w16QKqvdCP2Wa/0qVhJ0pBTYL53eQ/7
ph/wHLIclga8dRrRbgO/KRD8Mv4Yv9I+hwUTWhF7P6PFU/1GvehdAX4NwBSeG9mPhL+J9FmFsuZr
w3Nn85QkmA1unKbLoJ2V5nCrzu+pbaglSUmxQJaNivdg6B5vG8bHty7WWxPVpKQbBzX5I4t/gmil
JicUMLaeu/7Fm8ry6rkBZmz9PV2n9565/XOIXQLmLzQJ90FINuMYyqIwRRmn0B7v5PGatNML1XwF
dhlAwiQhQ9RJZDGAWwnk2xIbxL3BSiF8dxsIty33XpBWRxQY+KrSqPHi55byhSB4nkG0dIYFRBKq
9ovWnbsuKG9hgLugn/EO7js5mos6lRRrD0/OyY6/KwFtZxiB2zU7DJ+pGpmOA3nZpQVc23pKqGr6
JZkEoo/WRM+WjYsSzJ1Wad/mLOs/QI90O8lTVQI6r1iBZMkS+3xIpop2ajGWuLZrSV7BVwb6/D/G
lREK8Cl0x1oqxJjN+cLsGMEGO6P6LPDx2t12pWnHmEFlg/T0+SbSXC2vk5epnXQ4AIWWE/dWETdK
qfbNBclFl3yEqbnpGJO/KnsyXMA8KQvpKzJ7INwzAD0w6/Nxq7hDi2H0+dSkfhT1V3cha9Wco2WM
Jnu31bxnPy3pCuRCAKx2RJ+kxgmJtYFs9RlwLWsayU3PSdCa4+qUImzoqRPnVXWZYTaoLsF2MmqM
xm4hExd4A4XnAZuZ3pgMghTE0WSApM5x6TxjrcATLNCGuGGvmjRUD+K3lrBLCw0J9UHx4mbAnWBP
6vrJZp+h0k0PlIqx1K9uJ9ih/FrhP4i5ZUYY0i2203Rmxavx2zO1UB+7ef2BBe5TxVCXU0p2NQmi
BfR4chfg1fLWSUJ66GpITEH7JzHmy7aAze+ZSPIDjTxD9fDn2lS9+W1zVF7GozjWBxAkRBm/RoHC
h7XUdQTRldRZLySaMyr3ZFuX+DqDLeJHWmavUbwvkwmqZ79KfJ00M/4uvbqwEfj570VI1/5qpoQ2
0Y3o8ijmU6CBTXQR+dfhJuEraH+r71k3VzJS/PoPTtgsdt+TtaeYrCE+6CRb7q6xQ+AdkCvy1J6z
CDmP7oxCzndRJPkkzXgW1W3bLJjxzyjLId7+Dc3gujqYPv40UnmBch8wV4tBeCyKNSMXXvG/ubty
AYK6OcozLPkWzMAYg3HdFRFXIyQrtYBjHB5XyX2RIAbnxA5HRXidkTfSSNa9sAZ57E44DrRPWjbU
Il8TJeqZSzj5x/wEvl4sUe/7VZYFZkkz5Lv4hmk99LUlCwJtYtNiVHQDBQDGNV0g9ozFqL6mU7hr
I5ncGj2V9oRuzlW0Wgnqr/nmRdfzlYjJLH9W4sFMphrCrON8jhCrK/qTXuhZhFrVZOLzmAgVq+eu
ah4dHzVer2JrZVBdXZ16eDrlszi+evayZHk4DX1HVFk62JqzeQKKKFUsBTfkXyIhHaYoATCQSBHg
jL9L3t5IpaWOKDEViqm/MJlGyejIUCesF2h4KdrGP9ZzKMswlRUSDr32Dg1O9mB9/9ufMPqRI1xC
ggHEpHcd0ArWyYLRlSbj8oyPDesoha7zwaVoEXBhA8+ofQCCIKNafQcoc7N772Nh01xNRrSMrFqm
UEyA/2Rh9zXJayY2p70+DxYbkDil/B39dndJ9IEu0MbXKNpbkuJcEZ6NIjVdmKBLNnBTLv+F2mYM
X0AN7lpb4uzm4JwrVCgR2UlmCKI+iJZOSwAzjIjht5iSg7QmQRcXIlHjoov4mRJKggKWpKHjtsFl
lPO0aF2UO9G9cC2D7ov0UlfWG5udbL+PFVTlXrscZ5XeW0jW1//oqa6amInRVguKC4PBfiw5KXIV
4H8mXukV3jBfwofIsO2QzO4HOFAsnkDWQoYGc74FS2U75GV14KclmyKsH6zxGiEzX4auRoH6GpxE
8xuggi9XQsZ83U5ZzPnI59EzHYzNonAoiLLiZ0GlafvYIPTv7q0dJdIWNGWwgyc4QvYDV02pomDP
T3PALmC65JIjN37YoNekX05dzK2bs1kD6Yv6i73XAOKHxhbSX9SiRV95THxx9ObL6gAm7UvV6UEs
mdyVwxTkZoavDIWK/dpncv31p903wRnRGWXwdha0KbALYYUi606u8Z9gb5t3QdA04qDz3u9jQ1MQ
lQsiYnlTTtrSy0XaJln4WFpchpfBBpP6+iROoacf1/XzeprI3oTgvExQI5AyLUkv9pzf7LA63e5g
WO97QGNbuHMZmgXdJVIJ1IzVd2Hj+enpr1l+73dZsNpU5WnKaK4wwSnSAvH3QLGmk/uVCS1dGHoe
ktVFkOTJJtyP6m2So5thFOuyLNLS8R6UbzuEca6tXSIxUXbfxckQ6pUZDv6dBUDZaRHnxko3mMsM
F0vRW54Q+SzNOkAL3tdbbr6+ABhV9tIBwXEbK+EWYwN9ARkPbnj4bcD9fwDdgCwAOVdDjQHhAxlf
FEYR08r6XqzI78toxcrC0koA4W1QmUHJZUvKBf7kehtdE28AkluA2H9Le1NcHIU9dU2kgyZh9WRk
qxFBM6yqNp/3M9gep/NXD4TWfPOm9SgIPnfyxrUt+usAsAoioCcxUBmGNrdu/acBu3f1oSLbImkd
qNjbk13zODOgigYlByNgIJZKkWwGeT/Li+xq/Y0xw8BSqutvpgIycBYSzgaX9utJC6z5sgAqSLgr
27oRgbp7Vvxt9WdRGdyGjL8Cie/GDjXjHSWVUwrwjLUKQAjal7QzGrrJLd8gxrQ9hUfx9korBzoP
1J4nLVaq+pRMlT2tq5Wpu+UlXWn5EvCzrr88q6RqVlCx+4R2tCFZV6Co0jmUoP6fmtqm3/x3rVAD
AET4r5eOjKPPVPNQSIh65R2rv2zoZa/MjxRlwCDIGfoIdz2TrqOTbSNw2eHO6e0czsiYy+ZUw+No
uPr+OtHqjq33B+qhfFdql+TJ54dhpTV7DMGBdwf/hdCMzu+8zKow5+UdpK30B4uTHZMf2NaAKA2O
z0GI0JFaKhcL5lUp/APB2GJ54jmfzKolOS9ap17IpUaM+zArTdbQ/EibwfhcnPY7UkTY53r+OALI
RZ1bOGPygcge24ZZwU9rdmMzXastQGLwLEQ0eqEzcKa6eNEryjnKrVoIDJjlUkePPs+c9P5mOXC2
LHNXHNWeaLIC3IP1O71h1hhSdaDACVTxqKKlVJPlOwBpsswxfNDIsXaf5hLgdvR53Aa+8HTeILPH
CamID7usm4tbRHFzicEu6QgbrxuZZONVuFpJRh5rIQ5i3unEofS/kDj4xI3DkeT3gwlyOd5B5mAk
xY8zsLzhNo5e+ioKAs9Ne0ngVzSbwd84aTmNTbrcackNBTrczH38qMEP7gsxwV7g+O8GYYkRwzKW
/1h1qLPzn/pRv9kJ/SEc0jE2i+AcYGh5s9BEKlS0jnYMw79OeC3XTEqgSGtGRuWxyGKyeUWGvIJK
LsH9NEp1s8yJ1FQmRKK9q200zSB3fezyj7UbAOlSP7X9y9Ac4UdRiuNRXyjBz5sAy4WliMGNPmYo
KMJqevolLc7KlIUpViiiQP52W6tiVEuzBkLq+Hg7l+jjmUltIjZhBpuS0Ncdrmvla4Mj/kS+c208
nud9Rd0FUzu32kKnHGlXfW4h9IJUtLZfxl8c7Op1tMG97TA2MP+u0e0rSv2ezzEFT7KeOmaS53SB
6lDJzpx+idfw4M/soDlxj3iWmKq1KBlyHO2iNNoSczMXPlx0MVkckNuZr+/HRIfpzGY2GGC9Wh8n
Jps8Pkm1VF8JrOk4HRD/JeXKRaNhYCf7Y6c9iTsOAI3fojWkGVdCEafkvHD/E4hpqoVb/y4p4Rqd
yCu23kH+fZAvk6rVgDIoIT6DeDfUJLJgVD4+zmBBzkBZJg2atK0NXw9oXbnvUpuHIVee1QBmRWYL
MZkajHiZ6/KAiovqIsIFEfOefbAMA5c999wwty7dOL5norS+ZGBOjMwO8KWjkdarKVAJx/vLPKyK
zT551wNunUHiMBEiQ54pHSh9Xcr3R0OXUw2OCVA4b+FkCRlzgXECCbhzTcwDKRa8y9nsUtLgPYBF
hdu7naRw/Kx41DsNxFzoXU/0ZWtAFRO5HuIaUj33fShQupC8JikohZQ+q0Ix+OFnLkccbgvBaqjN
S6/3HLywVUMgCST3DhAAAdKr6uKDxzPoTB1QHSI3XQrLOayxu7MaHZMLMcCk/edyNJjNCxlfyhqN
cPD+81YN/oy41A9g/U9il8EjbIChlWZcNvORcq4nU26HxjZtOPd6HYiEe2oWFMVoAvhnsDHSqH87
PjdhDf+U4zIjxLG4Zjiq9+XGIIoQlWQYmit6UXC7nNhGw/Oa5CpvfIufV1i8GyjVxWS6bQb0Yqru
0zOdhQyOwzcj2VdgDyyXtc4CqSYfBQ9FpIQu3WHXLYVhXxtQbJntCjEnRpQSIJBwpOSWAgoWLAif
9uWXPzyM4uWpXE3MysZT0XFQ6T9EMQpHjLe8+nszfL8IT3w3sa4aVWyQAkGmq+VqQtLbYNVgfUCn
lTUKy8TdTkdP/sISkb8cCN1zFJV0X4yYGUy5n7nnkKOHPzQcKpmmsbiayCgrQOAjzxlGvMhDBZ/m
Yd4eNpIZPnhpwmsJiIqReFRpoQrl3TuF+Fad5ceQRBg5v0GkCiXRHdnc6tBvl2DWbiY3svAvKHVX
x+SmVBFrG3K4saoUdTzEMGl5JIC0KgTYsVyKpNE4Es+B4JG5RQEPGOyr+7CGkhzaLxLtC1WIoP74
cBhk2uVmenmEH8zWVouMrqj6sy28l5+OqJ4qyLdu2TZNBungOlCswtA2zGVWpqETSTuoeExvlxh/
rs0sU+7BTAzNd9MJ/fTUo1mrS0FVvebkumHCAkyQlabJgyk7we/lOANw26PUG5llOjHFwTRp1ERo
i5/svb1REC/bZposoVQ3bGAlsi4ceNiOmE2larR8Li37Yu4YztzbtedoiYj3az3hnwDEcwnR5VAr
WCKeYAy6oom0BX4alaK7jhpGNPptPyHD0uO9NUmwCh6Bch93KdO0PJyI5RLw6Q7Ogwf39vaFK20D
OAQvbKn9/urmEHnv6JHnxxhlhomct9jKusAcWTF5qdVmEQ3iJK5DmT30H/vNq0xZfjPXb5OZFe5n
ImMOCve57kVPtn3fEyBKUO5b+uBD3xNzxePTyPTKu3mXBPfad0Dih1ebifXGsaseE63OPazZpRya
9tgeVEpe1UJUKNkUGOdnXKYRvSDZIlWoP27BdEN3UG+tpGOphtjJFh60gZwxlaa9ez1x2Y/b28fV
j+lBnMfYOf1Lz5lHyk1dqw+/n+LXBYtkgrHCH39Lf/vgoreHm7uiwK3I9pCsO1mXzaujecDzqy8N
L8mJ1hf9qiBWeVODy5usyeIl9+NFIhQZ+RDyYHiLChgert2pihmU5Hlc4HpoHAvUkIahTVVcFZRx
d/dQM5Kkj3uUGYD6HYyZHgDoE2BbrukrKujg39gmCdWaXHFDXc6VctTs7K/HLkjOL8Xj5yvKKJKE
Wx7X5oIvBzXu2LrjwXHeccLfW3TZn1m3W6mi9i1N+BdQlnnJI0n2byRPmhhQh4x90hDOb1H67nrc
NUMtJcWVwQusWYnad5DBTOON7Wpu9W219CvGTvoINBXmY1eDM3UimI0LGyEhQd+uRCrRL3j/DbnJ
RrybcV7VuMwF1gotQC5DowxCakfPS16BCJUY0zLdVFBKYtivW8Q0uYb1zhk+GYkHtAmMnVuEh8jL
ofh9rEGQ3xeCQ4eQ4dK333NTNPMNFYEciI868zKJ/T8LOibh49P0qw0kwJb8dlfAVwohxd1ZJ5Rd
tmE4LZtAy/oDLimwxU3IpIEHUS94woFpjWpD2M9JBT57rYTVuJvF3hC1lffIY9QqErP1OGfEOfhm
v8N7rSTahOzgfo+ZWCzkWf6VyL9Cf20lWYSOnyOhfAN2vVvgNfNbJzhXnU5+wT+Tp/H7ChxOXPob
9UxdTYCE3eiGCopj3ficY5yDBA6DYTbxLGkEYGUoEEd1f1WHGnmgGnZLEoH8thL0qJjauqjajIBX
zph+Z/HskbBVJDRZLSVJSFORVhyS8l/k7/ZW6VKg2PWJtRnEia2Ldif/x3bTEXEZb+/f+Z4c9KnX
qG93x4Yl7+39og/84pJQuHAy0aPR/Q3qb3ykCREE5US3Z0dXsjk+gsK3C1ROR/86VhaolOWvyj98
0frFTMNtfdqmIFFd3pwCnbCtzpOK/L87bivBZ6MrPgQcoBtwnhjR/t0NKTmJ5dJMDqXq89OzLS5j
b07/TQk2D7hyftV4IPJrExx1X3aNR+sGRExkcjJyhjq2O1ZuKxMSiyo8S3WQiIo+VIzWktAUDWPj
qpjvdfwiWmjvf2ThPy1C4sLqSw3C7OF3eDWcfwc/SKROKeb1cC7tHRW+xQand9BW0xi3K+VynOtU
X6WRnnI9fciOHpjrt2PosWk3AfaiinYTtyFUGPWXLdKWHBMeEg0f+ZjxzNhxucXor8J4AZYsqxFE
T0aZJOvwbzRXoBQwW6r5eN48k4sEfP4XI3LyUajGIYmS+YxJunDke25ActGXJNUMY+xDMHZyhdET
TtPnjtxFV2V7iDBQUna7fw3ocmNKFNwzuFDqxEF5AgZ9F6B3xQG2l73xy+owHdqJhLBdRQ6OMUIQ
Zcin4ymTnYQVycyzxoWiZLmGspvc/JFF64HXgzxWcCdte7gAO8mTJD2ipoWPYq/RgOBFid5PpgDy
n0o7+vX/pfO4AQAWc78hCZqwhVn2LuAOSJklZROV1Jh5Qoic1P3I4JxUBiMVXghK+djEDMS6xawF
UXdDKkQgvXbtaRilza1ppDZbgd5Garpff9u04bUi6c3YYu8JpibKlv4c64lZXUIzC5WNpeU6rxAq
a6TRrQp1C1OjTP/0GNMIaEZjCuEROnS85mGeMPFmD80tt+/zXM7OBYk4WCCj8xTnMfu1RkmG6Hyi
LkntEKhbSfHxULUFwR24o0B1ouj4JtAL0Jq5yz+mBAa6fIqoG1k+2RCyw7apa3gxLBXO+tuDH00B
Ms66WgbcSpIGu4ykOUTu8fQl3DHTy8Xj8AkNNJ824dLborp5PPVq7LhL5i4wJIyY/SYsLYKEDFu4
tvg5KW1bp1at2b9KIwdQ3vRIvNwK7SE9ob+gGrzbmzZFjjjlAFLt3kPkU/Qd/jGZfgOtHoE5dwEJ
+GHY2EaHmXRCdXMYiyWdAtgCPwizamzoxp3wCTJ/hIG7qoT/dSY09A5W9Zocdxp4pcdeb8/4tq4p
ExFJshshH45WerLqQmgVcRTXBXqGLrxhr5JvbLy+0U9ufuwnKO7rrVPHx299CuuuetLlhgMD7UBJ
twOCzzZt4pti+i9yjOw5lpR0fUZWiw/eEAaqGee66PuweyxAyQPThHLsxbAkjw7fXZuXplyCr0NH
p6d0mfijgpSBwOEPrXPp+6kf3zvD0X+3SKk3qBTZkm3h5CEiBlKJpFhm+Q5v5P7vgMSghYuHJyfb
bCEHRA+2y+4BQKsp3YRNTEcVo1bzHsz1ugqWb46zSZLYuwAyOFgYBcvvYFloZ/Ln0UzKZuJjrW1G
yxShBjOJW8vH8jqtq13Oidt3EvBXa/Oe3n1fMswykjsDshTFU7+qYkExStcIgXi8QWN7NBH+F4jB
FhkPGDizMZ18eAhWVHrsuk77Pn//WJ+0j/6fUbjBC4dAwMYUevl6s179ag0RzWvwUzCM0XuMgFgr
7t1ZgKFFJ6tqf+mzrdU7ijJ4uDK1/07wdxGULLV17swMe61UyU8s8RSVfENi0KsjPGGXt31v41wV
gXpkibDiUtoVHYmTZ8XO/6HPcwklFGk+cf0Mk83cTVV/Su6JESGtwg94qfh/939rRqGWYPZ2OeBX
4VDXxZ2k99cq1YhGE+b8FIPCWbUHeW1YICtulIQ7bqP6d6KXdELJuxjbgCf23pF9Etj+R4pSW/ua
1IO54pYtHGMuilFhysIjk5b3YDnuovdKqMbokNquFkHZXDHE8JfsddZgg6NEXDYK7hF7H4C1Ehsu
ZIEBf10TXXA+A4qCmBGBPYdmESpaBlQzp8w3gmPkNhMc2u2eOFrncWzWIfmze0IAJQZPBcCv6Q8O
tTQr4EjbBZxp9cJQq5pJqyI8D5tQG6hRYwyvvoFpLDGh1WYLhxdJlcAwg3cUZ3Xz3MhPi16/ycFG
Wl8l4vDaHZWWVcnfV6WtmqHzZUD2lDGx+hebv91cXY4gopOzTX0ChfVcn8U1HrRtE17Oojg312QL
7NDod7d6qXRVfOyFNh0WAHbCDIAhuBrQcnlfxLyqfmeWIblGD62rc7IUzOTNWXtepyuPydaQv4h3
iySjfjFwJJkGJXvsl2nEuICi4Yp/IqRXlyv3Hr6AQdslJ+MLZVn0SSdlnfs/6MzzLnPautJZaL9D
KxFM8pyl+yOfsvobTBt4gc48uanNYBdXAOfAhw/5LvVdzp65O62dWWhzi27nw2cbiZ5UQY4Y17Qv
K18cy6eXKWUSY50eQNPXvxtqAg+nW0sPatbn1/b1E4uIowCX0VKWNma00EWg19t+uOiOl2BbWJ2K
jddIi3W2qFHt3WJhUqTjz/qQ1wCFaV4NVmJjKrwG5X5AMP2qcZz3hIUwSHT1UMAKIIrPX/xDY//c
MrUHFlmNY1j/NMQWXYpa4dycrAQWSgp9M7d2KvcY6CZn58hkST7gqdO4cBCVWFka/IYwO4+evT8M
ShvLFYwXDELYY+9L2HJEfO24GdgmfJXTx5O3+r96nAZ6XwkxieVTKOVv7eOGDag0IbmzqhePHw1+
hKGSJX17umBIDgt7Nw8SZWjBWMHpG1d2cXZi0f3/91yPRDF5dpmRqpq4R2wcVcBBYy6J/VBtvZCl
9AueKR87NwEW0NNPM1KK99EPzc98j9uc3KNTzXmM7GnylXQECAuvupqKyjRYeIrXIQXXRAqfKq2g
DQzTaGl1v1E4RCpIdAvHNfZwZDZPVwBAZRvWE3Ey5j7JWsfnC7vHabOX+XTdo33Y0wY7qMUbuLct
DtUll1oIRAX3AXXmwrI8TEoUgFMCYxdh2cG3ycZVLkYeUq7/BycGzjJPoaFUz3RFvP3EkSwd+KJn
b9mBx7fyra4XOwo9rEr30HrTnjcJdhKxf1l33Qd5AqVdQS0Y5wGoiqzxnQBatveQXq6qtc2S/iBn
o3mBAtbdOv+PJY/RcT0YI+8NKezoReE/kB53KUwUg2qiunEZT6Zxikw3L+7DB8opXAywZRUC5Lm1
hmvKtlie99DGPYH6NbwetQ0EHfu3XZZUDTRtiScjF7SinwK+UJRaQAsK9xGF4cfsuovCBEG+2I7Q
kwZ/vC5HfOE5aOpT9n7JCgSRhUc22gcFn3WF+yp/e22sIJixBiEJbvGhWkxiTTbLE+W5RECV0vpY
+0QZfh0Uv1G5yZ9U0UASlT0TUTzkTJ/KIk9tRQ+kyqilQTL+25iFNy12wXcr88C+CoygtQ+kU36G
RPdFswnT3I90lJAvEMMdLxbmTzcgrXNdqy+KjL7hrp/Wx+zATRm6ZBGPCvwmyKDcYWXAImL0v8rW
LVzFRFpn53/wEJVyPYC3JH0lsiDoyNZuLgco+OwiadXGwPjut9wCMyiGsuTHyvMegx8XBMvA4KaX
jsexBPu0LNY0YYwTWs+SezqPFykiUhiVZVRN8GDvSgPN1U02zB6jdAFF6Y4jJahi24ClmXN2M5HH
6+V1wl8lrTixttNLT3PXb/1C4QgSa/1KJls14+OkAo11/s/crpyGi3EuYLuZVeBtFn4xDzx9N345
5Uq6t8pyr0iOf0ATK99Tvsl61kmhILK/DsGrurcpAFq19Gt5rJVx5zKcGzlw09AzT2mr7AU8tddR
X9hbveppusns20VL/2W95vBBwY8j+ixfTRxZAXzhWeGaa1pM32hx3TLSlHXlnMWUfqNVfBK33QWx
iUSx9puSiwFyuVABcgc6m06i0mdiryoK4y8cGKwAXZFD7G/J8ZcYyVDOU5W9yYRS1qOYI1Ms5zlq
2uWgtmmGO7/tb7GTwisaj2DSyQFRD4+jWWmwrWZneprY9Ipj+3I0LQxr39LxHNwzH6q+J45IVbcf
hKgAvnx95+nDUXHbAnLGdPX5cz9rkQJcj3bJ7GKh89a66huhYK55TsLztLpzFFOUHxUsYBbSPiuJ
nyHi5lB7gyZBhuncvnNnU/EjnbiNbLWWqp7Wer/c+ZBTeVV/PbFoYRcU515GslcYSNgejcJV0MV4
myhNGG+dA44v8tn9LJomfIJ0hKl67NXg6VYBt9/WMwlhwE0AWJ5v21aEkTz9H3WESw7JIcud9NNe
lc9cp5Wg5/Ok9ky6Jx4tF817IJFtN9vpdhhDjx3IFchWCXYkMH8jadJ7G+nBbFMqJ7OwMU61tclO
dB0IZOAa1k3bMGZVnhIBOfQmq1Bk49v8+AXvzUXK7bKdZqwjiXYXhBLWYQTWl5vQNwv5Tj35lftA
xcKValEiuD+sD2bOaWhcfGaaFUtWeJ3lw7G9YZ6cOWch9n08oAxSvxqxmirpt6TV5yT3f6F8ee6K
Ma4wZuUdvpYHrc1KiR2e6CGkKJX9KiZufQ8fABejvP0QLASd4FLFT6wlZjI14Xs5JQtas4nWRZSO
tzw2sMsZeHMkj5cjcfmUG1oVIwcGEoOZl1/MGrB1GiGCCsnaie6/cNyoArNDAws7+N3JFhYcVRFp
fmJcX8ATyTno7awFdKw9LVK9irj7x3Q+KfG+NfK6lwpsU346VgXmGqxbmdA+9JdOc+5R5FwYZUmC
6GSsclKGBkZsYUxd6CVhtg7GQBIDqcZhXU0jYRVuNYbjLCnYpOpFh7jJBAoUKmpCcq5bma1IGx7K
oRWSnCIXqUjlCPrDk3cy4Ekid1OjixUmKBylPyrlLo7ywsaYspjMhU5TQwIwuz8L3O2rTu1SuwgQ
tO0c27mNXArRnD2ygWE8iLWtFPhfPAHpCw1bixFTBQrOf230XZav+zomfP+K3+yuq04CgcaTIIUw
7twqROlSB3QLfJ2wqVm2B4ViyoR/tfhfHv4HDZqgBK/5NMf0AaCXnVDtrfGHc2W5rJtYLlkNFun0
wzkz0NHS+fIx6kE/0Yt/kvHQgFRVnL1uMQbZGm6IvW6Z0IIOSbUX6CwNFc1P9yM4aastxjqxRRWn
fYGSTUom3VHVQfU+lWl6soGcFtaEghsAluj91OD8YtWJim8LBv9YGlfRW5NjADTJfoMMQa88qfao
3X0H4GvB+0TDVyFs12UxtUP9Y9Lk2AWV90PmkKMX55U0Afcxl+0OCfOuaI4R3+57+lEg1riWbP2W
74l5aBYFuqUH8/tnbl1pzERZV2pt5hTecTuwHLirn6cGoiom6t25K3FTsxhn0IllnUYJ7ysHxbgI
RwUt4I3YE73/3jXlOalxSySnkvsEgcX45i/ZcF3E9oCutKJcZn5k+vGklXi1Jq9dxpQ0kWjsvxOQ
0Q7M0oO87/ZZLQS6zgVnjZOsOfb//b+f7t0wQqsTqutSCX3D28i5mrzlwFM1c1OOnVP9JLSeb+mW
vE5HZBJWtrsZPwhoF4Z8H0m9P3Sd7xA012uU+V0DuAkDEARdwaV1DDVKFCRqaHHS06DcEUKFiKbG
Lp6Lgc1tOZLLGjZz7DlLvfTlr3Awx9lKo3G07gVrD+uXjiALH/DhLpm4B4digztt13y3RaGxl1eR
OElczfcxL1GGUGeDHMrL3Z6WehkkaPVqPtt6x91V271K/Ls5+n4kmgRVht0i/mIiuZ3G5NwTnHqt
PvSkX9dI9RpFm6mMJpKNyJinqJ+OxbQ9E9E5kw/XHndGiOjw58z2T9Gv5uoOkIUKh8YusktBHpR5
ic5jMxB7HR+dXiWjqApQhIew2hDHJJZxbQ3G8w3GPYAr6q0odVcJeDVRVi5RU0jiSJgmuaZqZhy0
doLAoVPzJ4P1YmLmF5EIosR/XXmAkQ+aYR9Mop17cUoYxGYM4XoJwh2BuGkBuaU4S3UYCTZgm0yO
Y5mg+Q7Km4b4PdVUZtpKQzQVGgEM7VcRxTtlVpL9/ljEDOuVyW4nvcngeonbvb1MVm6pcTpbOach
47b8pAbqDgRvkvveDu/iOIoc57emZY1y8rrkiMiR+N0+dfoX15OLvIS2F6Xy7Uvfd0ibTpS/Uc0o
6DzCCJI6ewwZ1j3MyYYqPdDYsRMMfrHhVoh8E4fxCXt9swpeZaJ0XOG24SP3yQgEOxLnm1qkTz7z
2j6qE50I/fpd9b00/FsITI7wITnLCBiAyPc4rTFxROeCR/VV3MLEgRZpydNb0zCdBWc4LYB60ugo
G3T+mjPD1y9b2qR1v4h1GiXN/4k2jlHRyUd7DMTPS6mcEUAuCFEVm9+chyomKq7C45v1fjQUntt9
Q+Q2pjtRfzhCj2RcoZRv+ZWkE2BoqUe7QsdPs/MKnCGFYBoMrHvPj+tblAYAq4Cf8RYYJMsQZbK6
MQx9GsrYu0t411sWFB7rDOrzfyKsn2ZDWAqHPeGJB8OszMajCaxnAx2m2KUA2vecTTj3xQfiUz/T
UZEn1t76+OHuDnFMR9wSvzatztG4sHufMKYaaCY/x+ZY/usqXrhVQj+W5UPjAepiMqseg53jnMAc
xKeodc0+Cmauakdh5UklY+/VWGVw1vEwkew9/qjh1ggAreibz4DP47J26cti1UXlCq8JvYUYwujQ
t2h/q3DFIV2yU4eaPfZJ6nVz+QzrT9NlDxyxC5C2t9bZh9tOT7Hph6QQbtVtI7dger+eiGlJdWhW
/cOPgk1rWOFhbMug7u9/wD0rltfOjLTsomqm4tZ5mqwP+xpVOyfNhCfUj2n+LxKYEED+9b7GRzjt
ggJ5bvYTpqNTKbClyJIsDcZYV+oWQksu6zmE79BghNKUrhegXDOA5zY+BqEQnb3vK6zOSnynWlwl
ZQHrc3JF09CohpW0Oo9e1IB1142rOEe69SConwr3rTFJT5pHxh4c05FsVimIM1fbXQlz3HNrOZgS
SfEymTl5+u0AnLQQByen2kRT9muA7Zzvbe/XqNyPqh/kMrbhuoCVFEPXpu5zmEL7+rMlzYsX2frA
3UH8R/d1M75X2lL91wwr8LHiW5Qm09bBI5BSjZtVI02Ra0L2MSgKVTr5JZ/US2MBZ9pBiZQJ65VN
wHl985mb2JtEdRoH0CiSUhL6Akmu0BVH57rlqkqDDPyNKcjlYdPbmsn0LuSKCUvI6XW37Fts+6Xk
AVfKzbHFua5BJle5Cgm+8uL01pC8/g+EPBBSVy8HP09BuA3312FiLAwV9dS9XBfxE5pxdnsvhHYD
9eO27fP8ACLsoWBZ1MjrYuxIGGpZNsyd5HBipBxnjhhu6/5wYkumVRp8vwvSwT799ecrl3KaDJ54
9KbVA+XAxYAELYgEhuOop3u3Zv4DywIwRIykR/1A7gcYVTgHx8bcuXdwJwQKCETSL1+68kwm/Eza
B1OzkMoIiht9xCdxOXNM9HBBFN/NFitmNpeYnLI1lGff280HscbP88RvYt1BjNy+S6gPo6eKYkE9
Tn+nDMT0gM72j79Cr8eGTpzq/IG1V8WCcK01+3Rm8yptF/wiX1lAAsodCMskfaF3e46LPnjWNYWJ
yByg3qY981SLQBcDatYv0vPZIZ6LzTNGRpNUwBujS5KWKNfCeI3v9H77/Ou0jeX2SIGlWI+oPC1r
n1ufjnAXbso6iuLYkNUIDVotK/3C2uhpNWIoNX7JEewu2C1ttESXAPqLHMe0dVVbwo1TGVOEL6mQ
eWCMF2p+m+3si/WcLSZrsPjjy5ZDhszZcv/xzbZCYoL4h9EzhGr452OREtMiQkeMr6s1UQvTf+4L
bTeAw9jUAc2MAtEjWkf/C95sWb2nxvapejo2UrhXuW8jBA4I4+53pG5qh3H3tlrIKDyR5DFRNvIK
Va32NtTFXpBszqA3B0yUB+yH/MeCJGmCtsucwGtqw0iC0kGBK143C9R8jbYZZYN1qZg/cz37K5+q
iUMVfkCj9Uv/k7HJccgk7JW1Y2ZtvhD7pAhgDC5PbE84JOUOdVGz2rt2VkxTTPKp0Cc7E9Euf2dT
eqVYckuzt/yWSZS2B9C+NLDrZNRLzKnMvRzVhIqowKcVTmy784dUWLEBu4Htv1XIoUSMQffDw6yA
WwQdW/X8v24JcVM2k4hbXvo+gECcKODsOmvJTKvj5nxsoqF/uJH6PXuiV1ehamqdCvBbGLSuCh0y
SSHwgqzUBn63Mj0Ngapsj3XbKmzgxPilFDDLE9iO2Fsxpbb06C1ggqyiMX1AVcxSLPltO27QnoWz
hPrZxcgJ5iL3iQesMCLwSWCQwFTj9JOICfihcIueoNGwh3gI51BaguNkWvak9MPXZdds9S/yHr1O
dOe9fgZGDSNg7Eom6Y1+E2IJaVVAYLSn8v0wZWZLvzwTDYRZiTOG7+Dbg//sSPsI9Aohogrrwe1+
xHriHIhVWHEiOfCk01Jb1JSQAGGyrNbgTH7P+VXjbSi2x9tjUVd+gnlbSdm+qoC8ZlzVwpa70rBU
iNP+IXzP8YvijS2j4RwXVMN4vNSx/CfwIt5+45tLVfDDMKW9uwocAQNpExSIsCljzXMcN6v0v14l
cqnaG070LIH9VnCSlm+7Si4Sh+37+kfWQe8U59yfmXcu1B49b17Y9biZ2mUAo4lvxTxyIlEJrYB7
8o2awaiMlpHdojvD00ReyK7aHPBrzvOV2ullADHuOcvVjYn+ZwvEmlFPAiRc1uNUz2mqCVDG1u+x
6RuSxauXnqihHv+evP3NYPcin70iZ4A2TRbi3KqJAe91Eeu4H8aXEXioX9FxIr6H532U/9PQ2AgQ
6Fn443tEGYGr1n7Vup7jdsPqDbPm9UqJpRw5Bwe/ibHwUBgk9hiq6IkWwnPfX2E5wV6vC3GC5t20
bB1Lw+Rw7QA4mrPWwLPnOBrPn3iiV2UAS1jurtGuEPHF6NolK4IjiMTQrbedJf2s/7x7NotciXJP
djqJD4YGkJG9/oKl8JLFXfiSNp2o/miXQDZuO8Q0JRz90Eq0hboLxbIxa4XzIVUiw6P/QDuEEWTk
bHGTScdycUq4GemftGNELhzw08GpQgyS/enfKVuDyZ36/zUGqRRD93K5BsIvi/uFcyTvzQ/EXbEZ
JiM1MF6NUDzM3+YnPLESOGyL+ApSaE16Tmn2OlYjnVwjTMWn/+mBrW1bx0j7/dm7jS7PeTsaZyJw
DDk7V4vLQHObt+KrCh9QpV0LZNzqZfjNzB4FxxV7x3T2Nr0Xo9s65Gb2whW8RBm3ieCKAgyccVf2
JSBdDYt32tUzTyeEa1A4b8K6RDcF0x2AfqJvj6zA/a4iFRkMpya/XMsUlOB/MEV6FnxLb9B7cgoz
jVyWeyuowPQcdB3/E8wWnxWGxPYglBImaf4C2JjHl8Rf42wZyLLQrjFbnobWr+oJfui0x0OtTAJD
lJomyC6PMhNBEXHOKEM5j0JHaiqLW0oKpBYFRd/x2lXpHjgrvtRC7t2ZrQP+AUYRPHgyEVcSbOCV
16ZGP0px5zzmF2xvDvK1HLT1LmXCMmJ7eNV6aoc3aE0LogNRDYo0Sorp7NsXGHm0r0I2oa5eajnq
qOHH3mzMmYq8xZfTOKWRZICj58LpdR8ZNyyB7Zuu9DQ5cI9pnMrjVikL+eFa4M+ez68weKSssiZm
tLEpnW19BAIGHhNJHPnpd6B96o5O4sg1CohFz4Yd8pvm7ZPdgLVW2wUpJH5oNsUTd7hEAM82NRra
93/g3wtIk/Bxy8lwa3FGQOBVYZQlrnYVcK0GeciV6jev7fUVQ4tFA0B8CHxGtko4RFEfJVsOLram
vATHzKys0BL88qeRgsOheMM3xSv8fYFZoSqEaNr3j3yZEwajCw04Wt7740TMDGk7AXeu9Zek8r39
MkhwgKfF7C0+1mF3IaFWlCU9hvzFreVJOa/vxPBO9aBXZiu+cfUv1f5wnyo9Q8nxw5H5bAs5hwdm
X61RRUFVuxy8Shcw/r5xhaEllWfml1hQBy8CcloSPrjUKzFGDGYGMMVgnHeTQJCpgLpbmVMKM9qE
1K/PSRf68KNpXyGc4+Sya3gsAq1WDewnyRjL0awW/v7ybdGYW42prJz5EWVgzeip6ujyMMH0GSD/
PiliQqQvNv8PglkNx7DThfoZnMUcpTNfaVhICNF3dm9PtyFrOyBtxwq5VQTQjypCkTQ2pRjUdHrm
Z1NsP+66p6imzpM5VMLSlEKttwS8D7ePaKjDeutnoir6aElj0rqEMefJqGp5TP5SXUJyfhOjUHY1
SdJd6CkmIUbXNGUuHH4pCZv5fSj/1nfakMohTbK9dvW6a+a9OD+X1yGZzgDfOvPNJu3hWYiKolKM
Yvpl0d75X2b8qrSMhYtS9tDHn6jFSubkHQRIIfyfZG17HXwM1coQjBLuBY16IDZr7ODGzb1+/7Ca
VW+1JZzvXNoAVqf+i2GiWTidTMtjiTKiEWVKpbgKSq+fgehs5rjCHcGA1UB6RtBF0/S9gzEMkVre
5gOcWMmkbT7PmwC/dhDJdJMAxqLlobcliNJzlU9SlsjCiLYWMqzYDZzvvsC9VqlsTm7G4/mbPeAt
gr++yAjmIO0CzfmDYFxeVfXs6nPCA034EPhcx6Sul82l6Ng/gqKELATAzp5rH3/LaZNJtAgtrQvm
wz2q/mcLIww3QMSoq97hMHyFc2sV5r9MoSsaSSSeBFfobnhjSCFvJNxLfR2IA9buAunV5ckx5KVr
qmPnZ81/XGk5teK2QOmxAySdxjCozuq3Q94v4xlva98D0sbI3P0LFMVK7xIyUK7GdScrrgpaufgz
lE+hdHXRn7YY77MoJlNS1L8DX8sUJzGC1/YiqU6Y9M8srIGbgte8YM+90m+aSzRMporZoulAU9NX
DkB5fnTaWva+zy2uwwZQMq2GUgIWFx8iv+BgCyKCd8a3zT8IFgGmdgjki/N1gw1rLPaHKNsbHnBX
/UIFqKfnG/jDWODxoBrulmV+WsyedEsniIkWT3FvPxImAHunt7suT88ryrSnrAvJQvfQT4FBOvtL
3VdUNi0K7ZWYslsYao4qhUuxlYpjoz2q84JeobylVIA7d0MXNSKC3JzCTDZqcCvoC4P6AShkZy5G
fhnMCDM1KYJGNYvOO+/V46wvGhEdvoPWjGMFwmTvZrDMutfc1+QhjNAI5pXMs4dpKBpgoBPddwBU
NS9xZvmGveM7CfeYQIZI9fESnAUT6v7fUcRJrRkIj+L+0w0FGGTq+crhjf42FDvDYj7Bu2wRU6uc
eI9wYx0j2475k0qMtQC00fb8+9PQEuKH6Q3akblEUzrS9th0P4XxdlJcrTylt59XQHkP5lf10udS
E2isz8RM49flIk6YAZN2GfQGPe9bgLR+FqeOytfdnNWPhos9pxFuo7PK1HZcWuPqzhy1WftgKiTZ
djhl9EPV9MFwJ4UvXM+99gbz8Bn4dJ2rAESCixthwgmeXzOP/r3n11sZj0Z2DdsdmDxHBRkaxp0h
lHIu2lWAjv090A/Byk5TvbjlwDS5eUoKTcS8abVXy22GXAlfm4IcV6ohlCYHC+BgvG9Np9qsm7Qv
xeVlVA5JiDe9g+jBKByUDgvRAW2vZfDL/bQL32H7VWUlbHfxOzn0wFo3CB4aYRIVtAie21+DGL+z
O8nQt9nZReDccdxvkGcmaOyFPcCsReh7MpHl3O+j3ahIzrXQa9YNI/ETD6Fwm+xuWK0Z2Vh+WNQ1
7DHRgbCBsRKhzZIB4gVaqrgxQh3ZlIPhf7gnIHHD9o4uvbjsPFegU7IOvZ15rEMH0A09t5+eBmQ+
H9lVg8gtuFP7MlqPlYnmgSmIYjuaKKQ7J2q+8JSUTbVQA9TspDL3Pi1fmwgg8Ns6wRqQ9Fov4HbR
u8eWCtY6+3c9dkt5z8q9H2IHxPYtslinfleuwGbPaJNbdXmogFFBLVbyqCDAwSbVIldF0SqtBKLC
ZcrW1Q5Ap0ssUOAxmLYswChxpLi5fii/nntn6z8bQ7gqcCds6/4MWJG0g5lpa6wrOx0+70pzu1d6
EOfXpkRm4MkbhwSkn0WGEWv2mLXgwyThqjHx8EqfwzWK5U6K7DkKOGkG7tXwR3I4iwl6SQYW80q+
p8v8tSZRLWdrkzfIYONHkgfdPA3VV+t3Qzdz0FJuCJr6FlYgDrhyQDzV7r6MQciwcyj3SKYVsuBL
NAKErO8Nngd1HRmXYpXHvajRQJQjece4Ip6UxaRrikazDWhqq9hxbucQ/ZIAjx1JM45etnkXK5LF
7jUOuaHnKfOtjH589UZWrDYtvz/j1Y2wDtGVPG+Le7lv77IssHcpJjab2FVcDUhg/FyApdQBXJ0h
GW/zVCsHNGf6CxJR42e0npNTasL9KKn5PfqyoU0iK8TN4xs6KXsukm3ShBp5Jf3eyEIPEL7ijrVD
kisexs1t1xtDpbSvziytfyIt6QknptRxW9EfcuSbUmfay1YR6hIMSHivXDx3DMLgKdh561DnlVZY
GLoji3o4UZaH7KWZddrzaiNk+OdSEuyYJp7BvzI0jECyl4tIjxj83pfP2NHVIoEdOcFjHr2JoBY/
2KBYi2s+tRbk4uZKO6J3j+2HM1rLEZZxx2LGja6xKMjiHM1XqiDDUkvJMCQKpwFV9vh1ec4DlFYM
YYi2xprvhZOXlfEilufF/OuiZGG2wK5GGXVZzUOyBgW8tS0PaNfXPCd8Meq5xCsZduNUDtQkMICr
tAWDkrCHckiGKoaozmTYtyxJ+qWIHNDQVdW/zSuXttGBSouAAOFlbGrq6bwfdi30OK+gKHKOfUSs
28JVRCmEP0naOT0/P3SEMFXW15YADtI6BIluR4G65FQHOLlqi/b4/2jXdjLj0kPrYlm9wujepcNl
Fz3jQ5BrBAYkdzID4SQLwdzl4NlBNGfxogFRZzb83YelUmj/k6pqxDOpRsjyHQ74E5UGF+HBBbhZ
3SLM3yMwNmIMvt7AhN9oDBofCpfYz9eKvfFKAnZIXH6AkdsG461WmpTIkWmlz+MSt9QeHLZFk9FL
1Pet15uWmJ8Mn/YnhaP2SKFK4VEPZ5Uagm3rVUPuuZl2JlES7RRBjynDqKu+BtSiUVHhJv9VMarE
SwnsWaegDCwNZAWUz6oMrViOM8H/pXGMI0eiYL3+ODh5KPfChjZYRAedckDefDACA2oQ7H7v1WQD
ivITD5vcIVqhlTxqJGeF41NAU2A/dZPT3p3jSUY7BJ0qScxfXJA75e6Adz/b5P+hUzwyDZ34UiMq
s9VHpX0kHhMd7Jc1zeSP7J+Nza7jHIvML7twhKbQObS56eNVOUatbDtZG2NY6P4vUF3Ai1Do7sOQ
vAQA+v8cl3X66PqOiy7SxY5LmtadtwsIZVb2tPLCkpxF8o5+rF7D7oE2f7VLaFwWLQBXSiwNIgsr
fZHqf+/0xGIagnYQUGEEA074IF0GjWlpzk0cjmzN7Z2NCAx7WqxKDLNLjj5p+x5XER8nSb57oNs4
4bpdjHo4F3ku1daQYDsPe3v2zXwur+nyGn2vwrzNUl1FkGBWhBMwTtG/xhTtYOb7Ptl6uHCf6kTr
Kw6f5qgdPVXetWt4VJlvr8QVSeolqRfHTBDf9M3SXN7vZ8uCnl7XMRaUQOOab2vcOpkfzyFAviMi
IOWj/v58Ys4RdgFjzxKT/AoNnL33fXIdNXikAf3r533Mqd/8C8hkXgB2EtzNl3S7QSBIg4CWDlRh
vBfLFj3m99v8j9wz1XUJKX1i6Zie0ReKHWZOk5Sh2uBFjowMduyEmf5oiXszzif/HnHznUwCL9Lo
v5XafyGs4Kg4ZhnkOIGxsyMK4Ps4G/DsJdrQprOrqd7evi26qHnnejEKM8/dQcVENMCza6bPbzyq
2diCt3Rh3OLyhMBJ8/oFRke9jA2NNLyVCwTCYVtHCzLqJ6KBStdFlYX+bUsPCWk/R8WGsjSKrsO0
EksMRy9oZnkbxQon3AruywMXXRrvI4P2is7OyG04Nf8ESLQ0uSg0Yr2r91juV3/Z2QUzbD41cw3j
j8oWsq5FajwGg6+ripZ/+5WolakhmcV09nWoyOcttmQEQUfxVFfCx5k0hzyuNnyQWHJ55wqGZenB
Mn6EC2sKZHqV2i+HQJJ9XOSDv6FF003x8lgQcWCw6W3Fm88MFVsMYS1ShcJ+VA+fAyzEDFgecBzM
7MjXWJcFkbcYmeVBOfOg4PRcuwgZPbn26FnrUnvIRbvBDh8zN+XJTMJ6PI34gc3BSZtJoc0lq0G/
RmT+ypHlDoHB65BjmjrAvIzS35cpxnYpI/1PpjCzckRzTBCBjmrtakCRWkFL2B92WD5fiup/JmDa
dsd9c62TTlpo0KaBkZk/ACKlN3wQmvH2J6ez0/V1AZQM2WXKfK8SUm/Tv59GrJ1rlBfeseS8+9e0
o+4iJaiBB3XMWfosEiA2ORHzjGI7xeEnkXEEu03nuTjJD/NqeDUURSaHWUri6w36XyuiEXpzdSR+
QK2FSxa7rqgKVsOhZF/MpOCW2NnGo7hw221qn0UCLOzssJEE64rC+9tKqxJ7VglAn3dQ6Kd3iGG4
7rHXQvf16EaJtfX2LFObGWzzJ4V72UbCNxBMeE8SpBmWXz3rDf6HwRyx7epmdLXveqwFJekrAzwE
YffhmZu0NzfXuvGBOLcm078/rzVWp42CQ2bn7cdB0OgxJUe2WkSInCH6u7LyWi4I+OVnHuIlC5sG
2qlwUbzLGuE1cQeb0e1ioQq6noMCghBFKP8Bhx8n+NnIY+ChJ5Ce5tkdKE4zjOcbQpd6vMUQpX+I
+0Da4EYFPJ1Iw5gTn8Yh0UA5ErT+a/OI2CsQbUDDcnFCbvXcNe2fQBUVUiHt+1vS7kknNF94U5cX
4XZszvVBPn58vZgMN6vZMZhjRy0j0wWvuLu97Lb9YPUSPEQKW3bP4eqjWSB3Hsx3UrtoxerLZvZh
udee7lrZ56KWJhCnpoucHASsQc8qJDYUhbflfnO4RbkMJTAB5GY1SpTLEXA0NzStZwDByhSU3l4G
026zOnF5gY+DqmD9x3uDNIEvhHqfYSmD73AoGSfnxdCs0iymzMaXiz/7D049/fGoLsSyj3H6BPQG
9iZ1QOVXATJGuN0P1KII5nlFHT8KT65qcJ6sINWlkvbWYGGkluWL/UjQ145RmBMRVv7QiblJqTEH
l0nINQqlmjHgt28NWCOEhYV5H5H3m3oBpmp6VbedvITAVuqbl6BeoV6wBSmHELuz1hi/EXCvPOVM
r4Cd8J8gSvFE9Z+sn6aDjsYIFu5gIzzSJ2YxG2fxOtc6wU69vLGd+BEDZFqTX7i65P0xWwpO6zE/
87b7awVfZs0aGrtq2MIBJKFzjlNDK1pMuJssicZzQ6Vaj54UARLduCC+5YpgOumAXAcl1/fc4nIp
nYXUWFkvyEx3ta4DxtKfyHzdRppU9bVCf0OT1xofV+l7EDmHsqn8tpcwXEDQ0TBrXhc8SwULEs4X
rydgYJWtKMh5rliKfAEZy8AJIes8Fl9jK2bL1YwxaeQD5WRJvvuXMfnb6VpxSclv6hTd45RHNkEQ
F1z33iHvrADtaNdAaOlfljf6U3fVzV3pti60lMANrdZNKmQd/QqzNDxdMZHrwTRndIsi1nv355/L
tKeIEanTVeBN1ixZnAcpBROv8/pCc0A6BZm1wuzpkE9jT6W1n4bjLmf2TDU5HcwXDBIyFO6V7PFa
9sCUWtk3P3WIaomX3JEZyGFU2gEiueAW/B/rtl8zkyNqm63cwFWjw3lZuMAOvzu9IXgobb4tatNb
AgEbySSmScgNtS3ONkWNkbkIey7e783gvFSy6TdY1/YRftmXLDEYg3C1R8Wjt2TfcmK8Wz1HiKDv
tY2pIjhNsw3ALAukpwu48i3jAU/qIJIpuLZL5uBSxOiMtTWwIs2jQOAwuirJ9FrbOKHeEy6aJlMs
8gVl7hlEG5Ev6eqzDhQ4D92I5+CW8GDo+8WgIS7NFE90ZG2n1fgXPa1t1o2pRTMXziHpKJKjkSm1
+vNdalkzc2+a/gRqH1WsybOuYqHufxfNIaRBso+KBFX0tyxqBsllEk+x+SVmzC8kD7u2JUpHJTq2
eQA/MpM1qpnvEbHJNMHntaxWMR2uKyrASMDGx8HIUmXqnEpVlWfTuJZ9sEsUIzqJbjQmKHn2vgEa
Prs2GyfBBdBx765kaFpozJnrliDdT8itJuVFJZRBXoiWfF2zJNNnNhromLBgKPokzrj2WGk3r1NM
PBcT5m3bdg09HITDlDFY+fBue0UXLRA7rZGK+FQhpWNmXFrPsm9+FA1PFOFRALVo34le697s4xON
f2S8etmru4cMDwoeD5OAAVoI9b37R2ER3JVs56bTx0cYuFqKFrx/4p0fUAb9fHwPZ8meCb5MKNz5
0vqv7Mk38dnddYUf9nG38mNW9I5Kz52HW9UltaWOx0xxmS22MHN2/PzEH5edyI9dDF0czDeUrZsn
vGx60C1+G6/6IbFZuS2YhmXDJzXo9+EKs3gqCWcVnWokOvHFobU89a/YoobtAlHATJaHVeJVA+jt
/FZrSGXJCnnvCSr7w0xUko/KX+z+X9Xa0KZJiqy6O65F5SPlEYZMn/ttaQaEPba5EwTsKQAKTwD5
KRVNBH0miC+1WBhPVGkCw4SuKtgHXSyXkur7+DFRRUbNIxg2SkvFx3kjeUK/ZAjGoT5P3e+7Zw95
EkqEGP8fvxKG354dX+mbg/l3PoCuLacd4uFJaKIDlPAdC7GnFcGr/yxnb4Hgf3KBpVxSsObcG56n
uYgTRofjNdZ+qCTBgyUZ7OS39Z9irHNnRDIsjC6+2D1Y+4CY6hlOZFM/6me1wH7FPdTNKsSn1Reg
si+ipA6E2YUNPvlUpEhY0qJ1TNZceKFKTQy2B55wQMCVszLt2fbFjdlfErJRH9qn078XwF/iFFzW
U0mam/I7jRO/BMe7mV2QGlzstsQGaz0IFSSyMHEaHBEY4Cdq/cHucByc5rCvSkFmi4JcjU/2yocm
SmLdx5k2OmLqbnwBlk+oaNf0J9SDI+rshwQ//uY8aBNdMLPp02xYCs4h1pOuq5KeQBChmkuTDI5A
sEpBknz10SRRZ0W3HUbI1LU7Bytvzk5/22OGBE0HZljrUQXPXLz2g3Nlqi+gFnhc4ohDp03hakes
iRSCm5wEu/VpJ5FMAFZNR06UdpNYlbsBWID7b4uzWrWnAs060df8+TCKy3knVHE6T309Y8lDONxN
53eEqxRbrRqAgF1UGYqkWvzso9otSBAf1tb324FMSXZHGOX4wQqt4wtSvRb/5u9TSmmxpGFxfwnK
1ebFXnThGfXohmi2bdCNMWfh9gyA+7QBkFG5weaM8OgdN3NBaskgC+dU/fw4qk435NG8iU/f3aZc
9mfh/x6Wq1lHaNzYQIH/u4CHQiPMOuCVR/VHNkgWMo/0c8qzi3tI9zlHpxyEfnX6gS7+UttVCdvv
c8o7rnnsIa9zkPAnSfsyVxNbG61mW3fKzEpp/FyHNLx5eRogfy4Y7y9xMPN4f/6F6zPRJwbggHal
qBc/CXslfBy/t0HOU9YQNmNGuC1XFXh2hEb21IGF9uHG/knzRHlER3B2zAkp7lmersV7uBYJVx/4
Oi7aKPxwK2AWKdTVLWwFpRKX9d4EvEGRcWdeyBlrGHnBo2Sey5DyuYI08LPAPClBK5Xk247acGfL
ZkyI2LkV0rTTb06QQ6FMa6seyzSwNO6vFj29wTVxv+eRLckKNRsuI9gS25zUdZBmFYC0RJHvIHp4
e0xo+xP0PmhEW9wWD4mtKz7ADmqR6Y2qp1JSld+pzkEMzQ+lw2PIpQPdit8UiPFw9muCKD00bHNv
ChNpq71N/v1Nh/6l1H/5GZU5rkuTmSof4703VuhurR66jMuGP8zulDfSwytuXrVUZEH0wHTd5bZ6
C+BTOv48H/huYkcRudMEE1BVjhWbAnK0kSObEFTRXNdeyz+OEdCnZl3tIJaIiQXmGuLQEtMO0mAA
pu9LfRAeR3VJJcpnSIe0IVwO7LfeyFoyN4p8I5mbNolRlv2j1MrovK0y+6z/gloTLN0YvU23ljir
evDXWL/v6XmHo/UmSwgsMHk/JBnHLUCzlumGwHzJmbrkK5On7S9f0xgwx432qS35+5sYG+T9eYM3
dJHixukDzwsoBSHRH58NVBwdTnlgLpi6ht2y0KqnE7q+gpTQeaL0Jt3CO1mEFf+Y9kL6j2V5JtJi
8IvazbqyDuNzudWdmx1Gd6CTsIHe2RunwL9boApJHvZ7+L18dcVCDhCNEaI2O5mY5Ye0OZNxsPx3
2O7XBDsOk+DD5jil9LIlFFRO0GPKKYcmgfIlHDwQzZk1b7EhojCsyFcP7kjPH5be3omPVCNfR91g
OJweB2LFa8QiUh2H5RSZ3YnxokIRas+qwmn1/tZnF/PzPOd2oUDLmpDDfvy/DRgvpsa7f+mhqY4a
XK9CNL1iuzRivum+f1o617ahBOIqpgqF9ROrm60FeqlSolZtyD91ZxsIAg9uxCEY3MkzR9NXflPR
msQWsYRbb3gXVzEbD0P37QwCc+XEnoVpsbEsYng+esx2JUes0RkQOvGhDFZr7i4r6gSY+B7m+5gJ
fX/mnAzNjpnhSuZqsK7UuqhDs32AUP8r868mGTm8a/tyR/xBGRsVTz8cs0PTiI+Slp+EhgbAP+Hh
FEyB699PX0vH550zXyminGh8gro1ya9P3y+I1yYFT/mMBEWK6imkLQtVPqFyq6g99IGJzlXVkUoV
bhPct+GurDrBQxtFscTegT2Xc2bQTSHaZg8jq5N6VOkUkg/8vdjFqE/lRKGYQrUGbtLI3GKwev33
o0g3EEmDDH6Ht4PZXgRnYYOaoiOiO5Uf6fks51JDBi+x/Oj2m3F7qMPSldGgdPdM9liuV7aLErbn
sQgpR4qrsR0Be6asTRYe4zK9CRWqB5GTpYb3P3tDCVPXusu2xi7z3/ElvbnO02cCIdHxmWO30EG8
UsBKZsWfG9aP6A5fuGTUvr8rLzNQUzwnUBS61ltGPSxgC1z9gCxXjrv2nG2PNcdl71mw2KvCle13
a6+i3Lqx4dqV33Anrq8v7dGnCaJFLgGm/KWIfV+9XjYuY11eI767h8mrtRg7r96J5Oujb/+krsQO
v6KO3drz5UnBuFFk32fooJgG2UAu/olJ6i322gwCRrxfUyC1+XTzQbeCXzG3TSKfxoElzqmWy8OL
rDUODXpUZA4fS/Gw08uhD2ft4KprxSxxUlxh4deK+cCQ7Qg7zKa3TtQv7jMFDyCO2WrLOa7e/++8
D5VsbMX8Q+N4ZlhYpVfzcCsvDWwMDFiFt93eS/Tggsrgo+I3KKiu2uh/wOLtYSbjfyWQJpY4lnTb
1R1vC5OjbikZch2b7zHrZFgFRvruPFxQHhHIqQFLiGQ6bHbV3IweCcRHdwKT5I3WoqLAh0rIT9/Y
B5M13d3BJ9Hc0f1x+v3MJ1Hcq/U/EsMgr018zNpn1oQ/Sd/jO0LICdoAj7Bl3UPiW9hNq7ruE6uv
+ia7MlLyBiRA/S85Vo1x92WCL9r5CUJ/Jp5rJyq9XGwpEcVu6GWMelhU/iHKdC59GNi37LDpsJCt
HHb0Y90qvAHTfejrpVrIeaBvByur1SHM1CG7zSWJPMkX3MMvNHkauZxLNwJ1A4knQ+IqIOxYwNmQ
Xv6kQo+rUz+crGsAOH9Cog6S5O0ZE0jXTnz0K0Yva4k9aVEf3jzH6+21tQ/yXVxIoCsFV2vKb+C1
RljdBLhSIyL5WCNYah3a2lA4CHEhB8VeBKrpj/pVowejJRb4kOT/WSYUk/4JKWAemTNDLhUAN0nS
AQVW74pR2y6Ue3Db1GIkF+Rkj+TYmtM63kZWsqyYFCYqkC7r2iALeOJcUuvabVZFGN5H7fo5e9Xt
30IPhSxSe91pG1MOxtPbhEG+yppOHZOJn36yxICtrg6s9n5WxZ7oWn+0D3OWWb4B88tXpkzYdUim
zxQf1Ww2ZbQrxA1Zmu1YWJfaBJX6QT1i3oKcHmAPymrEh6zivFvF8cIEPumH02kVaa211LJr0Yuj
PCC+kTCPDLwLEu519Gx9L+5BoZTNUK2wgtnffKERgUGRTjbJZYyDYqOHiVCdCx4S0js1cF+4H9Cr
xgoKb59fe+nFFAWqrghFHJGPTBxzjTIXwxxIdMh4RTGFBfeJf42RKVfdvnIu2JJxIEJfw05YPESq
DTwf5PrIEU9WCL5Gr6cUvSsuS2RyJCLFSy8+vhs+rYDyI2knJ5DwSKLyEdL2wrMHGADIzSeEDTzw
U5FWJm3R511EA7Qvv0OWksjUhoeD0zFwVKapyEE6EFsEkCHNDerSk6ojNEhjsQL4EQG61I3oTiyE
rdXsEMS3lHf6zBkoxQ==
`protect end_protected


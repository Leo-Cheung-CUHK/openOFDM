

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZBY06y5BSEA3vwLtCYy6nxOZv3rYFFgZv5ABjBaqtaItkwdtQfFvZBIMhBOgu0+1i4DhnUz7pdYr
Y88DaxXmyw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Q91nMYZhjxb8KT0ODrW+miquus8bIV0xJDXXyQLu4mbE2ZGK0HYqPk6xE96lKrNSpNViHea0rEyX
J3Qsb1QJLBM/4rnfg8PNzn8acqAN22JgnqyTntYQVpk0fARej5ldkyKbsCPgkFDFJQnDbUHBIcF2
clV1QCjE7A3SvN91cV0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fpeDNxCbq4trL0iAEhu+gbl4Rix2OTBKp+3DlpwRVRrJB8M79X6xv2dY4g29GTJWY/qcPCM3xauG
RxLbIsN70w9DSrpdJ31jxXSOp/N0b21smrkPYOGR9al1eBkfjYMFWbiVzWEKHK/6z705awwEunRN
qhtuKyDzs9JphrMi08O8ld4FYuGNYbtDOUXkizCIgaOdAfQTq0yCDea9z6uJ5sQUPwqrjRIroSnJ
mW8XvC4+hFTtIH4kcsR/hWe9eHVCVq7yIdgTrHznDz5I4c7+A0ZUoahnR5dHirQC2z7KKzrCldej
93tdxPQksB7VjPElshg8WP1MGrwn+7hvSijdSw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
No6agU7QCIBdcP4teTJDlwXV+g3qBzu8V5gqFUsql+qUP2ZRyYvAPscmGZyPnHh9xvIYYFmXqCE7
RRM/BcEtyrJ9GJvahRcE/doL0n1EHIOASw/MZnFHkf6gtqWvN+SIv29/H/UyUfhuDXqJBGjBGBRs
+/RValRovCLF1SU7AdbCQbWKJbpj9JDmu7gpnhPbkiKkLcd0L7j/KcvlPBvHLG2JvHXct9Oyye9y
FJ190Nne/diMvLsfTBKIzRzQiV/kj3aSYxw4yzuKLbdVZ9eZYqFHwhjBXrVIvIAq9zy3Z0JajEGH
8Eg7Z1uVL2BNbnB2qP4/6a3wYkq6RDa/mFw99g==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Au9tuW8YCiySVmtwoSZ2LqBsVMwu9uzGBs0i03rtA+ohnDzpS7/saWzSdnxtvJsmHKLPTnuG8etw
O+1iKknogGQAhYN8j4DK0/PmelqEJy8N5vwkQ/o6l1cfVFLfqvAMRbZ7lkPzco2SCT7/KjEJHW7i
5gy7tqPxnW7QwYv2vH65EVqe0p2tQ2kCHVUvvPaAZbeDzA1LHleCahBpWEI3g5wztTT869s7a4yn
1IeWyD5NV38NHHcwqubPZ09C1Vm5NLAHW7sEnM3is9mRkFnCh/x4Fb6Ecuu4bJYFhgmNzCCKgYK9
PEdkW2OgY7EzDM7ocQQuoE0+aHQvw9lRdJm00Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
n8+Js6UruWrTa5ioc59l4AeAloQ6ZDwzPNPXUOknQWFRecrzd2eOQ2KSf6tv5Oxix315yAoI88kJ
L1R7xZeU1dj4QCJCinzjHZXGEfUurXJVEcq84ofioKIpCyBd7YnxOq469vjhUCYiTJvMARwPVvDY
U+jspt29lk+k5/XFur0=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HvScITgcbiG4YgkXwlLAPuMki7p9oPIAapsMuPCpK/tVnY9llE0MvUk/POKYiMFRuKgzht1jfNyM
pX8Qwv3/+iDiBgwTwibzi053ET+OglbpoF/MDrRErGx8VRvmBKwxnlefbxg6dCEzjNwYuFpDkHVT
YZySWRuz7hA0uzRJwLLkvg9LoVoAsjHpp+GqlpSqfuVaV3IJzpIboKGmFv2qLj7Z3k2aE4HhZfXc
HclRJsWxw/CA2DK86EGTnPC71xJNT7pgY1DSHCglqFwF35L0FfZes57Wpz5Ka6YR9dKPNCocMfXO
DZKOoy0+Zz/G4HOrhtHGxgzfEtHjRq0ZthhxDQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 99168)
`protect data_block
VGPDfuyUzWKG7ctIlRofDvNiiirq2WwPjjIs19AOm0C70X3Wv1E0JPenlx5mRmLqQV4imWILDOUr
zRpclGj+qTEL65m0LsB67Z84AoviX64xC1i9hYsqJRG9v2tTxZ64+iMOFb6k6XmzHus85zWduREv
7IlDPP2w4j09yHPlzzHs/7pHaV3kC4F9OG1QAX6W6lNXLKvy3ITrqLBEwPe7mc5CBQLKoUX2LDlV
MYmCki3/9IDmAXkvqI1sD6+RMvc1gfTMly4xSZmtThb9TL5VjRHBpeQ49XZRwyX4PoGqXk9DpRln
dWqUCAfHJz3JK6wJYI7anGHJ6aRRzdKD0WWPD+PjJrs25OawCrCLi/W8Smo9qJUWZyBSA0o1+nH4
t2b+JiE7p9cGJ68msNwpq8ENo42ffcya4j7Z9ucSwVoA/FRHOBqm/Tj8QjxHNITwuzxeX+jVkZju
aLGmU6ghgnSH8sOobTbdOECBOF6zaPvsoPbsCQXTsUzC2Pg9Gok391Txpotb4bnJhV42oC1HnLIG
R8nh7YP2grpnsHFSenHmecOdh9gEWbGSYVP1MUtPsq1k00NfbIPKtfJZmoOC4jSX7NlDpeChNDBp
fHbCxtLMawyuhABWdrpgLUMY6W9ledxjnvjziXNG5rdchei176dKv2xjUuUQLIRvu2V3PuFaZAiS
aFtuLtwfM+1Wek9voXbYoB8ILQVt0kg+16HMq/QFPx7JdMjpaAiT6NYEyTUbWe2KvqdFG9+xOPOu
NENvwAq2A/cwpqEfZsZZsFLyzS7bIUFlKs6KIMHHOpi8UaDllFe+zPIvw4MB+URzN5+H0wlZ2tR/
51/+jqYL/QriIMA5EJF08ZmsaScJoS96lcsmu5d+XaVzL5zYZgLTLSMMANX2U0K0u49MjF4F/ZYy
1RIPvVtbvYrJLMipnRYAmmCayrMhYdVjofI1RmSV2ZcCHIzNFePXcpR/K2gb08IMdyViiEVzLTmT
am8Sjl8a5KaaL4NJx28XKoeh1nTpk0MB9tMd5+SHXywf8v7/37m8QGsrUn23YDGOefDkzdlgAJyr
121Ls2sX7iSgp3ke9soWv9j2jXpT98sKmYBF8IL5x8kzBAFB0/g3qXJanqLDbZf2QqmAe7I3qN2c
3Wmw1waXPOO+Vv9zutN+tDGRge8w3K/SfCbfoxosldkFVP8OFb46yV5EJi3HNOPhpqHrAAnBxEiQ
2SNixHIUqBUbNXxdmmByo5cMppBP20/cKj2AabCaWwfCZdtV6lR3bCKMIzLegFrqYRhb4whROw/c
ED743oSktjSFdsKxhn//Vkjy56qPqKEwKHDPAyK9qCifjkZQsXFOpB64gx8FNKxTFrC+T27ZamqM
0PfwmVn0Rgw8EYDYPpKtLUSlpMkhAnGw9NgvJenkGdHmBCsZmTbkFot1obWNStfSxuQCrCG9XG63
Np5o30WQZkXGTytz6WLaUOSlBYaAFr0dVivod8DtJVNSxjMyz52AhdgF+VRTsGmBxyLP7Ilum+9J
olU+mjYh2/UI3HxmZBaBRmFW8MnMfjsOVg/tnm5BkXaFThoy3CFgM7RIc9D4zt5A3a5hjODGsLMe
o0c0n+wP8Vv+d0GD9xJ57RnkmIwxJhr+v4PUdrFa3NUccodeM19/63ksqo3R+422P5YjTHOWEwTy
44ALB4+16aO9n4aAC/49TlDJxB98JHhmQpau3TOnxNE9ijpYKEJNFX2FO69G0DTYjRnAev+0CwOo
lyLuvrmoAq1sKtb/z7UFpNvnlS6hbsfW/ch0GLXo3KtI0pkD5qvohTT+rYnUPiOiua5gHJDDLBw1
AHs8Xk1z5a0N1FW/JRBKV6AO+tgWvuh/nGEcB4WlZ3hRywd24Av1HuvlCWaRiM41q+zFDwY7IWeL
901rFwi9NkikAN2GT38ra9a55sPLJF8eZwAvSF2ngLf39AlKV2IQAJHX3MRoWNpiy5W9b16OYNkr
34MhT8nH+SO332Xd5WP5o3eHgd6ndaTxbX+ZxOUaHl/UpsYVwlzTJBZHxmf9NuNZhE049HteWryV
u8YR4MX/xFyJmOphVSpa1+FH5tuvZlWuSLq51VD+XRb94QxdFOopa7Ik8sJO1GVjsUK+n4O4C6hJ
ZYtBe4HX6RfK09BcZDdv3ZhQ3bd1ACauPBbCywAEs9hoTfx/vkx117bU0rzxM2LeH21Q35Bh+0pk
ZWZzeEgAnXK1n4f46LsSuwuXCuKNSt+L7+QofaQqAlKaVhGWc1hvsut/mEaBcg1ZqXzPkxHhmF6Q
2ZOSPku2gGzNWM4hTVnLr4iD66/XM5LqWZ2h77VEiRS9rO1smhr6gRtO5IiJ+Njm+A2mRBbwZBWk
npkyP5nkpdUTrzgILAaFfFc/+zNzF/5SnL5krni9hGSes1D6on9aW3ft3w4PmPkzPkbxhhmFb/b2
7Efx4Ul6qanG2DG9Te7nxhRpa6iuOzslsWFCCKGRrAHaOKnSROOEBx+3p3uo+leQDRrrsjLmLJat
I7cyNMm5W7IdscAqeGdownqculW6JHnXD/we4eRUYonj+R471kPFbgONDVWhMAVw7GgcHcXN20w8
KUSjsa6CNZqMkZYi7/9vB0sIRMas9atSlU1hcHgsSpS8ab2YWpkZdgkzxSR5SMqkgvHLN8dCTUb7
Ythd4B4VG5ZHo2/E9+gIJKFvFupU/unjgo0dGQjjRa1Wq2j10LN6WG/xyMZsDhRF5J3B0eEyy/M4
ieB8qpLvvG403sKgV8zOWb5T+z8EyUh2qq/UdyRwg3WQN0qarMjUAxR7z/CbanoktQmG0OjXhY3Y
uuSPkJKIgaaD2iBEr6qbKVOd04duPwbpLd7SVon4oJ9b0ultMcOK0eZPuYKcSzLBEJrNd83VONRK
AkP/xj/yIKGhR0vUmotO6rKh6cH0VhjpS/WkV0h038yVdCXCQ8mX287nCfxtBkLJr3JM/ID9RNSC
EJnoAg1Zwmx18wyS2e24I1qxtuJG7OjNihqExvtYlTITTkwdecFfrMEAkqrlCs9okRieAsKyZGi/
6AEa3qaCkmYeCvvYtinxgDNC7aGJWB/rKxK/ylV6OnQVQQISW6XbUj80KwmnWy+4Jq4y0t9b4K/8
eFGqcp3xklqs7BapqUKdfkTRPdHXhE4UdsY4l6rqgMd2HjZJeNYf6k8Te0O1E6ZauM8G1HPDpF5V
b5cBLpP1bEDhe1Wq++UJx8PAigayXi+2d7RIoIyRIQC2uNck1jUb9398QFGcpwxkgn3Uy7WbfJiS
Xuu0xdPHCrvkXAfL6lejKga4+XL/+rZJlMPeSnSczkwYisfVUMAagZctPO4mR+NCnZJI1/uSjj/6
AirghCLYxL+0j9Onrn/h3UvrIUB/QJ2JkXZUd19uCiySuiVd0LKR7rd8XW+qh3ATPvivQoHkrDbC
YK2Ob05QKFXfxA0dn1n6qVpHwRF+Yh8lfzX8GZb75QRVYQ9imrVokBp+LTk3xIwzg1to9uaC74vn
A/5LfZQrEu5IbY29j8ylxkmCLpUhdcN4iBnj3SIxUUH/Flrw0uJPns9JqdQQANOVi67EL0XlrNVH
/Ellgiw6yPGBFuJQ0VEB6vjrr4wHIq6coGpKyAwP+O2gK/xNj49u60VVb1wH+f3ePzAmJq2cjY8S
rpDQE7QH8ZmhFYAGqKgmjGt+CCT35TLtLvymzBwFxOHn5AUhPX02GOIzM5/BL46rLaHPT5W4Y9bY
77KPPDpFc44GU7PKT8be6BNAbgqXpTiLt1K4oS2JgWI4dS675jWlATw0vP+FhIoKyxS/ROyzlNcf
RhEAhWf/S6uxV8qH41lvpJjUS6USkDmT3kDaE/lN5nXV7ufSasNcMfTKZlb8NEFCGTimyE01e+4r
wV18k3qkgVISNYEBOMtQ2dg3xpiqzmuZ5bj1ukk6niMrM9GosNa3cMmBckVk+OXNaCCJcR4N128/
Hk4RrFDSslbWKsdKr20aN1tZU2yCroe6OUSKVTJ5HeiAWqTzt/LTkrm0CataT0JhmVdVuEYa3hxo
qBZmbH8N3J4nujOSegtP91jOMNh8S1p1jo+bZBPYV5e/kOIwNT1B28NGw9hvWCG3FYZaAepolbqw
aWuPSxwkVD1AfdHcoVgMUBy/XzHkzB0AHEwEqMXZpcZ3dJEaXlK5vxfKdV9olQtSuw+gBz7tjbjL
z3FQ6MWNlvVw9VrW5fOzhJ+Zxn1TWrYAGrTzatUZMAs4CdNWZko776h2Rg0f9n3/yPOobVw5xDcU
x1A5q55Vj0nUCxuzQbODHf0B4HUAKiv2SzI0VVlYwuixrEXvz6HPkO5id+PGCl2/QMi9lH/Fpgp5
k1elYDgXAlinYJ8A6cR+y4yRauL7lVEkvHKAwWK1lEgWAFv9cRwq/B7v2hLsaWQwPurKUEesaFcJ
ipyUmtbu4fM8r1BkY2HxKZzn9L58bKQYYJ72Othnr3O7LLWMl3VmpW588U/1yExcNkiVYrIwIA4+
++9px+st9z/FXJ4/+f7XGQZ61hHDJCXM67NxYEhrF44vDHUogwHmuRQQHeBIIy2UAjt3ApbjtHKb
8Dw0l4sj+63AepEVqJ6FwGrNPt5AtmVgdaasPbnDJyJQLlskn7ISzSaZzyjq6n+kVNXwX6/T1VSY
4AoQdRB6eDuNHdjLZ8JodeBlpUzBtY9Fbxqg9qI2TF9spR0lZbaxjZFmT36+mcRbIjDab2cctvn2
e3uK8wRt3RP5m2MIOg9/lYSosJ3/vd9Qq+sFRVPBf+UDPBoEa2hbXW2w8naMUqXGMBi0WXrU+xXF
wcJ2/KS8N4XeFHic6Rq7iGfJ4hvxwWZjotrmVXDG1qvh7pn8ECd1ASvprixBbfu6P2ApTSPohNkz
zIvGvhWL9beaQPYO7XR+aOZ0FOgNBqsE2briH8/z/qgfk6mlmFJXkgl2ObpA8R1XlES5uJEtgTPA
/XrWMVPiPumzIDh6s/SBCUTNL/7zCcpg26ImIQspBxDMvd/CF+S23hP94PQnnVN6XFkaN0oLVNVH
AF1gMZqbk2+veqO7qNrLGtz6q1+NORfIbnN/1JYhORbpu5BOMQbZgflJB9gFjTDmzg5HkdstaAuw
yv01CxPK2T4IfwchAUhiFRp3ztvKCTemFkTXw4Mqbl8Ku5BkfxisxQ4YbwAqUeyQk2IL2/bBfOYZ
vCFNx38mfu+6aBLOFB9fIRsuvAxNwPYv6EMwbl8zmv9kAkP+X9amPPLy6k/rMuV70JShLmmM0Rht
euRdZUTOf5XWvfiRIRBnKhLjIu20IHXAZfLSR21Ov3vR9Q3e0cX+jdUE3EkjsFXTtyT9vqiiGqOo
xtmF9t5ocbhdOYSPOv4QIGhuW0Br/zLgtHTJHgAWc7yfDXw8iGuSQmM0rRkgG1bXm7h2fC5M9tf4
gIVfC4OhAlWYDTFbk+lwlqmovvoALTnfNEh+JUYcwLn9VJOb2+7B4nWLmZo2YXZfUmQ85Be+A+sM
sOnPrkrIqSW0aLAfYuhqY1SQB4C7oMqFyWS3bp52XOIIOfQCv8dBAUeIQG8ODEoYbHV4c94k4/Nd
fsUTDQDD/54PypFklhA+yozCYep1mlWeN8h0KGezt36ygXgPEYX0mPaCabINAiZmeSnfdhtn3hb3
QCxBw0D9ZcLISb3OJlIr1P3YYWSK+KVaOZcld3D0xR7YdWWjVtYAq9dq1ci5z9Z0CrI8s+2R4Ysy
JIOQEVsrx2fSZS5ijMKmUkLo6elRNfd7BDiS1lbRTD1D930J2k9oMmn6CvmEgO0fLkDu07Km0vlC
+gsphOuk5UARXblPQsP3Vw8T86ygbhWXx6viVu+iahBN6pwCyTcw6uJhTA1k8U7VXS0B/mIajwZa
mrEPqGLmBNNbeWuzYcy06Xhazu0px+mcF78p2XHtF8tJnBIZ5qxBoEdYKT/VdpAYl7JE9LO4QiT5
BUJHDgUOXKLghveGuQY+JC/hpebOq1r9W/S3M/WburmnYmT9RXViHCWMJ3k5WaWKBCE8ny1OwdrQ
zn4oE2M8B7i4kwZv9vpgg3HFDDO0HJW+ECOnwbE437AeqJr/2IIvYLUHDFLi1XY6fDjvJeKpmslD
Y8NFTQIwJk1V4hqJVOUTfW47lRLR0oZNEnMifKuZnYVhRnUpXbgkMKcpfmIgTG3oSH8J1ngzfVnq
P1O7WyJf73yWcHL5aiMOJ27nEtSFeq1ahntpYjzxR2SXU2FR7Vvva+p+SwTCWtx5FELkgk0+m5vL
uZrtvNmo4ThN14uTLsRosByk2EokARLz5sFRntHngKKO++xnZFiMhMB+cYZV50XRz915Idu7dtoj
O8y9sHTRoSgB566m1BhsTg8/2qxkFie5DSLwQrRWtUKMdmACkwoWNYT9XN+EsA7rI5b+cXhj2Bjl
oHTVf5ah7Lvp9+TXDwEAxxecATeH2/SaxcIGFnu4Jyx34CoGEdm5/9vQEqLQRefauKLEOKemrnnb
EfvmoTaNwDsn/djoTBaN5VbDLVBS3CrPhc968kBZdagxL8lJs4xT29UUpSgJsWO7YeOzYC98r2iE
fEjNuplJyV/bzH7QgWg8DIQBHAOhnCOAlccYX9M9yf6TIJtZzEnagoJIgAd8i/sHtb9NCjc8N07v
DF8tzh5WeuRlsRnstbi5tTdSHgmBVtkva4EUJPtDN9fEG/Id9ZnEeK2UqsJLx9CeFYCjgPQO7Z+E
CHmjnPVHLkVcM7r6ZSa0QCdTwntLP/u/xqpoB8omVY6KDTZYIa0DFlPbSMj8tuxK5l6nVeOhc2J7
5M6R8iFyd5CNkOP60jIzI1c8cuePaIOEVPdk48MAGsKqAI82kC0qA04YBn4GhISYRMuYHkiW15he
Tl/frnF0y2Nk5/jnnI81qpDisjj7itkQWuHSv+DK+7Pj7Ie5Tn9hKSIeMA+HZaDo3wQWSXf429I2
fskoMlZILfRsBxk+0R9bHm/n3Ijtn2rCVQhUVhjA5LNsWwAGCRh+b0a5fgBAk8CSdup+J7tNPBzJ
YVQjOFcfBAxdcHenfWB1KdsXsicVeKic85Q5QYVd7pCAa1leHH4I5UzF1mrXin+ARysmvtb9LLQo
MfFQ78vjOonUU/uSLk+30Q4jsMiuoNdTqxXn3CtM6ORhMHfuAc5qOhRcDPARIaqrelDJmgXYpI0J
6afYe7D18tx4gu52KJGVqZMcESv90rVWmHecMk4i4AO+RhfOEvZSil2BcojS2KKndFVYiaHlpRn8
QRn2BLlwPp69UH1Z0xFhN5vlQ+HIHNl7hkxD8tAysh0oY/D74j1aOPlyAS+sBleFF/ve1/fYqIvT
SucNunqihgvNECKG8sOShqaTpBcJ0XxCyMHck7d51nhAi9Ofo2E45Snmg9w8s2ZVleBZU6ZWRXef
XQMRjo7tjXIO5Ei7OxOnoS7FbNmXYirRyaLRJsw8XwKns5wSNxqJXFppvBG11ltG1zwadW3XaCwH
jycxDuOo3/RvHSK2yACYYzQCH38CVrzbJvVQPSfbI4hCnDkBE8hxB59qHmMedfYclTcoF8VlTHS7
/UlhzYJq2hwrAOZNKr4UHtjSHQNwEfHalKxKzEbMwQjURdAr0Elkh509BgvJ7b0h3ElJweQlaFQ8
uh6QuLG3/wRb/P/Sg1Yz3muOn3U5Km3joZh0h6plpz/qDm+d8+DAiz4FW6vaqf7PVcnKtYdq2lL8
Bw4/OdZKwI28bkuuYI7G5QPJQDvhscLDPTwZwhQ3y9H8lxjN8F/CIWpWanzN0lZ24qTmnnfU1bns
xawObAcGwA+VBgIUO1ctreWs/8g0W7jEu3/6puyIUJyfy1pWfPbEpTI92pB8lyBuj+Zq3brfL9pC
GjhEfnEs0nci9uZUa8lj4JSgquRoRZtnBIspK3635+yTHKgFhJmO32S8AncKymsWjs1CGlmqnCUS
90BiP661MwDsbEpdhFdNT5wvoczpXVSHv8UvJ7+JCs3g5URRM7TS2VFoETh1dyfbLiI4X6hFTR4h
s3+kLZqYACRFADtmUsSgaFi+chuRfCjLxbVzAfc8ou3kzyXilaVaw2jswPASqENQuKSflstLaxl8
4LSnZiZ5L1WYPVXvWDidDTa8J5dhEFLeNvoVGjsjOb93js6ZsByRSF4MTjy3hC+ZnUx5j/SWpMLj
hYltwGHtwMIfu31nLm8dhjSiv4nNUyh/Sw+/Q5BnsWoWwfi5tx8zvjbuxH8ZOBKgZGxvIUlFAOjc
dZNNoXPSor/bfRyC6Wnb6WUjxOcb+NpCvZYBNv4KNqb7QaXa2DNjQqecbmIjg/hfyb0meVVGIZX0
ZysrErP0UC7WrMLbcmgylIqYMYgjry695Ond6nzCocrftrkuSo81TV++BY5MHfNMfMgomWVWDMV0
yXurWaWpFhVbFr2ajf3DygsBYKJFFhoCCS1TAkLHmvYrTtY/PexDj8WpOvVBbCfoHhwKKoW9/blT
ha8FvmlVryDMBnV4AKubddeqs63UY5B6PS9f9FJqgjWtak0nHoT9e3i82E1XOuNcB5aJ+rAc2YTx
tXlCgUGW3DQ2bcusAsIBXLyLgH5vs4Zl1d9ShkQY0xf9RZ/7pccmaVZQ7usqmlQX7mbE2FIBHXvv
9JmzDV+vWBcQmEtmDfib3CvfuDtAceXsX4HdN1fNoP+Oyq/Np4HAmFWzVYfD4Ht7QJ5+rDTVT12M
jjTohl0ffJgE3sPO1/imgIzu4Zo2/HkecGtbgSqzJqm/axrjEpCpHT0QlEklZJaqxmM5DsQdLapy
QoLQXKxhEIq6Anz923QkijUnVjPtWTQKURBu7sYzhhj5b9KOES5IaKJHXSo9Rm9BkMVG7eYoy2AC
Ap2noCHhDSrQPWLJdIuZRj81zBgyVDSNJ+5KdsCqqgQx3RRMqVwj8O3j4dqYEtTE2IccfGMboYCX
W2VqwoXG90cAT3pyUwYs9mIPdVybtDdlgPZpIpvLlyK+6tMjipOf5wQ9wzvn1oNznuGjkwmWVjmL
VYpSrIfAn3hLYTZTus2VIcNZULXlSoF1WdbbhTQpZg1MRE4zTdPzW+DBs1O4y2UPUCAnqRiW9ENJ
Td63DuG+s33BRErKucTcxTL61uKLMt1PA/Ley/WMxnbT81Sd2KqJ5tu+QI1m2EK2LQTwS83oJgGn
yFyWvEb7SSeOanYLcqS9HBU3FhKrit/qwwYRr+pHHXNsg45tMTpXWohq4hsIIBy1xPTy5+3QLiQY
NvTgyiW1HWEu2WEVFe1rUTnQWr37+05bzJb8MATMf8CheQnNFtAa9YQN3wpSFcrVGCRe7LDX2hlO
qvcXKiM2tqxsdyZ3WHq1WoEBETaqyyyJnaCFZ3DqhctOw29319qouu6JZ0cPHHTU2qeXd3Ib3PPV
Mu3j05fM2yM5b8KKXzLyrnZfffMBjV/qK9m9sLHbc7kqoNY4FHE2lXb8gKMBveETKt5AFFK3TymT
Kh61uSoRtKrWBenbTXWkQhWKz4CM6KTZO5KGA/IQJRaBEn06nDCbzdbJsrk1eIDTiAJundypKXfE
+LMEnyAuUg8r3jt6Wr3bwqPZBwc9KlOIvNqtHDLLW1nXFfKdNT5M5TjoquVdx4KEJ4YZK2U7/57V
U574+D42hR1Xfpx/SlyPjIHMdaD7x32dcFVOGagiZBrfXD53uP9Kd4qmSbw4VpQbvm7vn7u51Xkn
mNSJw4F9+eFusb0Bi4et/uQWMJhLRl3KK5csUw1zsAbjm+9M5EHDEdneXOn8/sUx8FACya49Jcym
uVDb5ulA7bpxnKEo3n1V2jxOme7MuvTm2PwIoNqNKabaPR+qae6gPLQ5+voc1xwfBNBN0Zlj8SCY
KpmgtB3MyboOM1yIVnqr4FtU0M2HtBGMy9Hwra0cww0PHGltRvIep4yoMFMyKZXIy/YkRTWhtpiw
qxnHKlRP6OUfdCqDYXqh73bIW4ygKTMlYBb46h2MInMCqS1xa18tO2xgtK2BlODjcl7xEGQdvUvp
GUa38x9A9uMV2GnAy7ZJihGy1xot/pDopSTZJpZSeoE8pHHoYQ9nMrm/t9U7udenYL/kEC77ezg5
1S289dGzlW/Fwj8j66kUNhafr3x5hZyM6BSTN89Jpex/9G+cPZdEnnf5jvAQV0oykWq7eRDrf4rV
1QrX1+BESJgIleYVQnKzNucCfT+2ALEWG244D+KzCbD/sA76sDonVNqH24Mosfi2QuW4qgVyZKG2
bs/2BON6m0YhwpziPXgY3pX0rJBW8EdURXCyM/MZgfTcbXmwf8rA1DKGZvimywWbHFt0jCYz8+hi
sHXpVWyZ9K/ndV2/CBaYrr10ILBR3z3beHJe4reMJvVMwZvXRd3gV8ZwdGkwsCQLkJ+drZu0UcUQ
jp65oBoVb2k3abm7TcLjyX3Vc2dSmo2j3HL8z+8dl9UhFqYOHGv0ul1/zStiRt9lnTiuGXbXQXZ7
Akfi7/xIZR/25z1ednmufP9OkWtlEs1oHfHV+AsBa+TiPSm89indXB0Z86aRztohlxzbaKV93dXI
6nWc4Fbppdb8PF2nEGVyXCNU6KSNGL+uWVu9JqbSuUI4Yhjz1wTFb7Ef3FJLUfNLk/JQfgX0Z8bP
QHqzkG8IzUJCDHy7z6vbkGO+z4GKBRiBJ/no87kibkxg/T7RZgPmXZsh56c0t9slbavdDMdzDSzH
+lar//OjfGG7QJdKP2gRSPRkxqWUVLtjQnGLLOlHzB6gx5bPixTLxrYuSnmbxVXbt/Yj9SQumP0h
NZHKin+JM3xKsxhZ0lIQM1U0TI8q9D2U85uhHn5HUXg0u5x2l8i1E7fmCTKKz/MzXUtwt5AoX2ez
RMo/g3l91fAD6gCCkRVTWDpJa3L4G4TwqLjy6q+q8oz9pdy5xPCT0AGKJVPbxUJ+iYnNCTZFTDC6
SZ3umII1BFIcchJN7FXGT3EReDNeT3EHFsRJJD+YOqQ49uA60tekq2fa3jOArXkBaK3/vKSX72hY
XFzUk9mx1BV6evB45FjHCjD27Vu6PlmixOwvEtE0Ml4gVMcwySRCpbZRnhhDohN7bhqZAn3/DV4B
D4dwIpo5f+Yge4d4pd5lH5YGr24X2fQkohrHFh1YZCh9gZGbBIRaiOOJzNDT2MZVK0Ed0pGoSPJr
SFRlPqfq53oXTsrVP1bRscxAl+S2z0OmpiVbLO9dIADrp3eTbZo1vR+WQfiNfadr2g17rYQ+Zpn6
gLIkJv25BcVUvjsvVF4hr5MhzisI3DwOWGXMLBmz41Z8iYPBdy1TlLAJliRQUqAkLetwQzAEh/P0
O4e664QsxJTAjpWmVPvBdLus4PV40ZE+JSOsQ3SAzx4lFJUH026w/TKcoRgTeri2w4vLz/qmLmhr
Lcil/EqAJm2/Q6aGQMDqW729LBN+31/MZomV4q0dmCRXSpfXlRsYD9/+3YGecng9JIltYEaK2Q4/
6LykgbfDcrQGnVJOf6zuycvNEply+moAip6Pm0qzJeLGMQ4h3cORD9ajrBXPaVSOY2htqPg2eth0
dFDgadNFOKnwm3b2R2RZgWk3CXdcwCchxiR6CP3MrW4K35Zwf8lJLyK3JClZQXE47yjU+o5u972s
vvZQs6KkX8zs4dI30Q5hQAiyJc77D47JsxP5kR96EHnA2dwRL/Ef2Jhz7mK1RKd7ixN1n9XQ4Bgj
TowoSLQgycZhSF/JVA2sZVa5rbhsfRU0fHPmNcLsj9CLC5QYoRUc8ay/pBlzodMTT3HpRQUjQs7u
iVl4KC6JBYr+8MbUkjzaGjSAJ8qfS9jALTg12Qfk+HCkpic9uhiXJfwV7Kwr1LHA0W5rrckRGM5e
6FUckbEohBXNp8WVCgYb5T0YPoUIHt7HGKRPFy+0uw5JDK+rJjrlF01p9pxyB4za6+wF8yaQdrB3
lC0mvHFBDYETqWoF4CA3mSyzX3tqk2zjE2yedGG7hKCw6pl+zMK+Yx1NkiTMZ1D1ifa824lLKBoC
74oRykzENd5Q+zjVq53o71Rg62WjpWWhOxM2/xsuGmj9o1DCALfDYHIiNpdGJfKAmDUNM7RDrhY9
BiCGd+yqUyTn/TxpVydVfZcUSi95gMweCwff7l9S7CnbrIn3w+5Su6ef19XY0zTgrEPr1b1VAL2f
LWj4q9OI43qb3PLw7fHZG6r3hBJ4XJRk3GfIEotEKAoGkiFPjaIAgkQBQjCuDX1/0UdzP9oWUQVn
/karZ4CgGw1YHF/AzgOMeiysPugsAzHAlRXulFCUB2SZNTG7P1WKpij8YLnQEphhlYMdIJftA8ku
95KZHKREkyW+a78r3rmRH4diD3qODCpWtzdFZiBXjgEG9832YB9Eg73nFR7wd2cLATvWJzIHfZxZ
3CpekJSoL8LdAnTgYyy976ezp03VU3UiCY+28LQfPIOmDfmp7jiYkURVXYxSUecDeQ0yViJDb5wM
VxeQVRBacF8kGN5iNPOVxMgFUxBQLqPZcKQIuZc+U/ptWIhwO8TEIgrTXlhYXLacierxfjg5qXcE
7JLCyyGR4zSl/YMuIzBnm0CQUu/nnVithI94AXYPbNXkVD06fXHpoKu5v0sSOZUtT0TY178H1Q/L
KWlxZHX3Wtdd53h2GQgIMkuh2cMF+p5Oskvcb97TeIJPDLFqDYaWrH0x9dAl2+BdXn5RkOk0W99L
lmSLciDjPiHwAnCC7/bPZCxg061JqyHHR/W98onU7HYGQOuwdmFI++luOeQn9iai8qUedikKyyJg
FE8sTZEPKF8UlCMRhf+GnuAR1BcNQYjUY+L3fmSIiGj3Aupa++N9GErFcV6i+8DU4uiwY3oIWDqk
TbcYvki85fekChStkalFv2zMqdlI0EBQ0hAmmb46WyLcyeCduXR42QCdSmCfI76kP4lOgSfZfGrQ
y2CLqy2x4VvIbxoX/RiL+ZYgEEX7du7vD5kp59gfMBR1jcxYh2EWW+CPAjXSPn5QuaIuYfWoU4sS
RjlcXiPHGRvVuUkwjxPwjnnmKwtp6IrSdiSIXrqAs/wtvIpeaqmtfT4E1GzcZyUWT7FR/yT0Tpxw
ck5+yAp/1cKPENOxBu+u+JkkXQOqsddiCMlmDXcugUwiW6H5cFdFdWeMR5GuwaCrL5fr9uV2+jAa
hBcrNsPCKpcY69Ea3LjEzIyq3lxwCgj1N45ayjS9PH6sDjQD2nmE6wNlvRJbUWqNCnP3v7MCdVTi
0EaNiNQr2sF1yscSP1D9OJVRnhUr+6mwvXpaHKi7VTm3jr5i/I/hXff0ncr2Zny3+UKouq/qJWkQ
HvRB+IliYQpOUU9samLA61vSJotXxdMyl4ysvT3uAum+KTEfGSYYyk79d7ntSifL0yM+0/t0+j4E
z6KoIbhXOso9whRqg67QHOCh7/Zrx4kjqiPAzY1QZ7YuvknOI7Uah3kfS3PuPmEfvucaovhDhxXX
nbcUCTsCXdW4kwh1lC/0DSnR3q9VqdCt9ZoyNxHktGJhZFFwSKUxIp3OW1bMEpJMpWpaCGY9bw7C
strz2bbdsIJuKoHXDINOJUB1SL6Kpm1yNZNiLA5rgyKOT8Cqm3yYlWEX/OIjSk9QplbXx3RrD8ux
swllxCy+QtDxmINGAwmTvzDxidL/Onj5/FntXb8HUxRzbKKiiCLEcPK5l9DerrQNcV9w8+iBjbGo
8wVkTEYSP4kDLtgp4dcOWXUTM0uP2Sb/jH0hCBwozgXM2TTdOBJznQycSUtolE03p9AiI18sAtpX
VasTDKhxigxYpiOMuQ4Yfi5xr2REx2wW5QF40z9jDlHiwBsfPMGK1RKGC4MgGtlcYdYjCb6T7QF/
nUcYayfpbp3ZgahJuJm8/n3AYugpT6Zj56s6PY29j6FxwpDzTximlSJOic+vhaARv/G2LpDLEjtE
zeOb7xG028rLZGEnTyUEIdDE6JGF2W32pujI1RMakxpSnftE+7Shm8QDj+/xG7O7U7Wm4pv/eMPq
AoSkcJuN4d0qOSIFv3UsApiuNifDyJuH3j47bcG60pxneJW6Lzd90TedxkCSmbMmDydnI4oF8QBs
Q8qkPLZepC4joQS7VJamMWeGOaHBHbpTs2CaSpQM+EU55tqXPmnxvCul8o2DcSOdvo8PYGJ65pq3
VPi4PuDAw3CiIuHvBi9F5KLmWoQSG7mf1CIqbUbQe4U+/oEmWCWhkkgvPKK10hKf/SanxC8aQW/H
stGDhGyGVhYs/VYWrm+D4mGjmF2SKisLF5FujnoJ8GkdBDnjSRbZlg7AeIeAto14UYWrjmMjXCEZ
cL25okawKHD0Azo6C7+692CTORGFeWq/94vmD0QOlm7dNyZ5EZeZpSHRO3ioruRUMRg2C7PUBsSR
YnB+cvH1o7p7Rd5S4D7kdNnYaoN+4plg6RXoffAlR+fPs9oCtyABPfO+Z5N6uptMKs2S8gf5flf/
NE/9SOWBip8rwUkJj2i1Tlyqxy4x3cCU0sS3hMFQA87kzzQyHka61OBXPT2cG2UkGY/OW2vO4oQO
6wGpF7BUKEoF+CmY0c5RsAECgyIEoZk5jrFJdhOsi8p6pwH3oNs3tcVZM4ZTkD4X1qBalw7Mk1CA
QgQ17rdlNTNXv2PvlJO8fAx3WiOllbgZJhDrVdZUTrlR2geFdX6AE20yWV2x6P8VFvbWxl7uY7K6
f+dcPNSrKBpfq9wZXdo46UM9m9R1pYi+zLNYt5LVDGpupTcWo0W/bPbqnSsvaJhHdlYUM7GsBUr9
Snajxtu/aN38YhcIZJ9PGqpiIskBuyg7JcsZjGmUgwbgcKSGdkXXV1B0XOvtD5OMLxyBuMTpxCQO
N2IG8QmmtrIOuqvKRIFbtD0a2Ahc1YAkbDlzDNjIJ/W2FtPQ3mTLZonq17r6Hz0Hv0IUloW2wRcU
f9/YoLHSZ8ZeVEyWRcVBXOO7IuH9CaP82rzgLuhc69ag+KiUuUeyYGP/LsKZzGxQGWbHPWTYljiC
ytSQNFFJ4npUrvKFXygOHc0FkVqfJOGooe0DjDLG7XkMir5qNPOhRo1TreAot7Wl+EZcZyLuog5g
uzhM1WcszpWDcCHZAjcrdchNkvCWNucx9ELIqeCO/g1lP8lKyBWNhqrkWVx8lRf88lWkSqFE8M4T
PP0jXGSz5ajH8FuRyA8JL4gey17P01MtV8z6gm+2cuLX0rBnbPJDMr8jopwDkdFkeGATVVxk3yUs
r0J4RT1pQDyL06cpT+mOf0JMhB2MlIRGwSjD9qiMp/lB47RDL4DuckL5d1TYtdpKuMmd9EOpep5Y
mqF0tS6Fp/G1cfzuHnnbNy5dLOkXxUjZWGVmqUZl09+pyblhaqhfo9NjbVeTpP2pGSTlELNwNuKP
V48mp3CYZJmF0R97QkGeP5Bi05Tab47LA5OE7m6BS8OF4WP0BKeTfwgyBW+RIrHgXoESyfc598YO
nnIZz9HPvYtTj+eC2vVua6iTUCsgCa4jX/e7GAaLw6LlIpGM0YgSc15ZWsDAf4XWtU9h5T4eD5SJ
vzZXt9u/I8mjO9PEp+gvejXkszQkuLCzXaH+qfYkV96hmgNFh68qZwSYp8qgP5+fMrbwFo7wBob7
3897pGUAS6TMK1YJAQ0g+55uPRhqEHW1JPCPb6nuKxsjaV2YmVF9W3MCI/sg2F912XK53NJXYNEm
CtPZox185mSa/VoOwiIZ1KwpNo8SLfB4+8F3WTOAHFgY8BHNC02ojRAFkzWUeDIU5zqgtcMFLxVq
IbeS64RNhwjENqm5/+mzkVmhS5UY4D0czJ23ILrP6LseNYca/1/p/czjgtLTXS0SaxwUPmrk5MyV
VbZNPIVv1dvLVVaVmnFG36gTL41gpjr66y0ZI3o8qC13KSPR7aju3u2MvxS5SQct0t/s3+Y8/5hM
yCHzxOtEx/VE8grghRzHXQvbczmGdTcBsMZ7+2/SQUhMWRL5ThDOHh2Mo6wmRL+16gWBEDSfaU/b
NITdjjx1C76SuRemSncYNHNfXs4CYK9KkGtPBG5OWwX5YfzmFNLqi0SCb2sRvNyUIJipwjLgVVA6
GXzf9qAnWCVzNzHqPiTKGCKEEqiSWbV3qxxxoQEQieRDn4jnFH3/L3UrqYZD0MlsD58Av5DgzO32
mc2kjGJ3LBW/HAYiWS0DkWrNUfXO0iTr/rbojx0N7IOTr7Tkta6jaUyD5UocuyfCoWU08iSCb/M7
Buhmrat+H0TXsbLQIC/ICEggHR7YhABiIzPy4zsbIRJKPvNqWb77rBPF/+ayJWbMvoUYZJDAWjoy
dpfFWTzaxs8OddnQ0u5wCMPXNfUcVoHuYribAdUPjm/PL6mGA8Q5l80JvitSxVWUDHJpgHc1dRaS
2l6WZX3NTAGcGfBli+ny0CpdPgijlCB69LI8xqSmjmbFToE2GfuSHrmvXqFElEk9e7bqQQYnsMtG
ZIMnHevYWdKrQZvsusljMBnGNAdiHNZFMLTCZf6jijQMdtOFdD6B9L6zBcOyOF88LKx9IGz5XbeM
JHj/x6HZzGX1JXN2DVqf9dgsHsmSKRpDEKQCZOT+mZT8IKrRqz7FoY1bD5XAqZy3lIgQhuyJV5Cq
nX/pWuR38OgGPdJjEcdD+a82xyYyPPYGePsilYHQyU6wtbwst0KaneMNqp8QJbOAl3bGJcNY3X+C
8HRnCmas7kV6TLKqf0r6mGr/Icoho+ydkOT7SlJgHX7IOddIWPELzeSkwQCGSBqdilGOUlGfph8W
JeiNIOtEVL/Mm10nFk1NqYnZX7/YzbLRcpdOtvVGfL6kKEfDnrCF39BaXluPXJqjvFMPOInTL8xM
gJ0ovYrLiI2bjDy1v+OEfOV9rVwatrRhLJUqeKkDK+SFw92pjS137ujP9rFJT6euF8fUuveEQOfB
LG0PZcGcE0vijag75GYoxwDbAi8XjPEwUjT4kCYuaBtXUNfos2AhCDUxQHWDVoDsQsqJbmwUV+4y
Y0SRFfKcUVomBea4O4XzpyDjc3KgKHPSMUZuhPHrzruz+GcXnLrV6vgwPI8vdZAw9BKTxwGJwHAy
szbUA30cp3Ht4WnKH9w1Xrx54Shj9t38OHeVYGv0Q2vdxSmsuCcIM4ukurbSyWhBJMsjgbLMjs9l
JnkUyewF0bVn0IkS1dxeafhkwtNXXssJ2DEmuDNUEFNTvCRsClDYIJdX1UnHPorKpcbdvv/BAeBU
cRK17x1rJm0PLjXtCSh7hj/i0OI0abPq8CnejjWugca60dkkShqDz+nU9RzqnIoAyAKHmG8Fa8Mu
6nj4eLdBpLcVa94LEJa4xPt+tegPc9GYuV585pI2+kbW8QNIapxtCkNC7NbliswcGwiQ8HWevJex
RvzuBQybN9ucku027Clj4BNxvWrNSp98GIgq5W3cszcG75c5bxsIQ3ynm8dwc5MhPLwdBNuSnnHA
RM+JoHEuOyOL+FI0vfXz7KzKR9GunRM4YWtmeKmAKBisNZ80pzcDTvAWx/JcBu32tAsbv5VEAdxQ
vX06OANaNvYO7qiX4NQQCNTJL2tWhcfLeX76wMXT8dYX5Gvg55AjbtkyGAW/9X8Z4OgdNyRozdtx
/YVuBvPU8j29boeBkK+9ZTREW9VcxYCaoIdxnPLXb7UO0Ohm3zdRcgbsRBUosMkQ7OeGeYsHK1Yh
3j1dm2zslletqC5fCdtyuE6V1zeI1IpTn0qeMcQfUX3VxBloP2xyNTp7wt66WAOR9qJC85HrTOve
jfQPdCfJndy8fTTw/ut9Sd5yOobpOuVM+ShS/wmL1boaY7U7q2PZdy4vk1QvUzXCkSiAbxvkvPsd
cQWFBvxfqpXEWWsWNLToIJQWDTZwNmUhxwHfDAUdj+XZqdmRCZfXPx8hgYERHePWB3hyvT3Z6g6o
pykkfDviyNKgkqzHsAo8r1gJejp0avoHGhB6KIxj+xmYKd7CCFHU0SDfw36DOOzZDm2OlzquHI3k
D+ZnCmCQ2KxlhdL9aEuEGQqhspLKL7H+jixBcgV3jwU/9Xs4CPbkKs+YCOK6WS62iC7b8veQkhVz
v5bFPa943JhGi+FKQ3Jp1dRd9DC22JPCfNKRA0jVq8ITlDwnvPg0TpPohZpE9H5Fw6N3+PAeeBpC
jkoPtKmQ62qqRbDHl2S2ID1hN5WPixo0LP+YdwRg9Wvb0VxP+++2ky9oAeNADoAY5fe7UYslsOCv
49CdRlYdVoQa0ZRR7ZT43C0PHlSTmCnpsDblkYy85OY6gM/57kk3pXnKJnO/U90Et+ctyC8CNA1w
K8tb4g+nu60wZLVeGTWUMAKi8WcE6s8g5lWCBixugI1mSSfiT4Obimjud+ZhuLzwkDKEsCWAzL4X
RC62UcFjGTJUZPo2Kv3YJ75QEPugmX1RCCIWj9qrVbvcV+qZFvzDNUsBQ4kN86PWYLmIyI/BFhe2
mK04wQNDDcIWPOboqkWBMcxeFohTemuCIZqj8JtdIXgGq8xjzKPUu25u/d4PHjeksMRfuLHT81vr
bPxV0pEd5eQ09sd0fLJuW0oAilEa79F7Nc6f2+Ig+/LnD0zNBt//26SPogjQZMp46iDtKGc+o2BM
3KslWOImIWMZVjysQEmCwhQcvwmhYGhhn8s5hT2/QZ+Egz5SV4ZSmt5Vv0IK50EDVYnOKee/Tq7o
/zlvOUMMm67e4gIUsshX94rh/5PKeIkt4Cq0xwYsoj7PtQ24HzEWC31LLpy41yfT3KgY4vAVSg2x
48Zv+ugAf/+6zaiZIj9UQbKYadE8CBZDr9mwd8VXFiimFyx0kUx7dVPYgDxxDP/C9+FrogKMBnFy
NWZSGt0AAe9lV0edcQtHHnerYBItEg23MdyxXWz2LxCwq5F5/nFbiiIL1Bxa7AtelqBi4FwUngel
5FbwmmQfrfzhFvPFXxo10SFqfBL8VdND+ixpm9RUFy6u+ll++JIWw4kg4R9YnjWeEiTeIvAgYLmH
cxV8y0NOx7v4/MrKFYDukIBqR9cVNyZJcPVm0oR1MWymdvjyb112uxyDgENBFQATB3omiLrqrDyI
Ifjl3TCaT9qk4Q+JBEQBqo/MsNoNBMuo2mAIy321Sw3Sxk8hmW2uPs34MIFXpI02Rk/f43Bv0WCv
GXWfea7SRspTycyOlEdfJ3VzxhzJLfLaGg5zByDNcB5ZHvh5l9NINROnnYFSC98zuM/Zf0Gc1rbM
roHDbvIIGtpjTXM+dbZDYDDzWpb2rf0kHCRjOK1Zb3QoUHwMfXPRlpFQXS6JGKTW8Xo5b+w7fFko
CBWNiB4Hwbvx5uzLFIyC87i/Lft5ek+eaadh7Bmg2Xr8nPzujHGIi8HdnCZFZg5dTdrBkxlo2FjK
FgttDc6a5HdVRv5Btl4eJ/M0khk4jVCRlp/9l0dTAF1XcCQFyDfU43ybU0wNRBZlXe+1w1nH/22N
N6wxU9t2TWm3UbJB3PB+V1zCv8lF3hV6Gybrc92bj5oATMgVSQFK/kE3SOSMiD17+RmKCd2VnezE
qsrxUdXibjXUAO3Uh7niUa2rQgG3K46ciIp0dUOll8y7kC1BzVhkeonvnuSlvcmGY+6tvCVS0M10
FrM0FXwGEqdxASqpUMKlSkFoTa9xPZ20Zg3R8+IuE3rymBtmLimYbTiIv95caJJcR2FXc+Zcp2x1
2HzN4ifqJKEhYaK+Yz+goaAYduE9HN/HmG1J7/39a0XRonImVDh1n+8Sic1ReltVdsVLNoyH6947
/u0WcbqS4OukPwy/npP+d46HHGBnmaro9C7b52x1wp6BqFH6jd8r4JPiHwFwsCgMhsRYzOoHRzJo
m4sNqcYQfDxAHNlfhbnRjYIQ6evIpkduHJGojm7XrvZdvv+ICi5p7a/qw5ANiphe5ryHtWYKLUjG
HZLhemBzV0nSiUZOi3WTMDT2m/AvLhfzXD3wrogLvAopWjLtAMTN7oGl6d+JaqnzvXC4GPqGGVFj
+vQpbPZ/zrvtNZ2Z/sFC5EC4OYCMpp29YrPu+/Ef0oBYYpAvWAsmXv1RHV7CzC9gMLtV5YAu6JUr
aZGE4X4ZAZUasNERmeHOkUus5xTNFFhF5VD4RGl3/EuhC2NnuCfIqI/StAHP6atZXP5/qMi6rMZx
vPngbGl33n+svPciw41WmiSz9Orgw7OB8KRZJnnNUzPy+/t8BTv++JAsfxn8H+VDt9Hx6i2jL/t7
jN58uLF9Xp+BXHHyBSZXbo9xDBrItrSmFkQcUk7bVucJS8ZGbbsuNvQIuQUxz3+GQeqZKUjuHxNv
e+p2qlvpFv+JIJ2pOEk6tBBy7Swj++4d3l2HIrNw1Mlt/NoZ8FDI81z4Yux4ifoK2DYoxT00JOoo
4xgddKIhj4Att6k8Ek/aFdHk80ZdJK53Ydh6s9TLwBonReUS01touAUcRDb5d/nNCCSuijqi44fU
dXxWTqPxGO7p1XHKP8f9q3fVrDum0iSeyhs9OFU1H8vxs+4qX71s6MBmqvZjyYktflgiJfji4AMq
dbiINjo0A+rqKz0GZVh+nQyp6ObHR2kYIjYLHMqyh8DPS5mezfr5VrCLM1NB7HzWeEsCBK8ynXbs
6Xva8VxzPC4rhgDZC8cMPQeENnJ2m/Da+9Y8uqP9592JNv6F0wLobD+qhyf8y1K4Sr1whvF1X1G6
n+w2J5a4OTDjd15Vey+wBUC9z5j3mUHHceBm6X0iB3XNhvOFkkQ7NrUgE/wMDkCiUmVezmLABHaB
2g+kI6tE233UiD/AvB96rhJyKeDg6VptEIOa4maBAfbZKeMIQUgnXi1bpUvHGSKeDwq7jzTGNcUP
RjhAvE/f8bv1lEU3JJI262WYPmpO6Md1YsvJg2nOJZ9b+EJlR89+nBnwcY7EV9B2T0G8ezfVM+4j
2QKUdR1Ww9fv3IfE8JDhu74LK2MqUZqgqQkx1Pwm+lgrgwcMm7HV3FEvDjlDGwPrPzNLHdNFdmRk
hkDl/DOb7UosP5n3cwTg47tpEpMTu3/BZa6NA5TysLXCEXsa2h6z5bvl+Q5XiDvo06XB5O4yLqiE
jWBDnyQBbaNbJL9/xHFi64maQlfZpbnXho2Al+CguB5NtBbe/8kRSzCJ2DMDqpEkjfMBLF0+eJ/X
DsxqDTYrb51PETIr45i80B979chi6d2KYeGayLXjl4HFW03rGMxKJdiVcVKq2LqzVdZW2rpKC807
XwsBopxMfQx98xAFPIuD7pZYNozM8n6zljqO3cGtGPOeU2ZDb4jbOKbl+pHHk0e2rZFwsFyJ5pEo
42PlMJgvPdBX0XLMDMndGbFAvlHregdjOhV2xf79j8CumjPgd3IZrgJIaVXdJJccnQ1YzKU9oGXP
UQT8yo5ci9H5CmQSpIwztTjEd9XO+HCkp1/KeYC/nA2INQyidL9h3si/ZNCE6ZH8GFosAyLhNEPD
uGaQl0rcfvGZZhOuKxel5ng5waRY3p5Mq1buyocOu9UPaS4sIRFOsJvJzHhuuQ3vjl8KVtBo/491
IaH6rcJNJsacQCAslfHCMn1EB0HpjNAWKT4e3JFafRNjFzjJhUmp69CpPzt4n8yAsY01g1DhEdEC
27MnJLqKoH4sNHVgeaQh2j9UU0SgmeYRiGaT+dWFTfm4wMk4riv7MIkVpz28KutnXmpAbY5mOhuZ
eTNFVPh1erZ8T0rUwo0+4wyPv5AgszqruqHc5Txtk66t7bNWD/tWE6iZwqQVDEd5KMovrNCOXGgw
KXILhw58i4rWFAM5k4A6GLMXlb+JTCRf/F3dyJGR4dBo4kXEcLPhKktNKkVFye4cayOgnsN4A6VC
E0aQGMVNHjjPND3cdVGJGPPNse3drrKs2lYJ9IjD+0iuz1+TrHQ04Nr3TYvCcCCHmID5/Ikkgoqp
pnD+34mPD2sSBxWrqFmFe9Rr07kPBAh8s3+zlNfQqewqtQcO4Mr3FtLV2Q5TYyhiIKFN3E3ZN+DU
8n2RIpkz3Bz2EHEIWktWGrwkw1xUH8p7g9ThoirfKx08a853u94tDkPD+jWhgoyUPrb93NZILufD
87k11wfj6X6AS2twIdYWsfeZU3Y2VhhX2TSJ4bD00HarNe/jPbzZF2y4+d/lQw8SM/27kU0mJ2Qu
fmYaUX8mAlV+iXobk+Xh/ZFyXwCL7o7L5VrA7o8DNJdvgEoRp/Qy7aacmv5m0bg6u4RZFC44jC2P
nadR7ySGcJRzEeu06XyDLJJrunseHmVGVaBUOey8wC54re2qQaf/V9nJ0zrKzsnLTTOz5WOHEjBe
ZXX4sVlyNO/7LeGx6fphx4EGQHnopuv2NUEio/kUGJE4sIfrnV5W2jKOKAYwiC8I/dv29uvrCjV9
y/WvhERsDzmQTCuY2nWbwG4jETSV7Di2QgBU0D0dibMWsFa7XlTmH9DmcdKk/XtjKbYcyPY1edhB
d+rRrFHp0drBQhCDRMUepa6GATQyvCP4vNlwWUH9cMN24OTpxsxvE6bqnbAWkfQQHumoZn9yu4CL
eXkvqtZ65dwvC2zOBNBGGk+QY4A5hiczuDDYlpAgYNlnBk92sm5MkR5Ow6TCDOSY0AEJNdyz6IJe
9sdu/Z6hLqm/BWFq0+orCbVQ0+6YnIdQ1s6Xwpc0hvrGtN7t0b7SAwB23gV/2rbi9gQgo7sRuNTg
jxm7ZpucFD1+IM4pqWpamref2+hZVHGBj8n4ikCY26TAUBEuE7igMIrNmnChY5c1Du24vOZPqoiS
XZY286+3BKYheTtN99bKsB4ZQEPeIDDatn0GCPL4ZtYIueuuBp04JrMmBhdwK+37Jzj/kkNzfg2s
U1TDEfLUBPxJH6NsbWGB49J8JDEPqaB1Jhj5LPh5uBPYyaAx8RTszp1iWGR79nzwyiP0dBEacSzz
eVfpFISeve/TXA9xleRwksQywSeN3IPHkdR6y5aLZW2ZPXHFDu/TWwwiXkrwGMF9WTuFmFXtticW
Zd7qDCRMx86AIt2pX3/FCBn3wGyRaZtupkzujHgUryWN/mHCDwZu27vsLxObYQkfzP3Y3Kqo8ttB
Md6TlixD8D80qGQ6sZiuvq96vJ/tRjP+w+7E2bL/k7X7k/oXm1gqKl2jH19IaswWWEyKO3HQXkkH
IuUs1yJkayMWVLcMT0/xcbkKui2O0lbj+gLQ36dio6uROwetrgkWTN1qKxF9oxcRz48n8TIeK6oI
WTj+6gN/Q2+GZ2Q2TwjPyZa6Dub16QJPrY4umQL8vNZx/QDjMEjICzk9oapRSLD2KCvXKno0AR2L
f0Q1Tfexo4Ar4eIInRuE8N0OERuoVj4CNMfKFOmsuQZAp2MFrzeslM4B3oYoz0eFZFB8vCHA1ZLa
QL38VeL5U67UF3Wb4ZU/YZgGM80ckDJSEE0zO/luhu+SF9gK5f0wPaLgGtcfgtkNv/Zw8j19gMEt
jHy8yJtvAcgObgoJ/9Zu2N3WP8geG/il05kmonHPHfbOyjnbUMsFDFeS5/6V25DwiF4R2/CtP/DA
KU2N+qhT0VP++Sn3jfw9DvPAcPhk7wLsI3s1qcjxOofxAhaOZFu1ULvNw2LBmyAtE7oSnRxOSQN2
/8RGFKNAxzSHGyRlGtbDc7AwlbcFgjUESs+f52vosv14GQgixG4U7NX/L6IyvIhyZoJdbYS03f/y
lG6aqBOjOw+aCN2ZHTsWjQPfW27Pm3p35GBfoZ6YswA3JY7zzmzhwLVSSY9UADEkHkCeVyZ1b1bJ
WDKInjqhafaWC/XLwehf6WU4rcziNS6Kq8kFnXamJH/ww0nQWCiUbnOW5Fx7nwK9rpyjTj0c7nRt
UexUg5xYy9QHVGdkUOK1WiaI+L9Eyzyfmn1yT16NQKenoNRp+nTjNwHco9WblpLtN7wuJokKTmFN
ofjzirpWnxsw1huhWZ1sHW85AcSZ0hCHBaYgidVJ9fAcP+A90vD9gdx7TWx3FXrJw9Yi5IMH7jFA
twYRjH4RMs82fuj0tTLJsGXhZyQgRCSxBpRplaOScc6NnHc9FpzgoRQ0LaGbKMHeMu9+D0sI4M5M
U3Mih2+xo6aZbr6JJoXBz5HKO7B682rXD3S8TOkWDJGA94IE2rQo2Q0xxvsfEq+AjATZ+GhlfhYH
ZgHKm8G+Z3OM2UJo4IcjEqc/OsSpOEXt5MfEu3JwDvo2+QE4v4GOCQBDxCz00sTH1tkMcN0rxo6E
xQWLPoUMNUoQLSminRYIfkTTXzUakslsT6wZh5QT4CLGKroLKbDjvzPKBt+aC4+uiwmytaER0Zuf
7EEHS6Hg4CblltqMLhPg2hl3MpQ9A45n6SF27Wi/KzCVTwHB6OLCB0ZcwfC7X/nXY6W1FlzCSEAF
ERvs69pYnYokGLjUJjFj42oteeDCPdlHL2JyApqhP7fT6W6Ye1UZtQFRNVx38foGZ9dDHx9yQxMC
TH78Q2qBVqKaR5Ik7MG15euP3Kcvm1IlafxITfA1Mf5zj+1SjeLW24KU1kd1lv6nlvr1+QslFwEJ
DulZbma49u3zUWh2yWO+oUuHaoH1utdzMjE3EzC7BtFt5c/AG/yMSABJE9cBU4aO0wobQG9D8ppc
8WzYJkt8fc86S0ujWtyavuELtjtW5nQYTFOFPqcarbCLG9Jj7QHpaIlXbP1idCpH5Nvh37qm75db
Uc4GCnNcrvWzVAztD/wcOAoiUkUHV9iR5BP/4Vj7pBDWqDQlEDpG+x1DRULXyVuUNyg8UvjUqGVa
H0HnGIons40kZqgY+PZrZVC8XPS0DUEEycEwTdPmQxDpl8qsX50OwwqTLzTvVpV6lwPCDzizF5I+
L4v2i0RcZ5C+wBHLn55WKV8Jzc7qIMCdjI6HEVxi/0ojo+n+yfu90BQB0V574KdXfdlLxbw2D8Q/
PwAniLT0PsXvM5E+Aqly/k0FWkKoIhHl8AggDergysKYFSJICul0HKki2cVgOxjyKEJNpWL3AcDe
k4sSYtnijX3iQYGnY3btmtkRXNDsPFTApq5VIQhU/PJuZykHt1s2BbR1aO/ka5dk+YDXLPrdtzpy
W09PfHi+yrA+2rRxPdiGDxH250yF3JoGM/vcMiPd+azvTelu5cChnoSGn1kyhwmGtYXZW5Jd/JRF
eSvgTYil8tO+axjmQuMz1SeMGIeiAQlwgvgq/mMHm/CPPJOP3gTJg+vRgUVapxybpO0+mProhdKs
35lZGqCCQM2hTx0MZ6pCDoCREtqh839ZvyGtZE40jkd9HPoUnIAhOxPGEbtbY+3B/ODxKRBbAcPH
+oEtFwQVRAn8O8nJYBgPucxS+ieKVxVaCn5Mulfl9pY51xTEdLclAHqYl/k9eCzst3m68pDu+Zxk
5myQyZrB4corgbc0QesjuiT/QYiCswAXWJItdoqih8ROWNxT0/A0g5AW4X4nlQDs4ZnfVzlXb0HD
sVyVyjUrcAbqY0XwsjQHcZ/PfexHn6OyyHOoIFYkrBAis2qbBiJNkwNX64XKKF8Kdtcl96WTJjGZ
gIHnxqIrVjZtrKeO9ej8v+izNa4tq2CBM4M76r51LwSX/v8hlDCgV4AgXYyzfCzsp4i3Wp65IeXl
cS3DyN5/bziGCYAcgxhNJMrDVrP0Ivoom5a2HRQ+m4a2zsDxnkHY0DYZFNAdRcgdBxLu/cCRPF95
bV3y4QlCn+oLRi/Eexz1xk9+HFFsKHYJfNQQJr5Cfo+8n/EpOyox4+T7sL67YlqoMIoBt69mRoP6
VYygNpBaG7Cytq+mhv3I+xx/t7IiGciy2vHaDKWskSFAo9dKUCzWpNS/313UZV5kKtdlARMEyFzs
84+fnIQibzqYUePhiaH4yxfcX4KZLZZUm7YKPH4UM43tVNG1v5TQH3Dfg3cRfgTvzI9Gwq46ogH2
iZo6625MV5JnAvQAjEeGe9gQsZDFf0fe2eHFBH3M2z+MEIPRj1lqR7U03L9wou3qUfq3nBQuWKtu
L39juTsCeq/2rIMLhpwa/wD3Gb8I+0bQzZhqsp5uCEHe+HVRQAx9ILEZEjoDU84XNus/c3juiUqn
p/AQUzqzG2hGJtHPMc7OcQXjZGga1p7VzEQiOpaV06GfEcsHeqbBR/E27F9zyyb+3EvIkJGs/HCO
jKpSyKhcs/lEAD3Nf+Y81qz1L3QyEJK5ceJ/8K5WltBFYYNLlN69xR8GnE5OTtpd6fM7eeC2Sgvj
FkUJnljHUuqHHiTixhXinRrS5HAJ7tW4YA0QZT7nIiW/KyLtlcIPJPT26vDR0EZsOO2mIsdYnxsf
01YEYJigKD6/NpCgS0WgZ6dCFHk3nNwB/Ovuy7tvXA35tZKAW7vlYM2pLOHwwMBpFow1eII+GAcv
G0+/KE088m93x4IYny2kIrZce8LXPNCtlrEiZ0PSu3OLIug5qML8D200dw//fyrK7sPBCwPz9PGb
MA5mH0FoIOqxWwSp2tCwoVk5JDu94380pqb6m8nd/aJHaf1mtUGFhJcQSGX6XjillkpEWrx51mDp
Ap4Tv0WI8O4c94LW86b8qLSsSPXPJ9Za5bZw5Iw31Mpp7FrDz7Gj5PY2c4jCreD7x7/5p/Aanx50
IP7bIu/kdots8XAis+bWftpdGznf/QhOZAuBTgSkU8zLe15D1vYCPf8jYDQwqcuFoxVJbmOe3rp5
GMBUNZEk/X9CNwzPLbVkd61FsKTcURTOA+HGOFGExUyQOehaesjn/p3c8djkM56EZoF7ojzYG9LT
Hn/+63s5Qk2bDFNlu+iE5IuUQtIGfOuDPi7vPNCn8dk7DtM0N/F+epABE9BYh+eCxes9A/cuAeDm
CtoqnvHdOCxLVnGDviIjDc8E2dTOGGeXvaa4c1nxIOqsQ99/G2K+gEH6sIAizsUCqBKWJLYRrAFK
v7hLzgBoRHycuNn6P5gT+09juSLaKTgzKjQPOmkMlhOJ+OC9Rowcoa8wyzWpKQ+NuRZYn9xUyYlX
rFfzeydZ/5Xc0nylB6SV1NgiNPotOmP2zP53lN3fLwNb+fGTaE1ikcExVaU9BU3MI9ZFmkrCm4f6
x7tqZmBFKydIPzRTZdMgF//LT7tG54ZEyISnAiSsnfUfUHvi7teTYq78sHulcAUoWOSPFzqNFHJr
SDaLIlWqiK2uGeBhg2DZzPqykiD321JjpUUtYNuUZC0K/fWYmmkNDoqBVj2FFmRNUBc0mkiC5ySO
SY3ljmVaTOISlktE7W9A5mKHSJMcHPNt8TwMmnNhxremW+IoLR+Sg2fUQwmFu1bkkWMvFx+o9oHc
FK+iOwEHA6Qc6G3RtCxJXLHtdWhlGrCMXT/lbeiG32nBUFXC/0ofap4XSz6iuhH1jKafA6Uf703X
VrR7MOxWTEDHMDrO+iSkrNFJoexx4KbB0XQx1T5e83rtmj75fPkyLze7GtzYJRYjyvsnG3KMk5XQ
xJANbYaUMgwjhv7f0qRnW7gZSHi7o8qeiVSmQM/nQ9/LNC9OKymnJhJ0M31dhIQ997cygLwZyeR6
7rLwmo8NPbreGVfZObcdBQ16V+t1x1mRyMrxmMeDl9lXhYdZj66zMV4X74dbkbfR4rQdIGtE0YDq
aaPllYXpxS0jPpr0fMe/ahFlH3cWz2fWN0wB/bz1T94zap1mBxJcX5ZPB4uBifXD7zQh3Eb0Znq5
5ZqB6qQ6fO6uhkc6cvvs2/dypF419ra3jPZsSHrkKyI0vKuNd4rxvPTzXt5E7xcC/MtMTrbIWtZk
bRvKsF+Y+d4lCdkdGoDFPatvrd4v4cQ+7SZrj8GJrxdbE1mXiXfbhl728vl/10DNbDsUbADSGIbx
KcsjEmwP1q6A1VGElvG27MaR4ilkOIvivKs0SmiqyHwiFBuTcJwqJXwlC2F7YOaVmuAuWfJ71S1L
uabl1URzw+aaaHAKkeacilU8z/rN5Lp3A4Y7YdAQlkL1ISCi04D2P7+v8DBCge+jSLgJsnm06zLp
Pzqpd0Lqy3fd8M9IJi0zY9wbb9Rr1M+dtojpRR+txq/XR6KVSUT3H2Sk19kfQb2T40pXK21Jbs/P
z9GNZHfLOVekVaMHva+BpYYPETX8hxWlgZFzmKGx4b4Fnys0aF0ow/GYgh8Vk2ZRpVtkjKT7sWk4
4sWjt7LE3a73gvhPq6QQw3x+tZzPoxfCsQ+M3kpTveiVAoHX5f5kr+anz11YreWtsfO7rvSpsh68
G6j4klBRWtx3km81G74JuBrFsBgW8LmqIAj3tFaDc8LmKlYZHIUdkS1SW7gZ/LQKp8O78XhrWL7J
VaFGhOV3OJHsUgVUbQZYNIfDhXcvgNHoo4cypukUB4Y0iq2rQezegdHL+RrlJ/og0j8CeqlhRh1o
Lkac7PYiitPsY/onHwlb2Ghl2QMDtHnMPbfzJtzzYbC/bVg+9IeulPgg2RjuJ8HyI2CIE7WUNZdt
efHhkTujsS/8CPZvbq/tO4QoslrH9Fo5Cr2Z/WlFQ9nOjAY4XvtytkzCpGGarg/AjVarc249dFH3
FVNpyPD/qh742X1WPC9f0WjgJVsrEwjiQovD+hKlW1QB5cEtP7xltOWmr09C4FSBWBJlS0KR0qLq
20445ykbo4F/dLI8dHy9JQyeKo/+0Qwwso9/Q1pNIJ+NTpbS+m8s+1FPgq60IDuUFI8no8/FVcne
vdhOwU2NpeFWG82SUi4eyKJifaVX7NSHOhIcgex0iyW67K85y2UFCWGR15nIAstwPKOIc2DXec4m
Rayp/59Za6GKjs1boqYrO3tkjmdpLTafK/zwVYWxMpMiW51uVJ6iGfesMNJyn7QcpTb+ral1FkvB
tlFW4giy9p63b/FceBsIvjEMbdAsMsoeXn1vihHuQxupQVjgG0TY1X6+wXjIWvxwfwgvCto/agzY
0ff+XGT16CzSOh8jYZKGR6TGBb2jAx/0dvEt7+X5Qd3yuLOuvSNNS2buGPY+7K3LVZaAvlCAUHM9
HDE4VnBp05wsGYE+BR7XIFPKky7ujWmXvNTrytQHyRiKNqeeaKofqT+28r1vME1XpTnKhCu/GhLc
MN3GHSOvtKFre5p3w8QmJV43NXwpt0zlbh9Oy6rHUtSIV4CXmADJEpR+iy4Exku7E2pzdlViUVrn
ZvBifEyZ/C6XM5SZ1xetFr3e+Fj6Tr4tDJs58PdqQp014h0wr3xbwaX1XdFgx2qx+bZDKQnVNxCs
C7+GGficFx2k99ohduG0x1ybeheQsayc2s+Tjfb0rdGGxKedCgcGsCmDM4wSf4QNrvzfnj9qKmRG
4ax+EPtJqri1beW+kKwKSHu+AbFErbfuxEBIQbGRKsI8KxVpgl8niwziCLrQLxjyg5GdWgxnon7/
DcMgMxuKx0g+JEhSS89E4O3n/+V78nKGkWo3K0cto/8QTFXbvOcm1ZyQwFWNsUVTwkkBHoL+OUph
/duc7a59SorBpQ5q6e6up3lBWMEnRFCJMkgc5YUNBk0M3m8na6v/Hj6sN7VdWQ8Qf44vDN8aW5EG
o6sQiCvrvomJo/SMCQne2WtKFgl6qYVou143pwGuvodghVrjZGGseGr+YDpZZIzu/XbPIM6GHUlQ
t+5XnThsw/Fr/L7kDk5BerLcMlwySsAdHoluk/Vo/Lt1bRmglDASbDQBMrZGFOloeflywoP6S0S/
1VkExB+CNbVk7ujwdZAEiOridNuV3fR6Ifc4Q3+KFf+pWr6Hf9cj02inDCCApfLE4bPQIyT0IEKy
jvRbUJTGd8LEa1Fkd4An5x+yGev5OGyj9awMECVkFCNavuhB61v0RclIv9PVsO/5AR91xvfKN1wa
xGwy7/KNnfHzypeG+H7XPWDiwbJ2i/uS6j0YW4Hv89Mu5t38/czgAbKBdmYW5i3Qez0gH8xgxrlJ
yOeKKvWwllSGnVJ3nIqesNQCYjspvAXVXUPG8G0FaQRkZb+z3v3ZvGv7wyHXg6xfweHn5sAxMN5i
NJXLxOalm4KWlUuRC52TuLDLqJaDDwICzH3e7BYy5DfD26UHFnvtun6hYXRrkvdgsIFQb2FGhFzE
cQG2A7Og1b8HsqLx94+ACvXTstj6PabMpxM3nmBGEoxn3nZpFjgs4BdOOUuR+srKnpIpEpHTzocy
GN0xeG6ayuqy0/G8+/HkTfAX02se2fHsOVAD8qV5Cxbk6h9OHWwpHsAcET995vXt78k1HRSnPRlW
7J2q5wm6ne+q2yn3CddLgF3q4/8+nkzt06bhb6Gh56jRAEw1HZY41G5qmLT9UubVlTU2K1K7GiEU
1tjgwsOwxMyFqj7Q3p3JOm0wbnDXTysXTQnCBnq8D5+05tSlzwU8W0PEVslRggfGxG5Qjd7DaTqC
p+5dDEVBdDXXBkX5mGmJqdJekpV5Toplf/bFtnEkm+eG8Gp/YOFulnREDOeX5JMxnbGs4hwt5NmK
Bms9abGFVD08b+xFOjbvuA+mVl+rQ+jLDTLMEwxPAgIiyeCwjKQgxUafy8dmdkZIPUMJExXZy0cY
aulzdkg3heMD4l4Cy8vBWk59qFEuYEqWKg4t67twU0Y3x3ovKBAx4n7TWTzvI/tmeNjDvBWH98LE
9GUujjQvWlVcvXF2iIfmGbNGfXKPOSu7NzmBEVKcPaAmHRc/oCMtkoW5fMpFwa1Y2rYXucia7N9E
ziNq+koJF3E0OWw0LaVmW1uA+/DIQjIbi7/y1i7Ll1UXyZN3SppmM4FkkxpJROF7lKjYLYuA2tRo
gC+5hovmL+GqOkAMK2ig16L08a/0wxIyxYHg/PtP4SkYz2Wq0/XE3H+2AXgnpp1f46UIcHTZK9pB
UhaBgDFyIgnVJXwTdDL81KsbFIL5XWxvrjMRzRmtDf1LkyKH7uCdJbnUuvWdhg4lvzwDycQ25W9T
SBN+LKV+vkCjRu4NczNFGA8LTPR1Gg9zMp9jUUfnbT9zWmw4s8d/XYcwRRJSZ4d8H96mlcrnQAsG
RwQAKP7WNomgPO/7an5BsTgPSZhGP093VOZoXbWH26xya61yyUURj496mxepq9WpZt/Nhs2Atir3
TAchGfA32fCeh8TtuZvgNuqzo/AB2evL61ALQb6gDa6TQge2aJ+Yn7gPUAcxBNFCgxWKqED5/rxR
j31oa3iATc+vF0LXn8Ea2IclPPXUA1e/33NmiroKoQcCGu0L/jfjj9fwl05GqAOwo2IMf9EBiSNw
944t5RoYShnCaobG8/D6wshMyocHnyJGBNWCQlqaWdnZY7AwHTvcI74I6WLkTYlGJKOZ4iw/edTr
64sxnQIMs24TdTF+Xn12RsREwzhDM4uVjHFBfBzrTDn9fotDdoD+E4LAEdDuMNhZpS3/4hqwBRp2
D/iom3HwySmV22h3cJw4HGFveSJFaEOh0x+IPcRGpvR0f4XQP1gwnpIuqhzOL7uq0FvLfLYVOm9X
cWC7lGbjC2pQDDDM7TdB1euZc1MxkKL41rwQoJH3Oh0eT34/6SFlhizC0fXvsAIm3R30JQctkFFN
mZlI0RPYtlROy7eaZ+Sl951wKgBnlTi59oKsmSkOGWHEfv0WYSTL6ZF/wjBz/fprd0Y67dmrG+oN
nS8okNWJeSovZCJwbLrhzWEndD6jzPNUgT+gB7Ay/PMnAu5l3j8vP07Wm9mIRQJb1xCJSPbvev9M
iKgEKmcitqm0lzVX7zogwJG77EfRRVC2ewr1EBNejuIG+16gEj0WnsLinUabWcTvauzvbqjtNwEX
ldvJzpd1k/KHMRU98ZJz5ETB3B8HsZSItXhphvPdWR0Ixek34s+MynHob/kgAYRnmt+Kd0GCwoQC
3b9EFDN0s4095KRwQWci6zai3OfpZ11ps6sxahItxsqEP9PmqVTWcqFelAbec29kjfB/t0bRcvpr
3oizFi/sRNqJ5NJaWnDl0dhAwb6ez0sZAQ5wJOgcQDwVrWl+jxDGQ2k6YrSPwrKbiv4CNO1qCsSV
9GxZwTn+fliy8PnuUDuLuAQk4W5MTFBABepXdtDgxv94lpo9wjhfWn8rmS5jDQ+GskpF6OJh6brA
AK/wCwoY+j470qDim2RWMJn93OQ+vxzIhlPGF1+c9PKHLRHs/Sb5WlMXr8itXP1ZUZRuTzGdltDV
WzLbWuamTmKvaTzmnjBK0/ijjh1YuHyj8gQgUHj+iAnTf08URKOFIYEzTWJOqG6BBQpOZG7KgMD3
8EG6zdg9bP5R5793fYZPupmZtdRt/Uro8Q57P+/E0F04cA+6SZrDHaxqFqd5G4jE7HNRwDXTfrZh
8ghfae41YtJ9thl87DlDbGGyY4zjN6l0Dnni91fVPAJQKR7k+liudfCCra2llzaPH1iijtsGO/uA
blsEM+qnGIK+eraU5pP+yICv490bZt+3GthwPWqq/HAHUNfTrgBadEM6Pr17mya4dFYENiSZUcTa
HxPIlZ0cnYZi0rN6kruI8pzBD8Yz5kLLA2TU3/JfTtugpmuQwA3lG+Hu5ltAlvhigCrGdK5H6/2A
gNR1h+7/O9gIYT8KjA9PGdAWq04hI+QYDN+fX62xGR6y9gx6NmbTIDVwIIR7s6llXlw39YTlxzf3
77mGZmScHvpN3f8CGnmPdGr5FLhdsdSPPhaQfS4dWBerATdQezoePTGPbmJeWF/Gd4n5gEcd+2GQ
GzgjS0piubZDq23eDaTOJCEP5gWnu9pXPa9Z6KEfXZMbnOqxrVoRFNZqx5+1Ye3jUfd76dKG+yLl
95BbS10DwRj4lqIDr/iZiJu/Sv/bfklyQjfjsshOXKLE6URLAHAUY3satT6aUHh/eHnfz0Q7rBhl
wQEcmuTMxVSOpa9KvNoiGuzurgtVETNGzRH7SsnRKY3s4FVHJ1osz3MMbQc13eyvoOubPsASNR6Z
1ETrfxvgBKYSxyXnd+e2HFM5+a9WKVNXXMdO69rIBvSPKgbcdFpHu0LaIM+We6C3s6zXQ2TVSk8C
ZVReiRj+BTGjYmOBBqrvG1m+eHvsLYE15wtwPnds5CcOuaYSN7FsP1dfX0WBKXD8saYBTUd6ryk9
EDSGKCEVrEKNN7Ripbi/GAmn3Tr47IRDxQlenG/zRjQjHSiUA0h7vNSirG3bN30zwyAPI+cL1mvb
V5g39DSszFTq36RyWISu2uEhP62+imzguL/yTp2fzSTY52kzByaXHZBRxfZFlwn1629AMQZe3CV0
X/GWoErq7M2HdCVlUy2wL/KEuC3igdgBHhigJUgQ+ZtFujfky4+3pIu5d+HevIstpN0gSUp/BVPR
VDREBK9jwGKxe0cYxZ7sgr30dUEpWhZkFAncf+gPLHFJj3LwBPiowBY/fuz1kROa876bW7DApM3j
t7sVddlU6Lm9X41v+IF55Qr5913rruME7M4O+LbRGXAklhs/FCCkqA8nORz5xG3Z5JmcsS5X41Wk
+smHdzp+/r5Tv2p64zVxK/Yx4HlljV17sD93Gy/+ka9hdLoIoNXm+6QQnOwMQq1JEOjNgEdAzfWL
MlPXxFkQ6QMLyOQsM9R+T8hKqdEF2moQSmUs5lN8ZG3frIHICOsVymZPsdadm/Np4rn66IRkLsx5
I4mwx5SVrXb8iLcCUhUwIwQzqP+A+lwYsip8H0I7AZgKrt8KgcQ8vG3xJkNXHRtQNSAImSU2U4f+
rw1qyMQ6E8t60NXyYbvPRPwlISdYxhfUovoiLd8tLwaPa3mhMdPzGIwYurVBnVnRQWm292gPk00e
kLVA0obJRH1MPdvnP00sfA3GPIKyYWF4alwDXmyJrq0wLAp62f2knZqgk3bL4WnmKQUWl/2ypKYu
pqTSO4Gxlzl728VMn29vRxgxluJWqQ4i7oTuxkSJc8IT1E+55Fi1UhmcWT+Li8h/Iz8dqH+f3jxp
9nIUKc8BBdrCG8dagg8sit5U1/4H/XChEvAP8fw+s80f87UT3sYU4MuXpKxQnvxnwSoVPoas1UE+
aVK3Hw+U3fsLhyRGblR5feg937GoUjZUtcdX6DrCZ9wuU72LHw9DYFOiWlZX5XFtvNCNb/rgr5R0
7bj67whjQgKaTz7yrwoDxEm1VMeDfCc7yT8BT5Xpw884JvS+MwCQycMofKbSwOW7UU3DQ2BdfLIo
OhUA38fL8xsg53trzJZ3Zfvfvirbv+YE4vxQEZH7yr1/tXaqA3fi2jB1KaCZ9YUTZBibT+eqv6s6
xiIbRXEZ1OCUDwVvKBGxlIoO5833wG58+KtH78QsMCQRNxsv5qUEhxMZiYbUWlZbE7J4fVpYPTom
nOnTlp9rKkXkULrcWub0iDhHb2H5K9lxZmZtOF8yQg3TR2qn0SIWtv1vFxvaFQ0m7D08MmT5k7b9
c2WrFuFFLo+2EbQRL35tf40tT4QCWTUOBjcXXvEnaw16vOf4btqgFvEi6qhvYZ+olDrI6ZvwTacR
nLfwtzZ3Z9oUcqszrj4JyO0SOxkLSnNrNdFpO/hi1mQZJiZggVVnJ2Hbk5ZTkJGve8jKimePqzoS
1ilanRYAifqq00Vp4f39SCiaxO97CKJu8CD5+QYR6L2r9evwMvAciU2QhiRLdVjeBpMgY8xLvkDL
K0MyianLtcupW2aQD5TJjr9gqHpmR+MaHGeL/7l1MSlJSZ1UQmW/gmqzdKRePBaK2NCA0dse8Za+
PgNfZNSKyVqPr3r5bCHRduI7JyAEc7EFgdGHOAQddQQGUixq+FkIRnmV908TBaWaWH5hNkd6Nctj
HlEw/1HDRbLLaScpKX/w+HAd58a6WBAU1TNAdv+cxa8tDx/1aM/EqXijr/RHh9x2JuRMQkIqY4RX
0OznD1vBwnfMKyOo0fpAoHEBBIHHtYkhJ710Fd0+YGTpRtOcpd51e1gHdhW5ODd70AOZuwI9FFkB
oLs1cacTj0CgosetRHs2PMD+L8m+3WAD5d/DiNoW7LnLRp/+2FdJWYktTmAXQpJqSa178REN+5K+
GFCVIcLYecSjjsM9gfk1ryMwQhBunCODcBttV/7h4kb8yWqrxfv953T0zDrz5gJPQi3NfwoJAnBU
6AaGFAczIidK6VX8OVoQXrDaHObJ170LoXVoJasgKNWIVAeADELobNUPvBu1qd/D75p6+UWPkeIQ
QFk74bQ8mLxt6JzYt2Dxw4A2qixXt34Mn0Wrh/O8fHMoKF14qq8dCnSV/adRq5w6+Ii7uVmFgl4o
dhBmaG9vivTQI3roajIifMOX1hjX4BfcNhcDz2deb7Nwfv0XPNoOYLcKtbX/YhDljlrC6qxd0DyD
ecZh+PgCZc5DrbtNS4+8fZ/sE5UdsXE/Ma8/t8jaIiz+mPVs0aYZSuYzlg1nmxrn3xQm1ijON1ZU
H2t08g1FWSxu0OhtTeuyXhBv50I/Ohkmb3HVnixMJNkE0IvUO+jBY3M9N1O0SpN8d2h0eREAes2z
dxlYMZEfm8r4m8EkeyHjmw/2yNpW8pwvUtCufAJREBJxB8gHs5x7fG52WQXrKi1571idV1bvGG7t
dEBXnYSXGrlwKPNuvp0BZjApC25knehb9IaHH602qGdYp/fsur5L1sJVoBn39NGkMtd35OtWapOn
Bfm0KdtQrttg16tW7Op8ANgr45aktSmVIP72aKJhOBdSjArcPdpXBCmatp6A0nUYuQAXbzIR0yEo
G4uUkR8F6hxvRpVqZNEypDSVWFsWX1aKTpLd5K1/HsAOm+lKAhW8Vrmr1QK04HeDX8yp8d6EKIUn
uo0yOhWrKESGGlMSrOiKVQfKl1pbWWYRr9zTDIyzd+qaYZAnhhkZdEIOs7/fIOmj5CYVVbXOi4LF
yhvELIBPFzgr3JEYEeuY1nTaFVCPMseFlisa+SXwbHu2lb3UCbcK2j+/wLrc4McBIFPZOk7/jbMy
eNhke80U2knoAtikbBevbWvFCE1c+2Xbw1JJrTiZVTkAeUEmrdhxUEqUmgwwyaJwUzJ5otlC0Lyc
qjodT9vmpuM9F+895ohA1ctOwUapCQYZDMQX9WTIygn7Il+j2vWgCQ0zQI09yISfVg9Xg/OwVTjh
CjCH/9KxGg+nhCAOZH1Em7nr8EnjGTfKZPizmYAvdQfmXcc5VSFw/YB70WnWyERTi6Y+vbmUQGtk
U/jNdLfZWl01K+KzEpN+AuthN/VhWCTweH3HybY0altsGh2yfh2X3/nQfYjLZyBkO9wdoixSy69+
eRQ7w1s+HCrgmz+XXFg92SVBzFCah/ujsdcgWGbl7ije++C/yqqRJfCR28HeZuUunQdRheUEFHL7
Qj/rvHSGT+SYx6Pi84VOpIsoNQqtgWGKT52YnoQqUf4BeOE0IxxGHE365KBcIWQqSJx/K/XM4Syj
/4kgKdkUmlu9W6oocVD8/U0XOx2+f8KAMRvjtnXV1izgcYD9THs1b0VrxjR0J/6nJAg5CAhDyfJ1
emurU7RnN0QAvvZj4FFuxbYkW92ek8pl76FWTFX9dW1IcYBd1JXhauykMdfMYUQ9orZhkDf2m+Bt
Ds6YTTfY75V2AmbldhiD4RCBJ4NqTR5tCuYBRzLtp/SmVlBEMY8RJu/UdN2u5rDR3JLtwxtYocoy
zIgIstIXFWB/5TD1ayQkkAfqrM8PESgOqgzO9zWEJZYk5XlwKUfM/WmqyhtYZJyvF89s3JyVIcWF
lDlqBbVcCSdsDu6tnV4ZWDCWbaqG4io4HJSnr42JOtwrshSNG8T8FZhzOgioefwlpNcCMDfIThtb
gg4stvODHlG5O5TjXBX9ZFF6aT+86Gr1n+UkuyAdmoQj4ysPyC+HkM+IusNrh9PQgyA5tvdlyDM5
8vHmkNqRzBfZRV89/0NlGMoSDQdPCFBN47MjaTMZcySDh5Gw3MEWpk8uqy9eXcpFGE/NWEKFMFbK
1gXrqqyvHt0tpyv2FZkRgsKXcHGrYlG8Z/t8MmLHpCwVccR7cg8q04xw9OaYZZcR9GO2euR8wXdv
pDvvkU1jhEFEKpTrRChcMXOjsvvNA79+uTbkQX0pnvQfp0VuStX+77mnT65fo/lD8guuE04+o6zZ
kd6Jd1JTLmeTJYu+jllqAXO0NhnCrRCFT4ZYiFUhFekmhkhJEgBW4SdYL5yC3GdAFm7PfD8S+utx
hXM4PylXQGILwZI4bMfTTwqoOUsN/aDKKDqUu5/qjg2MSi/4yB5P8HOwsZBIONLiNvzG0pxAz/5S
EylEOyYVRJFpBfl0N0/B9+OfZrJgYCixkMne8IPrxgrrcJCcMJQSqa8Zv5JS4UMCB7jUu3XSzabS
VEZMBGYSElB+KLSAQt9tvEvnXnMLOhZ01js6CRQsOSMcLRB8Q0dPVHUCFwN8RfYFcPydfL9Y1+qq
zjxRiRcpjtYWQLWYVYtuNurqNkozF7kQGkH92AwYDVRHeGCTHeV6KdYipG4/lFO14GTaMgeyC3bJ
rPJ68F75S0shUQgNRlzw6zkHrnVus3dJUfBltPnuJBu0MZyRNZaM80/AmKegUhb9KKuEBEW6rLlA
DCIcQyGjUOtuMCuOCqieMpFaib4z+IQ2C8FVX+/zSI2E6lBPYsdwKaHrFUBOiVsEhxuAzUYTX/Mz
UT0TPHoWL0W+ReaWDyRMcfr7EhDR9FljWgLl3zqpnBEEw+YwHJs8nBI8nOfjw9nfnoMuNIUJ11ra
QayiNNjlKlzqidlI75cwx7AVq+dU/axukircLEKUJrHpYgnaaDEicjFd3Od4NDJGSTLDK10W8mQC
YgueqK5AAlpaJMrr1RpvN8r9Chhj0nM0lXFJ2PN2amqsIIPcPYNb/EfvLxRNQfP3OBHuTHrr5NUQ
ncMpx//XpAWxFgXgDEitWESu2Bu5R4ZaX8kt9XaLx0emwIISfTP5ZQsBjuoi4hWdhJ3BpHXloy14
z65e+eTkAwXFjdrfkWuZApqNMVJADs0apprT4TE6bdcsZeyMgyNibPtdBDrrW/EjuJECl3OefgzS
0IfarNGAY2942Z3vZG4bl446/X3s4UlJ/7G9FgricqgDyS0CWh/Fyh6OGpZIRq3iQmGFIWVyRw9/
4BkL8RnsfTPyM+P3OJtWJIwSNV8ZJYRmVI09LEhfb1lkpBPgCx9MzWIz1kqSPokcerQz0IBgQ8dm
gaaFVFcvJsfAlAqY/V6YHtqlldlLH7w8H2dlPnBMKilb/Pc5XXvTDS8Xm3RvleC29VtxbDTh+Aqz
IS7zFQVQxvrDYa8OZWGMNKah4URKujWn5uyf7Ob4G+LyiTAeSJFRQCnGT7wpHyVKR8Idx2KCrqlj
Ln5XmbFqUmu0IQLUInWuF4bp6U/Pt/UYTdpymwj9m0b+UBuPIPerDj2wCXNx0FIKQECn2bN+bbQl
EF//TnSG46w0MkVWf7fP6is6Auo0iM2umUBb392M7/UNIYbr5MAc65S10/Y7Qkn+0CVXt3Tetp9Z
JxI4jl7u1od2/K0MJbEX/wCFfp7ntQopBTomeNu7J4DltFEUmYrQwtEv+nZoBpmIt7kZDIXERORA
pieUJTQIvK9fTcRjd9luD0wJrmX8DAffFME4X6W74KEeBZMFFN6m8DW+ranI9G9d72SmzOfK2kj5
2fWW+CAi3NR2Tt6uOJDcTj+xJqr5zW2zWOFr0B7lS/siwQRr92cVA7yojVAXnIWWPG8McU0jOPFp
JqRa8gmiLSUW/TTz6fd8K+gTvEPrMg3fxKfssb6zbbcaBgS26sz78PLC7bsDC31W7aR/WhNpAVZD
ngyuCyrqMZmNJP+7mdGFF8e7tx3BXU4xY5QWYMYSTRVgBEyqqHmGIGT5Bf0E19USDQVVF/yE2Liw
0ywpLTCXx2q0gTvMEFkH33/qAkma8ndCZOBMDyM+gwl8jC/S48DuYxtGZV0mIXs25RB6AW8NqVP7
3VdpakgjNUH9+usWC6EgDPBBWJ7GmocR81kWZypOqj1/3sHGGyeB0gKGJ94g6F5HDb4nivZaiUNN
36bZsB2idGk8aftnKduEQgyTlK1fnn9ybhKEr8/gt/ZhB6F0weqEosg82XHZfgpQtFeHWO/ZkVWZ
eheVG7smIfzlSh2KklsybxWbknk5fQVOgMkqUsyMlBa7RwPtYzoXKIiDkNCioNGuQwrGAnxYehNu
Gb2l8fc2H7euuN8QJiK7MfPVm8hXquzggF56glLgA3+MEroHJ62vEWran/1JS8m0JezqiZMLA10T
a43hJGVU+5bpNyS0rS0N8PLMJUK9nPBTFrPNFyCGkebxRF8tE66t7nmo2z76i5/RGrCrlPkX7SfS
lTutp7wRMgTCDoZMbfUp1Vgmg6e78bBfIYYfUG0JSgnpJMepU4fhUJ16GyHboc9nSTME+Zbgvdbv
gYSOKJu63aub7P6PbUKCznmKUPt9saoE7o7dLR/toiPSbgaWjEsSvHk1HzGJ3kDsWSffiUM6GNhx
lu6vKIBRYVRkhCinswztx+1GNK+L5lbe8I4uvK1eib3HuBhFB/v/G9973bRBArAxAnv+uRDrT06O
i6lKuv6zvGYLCAexK1vy0//3AUvDG2SH1aqktr23EN5JAl7k3qHMUuLwWBHMmc1rVLtCE1cqXM+0
XrAdrQir+PjTC+uy5e5kebsb6VZDqtKcduaagShimpj7Ax8YgnmHseS/6DnuHCblVrJ26j2GuuZP
Sl2+qnNHYe5SIDIFUr74yIzzx3hXSgIQWlJl+1+kaXegu9wOlflBQH3XhI3zsJuaQaO9202Kc7TJ
HzN0G0ZmdDbpZJvz7bn02z3XtWeYNPj/wYT3Ahp/8igDaXKwEsDxn1qqOK8ssdxJkQb133OkTRBC
dO8/T7+8dOn3sgoxzDXvgO1UroZJYBesNfWZmvv88s5tTk8lhYiJMt07AhTvS595Eg4ABBaK6NDj
zWIt6aBRDFX+dR8z643Y2Iz1GDm+PWSA/P+Jf3OG5ZOZqp2fIch/LveXDOxmNPnJaC+PSWCQgOzt
JavJn6aGrhfnFgEoZaAmrf+MhEl0LBfr8FHdtNR7IW1RSpzD1M/PX6tczwbUKZnZJha+cYgKwFWy
L7VSoWyne8Cruw7fUSHId1QrPDMZ/wYZ5GDybJw7jNa/ujXtO6IJppXXe/nTWPQZ1U9z10ayTYzf
yxvFQaN/UfKGr6H+BVTFQIU4iTfYHInUeXOFU6g6PMWuja83eiJb6iymufrG3wRrD0Ha7UJvItHe
hjbhv7qf30iUc3e+4zy4yfX81ktwbshp2qthJNvnG1tgdplON2JkYtKtyicYrPIoDH/q6naiAWoj
sqKI83zBDSdIcp9GVUJ++IcxoAhEBGbyrObhmvUj0JuQvfyfnfxKMQ2qIiU187eFGnEkjg8zy5gi
Phv8W3sjlYsDrVO1B0sK4JofLDlmEZu2tt25GWKEbKRfI1H3j/S8zBM0e1R70wqY/zPmkq/cD/ND
NdssLbWKz0gnVtlG1w2Z7M1FRnHpvqdTA7aNdNmkq+f7FfgfWH0kadZXzURDatzCW7COjtbobvQj
eVaXhhgZPLwfxPXCWjiq+SGMWC2FowXgP1PjiWg1BlMXlV3A/l+xY5IYbNuH3/+xuKS3B5X+K3TI
XZ5Kd5XCtJiSOF9rxcgXXNsXqSJ1Vk6sWV5gyKq9rHWjzXOo3FrqzIog9v9VpXCSMYRMT4qlEEIe
8CF2bfuU1enORYIWU4qJY2/zY7/oz6cUQE6SptvvQ5LE+YnHW/S6MfWz8Hl0Xap02beUD21LWa7p
zMugblTz9jlV0QH5swxgs1H0TkiXit9Rc9FuPA3X8TOYkA9yXMPtiY8jWmdlSmdFDEj8VVi1vjIk
FatqytqMzHV87naU5adlLtJ0OePJcSRH0zcutvOvsu+9v1RcRoQGow/lIlgeVrbHWuG+crmctrVf
aWP+k0lU6MNt+6UsZREU268gEKFZaHsyHc5t0rTK+ZB52b6FIu2yx4FgZlDWmAZMm4uhTnI9AETd
j81zDd3tWNMrCbVXQJqqshj55IpTETc+ABtCSityyT9gXHy+Fow1n5h1Dmi4AhvGx21uhRT9f098
QvR6c6FSR/nXUzMRtjm71XyfzeMeT0QLzqeIDokyVzyvzZDh006nJkXq0jSXhgFHCFJAmouA3PzF
pY/r8+LuWPeZRGElUGZVNKYD3LojRwj5XbnyJZtvsoQTXPPpFHG/lvqihyw0u8MF27UM7j7ry4Hk
vg0c5i4WvHDvkfvKQzG6dh7i2N7/1Vpnf25IQ9187sTG+AZtSkvTPVGonceNI+/Y4gZH5tkmz9Vo
UipgFKbuTIedNRn9rm8rTYvxuSnu3dCP8nF0XUfR8osJT92ZntRzfXap8NzTJkhZMWh1U4pcz0Nr
RUKMZH0+IY9XztYIXwMf4ZZRkXicKcouSfBqVKGLVgx7Uc2HXZUtWQIPExgEmh0Y+0tveseMN/Ze
9rpBNLXLAEEuDvfu7rhVkaRUCGIAMdJqpzGrX7q0HkHvcMnZwu+P344CXYZJai36fziqpouMFkza
JG+7LWbunoPwgihO7E2PRvpVUEL8rY5UvSfIwrW0KhKeELJOkP06CaB08Hn5rD4gV7KR51J+UJpk
URgOauec7PS5EzcYulV4b5zGjfyO69s+N/bpknwXILQHGlRSplKpbPfr8V7WDUFo+gwN9aL3P+95
VXiTSEEZijwZ++qfQ/LBc/MCOOUOOlLyVsR2EnTltMJx6b4+wrw1PrJTH8zEpp17tl2d4T5J/5oh
BCHrL1DJQj+TGmKPgkj4PlUnd3Sz61sHCnzWoyvDTt2Y/VbGpHrzyZAGt6LTRM3GQKeOJiv/8fQ2
dJ5u07AfG8zG3ONg41fNDMfnR2Hic35x6g5Fcu9jgL9+px/e7CgCZgqLHcsIaBdR+bqOf2O8GvKp
uPpAbWSG1b7sOj/kBWSg0HQchGIDUWg1/Oaj5e0oSTKGpPHwqCvH0hLNZUPLz4UCMSIr+I+7EYUn
to0V5nGo9HF2e9ge9A1a1zMVa82ZGv9d/5z/VVAqEjV2Mvu/+8m9KfNtpbEIsVoaZLp9XSXOMVwq
djeoKWSokTfZL8W1NiDjle6/DQIoBZxW5LSJDTgHvF6rs+bfN3hYgWMTyAWt/y11FDHYVnd9Rqt1
bMJ1YATzm16u2N4OxV1+TaAoSnZrmf557SGc8e23EVhzv7JE06H2v5EBE7Cw8ONE7UzGgqzn6gm5
y8jod34Lv8F0VA6jSSZBO0bVE03T4vuKc14iAdMMngtR5MxSyjMx/D+LTyaOmRuhUAFsUM/R3gcj
Ow2u+OF4aXvwecDKZIw+ur/VTreKME6l61BtSjemxkoGVvYSSRDEyqdJDguUszIUhHNZOQz+tVoR
n4Lx981QO21xkNwghbFVs06te/+gMOcMNF9hcn8OKBWFOx4pj48lAdGYnUGivNj/Fe4+dDXF0Vxe
YqKK5zA4YGHgOozCZa80SsZlji5CN3sN2YpcXd1VynzCbI8ZLXjGxRHIRAvCM/cc4uFGG9bRJ6BR
ReQnh36Sfj5zKj6livaX4NLeMIU6vMvwdD7ylmUOm3g36/cDbIlCKXrN4NKdneitwITZaBfxyNyT
P/X7pgO+Flcf+AALKd5BOccGsVTNyOLpf0DEmelbQWcmIa27QaZlmKjv4RPp+aXLQiMMXTlTO6HJ
QMQikNxfW7WDqEC/Kpl1QN1Oqvb+4nNz5SgwBsRUBYZtyPY3cfAlIgnAvkazvzjxKF+9EmacUXIG
GRoAM1An2VV7rf52oWhQur+kaeyh7kcLdD+eKSUuepSNTK/dyfO4MIKetvuoT2pgOfjZg+3LsAa4
6MUIGHIKkaKw0cLg2X+eb5fPb3bf89SZESteei4ZeEa6usOCs3FLFrErGeTiXeeh6L2hwp1blO7A
RavdUtfSyGeY7B/0VxAEIkXmMsr22l9gu0GpUd4+JTQpNwCpcclrktagMQYAzOstP/tnwYvt2qJL
FFmRYvtEigngHCX299S9hlnLn4IWrv0QqxvFkln0DKkXwDzSF0uDulAx5fWusmUtUHw9V6B/g+zI
wQ1L7ltG5nwVou22QvHPBjaqSMz9WB+4OugwsjjgaBsnA0NdnwwUiVOBsPTl6LS6ny3gFUp6zC6h
+uNmOrZeWO0nrr9nMF8WxRMAHFIUqbSN69MrpVzeyTQOJVbzmaoJsZyD3TjRSzCvsPePmcatJtiQ
jd68/zOSlBjIjFoPg0fqIE8JmKYgkG2A4aqqlMZgNGbuvQnUKhwIxSbtN3B0oWaoy5tpizZC358t
gCZOY6kXmVAX0zdRJwSpf/KzjuHn/gYpLCcr7ZY5MJ0sPRmttvQTSP7c1J/Zoozo+Kd46hOytQw8
racZk7mTB8NkZbbKkQ8wHALCuZfgT7ZkpvLHjTg6rFS3sqfKes6JD3L8xmvVd7ZCCfORCVOn12Sk
AwyCnyCyFFa1R3tJZKASGmqnH7t1vszDsr6IYebCFtO/pyH6sxqn+09FC7QyQnyei2NxpseYmAp3
w/aU2IeJ2xYbhUOcFRay47Q4XK7Ny3jzwL350UkJfE++R3Milq2Szq0U0FqH+UJYubJumsZYmwDe
0sra2mnq3WOlAX+hv8jZxgtbWsZdT/Zk4W46LeHyM5mxxBpZDHCoXIupXTF309feUgZcPPEHz3UF
2Be3dMZ2Vn58dq2cXKSufBT+NM9d1iZjMecPUUpPGNeiRCjhqLl8ov3GIMR0bLr1JAc0TNCZFOob
MbaNTljycJFCK82zQOcC3xBSUmD+eJY+Q2dkH4+KpSz8ZFFeESvW6kKPw+ssLqb/iRYRck2Dp1ce
XZsXfxvRcI5YvbvBVQ6f4LBTStv2BTeO7xeJ/Lgsg4yPPygqbK6ICGKj5NjtYaxGdUKfNyceRxjS
9niIHHVEtK4i/6QswJgQp8gpbTjYnlAyNZQzHVfKlrnkS3NztwB7bEVpGcXlWn6POPi9dOYOQvr4
U6f+ZK+C23AqGGA4/x/xrleKz558AISSJxO4pWKa/gmJsw7noA8cdLiw3oV7MzA/8NLMt5JRnixE
8Ofv84mt88+zGTOkX71EMjpOusmCqGFOQ4b6HaqaoRKDr+haTHH00cxww3QLU+aIrXSONkTN6+HN
jnfjiGWvZki+yi0r3DHLAYIzIYIXM0pqeVPLfpPd4psmDw3jd1sxGsz1hu/HHgxUd7UGYWMG1Uqt
Qsgg93qx45c4LxsYwsnm38Mz6Lr52qSRyQXLuKS7u4dLODPjY0KfxtD0eYr1jRwX1syoSpFz0dwg
jK57GWqdw0Y8RcKNqFxCPiu6TZ/VKEv5xfpfjB1fiB3oXZZCqcNXmmrbs96tnpHqNInSYkfZsoOV
SL/v+DgDQNdRYmh+LwzP6b5Mcqp/urZOmrTJUNonC6OI52v0maP3wn7c4tlSV+5Idqe5JfgHQ9Xy
rC9DKcwgeliIZp9zx0OY64/DHn7qUG+pmevYBRLlIZWhJpemCkKXx3usuBq1IvMLsw2CaRUUXDLk
V9EMS9/mx0cgoAFU5k7MJxheWVg9zrFhiGO56MKZ5HKoV2ObvWgcoJP1zMcNda09l//7Hsc+nbNW
PIigpxj7E2QKj9Umy8y0jXxrxk5QawdQ8EMdz9pbuLRsvsGzbqAYNMSEfdgR1hJ/nWjSP+O4vCDg
HOiaHuJXE5lTBWm3hU12cwEz+qXv5HOtciMeJ1g+i4HBYQr9TK0nnRSR449tgQgdSxTZOz/b9pJh
fdn5qy7F6GQ9Z6SxwonQbr1coyPeoANw0T6WTEty0Pfz16FuUpHCBe5tOarhR+kCh6hACtkY1Qgy
2sZ/yjqxFdraAS1UcRq8DqeTqm70xKdtEAfH6Jba4ARaWUOAfTZjNZntkoIhc09AOzX1+rpDs422
rw68SmH+yLjgfpdEJtxumVA/GX5DYLW+a/ICU5doZrtD+5dkmavdc+tJb3049y4rNdjT67TYnshZ
ol9lKZXh9inivzGbNM0nt2Trkqkd0k6GnGpCxG2dk0pYTkUOIftFJBUEDLb9KMZLp1yoRC/zjmtZ
7zmvsXnl2teIUGQs9Z3T33UaRHcthuzNskyq2cefw7pL6THbbv06PLOOl1gAMcACh24r8GwIGsNE
2MpDdHKxHw0Udb1CwVWAvyYxG+HUWtqnO8rneTAGgLdK37XUGIWxUehkjGQF/ZxlvDY6dsQHpG85
NZQZN09+LlN+iNefTCvNieGvjnl8WM19bK9894xBp4mHNCT1/FMJQF8HPBfbZ/jhmoEiew63qwlV
x55Dzjg+5qV3vSBYhal7u2YV/Rj60qGTGRcStSST4KE81FHLYOQvK6G/A2/1A2Gt3aMHamf4J+WQ
Q9GxIJ27qCNq60J6CsfS7hXiTrIsLfMajEEAo3fMGkdkoHptF56XAjdZE5cH2v/7Xyz8aKpMD0Tp
v1jOSZed6Tv9U+8paHF2kN91l+FP6XcW/9jNL2kq/HBeZlsoA4eOgs2/YMBcYsh4b9RDJx33LHzB
R9nzDW9XF4FVk6QafHVw2SlZyVhN8ViiO9Kyy6SEgHRl1Hfcw8GOakmKrnd84UyYemeLEbIDZIXd
DXNWFHMwkzFhqWpUL4ceoxvLr1DWRV+5DUD3SBy1MuE8WYpGPGd5HJ3AE6BrX5HJw7g5M36Rw7xY
RGscXrq8MixpDWJGaJRqHoCQR1Jrrq5bAaFsBMBIvZZmkGPAwRrEp9yFx4Z5colf5J+Y9Ai2pre/
6kWfVlrCgHZ2b1E6zk6mi+IrtO4mYNZzyv5+Dg8F3NTLku/QM6lyPYUKIxhni58egGQTnxanKF6j
xGNnpK8zDed5sY5taI8l1QS9LybAjLAxJwcvHyo+IoKlDYWtB/GVxmK+ZQqmeD0OgJ0lgMEs3F4e
GNfkjiv6lhMSNXe7L0kib19vHLyGMGNVWr/SL7f0BwgLh9GbO6uyk1TnOpFdkpKKkXHE6PpEXDaB
5zkhKwAeXMylv9fcdiH+74Hvr3rEA6c2vl9Mbc04HMPDf9YphTvgFHte7ngh++Mbl0PCCWv4iNd2
V7AEzVhXfJwAbI8tYMcMZlaNU+l8piaja0hflNsZ0iGCOABT7uvyOdkCimqPyZApGAyzYwN1YRMA
z24tS5zj+HYUaTMn8DRdfhmyVDD3r6WPPFFEI5O8r8BKfNINNYSIvQsNKX/LZ2UEQK4QEiSspxK8
n/sQvuorbBW1PPHBD+4yyotT9gEeASxrvsq9/49UZOFLpkDW9N7PONqDnNcwIci1uCkyBwtTE6Y+
hQHz01vOkWesPuUOGc8XcguOwLgcWxbbC4f+6b9WDUh0gg0DG/KBnBOhL5UPHsF93S4/OHmUKy7h
OdgjskIb1DBNeiUatp7tBhclV2uStIQXeAUoMP1EVBNJlgWLTTtFAULQZLORuBerr7fG74QXTuR9
iQQc4EIV3AzyU47c5JET+gg1dmKlkeGexmDR5QSKCAIRZIiPHMeBZZo46DB77SHDuffB/Xs9kU6D
PFqZjFJXGTJjU6EOBsbh/trimAsltRqeybkeF+MSBaRY+9Ld4+uagg4CJrLWFGeL1t5ieHDnQEcu
nnNGDdIhPesDWfNOQ7NcvW7ou5407n/GDOFP9gF9YkvlRB+sigGmQ2eaJoItwhiKJ+zeHFs2YYZT
syDSvYIJokbzBJEyS0nHCDeofJYCwxhccKkRJLugfEFZG/INNWIUVfQWMtQjLaMXWv5dxwkgFqCo
js1hFwBszKKthfY0priEU5uf27BW6EzXdiLBbGtO7wRDJFA74dmJ2L9r1qjwYhErt1PH3pUt9xtg
1v9idVDG+lrMWSeHWJgEtXgXLLQr3yWDOZtCRZMawTOpasgI1seNyo6cIFs1YWXvszl/aw9GoGuj
3GtOPw4QCNgl1ZkSqhOKNY/dvct2Ylb5TQES9F6/kjkaLZVMRa9lZ+j+/WyI421eJ4JFMjziOaaY
uZ8clf5YEEZZ//NivpHqkoEkx3ezYXwc+Wgc6YEN8o9i+G1Fw15jxeHDW5iXurL7CCra4rxAz6c4
/FvnopcymozK8iYcEjaGfaIJaqguqpqcorRzk1wE1Kmw+SM5FFNMswY5WxAZrNn9k27hojOCodeL
coUsVlveyuK0/S6JJzLyb315Eu8tTMmVqZANIf/RuvvnZVLWThZJu7OSoEcxTKznPQDRwlkGuiB5
gnQ259XP4CparHzaDzhf5WnveeSok0TSNMrJj/mQIpwQPbai5cD1Rrgj0rb2Wqy3RvzRhvTEBQ88
Al3TdpnF2WjeUVel6nkNpPXtlNgV09GxhLZFsILa9lERmmT9vTFVMVqYr5WS60Ru7Dwezw6R08BL
Az4FSHpw2F93JjkUpUBoH/U372wfwv4QQswQXOcoYywOg3g8RHOLh/XQtziOuEo8chyjVJRwjHfb
3VvaZM2sN+8kuTFTD8nV7RZbn0EP1aPtCRp52NxdIEfweRSgjnTHvqN9/tH1fY+DyDhF2AJMzzZu
pGKXxn2ebBL/Z8ratrsv3u4xYvWBRBDQQChDTpLxOyv7izdchclmwFbha8E5FJPBdXquNvqiKen5
moLIH/EoU3AuT29uZIEuq5e6+c/ez3PZbf8W/L6QGoHiCjdNTvWywhZ0P7XDIoRygAD6iezdvtDc
Ff/eLeExol2GEY6Tu0w/czttWgsMS/nRV8eqEPE9hf7e4+bRGoLGrzEt9LIjqm7Xycmq7pJGmj5G
Eu+GY9csseGRnXTe1Ix7hRuKdl8T4RISMYvE80mFfvg+4ZVl4Z1zfgiLIPq6fMD9U1Wp+ev29sI7
4noyElwNlDUTqcbRhXnnpHUmJ+s5QJeiduJSAzGQbCilQ2vg2+selbGDFGHJPTh4jPnFmfGFcMw5
QeY0SQstqSfI8FG/u9y4Byq3kl0lqDmdLyiH2VewG00B0llwsBw3K8PdCs+sChvWpDqtrSuWkno+
TIUgsn2r14KY+ufNnXIS+K5gnVkjjOpHwdpduDPfIn8rJKZ+QJMqi4I8d4pzWHbqgTklamOYopH/
7JT/lIrR+rgqM1O91QCV3ulc3DiINYoca9/9PUru6qz7jpemPHZ2o5X9X/zSVHLIG6oDQLp4/geG
BrvdSLor826zN87fVbQZqFJ75rrtq4rS1kmKPGrhUZVdDmV6DPc6VJ/8dq3d/GeoWJH4GsLzQQnH
G34Tpbfv9uukbCgaVD0omimqmOzFw1IfuNALfqapfvWOd15Ci6DAA4ILKYEOkuNCzXFz0Up/vlKN
MftJei12us0OXWfSvvpoEL3MHDiZ/mlAaudGbIwfrPCigZXeF4PvXSIGTN/NRGgNd6JQybHbVfHM
l9vgtKJupvJFDBdW9hiCkCmEpB6XA0Zs/79Lqx+KZPTOkaIAXyKcLk7SdquzoJ/NVE/g/AyZ1Zhw
ZJ8gjpME28T+ySQbuAlwhx90Q3+TmTYLIDE0V7TuY5I7mT4hekjrDKn1wuPblNf31Y1ZwIUeJdE0
GFzHx4ze2PPDhU3phEZd8rqoe4Dz3FDfmau6qrnKPOYYwRiAe5khHMYNMRF8eWIEpBCQGCqBGtUF
kLEfsN/fxl6pCG2DmOpOSSYAmO/iLOa41Wdxj7zlMNKXYCtNroumKDgMo7uR+McEp3jP0iO7CUth
Rk41tvvkZOTNmLyb/8k4biSh2kJyt7CRfptA0jTLeKiz5jD7X0rfT1UQTMFeIoLAU0dxYF8uHwDQ
boctkVdwX0N+02/IpcQfi5BH0fU86sLKjknCarpqCGj/AjA2oVm5fngHxIcX9DD8avqqtGL9kNrq
wmGmq0q+O2SWMRaerrTroxBomVqaq2yBqwsdtzfEppqL53Mf+EC+iSDhl+WEQDojE8NYPUyO0hi2
D9pjq+pyyB4zc6w5Pvu/wdZ9FSIuoDkr+QSDdVgLdAuSh0Ns/QrRkwz5K4P0Z5GWpSemzO2W7aEv
SWGQvCyr+1zP2lYxSQpzpFoflIGr7NyOnz15XTCgQFhWHiEn5EpqomNQNIiUxLPWbCbpkplZOFcn
duYNbqUzUaPglUX2sjLUqM9KfKqj4nbiZhQrhmzlIJZq+IIuh2wREtVhPh0AKIUq02MWmzO3Yv96
y1U20VlEB055ytf+xEzNra6voern7jsrBi81fEd/Mei37++jIF2AoasK+6xFTQrcBlQ69rppabqj
KELbcIEdMWGVxNyo34PTPlG1D6ZRGXQV5wY/8Vao/8laZIhK1itrbKSNaAMuLRYgcm3B9OstgUVI
rHpUzejwW45EXtZAMill5YgM56HmFrvKp4r+/Oq+afr0K0WZQzdGJpnhS7OAF6m1psnTsFRx9FvK
zF/FRDmQiDR47o/BJLC9H63aF/3Dpg4geZR6mnKFawtVXV+1sm84N55gietuJd1uhJa8oIXtHMW4
o2QljG5z83JwTBWDsvxnc7ZyB4XmB8ltP3rWZmfRZCAWUS8qn9byowQJtnZtHWGo/wTJHqi8+e34
acoi3BQ14qLNbGvALdopw0HJCd2Us9qONSLBhDguR6zJ0lBw7aWWzLPWpI7gNb0nkf28S1JsEsMY
mmemENAPS0HIpaNylWSioL75u0YUPJf9BXnSG9xS/o/N0GnspyObwx4je0ydcEC+5DixWYvkHraT
cOgvWGez9ExzOnFpdyMk+SUz0ZOv8Gl2V/p5CZgfVOQDO3XJxe6gY0C62DCSvMLWip2/63gU8eXl
RWCoZFMTcVR/uDDo44uf2JGZmm350tgPZw/KeD7HsLe9OsQxIaoG2MWJPqsD+mkcRJb/RIHQwRVn
XBQLV01XutghUheQ1sf4iVB09Mq+5izk6N7vWwvIOw1vNYn0/DXwMQxpih6A7qG7o35DjRHNGIw3
wa9XxLt7QaAHWpNAcRZqSGgzvV7eZcLk+wyFuaBX8ad618PpYd7Cmb0+PllICFeInHPSq7wFU/Ji
NG3PsqkiJf+Q0Fxfj6GJYJjGr/g5uZl9GXgCe2Qfg28qjn2wMoOrlDoyDI8GVS/W/7E3ehVTAXmm
14z4+1u7QZJJCKbz8E1cvUutqNs42zawHK+YjlW0hum4hRfdY8sl/CTH0/TQbuSA9ujQy3QDNiqD
2jp8pXYDAtx7voW0KVKm1nm/6c80f9L0ChmYH18+/KZoI56se+Wc5qy4hZ5TA/klilhMeR2Yz/Z1
5+OYYwiqojiPi6FedSA7sEXspDU8EgljS8NlsTHoS2htH5nbRJK0jmWAsWDoi12T+irovNOCZx8U
BSfE7vBXuO/eaMYzZ36FtcJvUizehsV6up74VQAj8DyQiKWUP0ohN34THgjvD4TI7RlUHpZu9fMv
m+awtM9ynBfqRotv3ysXzuY/lZP+X3FgbQu5AujDwWK2eYlPVfdq4IlLydb1AloA5wv4sPlN2s2v
0hhe2XQAiiv5NU5l54B9gl9VdxAK0K+IctYyZ6hJwRMeWcMUBGduAZ1smn5rugTG0KWDWdhPwbht
BPlDVAXskkW+CxMFJaSRAAa/NqbCwnJfNJQo7tH0zJYQulKPgnMYLJx9pqWZP+UG6JV8yJvURGa3
+LWVU+RqbXnkUdzySARSGL/XPVXAGtjCcqANu9wu3TyR8KBiqkOnCcb2pGZSlIYyijqDiqM/+YHL
ur7eXexpFcAkiBpJXKHCg66Aq7Gz9YoDtcdOYNVCx2FpFS5wvbeMcBjcbCXhnUxIIG/gjtwXFt1W
kHhmDD19KsQnTu07SW8G+4YBkbVkxHH3XTKkEFQNhCN6vC/mVrqE+hW8NvDWmpn91rgi6dQPjnRG
7jPQ7kf29bn0LSzCiQFcpFiIOvjgpuf5wRT9NWG5mEAvmxN08q7IGy0Nd7DJNaLqZDGh/OwcP7s1
rlQZmmjUNV6igGzKU1C6Oa0vh07yL2x2xwBLF5bsV3ALvvqu3JCdx+4cL+L+QnhptRCHknXYIMZc
a38QW90ECg3Ok+yJ++cgEIUmKsMi08mF2KYQSIj3atOONsiS1SWbv0Pztksm0lXYgjE/fYm4oXcu
0MJO/oZ5ejpcFEt69GQ6Bg/BkV0Bbnk4idsY0oEbzrFwpTD35yjjNOa4HEozB+LoVA5rxw7Ntv3Z
EeqBITGKKlGK6/z3mmNWM5XmtvfADNvO3C6+I39OhnLzZDkME8jMBEUmwbtqAWHMIUeC1bl4D8HU
KfG7kMJvtDUB3ooRXtZyFcc9Tk54CJLDvPhcbsHzTNfsxdgGn+hUwhd2SGwvIZMolQd8IEoTfiNz
/pDdjKyEASP1hjPLuviCRzwHkAg9Zg3aNBxzwoqjIPo35tY0002MtEtYBKzyqq/7SVHDZTNxdu/x
GgT4FY6z9iLbpAznZAgcWpjQ9lxNbk2hfMUYoXWO1OwI1my0VpBancXXM40u4SqCfHdJ4gsFirOE
W9DSg2vSL+2Ai01sg7YXB+2a9zBPrfixda/VPZmGfLGjFCAQ/AfGy6nKwHzeajcZZggHLglPUzRF
RhHplMVzphm/EjwyhKCzQth4wOd5AFkXORYfQsYLTkRZCpb8uIFo5Ve0fiyrZqg6njPEuXiKgbCa
hweEICPkX0ypQKoEvinPpyMWmf/WIAK8/o6lpAFr1ELTjKQAf0ZhO0SoOizXPVld00z/OONFqomE
D/jJnLSZ+IiomkkCZ1rpl1sAfFAAA11fNVCnX3skG+4pesWyirwV24aVWAlDJQw8VxXAdTtDHHsH
tMUFx3UIK8YxSUElE5EN7XB8Mc24Uqb/1YdQje0I/d2vXcuN6INS8NQWXLSmLJPZTiqKMmA0IiSj
cQVtxkYlzb5LiQIKTo9J30VwK89tY2UQLo2bB10+Lt01SY4H2ys0YpWcVzk5HgA0IxGx/kgB4g1L
HDGghONwcSaS6bBJCATPu9dzLkr1ni4vOh5o27WDuEevUnIxj9oYftuFS6F8Yc1TkNmfTp8yDopq
CQHUUKr5SGpnGjjUBE9SGA6gLy0KrWBtg5aqR/U2SipcYLafbj/5d9FiCAQN9i5Te77VksH72qIK
GDz4RspaSocqu2fjiXoT8i0CB7rdcSaWcun9vU2Sn9oFt63bd9Z5Zv7JVFN6PSICNJI/akU+csf8
ddM1UZyHNE5NDoov7hBYMIcrvbxQS2v4/QTfPs8Pgm4B18beejy0zfwirOazZHRFU7UkYdehffmF
Yc+gNzu88jkjjeDUCeRC0enMO90ASGRekjOzyWh9f9jWszXQzHox4rU0CGMVtXs1s8BdRYVNKkug
Zoi2mC7oxc4D+xkgJCmS6DG3XLW77LsqfrniBwadYAhcWKHOa0ML5xdZA0nk+y5nXfqjTm0GXOxC
boYcazjViELI8FOoHK9rm0B909McZuW8CE41wZu+c6u0hhjRspRfKGFs1kd6d9s4lo/jFLQ+d+SW
qkm8saC6oaD8rW4sQ0G742Tq+ElRuamfMUfoMx+C2I47dYZ5vh72FVcm8xRlk1vEF3SOIROZTlyD
WJPonNSGFsofjYpj9mGVTQUPe0NM4FXZbZqIV4U/CA40pdrKhkWeiizGkQ1CiwJxxTSLjjxBlwCF
pC1O9vK5SgANSVKkhIYVYLH5U1KWml2ZOduc8Gsu7FbJ1XMrEV8cSaN96PyhY9GIZ1PR54WjeD9s
BRue5YKuHlVnnl5IpRKjQI9X45mWf/s4P85Zk0MlU9R2084aUPYI3ZNb/zeEVWyUkKPRWy+HbSxe
oBsvxpyIuY114rZ0iSXfOErqnm1BZYNQGuCnaQ5P0kZLPtmhzV9HtU60kI/xluXuMAS2bBmj3yUt
PQae1kLD+qeAzTWSjMgGW0OcF+a3//o+K/mWI7QSTAY9yfssJN1APSSX5JThvGDUNIC2anI60uTY
ci0DBieFh59P7Rjm9a0hpODBaPIRpFsfXh6qiqRE8XZOkmCWEgD3Q6cQuskkFysg805an6Rs1L3p
HM2X8L2WUCTnz5nA7AnDNPk1ZVEGlu072p52+WucZdXUTxz2yRiaJeLqVuk3M1c2kd3JicaooaT2
EoHfDZm65ABlM6jr0TSD97OIcM08A87J+0ljUAV0jefYZAtB1N8GGAYMQbxWFrUqcFZtnmv/wwBC
0YeNCKESTszgCMb4e2PIJkCWWOv9P254viD7lp9TSAstpuTMO9/43KwQuVfT4CeYsXe8+xWKER5j
WFLwXISdIq6WgvANCqCdKFJecg4Nntk3B2y6NqEEasB94/hZFMIBPoH0UoCZVA8TfYEF2Lg3vScG
T6a7crc+jqXXY10ZztLy/FPz1L46cIdD3qhBypFCiFoI2nlyeKS4nEBUfikfWgT8C/tU+y7qcIbK
4+dzty0L5FMnk4wwdQGLzafCay5IhkRaDmDqCCKWVi90aLyVKAi4sbQ+/5hV689QiuoT7+ITiE21
0tBP7HQxKxO9g04Brcs2/wm0+eVeK5gbWHFMXhj1udllG/z77k5nF8tno/RAmnb0hDzgXYXZ9o0P
36al886EnhV0eYwrtDFyWo77fVDSJoRvWp9hylq5gLvd5ov+zHp+4NMcpQN9OMXhjfYHSHjMxlMo
KDFZW0ZcOAY+qbijsvG792YmKcwgFEa4JXz7YPZET+cZg9fcct+EryUx7ns1ZyizUeKnt1kgVTMj
X65ViA1QPOG+gTew1eIEYWqJgsQoF4SVRHRjf1OSl+bsQWnTXXIRP+TZCAbYSgK8JLAH3HiyOxti
9Sgubf4SbLVVu3R2rqkCPtBuAsImDmeoNVWjum9JgI3kHj2iIjm/bsUiNHsXL3dYV3XGKtJ72+Q7
5S401TvPunqVqaJ2MB3KL9vpbaXBtqDNWKRKQqe5BRZeMKvnh/sYnTaZLAFSnRS02h+bjs5+jt/n
X2jvnJnmgzczY6MmFjWHffIXtWxbYf6D+UYE2y2s/vFP2qTbSc1adv7ZOoZh0jBOhK8+bj5Ivr+d
D59mDvDa8mtxycUKcW48EvCqacZxqvyhwd34TR5uWuuNvHnouMcE5aGGYZ0wmOrIhn4ROzlT17M+
cLOZuqkFVROiZ1ViMzWrepfqNeaH6ocuBQNctYcK3g1kRPXgpOOOeieHjgzcBpP1WJ0dYiAhOSe9
GWQfZWl1bMx62U3sqP2V/DQMaRiit40VQFqsW8jOobXy6ba2V7mDmjjLHH0O7YsVJgsO6mf8C4PI
/vSLG8CmknY3YHjbWYRbf3vIOGiKo8HeIFgakgW8m9/tk8KiiEtOdk2n9zsHTQINF4FcypeEl+21
zt2u2tIgfGAbgk4MIV/ABtdeoMeJu/byFZT/G2j45rhkSOI7x5gjIbtA7IyzotkjMD7sBUNfVDaT
1O5p69OXlEDUOxabVTnC+xvj5xDt7uzT/LkgGHJ1I2GzKvHAwZGn1YZ5SmzMESZsmkD/WIDfjC07
BcuCL34qosswWWpJSHunRgn3X6voD+f00d0xl/luKtLNOJDzGPrcqUw7WkhyAPBwqVJc1LVhaCAX
Ys7nfS3QzLLEl8rcCFrI85mcAeZsQ1HfSgu41oOcmG77uZpCN55ZtOTwagIt49kWdqQpw5s2dpGC
B9P4GBZOCNm6Mrl5+XcX8jOVyzgA7/uGb6h0GZG5UtWBG4wP53croOBaFbwLEh16xlhB54x9BLC/
pHcEId+acH/u4BDJ15N46Zz9img1MXlATkzff0itABRy1gIZ/qSOf0Bxp0gcZiQCwuT7nmmtAVwY
4HmZPozQykgiYYT6VTGwWrqh4Vs2EW/n5YbZT1q42yYu9Js0JmJ6NXAfA0DDKEutN5/J6arrgcem
8tKnZjHOJVmoXcuZn07ESU/5oqocNyrHXDZbAWPaMxnivPIs3zGObhgniXxy0m+7lt8whXKfPSXJ
gPf51RNmSEzCs2loRmPTCERZk9stvWvSHHPdFfPnZag5JEOGzfhD2DotLkRL32+7WTwtjOqQVgaP
6E2B12JqtGyQbtzyzd4pq4Ke9upsS6FUKA6WxvyjPTBbX9jlRcPv+dZI4NGPYhI5byOHHorOKsqT
8qoa5sTM4l3HZeorePFItLWRI1TLafhaj/tXDsptQ0caKJnyfznAbVyU0w2C12P5cC1Svhkw/GgX
RvL4tI0gjz8BkHkDoAX0jYpbJ0KkUB3irwF5vWKsiUsH/FQraUYRJfrhFtmRT/4Fo2n2n72CVsff
Zl4I9+0MNnlomx2/ER0dRs/VTr7CBQssBaHLO7bhMLe/adWyrSiW/MBXTiPT8FuS2m0Yr3joBCAU
k+0rBhzsK1oK/03+X+SBxXkO7HSSh8dqKQCbcsRblcPaPwSwyAGG8+2NoygnmqP6368/36ff1zmM
+x45AwQiTf8h4jTBgiGG/cjw/XVEErot0F0kkBWfCuzImfhVWfJ+wOB3ddpdXy60fXD3RXJw45kG
GXzGeAV7jC2ga0/rELWOxwivp6b6zoXPhxqOs4ZrwatfxRHd1PR5sRUnfJRzMT9qLf8/848eGNF1
GqLgJXCf/FiJXcVVaR7/7usKMNM68KPu7DYaK1Gz4FKtToNaKHOze9UqGN4dGGaMfAAm5i1/jaod
FwgADUPI339WYRPLXEhmrKH1hwu/MNGqoZi7TZEqkzT7Ef/49ChaCdZ8LoaAI3qUcjW6ncGv3HPg
TolVr68RrvHr28HaVtnxnwE1OMbujl9jMiS4P22x/WCW/wz8Op207lQDryONqKSrkJpgRz22AOr0
OgqTIMughseq2Z63NxFrq+1AvVu5POwqnNfmlggQOgj68c0+Zoyt6Ggrt0nXjR+9SdfcIGI365hA
5Ze3IFpYqliQ/TOViINGBAI1Niec3bu94fbjy6V4HKhSEFBUCfDT3AZpHK6+6vfpiinUn1ONtJlB
BPGI7SLvFD2rqIGnigO2h9+BEj0RhKwN7U+xbU69fEtus58opojr3jPRzEFNyQ9CGbK8CHChBgg3
FI2/OoIcm4PkSohnLFyIqDWQArj24SZU57PGxmRlADrcy/EIZOP3ArsFbcNztoX6hiGX7V7Ul6n+
XvuOr4qnAi6qSFiZx1Z8QsoMXcri3qLYPV9yD5K/RsahmO1mqdo0OzjJuk/vF1yiEJS0HiLSdaUL
jD4pjWfp9ZOl0m+VXH94dISZkh6TKNmyTRYP6UV3zGg4wxzBhessXZCX02Bs3D1UUspJqXq+ImKD
/TGKGhu+mGb2lrZlr/kHXsrKyUu5fAwgPPoJCiHojc7wyuBe+v4PuvbdEh0x7Ta2NUSCIHWeUZVn
h1ZtF6lGtuZPd34FPU3S/AaHWPCXc+k9qrN+2ee/G+9E6ARxT4KcW8Bu4lywCWwTQMEE0FOJEcql
jfmEs6CC9I07A8fA3QGoRlyqpB0gK+clBXEJsdfeWjl5Zj72tsT3f8kWr05m4TYmzd/sP13wDgy6
A7OwKtMoWIJy7nL4az2fXdECEaZC5rLltBrWg2cW9LiYOQv+gHRv8WEXoO7z5C91zF1kBqLi5P8V
JTL64p+gP/+p5vNtDGbQzD2A8eWXuZwvUXnEGViKxe4vlOAXHvHTEK23Leio7WZWdkmUkr1hhvsk
uwpCHf6bw+Z1F33DEOeFfdlcKnidBIwkEE5x+dN5D6uUUWDSibncMEijo7LWO9iQzHsBuxNNdkn+
oLoXqeiaGOE5f3voCBbL261jamR9TLP5mY4v5mZNuIAP5MvSJ4rN+YHnSvgttaJFXRMVO6bV+LV1
7XTgPz5fEl17MXkrVX0JeII6JsUC91THn2TKLcdBMvNdU7ad7h3ujsQtZOCXBs1dcvpYM6QIVo3X
IZA701f+w5Xx9C8Fj0iGkOZ/BXo+XiGlkvCBpt1eYq4YB8rcvbrjJDUo97goL8YbW1u5rnCORKp7
zPbs2973tpcOlhgMypHseav/9g1ezE3gkrTly9jsxKHlEeS5EGH+8Wz/qn3odUwAiNkgNvMLWuBm
qZNrc2B/WBtnwHTtTlHdEY1Io3EjB05bMDxqYIzjRC2ixMjEG2LGjn6hP7A7U/t7Rr+AOmEivYs4
ZpIrPPMBjDqa5AyZ/t2Y2XGN1gogZnzSR/OdQ/2JKWkbYvcwCt0HluN5Miodl+hNGIMD6t3CtQhq
U5/sgT0X2uMEyCvKY9lnR/EB6fpCksi7Ffn+4irhDV08CZqQYfeguZP/Cr88gvPH/PIxI6ApgaGk
rX5EZHox+O0nTWCAW658RYBPgKciG4jmUUcTOQr0jSkqi+ZeYHptdmsi70JNsaTHhfHFevzTI3N6
+rarIBXgluOB1iz9pkS7al+tU3sYRh/Sr09SBydMEj7dX8AQD5m9SXYRRwL4TWqJuJpZ6IkSXZm+
N5Sl3Cbm34Fe0T188Mrqq0PsbUbsYoyxdEHr2GelUg6wz3Rf6XkyNp6pURslkUfj+mRS3nW1FQuf
kKkRYsr3IYE0/ANgGINmwOu6scUDmcXMnsIgji/RQ1D16IZ8ebr3fWH6zxW/AhM2OS/kNK3KkdpP
yCwlDAiEUkDm33h+OnUy+FPw7ON3seOdz2gN3t1ckNGtAJTNljtJCSvZada6ZWvrz+JNwCtJympM
V3sJ1Gamluion6kkCN5UqT/R81oOJlYo7xwuTilo9XQR3Qy7bEL8HoHV7aIM2bVu1YXFVNao1iWX
JWV8MMUxWFLW5CIr+OiELtvRp6QFjGYHd/KTXwIHbMIz002VcNPZMNahfDLx4Tw67WHU1FnTlXJu
E8+WMrNj56c9y03DRpFbdxkP4x9SVsl6YUXrB/WqnJ5KiacmPdNsxWurvoTgci8lwzEdjnJVK20n
TV2WAF2IvRbYdlKkJcO7/Y0IvAp6nubp0bbjwrDtRApEkb/XPXEmBu0jyjD/XWYi30FwvHnWEy+B
XscyLGNKSfDEhI6rhanGeC2jsZqQUB0G0nnDtv6Y8Hn1dVP+XKua0EX36AH5e0y/SN/LICMOvTpl
qoGyLnSwmCHtqCzTxTA5rr4cIV3D+8Eg7n8hjlzbeqogvy1Yr1olvb4XhoVtT22eKTmBBj62mttf
z0FaGMkmNWmkfcdMwQjjIWl/npakPxXPaJ56CAXq2AjPmvqf05sgh6gR3mPHYAseWjSdR0zFLXR0
E7FVP2AwImVvscPUKAne9++h5QdNe1PYe9LVc0rK/HVjAfylKhDKggoDya4mxISZBrn551Vg+x9v
cgr4JdBUWI5dyYJGH0BX4ah9D7lOzLGwxL8aaJKVSG7BEkUrbV3nmcV7wb3BZzaEm0qHRxjJGmmA
VlzR8vpeEySnmcXQMzpWdK6L9B6wAb/539UoPbPHxvR5j/xIYGs6q3Wbn4VK+okCQ4YSZM3FJp2W
J2M8sxQqfq4gTQuOYRyF0tiFsMMSw9Bhia6C2Wa1+8SWZ8VZJIjsi5ItCoQ/EQ7HctjGA770mY3L
wtU9EbBvG/TtUtRZiZ7WeN2QS0Ed2N/BLEe4LMs76Jy70KCxNDOMoWoIw8ufU0+ObP/nbMDvo4YU
89wDecMrzjUYFc9KZua75srxp3baWmQK5CQeEJYdhFoc4OF9LrbgZTgzjY4nr+bzzu2bFQj2MgIN
1idDsHisQISo7kZAhC8u1/4vjrRHyAtb/vWmwQxi7jzeEmTg+FIiH+VeK7P/FuKPIxYn7QwfPtH2
8qD+9HFL41mSpWn2TrdklA7XbYZMT8l7EKpsIlBRkNgSdW2lSa/RvQaX8dNdzThlP4OxpKlzQCXn
Kv65qCC6NS4N64LTodFclwVNH+SlujWKc5R89t7bs/0npm7MtVKRRGlSZgeP4kj47aMPG1yhMCeA
9k+T+fgsy+M8XqiiqPhz+eYfSrJyjptNQNbbO9uBTbe5rSUiR82PrBE+PEu60RH7pGoFFHXrVpnL
EYu8T/acRSXiC5BxBhB2CJPzyua3CAogwE4VPhYeORhAHLxoPP/flSoQ5oOJdbZlPDvmdy/qPufM
BFwdX9YIsKtIB9btWLzHhwJ3rP9RUEUNsEztAa/agVsqqE25uGBHc8Oal1FSJeoU6Q5horrCmwkm
4XgsJNoDKMuInoqpWSkoGxTMNKnqBa9JLuPcArZW19bway0jLaqKGrOG69oJx/ibKJpgbbobp/sz
hjDySC0QcEJL0IG2IjnywPuWI+xcUd1cZS6wf8LeGr0jgmsiW4JPPGJcI00TF8DpdDuY2MO7US9A
DAQAejrIm60POVDnUFgkuexoCan+iA2ASOZcj9ikXlYAVIcOU4GMMEbz/7blv2nXrx33JTbJALRX
dFruSWXMAvP4PaW9u/+/ZoN24JcgdZ1CJueQ1AqH/gns5C82i3IfjPHKH3P+c8xJgSgeiIp08tgO
ZFjOl3Z3+F26OxvVykxeZrjOLa4eAR4YTDpBqTuoLvMNdW/pMcgJAHn1sVXexVUbmXcYSptdhY1W
TxWVjppJuGeLyxF7+EC2oYpgtpwGYJe2LolzJiE5R8HQot4UkRBS2qSgPYylIKv2cj3JM7A36IwO
nYtaBW5qi5UGPwBH/4SLA3EvkWIrDhQmxVmihuSJWO205hVkyWmxOEO2SBOnfiQ4Cio6jK95j75R
tfDRBnrJ6JlXRVf2IIavV65pOg3iZtC2x1DWb6GnDOCifTX+L1+tcMVzuJu59hRA1GCUWH9CtYNm
7NJywS8fJwllriouA8HItcfYBWnXa2rK5DRvsyDIuoZJIiapidmmTst/os/UkngOgz40gsRPTISu
ZKh1jSwnLghHBgUccrjVGX3HqdWbMkRNsuProjqzDWNfkjDmrkTa7F26tZL0fpAco/6BheHJ13jm
ylmOKR+ZOlpwmVbNv2xyvr093ejj5NsF5PR1iq8fzJg78kg5QeVkVDuEzoK+ORrnXPRdEPOd4yCa
AkSWnf7VcWLRy8yYM5i6Bpn8EckiRkzTqxoLBCDHJftAMoGihwMNaW+aLZ2XfCXERjN04gbhFz+d
sXyaN7Fq6RrTP0+5/7Byd1lmODcnBESEPW3OcCmVy40EcoHeiqfPHCWL0Mt2ckkgHFSKKlcRRyZH
gzcLn2Q7tSVlMyNYg+bj3UScCWIsdl4kZhLgIFMo4KjdkGRTc6uoaA+t6eLKzPgYHbWtT2eWYEQ1
wbygkMUE6tOsQkizTyFbIQYWym/nl7RuRM6YSzK+gSu9ClZ/dz6dSob8JgcQiQbxl1AFtg/VAm6+
2R/NUIQ3w6WdCefjrKPUzXmnbcn/WnYqAGT41MvbLU2GbeWFTvP+Kal9AqbfKP6L9VPlorQ/uWkU
lNwcTm+XT9beJULZP5rnTfTRoqByX8e2H7q/wm6Se/I+8aGPQEBxS/Df1EK5ocqo8raFmOuBVPKb
WEJ3n9E64y/RQwPwB+OKXGVgMyy9nYf54NaW8sDERoIAAuu6v7hcPZGg35JMritktchZylgZkPMS
kEqLr1OFTDFlJrAifzb07++n/74jh9Z4RS7scJ3PywJZ7vUyMwhH7iQo8xqEicHhL0DivFaCFWwJ
ACkn7yFeLqTNtpFqF830c1WsPBqxGk006sHhB8Vy0hUYyU1+GWinMBw6WWj+mrJidIQ+VXqfXYJn
tEJEWaFzhs0F8G56HRmXvDI7ot9WjZ140cgkvDTwd+JvqSo+FSynYhZFZxpbxcDiV/DjsP/mKcLh
pY0VMneUdOgBVJ75ajWIa+XX2kiaEy9PmWGmiSFBr42wwOzQTjh026V2TgHH4sRsmBKSJ23Qccdt
rEKsbNil8Vt4RMpeP8RL3CBdOquSFV5dZ6ycIhRFOlKXVvmlcPBHUl6abtJNPq8SJFAUWja8UHx0
xwX7asMfGW+iGFWkZ1jj+4LDae85cQZnwr6DcE7tu4i8JKgVUlKbw234J3lHf4+TuuOa6+L+tBKB
WYqGMjloLX++9BQFn8M4PIxqslUgBOtOG/srYcvveCD6fRcYGIsTelokcAQQgYXV2GsQrs0GAq7/
8DeYEVkRcBE1vM05uQes73Q5ZSk2ElHi8hO8YZygSz5lUcLIFF0vRN0seVYpkY+7nVuSFHRron0R
9ioLd4AdoidSj73sdyAGXgM/0oDjSCUfqngTTM5v8URYo64kfE0Gx7uBE8ENo9BSypFs9lgaUqwp
6XBfPTdxAvIAFz+UXZTzxAUHTUR6Dj9yYm1N4PXtNDWOatQkjYHh5aewzhK2/7De5+N5GGE+quYg
pqE2sAsA6XcexkSqUk9nYdBHJfKpdcg+sEivrWhYO2ObIQR44AjPUvqfPX/PLxjgOFxxFm8ZZ0Z0
7OjrNMsVxvvKNeJZRBXz1cUj2LoePY1F6Z+tg2jm6/AzRGT/x4yQkF+Bq9TzU5ukNcboDCk2A0SH
nIR5kXMCwLDLcl1YPmXvWjDqO2gJ0wXDIyZxWByTbd0KkSVL7haE/dIs8gFz02Hv4uj+3nbWj2hm
WkTwrwbjjXRV9BhH1zNKrke52LQPI4Nd+Yc3s9KKUJbT5RtBviL07Vz1suiXrW7e8eYs4zPstdxC
6ZcBT2wTHDTEnUeyeLgWyDmv8pwL3lT2MLZ/RLj6z02mfzTOW3eYNkxx5XkAvCxcevtjYahm/r39
ZTkSnTdS8Wy1J3S9J2tjP3QCezcZ1YBBYdNxlFTO+3gE41cBIxuy+ZVlNh5pUg+1vfVZDg18/rWy
a2PSeJQKBTbQ/ykq2SEmVpXEDUHT0e5yjAE9tawA7+4IXQX/c97B++nNnEQ75Ed/AsoydavcFbWn
cWht6I2eMIGt2MP7YaNrkLo7GPHMVvu9sT5pZHN4y+s92b7JDHnXvosr7SDzq37injQdcRPwV2J5
nbLCVA03VrLUI129Pkbck09qpIdHz40iu2HLtn6xmzHZqpx8jDNfwrvyVa2PTcea2G9xuRNOTFvx
4oOom5bjKjQ/eG1nZvcERB2aarlrtJOObshLazEu92ddQXsz87Mxe77kXvWrksA3YdX+pTuFLb8m
8heIAmk2lw+45rf8QOKzmcC3NMemdIrw/OPKi015M/v7z/cOV+k7LSbuOYLjIrO5gChK2/BBSZ3B
wg2FeMyldviQuGOARWXbpUjXaTYtpGUnUUtYk+rmggAILQE3A0yez3NoYRoFnOekVMMj3lprK/QR
X26L6+zL2wLgG84GC2LzlsMG9+oD0GQfKEICqiIlefyWeTahdqoDBCHFCpQMJQ25fYNTK+ADNa81
oAbscBpa+Kk33PAoZOyiJ+CT+SYEmatw2cWF5pFrWIJS/XnfR6vy796+q3eBb3Fhf5u3xGw3jcjj
d1MtuGqR1AGvvIKP0gEX8ZsRzRZiHX+ct/kSCHHs/HS2j5oYx2JUnlHaXB5+NhK/uRgWoWlUVklC
fatuTODwn4w+YO0nTHaCNW2jYMdavA1HdrSCIc/7487PU/f7FAiZAVK9pi7u8+i7leNzTMZjQtXV
qunddVWG/dpSL14dVuXvLm3vRRVRKDqAILjudRihTIoa1YarZqPoa3+lfnlQiIUjVWRmKmlAx94W
HzYzBMeIx17ckEBOIB0Ls5WGUgTzMnUy00ptMRxK+VUvgdXyrEwj2ptBcZcrXFQ/zk8+zNHIymLR
150RYdX6k9VldBss+lWjSUos9oeFSCgWoWRVNgXuZHnPxvUhK9l0D1ReD4H+DiqkdBuCWHJeOy6C
K59nCAjqnakWXXWdLcLxv2Jycfas2NxmqirgwiCEALc8Q1BiQyw31OrYdi6P4fqVRAw255V+iFeT
98G4tc+ElWZrAsxMPqNSGzRcdF6KI2QkIMIRt0niZ+CxnH775hYAvFX3cjqNCzWs/MJ2gliMJbEY
pfa9odU4n31C2yWNojOOJ8IUesnAuOsbOnxZBiSJURHkWfkJIAIxvX+1UruNRNQdABq0pDJIOSlC
8u6mT/ixZagZiUiy7SRlex2Kg/xqY3Rbxgd95HuKJhi+4FJvvdNoBUSODvR8TWd6NjJ3av+byyU/
W/+ev6AnU7xCEHxAbLBvSNhLqw9TAfcCBEc38+jMOJjdI6AdIN/C5hIKBClIaris/CGT/XkGR4n7
/eJH0pqpqfMg3f87u8UgxziTr+yzX5tpnf4XVf4zaNmHNXzCUiiIIy/NFP4zMc1Qa5KXmVEBFnws
SFGROeHq0hlTawe3ccda4LV4y0VIMPTr4Pg1FKIKoDbKRGaBBvu75cC4vTto0sYH5IckBA5yzUcH
alqJsGx+ngA0PZ23EiaUKHm4t1v2Bb2kHFMgaPvuEILmosiqXP0ZcnPIbRKMdCMbpTbMPmjv3lrQ
qSFnXOAzB1mXZgAfav6F4xkKGkTJJ7zmD7Y54+V1xqS6eE8Z3GS42HqQxokzqziVhIBbsy3YDbeI
gLHRMasaIWgZBhGaO4DC3K5H1e6B9nC+yBk0hoXNzQzalvDvmiMmTCqhBQ+N9sWNqUE1MLn3lwz4
o1zdedXRZJUXVyVL+arjYtHRecM1OchtNPVVv9w8ndrbcCllPvxvIRnpLVR3eJfxqwnpKzQmEiwJ
29XUUrQnWMdsMcMeOZpZaMp9XOb/soTrD8NHVM1yVwUQOCvM+3IVrqBzbr/BhBxQEWPmbzeQj9X7
vuyn84ZI7Sb7JxP0EF/IYihcXybQoJUTr2DqiFL/uNpnUI5FEb2AkcASTy9LpcX3UxtZGvbdQRtL
Sf1bIO+hUrwI+LBkY/5dV7CixVQb4szenwIA/6D9V034a8ECi74PWhCdjtVlBs3jzi+zDbWBhAXX
Q+IEEjdJ5tgmULkdSwErb8P4qJlqHBME0zqd2TvjXpKHZtp08+/NFqnG4bws6KaaRA3GhjwtGDif
lAaQkSHcKKPiDUMwjzb/YSdPCVuHu3Kg7wWaBim3hMJDXRHA8fRP9Frz3WdrNNdwB61kiHaW7SMg
w9XSqavSzbd/HspMiztHGw9Lk2rPpY5jGx5U+iKqE1lTnVkQttV0GSWwKt6HgJ01Kqn7We+ihwws
zXq+wU03KzQ/dGoX6uJSucIMoa//DLiTOcVn3ITSlxaRa8rPIYPSKwqgHu9vzmnVtQF7JrRqq7Q+
cy8Ym5Q/g82MyF/qH5nScXd+OqvPaNTBsY5iy7DpkZ/sSU+XI6lYuy8/A+hR2OnWzKdrEsMcHfzf
7zHZNkPjsEBrU97Jc1CyCHX6Lx5Bv8vuPFteFGrxrqgXY2fUB8o8C9D1bmyB5r1otBozEYHeKEfl
g6EbmD/zPb4iBT9y3qHYVFivQv9N13nRLFN1OgzeF/zv1Q6B/aMJpALJT0Gm6+2GUv7J/IW5pQ/n
4v5hO3gJRAlW5nDJt5z7ENgysTG/S3t6C0RAq3gp1O6eoS/Yax6ucxEt4CFTvmz8DJwrI0cl/6jF
q90MEmhNYZ6QUsYIwSHvlgAL4skOlyTpwcaLwoYOhx2PdJ+GD3G7mWm5seBR+Q3/mz86XlP8mdo6
1/5rbnSM2qHhVEzmOdWV7SdBgVosZgiXodjJR//bXbkah4cyzs/xueUaOWi7tW2NODw2yL9SNz1K
SkuiVc9zr20M3GWKghbBeSKgyMJAuOYkUTpjuKc7Y6EULXEm/MKjX3m2LEqZvsPKmXr0VKutKWjz
OamN1GKE30qkPCNodx3h/Q8p8JvjnLw9cLLO9+/jqlbLsFtetQu1rX+IJ6j81xx1tV14DwB8H9Rn
w9M3RCeUb4eB/YT86GHI9RvUee/fQXjqowH5EIfwnKTR68UEfRCyHhHvobks3QLCUX3y+V201SeC
8Ax/wXCkyOEbWYww5DnhLQp+yTuBuZfGH6d4LMo73nPDx9vnUYEhhR2TEiGCY/fblgZLP0MKMuvP
L90WsaGlusv1ONboIxxbltwV1D4CzIh9wRD6DdAYjpCdmylXPSOEzCsrLWNrV94oItkNGpGqQTTD
MKagPT58YGB9fD2qTwVLUYLsTK5V6YobotMIOe2anHKt+P8Xq9s8OHGwL54Q9cdhO7AsevU0OJ/n
U0TiorOiUI3Y4Zq46Qbybv9PPdZWBhY7sH1TUQ7juVReJYedxhe9rgfEvA7GswpMI9Jata7B14qs
Dzz/4Mq8h5/3Sm6TM7qlRcb6CEIj23y2QOxq1P6RcQlGBLIXqjoyPnX0aKzfROtxVAlMbUOEVaL3
QwzP0y5S37EHW7SbEEaY0uHdiGuXMqufoW12DYOIpoxNurlV90h+FnNcIgTAnvGaw9PeDzueOCjl
6EdWzuIqfVCVDk2q5QhyXjrVE0kKUON0g2PlBPiw5mUbFURV7XSmLOdI7iAtPLchpkxk3zQdahN3
aeYRqWkBZwQhw2dvXr14ySU8VvgkcrG4cSIn2YQmjqbfrgarBd/8KA0FnU46EqRDcRnU8zNIJHEZ
Z72D7q3wpDNvvJCs3GFOB9U7yKAambICUhIEJiwsSVo6GMP25ma5K6RcHteexfkUYnnAI2raWXK/
/SrxpWu979bzaG5m1M2h5/v5LJZxnwdK1fw4EnNlw1PfcgP3J8J2rRXJHaFoPLIiu+yHmas+CRNP
laF9OJZnRQZXCbNi56te+FaRGRXbgHe2WVuSto5u8xRieOfjiWQtQiNcqjkDRcK7QZtSGclciFgI
LZffuvJT4AKYrTx47TuNEj/NGoChW4P4WC/MU+cs+mD+QG20PsDxxVr26veY8G5QHqdHhIJG0RsZ
sy8NjtmJFNT0uc1TEh6eMPPvcZeapzpgBQslaakF4N+iOlGZG3wXEA8fMeMPyxb+gZSMef++MYUb
UgJjyPBEuUg+lDr2iwRySL18G/FFGca7Hlk8ezztzUCMv2ZD4y6agCIf5xMFPnNuBcjQfHZKeui/
Tg3sU6pDcTmzkE8/VQT0JhYBD+ZJxrRC/4E8D5HQC1kZ/PzqF+qEF8Nua0ZdPbNOia3zpUow4TIU
ema86HLsM4V2OX5rQu7LqscyyNLwYFegePUHFMYNJ7IkltiTkghUAhhMwvIeu4q/7gANSQ3fMkRy
sdDnItT7lw7T7sqedZvDCFYGgGgYzKDTh0E1h3an0z1bgmHZ3fHIGW9pcQAUYb/+ii4n/iMm8NPI
XNCNiirVWQPx1jbqW6wT2NeJq4FcadPu8i/DQFxOxoIjRmGm8x/DaiFcNfeslWphVNU7wI+6ZbPu
LLHOWoxIisc8XR7QY91JqH/LXX0Cgvxs+zVyezjxx95HPJ529ioPVdRaavQarLaAXubugJ2rObZe
5chLOAmvLGClvpdASjdP4UUDr+ECtbTryPl2DbpEqSxGKIyz9BNRPjbMkhgBSEMbsHfvf8E1zBa1
YTb9pjxCqW05Fe230Ef4rl0NxMerQ2seiECGQsASJCU2iBqxtfpvk6XiUVcXPfjbzRTel31bih7L
OCpoMOGgo5Xt8Zo9Y8wPci/ldSDNK78esmXi++slLb62SALPqOXc9fJ4gqhwAag0ox25hjpSi921
fkSnqF261Z8N0NYzxL6iK5W3XiF4ro+lR6nZRhItvQRv33pM0Ln75h8c9RZoj4gMXVT+vVXJmY/t
DloLb9keMloW3Vj6HmyM8lLMmZWpn6LUW1mTDJK5XGg4Gz/5Leh0RThfGGi6+AlrzB/jXM+dx65y
SExjPKp28xxHM8qHgcdV56NU1syS+v8CgHGIbnSVmgs+r5cPagtEFr5ksTR4U9kTctrlOxoNNoIc
xrLTeKfzxENQtG+wi9b9wadC0yNN9eQ1aTl5LwSexQwC46xWespbTj2E5ZWOWcrP1W7C5/MpTEhZ
NZvn/rpJZ00NLDUS1n3rlUedKKtzBg30YADNAZxAJr43uBHArd5CnS7+jjXtGmsccP27BURehDqx
OidedNRWjeWhxIwmncGGSZCyrktXcJNqE4vOCslMRBWlI0BUzHoeEDpvp7fKEI3mTn54fbUZgVhG
y0R+5dvRsbXIpZFPjMBWOlu/cjCMR52OAvsjKorNL/6u/F38GQUXzaCSRHuUMudN4IzWtB+F1c0B
oyciHO4YHprxE+ti5hx2f4A2uNpIRFbpEmnmL0duwqKGUatiueyC13v8T2cr1XatZJR1y5phlAcb
0wIfq+809XhIw89xGAXLatPVXSKc9ISG3tfxt6BKQb/1QrIMBC6XsCcQUPUwow0Az2g7UU6IAhSX
lxap5HwAj2Z2ae6mn5kBKpZvYjusLJgGyEpv+qYL0nAPnO1Wm49j/JevInzrxKdnKeRoRkFp+0jx
+t6oIdZmyzVbo2SyV8BNzaks0835VQSklHVsDfd1JIhlhcANHKGN5D2trdY9h/I6Ds6r0eJm0Lhi
iDeemICXSiwsmLT9KXe6pC+4z4TveFiQvrU/o1viiQRzu7UDU1NWQS/txsYuVCgNmC3sEL/R0BUc
f6D70QTk5ybF74mzl7O25jla2XF1y6JlKWPXHpZGD699EJo69wmlwpJcCR1bn0HSWOBYYn+Yq6LA
/+73n4214H0l8jlNR+YvT3yC3klqqin595bGj7bkgtK9iOgqp2IjWzUmQjB6sSqT5SfNKnFDMu83
2VDTcBQYYQo2JEt1YseKDgh8J/OF7JzSaHudRloax2WHjoAd9am71AhdnjWXrv/RXRab1lz8+d5z
BAfpSuycvfpJ02pwpE/SqMdndmjjxMegdHkCMdgZSo4FTrip70Lp+RREvQkrn04lLizDLcLiA2k7
xct6SWhHUi7J5qcwpK4cMHWSnOX5tCGPd0MruX9xFJoATH4LwDfR/oh30er0XLGv8RbuGSxwBsbT
fYJ9sKnHg2Upl6w7fQItl6bmmYqgf49Tdyg7l3IZocQ82xcZ212+YiZM82kYajFfTqEz89/8WfUp
aXDHae/r53E61h4xlhg2EeSBsf56rUJ+j8hXMni+8I04+UeyD6SY6zBdpuK7KEZ9HpEg3rE4p6xJ
BMuQTTMGp75Ii7Mx70TeMZLik7VvMfdNE49cihSw3CVIa+aOiD5+wAUmDq25KETcHJa3hSWjV828
RIG2uncQ2UQkg2WER7xce/xFHiH9ppWFVMREe+Xf+JhfM6hm+lh2XuiYau1DtkpdvlZAa/Dr0Wnt
9tv31va/tEL+kGTJ9tFdrdiMjBriNsVakv2P3hg05hAvpXIt9bVyZeotQC4Mo8yiEfjrro3FYz+c
5WLAI2VTfdw+TByaa/kPV+6KNoSmoB/M8dyyxCX1HTLjVoXfJ4emNdrTK0M4c2+JLAQRzQxFod57
nLtZGjwhOCfN1NTkxE3Kb0wTwtOFCFYILQCl73SskHQ1pAWPYA+vmpL3ixPie4PxCPqQj40cP30c
EsXad1xQJ1NeF6BcLN9FaTeKfAxonhgn9t8GecGPZaWmnhp1EnqnduIpUmKItHgHPjf7GnqOVLhr
oL917+mCK6s21x/xLPQtCDGsKLferkVlKiTCEXgHxY0HFFmsDI2jaYyA2mfP7GK8c+zYH81tjZ0V
O+ckb6Yf2g47eR6RBotTApMp4YXyDfbx2lVUxR4MDFmvlgfRPs1SfLFMOi/15+5HmHv+ScoWaemp
lmK+lHAP+oNUeTIkUtxvgGAraRJySqBakDQopQQ/3v4Zsvb4nRafh67H1iX1mbjAhsSYmI9CJENQ
+m4o1UpdQkMZiCKApjwGnXkxboXrKDXe1MasWMEvjO5r6NDW2MSz7FT+l6cPqDP/mu6EOUcPEhro
H8aGXy1ldk3DSJ7JETBVWK3MQv6GP5pRTM6R3PchQStiDAKLsK8Z+/eu7yHwm1KUy9ABWtIeS+0B
BBuofH5FGegiL3BS2lJfUfzPkLlsl4JldDzTW09kMCOgdrVg/aj9TatMA+60fmPCwTV4b1XtT5c8
l3oyPFYKSrwfPxvx9bG/SQhfWRi9F3EdGC3jJWQ3m0g1DBU0/Rwobmbt0Dt+fL+AFHSzg0u6VBfB
TGOHVxHGZDXu/uK41ToWQPV8vOfjCMcOhHhTOyHdnNKQzpSJT3LlkttHsF5H0v61llwuxigGflrI
G02dYcERwaORmB24CpVIXFhwMGj5g8evnGg0WfOAy6QiPXfWD92i2Z6ZRuZBTdcFmjRkERfHE7H5
AwK0Cr7tXjoi0VSHAFS8K9t6WLj1LtLaACjJkxWLJVvsJ8fs/Zwzs/MIwJMWsUDto+XFFx3H0mv8
bI9F0djy2cTa4Nr3gt/3NZaby8bw3nP89/94ywQFePBynY1SoCF2WSXctIZFoJvjNg3yBDPNLwtY
ovn6BnqN2dyVqlVH/SwqlvGBBENf5kuQOHJgRlKhYlafyaQSeckmRRIsgEUdTYdUWuY5DNffGF1x
FTuxeuUBsK1I9/RvLKYHGHoIU6nEfsHYF63wKyAGKw4TjR/7mffXqp6vy+lWAwQ46FDw+brIzov5
Aa51KQEMziFDH5SVz5d+IVfX1gnNQQSabeHmsy4vqJMOefyuPi+n4B31TYAN1iGX0c8Z3zStOn7q
doS86LBYqo7phTTi/zHx6zScBjIHUhmV3smQOPnGKt5pEy6N7VaE2twuPtLauDfx0w/ptcKNSP1w
w0wSyDn8nCkOgqpjoOuTLXNDlM81bYaEigIFeA1TGjEwVnM1MgBcU4KRH3hoeM7CG9aT9pQzq1CP
Yc5HGFXHUmzg3sfbmYGFHNFQ/j6gnqhWpVKTKoZc5EgVwlF/AOfZTMqaihbjmh2o6Gw3Eg1JVMGG
PIox9EvcPI4RdTsLiVdttwzqAtbBsIR1UcqJXjLdIq7sJUcSSLsdbb5VxHgYaTC7O8FXwkMffGQq
n8qCX3kgW+GRs1XfNxdmnTact9GkVswiT6EfMp7tKE5V1PwbDfxF6mKxZOkcamWFp2+z4GMbcCJM
95baes5b6Orrd/7J+QXdeTlIbU+ZdB9VO9yvVPCzKGczh874Po15IhTxWMuxMi12GdtoNA3F0O0l
nbWrf/O9Z5CGYX2xB6T1TZ63Dh8Ev2jf/n04FkPqE4conYT/oOaRFTQ7xnDQBPwuzzC3tUg2RfD0
rpNTnDi0VI7P7jJFMszf08Pqr9mLtgpcTQJ8Kt7MwRn6BMgcWwupDDFUYwjSFm5ZWn1bHUpVUQLY
N1YM8LT9kw8gPmEwSxCJqpE/1QPzOEFs7WadnrbXveAmS2tZZFo6rWFK86R3/4T9zPSnj3RavBWB
wb76+1xLbd+OT8BUPpMqeZe344fTYzqIFOv4VCabNyNYiXEO4rqINyqqWDEpBwPRaIS6nwxzcJGI
qeV1pPeUY9hfwI2pu3TxhHqEkgmkYZwLYJ88HWT8Cm50WoL5hTKeGBHviROzn6kLPQOmtXZKvhqs
Gf2QxlrcMQ7xbNcggjZ4BRVdS/Kk9EWcJxowMK+IMmz4FTz4iXHqhVqeCSTQMLLujeWsu+vLyuRj
io5e8HqCRjMF2SNwP5Sm+CPwjHfWH4hUcUXwT1rKA5+ZjUDhkG2qimYe7/PDHBnJ8J2DdaFziqbq
WG5mXq65hdI5sV75KLnzjKFu8iSStkefgbWb0T1USnbooTfUvNxZj6DbzSGHkyLxDbPNxWKa3Fke
UOqiB+MWlRYOyV9qvX11sGbY58MOaWsrgj9Orl9p+/ZDAR5/NO4aye1nznq8+IW2xGOT3hA4heTm
Z030qj9AoO0EVm/0Pz70actqgr6eVE8gfAMirX9A+s9KYVKt6MDhMGthlldFK4Fxl/dLdB+b9Jzw
s1v0HvsDD0qRpeZWnRI72dIPn5SCj25cdlenYNoceQ5HX0blfZ6A/Sogt6cnz+DhiMst4A8eDF+R
bVhZjFSPIaQhmrnEXkRNQHQk1V2d0HhoBWQbKAQcp1fx8AVXmIrAULWi/IeP8UzYSuL8otctimXd
XksFICDwGlMsDr3MYOfJtLwovVnLXxtu6bQDCL7VfRw7U31s/j+cVXEp6Y+Ksdq5Tdo7ubv+VN8U
urHwZU5Y0mOvn6hQ29oq1MLMmbWYoXJ091GmrCrOPycJZNgQ12RocyxR8toEWIqEJX4mjk3vISDw
XJNQlt/YQCsLbOp2zSSzKhRTued4vP3ub+C7CldcdmQGfqwhrEJw522nRXDtfBjJhd8Nx7kw0cF7
QN1GlL552ATT+vTJkOTjaomN1F18Mqt/tjIWLZHEboHOr/5j4orJGVNCDM3ggzRB13SAtaqbBU+K
FaQ8gsYwChMVjtMvdUTVJtme+23fDPwE23xcaju5LYTOoUxFYTKn3k3nrJZw5/QNPNe02FMJqGB3
Pqhm0N11BDLffytiuEJH4iNpXmMOkO+mSCanCzhQGGOdeknYTX8mUmD7QszW2coo57ggtoGfeUCf
+Giquy/3csM+xoUF3spWyX2Nl58tFltf0dP54/e6Ipf/tnVCx9rZor1CfDEYEOD08kFtatwPVZ87
Uuwz26ADFSTZSIYXkefM7z9kTmmyFcJ04jmJXT1M0kkH/lSy9Arvz1tltW/FPgjR4dCcx1Vpa9aH
8E/Sh4tAENKh2nv4dys7wSnmWeEtJmb27ElFhVAa1sQM8ee9jfDfavy1bjYs4S2nFKNmWvbQjM5a
S95Rb43QUyBmG81VMzYylr/agTCMPZbPfGkIw8/RtxoqWl33KN78RgM5mThsPwJSewSpSKpRCakC
1GbnWq/40mzPjDGXxRI3rVFx0tzx5AdT3MyLgPL3GGkwaxYMGjT1oQnB025usSzY2hfEPNfgyG6n
3n/V9VG19k5J2tVhKemxMMSyhB3EVprTZUjvChfjQGMaCpd0CLtwD8QPVdPmoL5R6ef5WtZ8h1gJ
7hdoPbssYkRlSoIq0n0SY3nwLx8/DMDp4YROorFpGo9LVIRhlv3lPvi5XofWokZQcHzEYwl81MmX
8+0gS71MXf7yx9VntUSgeUwAs35fkPZCR4lYSPDs2QhzO8x61jGCEf64ELjLkS3oE+tfGXkx3O3a
Y9wAz10++VknbDuWDNxLIDu/Hd9q0+uZwPW9Tn2hG/ss7vgnnlfhVOAVk7UPWx1BxZwA41plvOfn
f9KF1+mpsKu6XFDstlXqKeoBFF52hAQsS2h5osgQIcWPBVCiFOy4oK8FahzxKGrxKiJjRy6Uvbey
Odd8WAiNoKO5WYH3jvA9r6hRV1pADOCwpatzDy6tWKswDQ2zix92KhNDG1rgzJ6RO8bNhKs6SyW3
QThGUiA2E3cnyLUJVJPgDkEYmFS8z8Xkbd8wKfVLweG43z1filJLkFhfGV+pf9a6LjwXJTCrF1pL
3bbL3nn3jJdq7VJ01/uXtP2Bvu9g3hD3TJgCnndyMZHuCavwpdn48u0UDhT7pDJbZcRF/YD84WL6
91fmZYgIzRjrZ64NATs/Gh7pnZdM69t9b0Bzh8PgGRQ3sZD6J2N4jsRjBHmW0WklOuXRVK4cop0/
Cla2BPmV/6YsMM16S/7Z+anY3PINgfnDpHsj3euSAVFbcSnNvrecX6umS4CzPd7HYEWAQ0LlqHnf
5msHwzHSh5j/Wv13oizZ8gLpZIUBVyZ6p16N29+Y6tkdr9YcabWf0n2KkY0pJ7PricSBzNMOX6iF
+kAsIGqN/hztrZNJ+GaVHuyBLSQoOOvshfJVtMZ++sjdD+mIkycoMyi6B0bXmUjBsg4ADCdduN3I
Jgc85kY7pUMKOgRnjbYzJRSBu2ppRU/WnuMlcPsHVaFAGeZjiRoi6qWeUD9nTaSK3SqrZ1Sn7qhp
mPK4M1UN3VS34hnzZFdTUn55+JZeffJpfFU27xnnhHcE6U679vwibzaMJTATmDTrmAZ5e5B+1fz0
+Jnf14c2H9bieXkDHXJAwrJIGTLsW2dJrf2zMIlzwkMnVJX5EndPSvfQfozrgdo0/MV65Bu/uZ8p
sI1VjBWwtxnMCq9SB7y8OqSuL250XmjZs2iEcuxJ3AmP5phoMBQMBpIr886uBro3qdXSfWOtxsdG
90rXrJxjH063tm8XltdYTGFFzh882I0bF+dB+g+3x0aRFP0MaRCuV/rAYB2pNqcCC7sjO1ZHpCIo
oEMty1Q0qMogSiRBKX0qxSbiPLXYHsRqiTPuYA61M1fCfEBpWZA9G6KFb9mUTZ3fP7bl6nCp9H5w
eA2BLQiO3xO0xID+uk9Kto4oA9ax7p7be/bsOWdpvW+jZH3w5OVyInhfXsCf0qkjN+iDevUlavTu
ViCSE0WP6URwqdxg3DQQBjZNRbiawIyyEHLXse+hZVM+8IEx1VHB+L3w8Bxw23uKqhnDYgSkY5Jw
6M9u29/Kn5u8dZJcbAvvy+inRF8qr8bcMu5KA67QO+H1HweSrDHI/xk3a8HlE+nEFikYwFh7msYp
Du9DmgM883GfgN8mPCdWIk//7po2VT/YqG75aVjHKWIcuhtT+2rSnkNVPaz4r5p35EGRWEktwmD3
JTE1TIdqEE8lBnq7LU0Wx3/O3sBJJTuclfFErUjabTZj8tGeQJTIFqjE1pu8FlUqN2MTNTDCHXRD
setFuYdcYm66R+TvNlHoFcwMBGb+bRwqI0G+ysaAT8Ur+CgD2GKZ9P2ZbiTess3MbG8DnLnrgUAg
o5LyrxI4/ahe4bZuEoshYmKVwvjS3fGNzIQVOwkzw1lanSUElodKz5cSL3pt4h9lO2RDy8IZBsMv
3v9pdvIeQFmIyCsN788fOcLq4mCkLSiOuRaiClrgzY6HurWX07RrTWd3uW2OegwkxWEbzoIl3T/+
tU8X3qQtmIj2ogxW7iMGpqVRCGM0ZQS02Qi1xSKiYRxwcU0FduIXZM4/404FZOD0OIAYEGyh5OR/
YvCM1ZEanZpMlX4C3o0sxa3JhQgraBeqlJd7MobOW9HJp/HoBEZgAssckU291/RZPSurb+NAsgtZ
0vsmF1U+dQ1CDzVqh1w83A57MImvmcps1c4SYXsCGRzuPyY2UbzLO2qcPMpUDBU1zIbzaxiJ/+GR
JWqivWZkbRwgYcRyIb2uJwb4pha97L0qI6Gx6bQs5t1L5tH7p6fbINuPVTNNJzbFgyTQjoM0DC2z
RysJuverDN39DRp/zGiBXgdYWl2Z0Rt8ziE00hqYGCSNMCLhvyqECrbLRdQgVnkKwa1UKqN0vChf
zzAT3FzJMoImtI8c5nIi+2oTAPOJPfpTJAVACmbe6Nyptj1CSJtkPV4ZVoTr7k4uu0Q/KU5n/SPN
UMsliSHr7OHFFGFfbV/Bzz/C/ZFhCzXy9ToNAKJBdHSzSVJNtKA75GSCMdv5ay5vCO/K0sXxMqsS
817UhMxGDrukWefZKaXseKMRKoqm+bQiV3468zDHg0tUQq38EfKZnMIfILyjDWve5lvlwADeo+SJ
1wtqfvN5qxafclSO2imURMbWvNSE6iSNoQKqUkaHSkjGvDRtGiUXvk/ggdRwBwaWA+dl8uRx9fbo
VuYWteBTwZCN+Shs6BepkCe+D59kGfSjvPW1/ztqqAiPAkYHqQEqMrMNH0/YRSlqtfxF7trWt8e1
M8uwBeSiq/iy+nCCUjdSd1sOTDfZ8G22gZ2ACTDJb/IhlWRVwCPGgrbuuWBGT4Cnk+9cMcbx+D8F
1SBNYxg7+z1acluzbWeXEst6xZvADOzV26xh6nn2fQD7TO/ZyvJExmJ7K24NUP/ud1RUFPosUlZF
MKQokiMGCwpQVdehrksMXI5hYSmru+tTrk1J4nN0HHggn1t1VC/4+45N57am7HOn9l7eoKFfsuZF
rpGVtwxXLWrzz9Shhw/BNkR7TZhFPNn18uqNN1BiEhXrfDzydRferUUy/A3q+mFLti151Xwo8q25
jFNTgSHT7d1WbP/z0QnveHn6PgkstQ9d4QQVJ03XH8LHOvVx6B0bbOakuYPgyZO25ZZmX8M5SKbk
miyRzuH3+Qx/T8osELA/HKbvWVA7X/rrhOt5gIkFpDpYQDXD6+n+NljQQ2ON+T8MppYq+mSDnmtj
1fLWn8tHuED1PJps9Z5xFtJXfPfqc4nhRTQSnIjLjHwJkg42JxQqtpHhm3HB/D2A0tKG47Yat6PV
mFK8hn4R2IFs28j93V9VUoInJyvORsWh7IF6smPvWc8X8zR3eZk1QGqjml43nUQIYFa7RJH5tAam
kfer3fy9xtEMjlUVIoFskdfZ99Vjve+9qhgSbSvhd/PeI348Qkaptwy0hjUGhKIm3VMt63O/nNB5
eOOBuYzyVrQ/aK7uC4thBLXr7oHIPX+AUOcDzqgMokq9QH8KDJvt45cQf+SWhn9olfX9eupoGFIP
Mn2Ybl0xRrNVGYnYdBQ3bwL8eFg4HMAVFHtxvZFH7J4LkrS0810JEk0n3FtOCkbF0byTAvunT95R
2Oh7Jll6ZJfGZ19bAuuETW0u7ggA48NQNBPlKuXlkbP/yk4tEYrou+Tsccr55ikVIrko0VaXQXyW
F8VgxIP1xAa5xv5cI7GJc8PpSpZ2/HbtHcJcpv2YtvQm74yptDtAycXSmWOrcQ88/9nB4PnvTMCO
DcIjxHJ7IoPQQSO7NrK7M3QZo00p4By+F9ESbBygHLKxWBpbRbHs2gylsKhcPNstWmJtJVI1gcuV
LvaBCxrpl5bRZJkRDl5o0tHk5sSqJsb4/kKOlVFElmozUp5Vfw0AfSsA64eSStCGIEUm2s42JfOI
2twXUntWBeIGxpsHNQ90gt5rofum68z58Ko0+RAXE1Iz2PNrBOFV4cq5ckEDzcJGzaAA7ZsKTPnJ
NidiT1BXfo8z2Gloy5xrwTgL7mmi5KAXnU3mENLtbWAuLknG6k+I3q0zZSCEayBWNZzhWt6F5Ktz
raJXasdaznfsEYduw3hRD66rO9E4j0C3waxl71/DIb8Hj+FAlTKsA//Rd8Cj3ah5eqpCPs5e7CFO
5hdl3Euo3zZUBHCIDDi50UK6rMvEMqTn6b5EDk/FgjeT30xnGJIdFH0svbAbeMQOux5O3t0s2tUK
UDvL2719lZouQCSYhYUcT4UicTncCkAkV+/QBY0NvUaQd5zcXqzrizlGhh7LU3fx2LjZPDoG+3qI
bCY+qtHb9KMvi44au0PAcu6jh84by7wJ1SflERIRyCtr4Mq8pzbNliNTPwDiY+N+N41IPx9TqLtz
7gpdi+MAALbhXinZPYDM1ivYUeEQn710sEtgoS+JKcSxhrV11sKD5u2e/iGwN2J3E7aBCJxrNs9J
r21xKh8tDpifLX4KL0tzf7lZkFmJH8hactJnANNOv+/F681XQd2UWuQ4d0rIbPOb6UYA1ugy+gLm
991mM2xSemMULH/ugx+QD9RccFMesfEt1dCWN/N71T+6iONuFjXJQkO6rr7O0fcK+bTuEH1aa0ov
PVxGxeSMefSn9gbQfTJxMYe6TwQ6VPdLublIelDTVHcloitRKDcc9JOWmFBB+thy7GJ8vx/FgSsi
GYkPAyu30OtNMZcUAZo/XSKkN9/ISl9kwv3g0Ac9FMHTNDV45WDMfYoFso0PLnBs1X77xipPDwJl
rIYCP4lZClFgnoFyUF7rjKjc4QqwmZhol4vXqXdy1oPe69+yScfwOSRjBVUGnHhlsrUkbb2YnB0C
9xHCdMFqbj8nruy7EnjP9/rmTORK97jY7VjovT4YjxqqjyYKZnIrWdLynekYZ78oYgfVbXQgUV3c
4GjSY3d5/SXqMEJIOIZb4C2sT4e5xx0EyD5IAVnWjqztp2BLHi4uu0LnH/7cTmMXdVPrb/2TJ5VI
QkVJLTff8MbE1DII29oJdvw6W1BHO/RZy/Srz3YZ8Ryfqhz5+4NIIgxSDvZsSLUzI9vB6WDcngcG
M6CQ4UIbw6gGxih9pSiFOEudrew/BnHq5yQd+GF4o6ur4IrZTell76a5xzQmsqdsC9hEaHQ4de/S
YXhhz1pwskqJ3EVJRskFWv375o73z6gMjWaSJZ1WivQRfHg2dFvWm916XEbNNTjHuprbP6sJ812H
2UJcotlMqBe7x336zqQPkT3Q/HpXIC1cBJ4+yzS346BK6hufFwbBH5LQ+qEqbreMaQmJmJVLhZ6K
0DMXoYCzoNUcOY5EgqrtjK32+C/Jn5ICAz8pXi+XYlefe8iCPAkTpYQIRJWT/hiH2DmQCfY+B+rD
XVTv5nIFJiWlYJbgYTXVeZg9XBRLWLBxzBse7RmjmFwQ2F+f7e/rB6PxD169m4Q3vX4mcr8vmOgF
bCds8l5AO3/gk23hCyU5Gx19rG3sqaLCkPv+9cqsnHRQ00pTqLrHe1zZKvLu/fZfwo6S4UKQX7ON
v1tNyoZSRpmvB7YqmjEkYIK7u87lUx0ReA1kBo01W5GCXYFx2AZWO0/JeVBU5fnEhOwmlfKp+U8H
GktaHhmUEqZ/NXailjzcFJVeljlXS2FpFa6pOBSJS/BX3qS57VXIY7BiWanNP7SQ0ESDBtMkEuv/
bN0Sgi6Gm8qpFhwbhTc/Cynj9hzYJWWFVb/KbrS9jNJgKfnb+rzOE4XmCI9zHjY6RyY2qvKpaZkn
GQ5HiUn6JLgJ/G4z3E8SqVLasTwHbIo6xGnFbom5jV6ZpLng012MQs8Ia6gnqWhkpIPB3Dcfd2nf
KEIlgV82+2ktI2jx2Mgcze5c7/7kMdvH/2XFgzc+hRMMnN/jVGfKDZqwlybLanFNcTVzQXWOBT1Y
2br4gtzxCKoDeJh3AaAF4Og9Tr2Zily5wDTSgBgu0WSTgKTUMd24AyDf4Sxo3gpnIbB2y3hc6foJ
JnqwD/DIqNEUiizDxGWop53PDaAuDshwof/pGX5Q2xXScROhcpZowwrp6rjGqLmPXG/icyHZlwEp
fVJdECv7vwOEe3+tn/7lghAAxRwf0MhoUArxNWf0cLSITDv7gFn+eNmgw9PjQ5OXVopEuIwJiDml
E9MKe7nSwXFb5GQCYYTm0xvqcakH1hSMksz/VDQFrXKKuwYwL2eQTUJXmsm9zCs+QV5Gm0gz6qHU
eQFx8iI07OPvo8MszSDw+QNufJmR4+Ti8GE2uGKmmBXdiPiTU6J0uS2w/B9GkaUh6L2TMzhdd3aV
79SKngwtrE1lOqXka/Xrid9grMwHP+PBvQ6vDFEehFr6q0nd9KoO9M3SH+atbIhE77TGCTxvoqs2
Rf7T8jrZcMGfnGbfGn8E1Is89rS+ZktDXIj/2hmWlZ0jcx+5tF/uup4y+sVSils0FWEpl/Bt7QP3
GnRwwotBYMF/MfIvLUby37hiFMmuVS+4Xy86bURKLeZOT/HvbwJLiRC67EQ8Ce7qqWrzh75txlMK
e2Ov1nAVzCJnAr13QKCTp3dvOFppoC+RkAnZonOfu8j8s1Cf6EG5B98WkfXvGJPb20wLO0cb3sKd
iggvW0tzz2pvD+7+gb9apK5wbSghwfwWSIGT3a1yEpiRSyhsrLvCZxuYWoJ9qsqyJnViGN13MuqQ
NeoqV/+zC6u19jDAYxO88HP+CFWoaozmY5+ZwnJ5d9zQ9KyLu9JnZi7XvjfYH3jsYuAvYBoznO83
AwS9bp639L9z1muxWYhkzzFDNwAPN26AJ12im1LteAKWH4QrcJLrM5CbBRNxDDjTrrU2nhoPxO/3
/vNEPc9VubKHdmCTkr9m9tlVwHVNcW0VGalozV/GIwZqgZvkOSstha0PsRdUcPBPg8E4BGqfW+K7
tc7UAkZlbh2x2Z5ch7zyOfQIXBsF1dYFNi0ZUWEob1lXPYYs0RO5RrpbEno9MI6OPiyUKa0pzjhz
T9/fe8l14yFf1CNrIzJY01HeXmhKx3DkxtUPqtrRbjxlB1hR6BHtWvmMwrS0INSvih+SpudfLCsY
lmLtl1MTFLeNheQQ3H+ympQKX1iBmaoLaxnpe+G86d1rLsWZKl35sPbZNamkijP/q1Pw1BjsC3FA
eitMXBrkvIQPWoBIHPtb7mj2ag/ZQVUmez4l0gqgnrIaqcaRGRhtx6P8dkrF8Gxv3n/b/JjjUWO/
Do5X5+LVnR+T5dXRqVR5AhNMI4lexE2w/rd6LW50PVE4khMX+3QdqpeEnEzf5x0i79W/NzOE3jSi
r90EZyFwOxOgKjAnlFbdLLSXVJyYmGQcWmkufAp2i10+F+Qj7aMn370NVibhT1iyTUUFZRrHZLGZ
GJ2UFnPUJylRVI8Co8amTDFfoG1fFRFcDZP4sVcqlrnnMS+ZoOwz0rb0R97uhkfE/0tOk+ubV9sO
FAcvXgYLFfpJdHdiQ6wZV3ZCDuBxy0yJACGL/NmgH8iziJKruE4Fc6OcM+B0wuPrS7v9Ziux7RHO
SnhSw9yEDJtNHWbPsQSnMdf3AvRQpEPTHs+foyHyX5rJAxSeaTukKuPHjr70Jl9tLdLdOJwRzXO1
kzAOwvw1p0Df3VcF/LezsiurFJtX1cQrxU74cQt2QKbTiuKWXlWmmxaXmoTirknozHOKpWJW13dn
6oPc2R1VZtS5CLxCwjNakiYBHTOcdaxP1QcNjuLEOW/0pHI8fYa/7fdBmfgwa0om8DYCT+17VvEd
LAfYw6pqs5RLLTmKqjYVpoR61CJSBlJp679mSDgD/XQXhbYmHBuHI9RhXdJ4f4DDCVCD1jI1qvtt
qH05P0Hoky11pfs8hBe1TeXcX6TOvf+g8yNkWrJKyf2pwfZlXzSCbKN3X19vy+cRDS9vq1yyGB6/
cqUUGBITSNKe9jxNmBvnZjVn+D12XEQtcTQ/qg1ZErObytyfzDwqNGfRviY0JQkELC6vMcqHsdY7
ewK1Gls6oq9tP1ZfwOmPoehNgNb00RJMockbDxPvU0J1q05WF7qgngj3ysYK4qQOcWnFZOAu/lvp
R1hAFDBFEF0QvMqS/wJmsfZlyeFrSm/A5oE4bxr5RPO+4QkxEzSs5DXNH+7RlfHBDb7rPecPpHWb
CoppLmOXY/01XHmnWBmC9fazchzvD9lyC4R/u0a6jcjHGMfIAngoMQ/poGnLegD4zoNlm2mYInlx
3Rni8YJApbsjxoSfAzyws833iIqGu/c0W3u6lIR6PxXtvlCmj9hqgLKUyHof4bdUo0VyQgEG+WGG
AxtrkRDl/RoH8Fepj3ZUVxltmFVNj5k4HudxgEp0PAcosPVYLWYrxthqe+NBWJ7pf1S2VOfJ/XE+
xAsbJK4Dsnl1tR+slt+qOZFuIi6m6GTx0bDtRJBpr2eawwOmIg4g83tN0w6aImV8aQyP4VltXXo2
5mbxHFlPEjzn2fUiS0NMZGDsV1rN3YDQ3F9w7dDPwjQBEki+hL0g0KgcBWpCjXKyksVayAziVw/W
YFx9Ih5R6ojVkXIlkI4ufoCMAcqKjguAT279D9nyytCJGezhN+SMtux4Otl+jmX4xiHDX3Kz02Xi
5Be9b6r0N/Fm6ysGTz5SY+gJ6RPk9Xxypr45UValDxZOFdtFnE34a2Ir3yA77JTyNbV05B2EWr9y
fBZBn3yDs7awZzMerflp8MMA0//FT9DvVhMR3R/1kE07n6YEU8F1ewi05PqXjy7v5A0JXvPq1saU
kZ+OaB6YScY+/hvsxtyuttWa2Ylv/2H42j3J7d3N1Y5xpqaSZpDDT24D2XLG4g5AGQirwMG2mDam
PoOP+wpsJfmI/NEcJdc637V2cMXh7vP2jEpYpkVRLhkFcY8+V1ZcMelnxzTaXEItseaTGuzGBK5T
gZEo9DAVk7gH5YGTcV3fKFXjQzpOIO302IatvCIh8Z1pmfLHLahr95dAjxFZxRs7AJpXq9EPMmby
iMZGshin6Q1FyqmcVz8VBD9mLaNkWq5Ml/hw6Cyx7HcVHwSPamiludbbuu+pW4+/htaZwgM8RT2t
NnLUtZXOWxUHij4j0KTQHXvC4Swgec30dp6rmQW2Rw6Hg8b5fi2Yh1TJbSsx1mXj5rQ3WPjZ+Cw6
oNHfqWU64F6Hb7wRA1N3yIEh6vvthorr385QuFmfHxqNDtjO1ySWLBRb8tDEYkTU1wHnsuIs1v/t
8OjRGZPnCNLdamHnqqSkpuMIGUQNWlPPBk61Kpc3DjoLVlD8KJbWPvsXzSXWBDeI0+pF55ZkcKCl
8pCNjAKNsO8tWmF4O5R4D+RTUzrt2ukRz2nonxGJjAK2Uy/n6FXHmP0V5tGNOz0ySuozfzkw4cR0
CqPlCX9Rr7VrG/fED6d2Y8KFFrLx6Dhu0/r9DA9I0gWLdcQYyQSiGyhsnDjmkTdP45ImUNH2ujcM
fFv3WtPrS+WjJgOA/pM+9IWO/IcNv9SHamrMdgYNH1RGhPGXRROLoIzlE9YDfuPTYCyoL57q50CP
HN55ZWVEhP1StxPAwarqJMVfpNHCWIvYPSDJVjNlpSYJRlktBZiehOkC2VPkCHIc2V160pnswdX8
u4O7k2Xocq6TTlR5qxahw2zoT/mRCqv1qBEvE8AcqClvzQFalagZQ7o/HEpBlUczF4/oLiI01+gk
vewCnOPrudS39dGvmIz65LlM/YaoPEIW6WnGC5zf9Op1GzySFT7fiQq+gDpoUqWspl1m+0/8AFFU
gqgwDyLmPfd3ROan1eMC5LDoPx7cBa56Fe3owVOiZ/EfoVf6qYKbFTzyPxmWPq7sNRBf66EpiwPX
TzO9dvywtdMBpnixtyzD4wYt/Q3Mz89d0HLwYWUYIq3EaIhX93zR/Dq/Urxp0xmCuRoZV/0SV+9t
o9duy6TCSJTvYurdn/a8vTGydjrIv8w9TxZAGIVVfC92n9iDOMxFsMnaiEOn3pDD5U9w5U913gb8
7H4/05ncm9H9e9raG4idEJP7lDBEqHPomdqujE9mMMoMFb67TeZccL9KrKpHvA3QJCLucub9wbBs
BI8G5DF3ZrfWd1/Tu92j0kgidFWn92r4hlYrJDNJHD15TkBXhj/gDdXscKWw6LhAvzHKj/4GTGdY
A6CtSXQ0E++kHbIdrmyUrx9FueE+lh3ND/a+eO3QwoYhjNQdnveXMZjS/rslY4yFOYFfAqXejbAf
Q1Fu4jS4QpAVTXUo7+T1XIygaatwHb/sG+1t7lcz6W72P0Q02mLvzG9IMS24PawMPslvR9R45SmT
9zmbEn3BId/z71/1s8D9rjlaaslmIVGoDSBbsGWS7cMTgbCMdUk+yrHaXuxzJJ7qyk2jMbXltvmk
hO7nM/lBh6RscRwrO9Tg2g7O+ypibmDWJdS9rvXSQQ3h9jQiKAfmazBX9Ja5AO/SEWlcDUDmtSH3
2iM8vHTnOGWBpp4+yXvTYAf7TBvvUeK4DQTxJOB3mYp902bWVHIZ5AhNbPN0CyKgVQQ/kGCJKolM
msMEFLxXAC6jiNBTeGMceFC3m5uoZM76/O5pG81M1eSgzGOwLWkuySt6IDlz7jBUCPQaNCYNhxSf
oGqohQP8gBLgM7CLPvG9y8VMchrzyuz7H8bFm/cBMbX5UAuMpk+oHCCgOWuoZ9udHL9791yABEKR
MYiXC+sEya/fqhR6QhaD1krlT+j5GB2eAqe4Al765+5fTxMmlglgGABm9lzw3v/aAM7AsiDBjsGc
ZCcZa/rABtFhof9X3HlxM7nOU39u8xCEf1uimTWMRXHILBlp5Gf6wRCKqlZiTGXi4+MVHQPXYv5n
dqf/Dhtq+VatpTE4PlVGRPCNk9BPK2tcUYHtnGwCUXzGEO36Qqh2qhiqmAXWwXDpgQZk1KWH3yzb
ZN+0YfoZKrO9+il9zeK81YmhBu6a7srOKueNYCEpVRwbmcmKsMSnn2Ki60FOVkUMTn1b2bfiCAiv
LduVbP1Y1xMDm3dc494ajDedGFi6qj6V8xZsWEjJFjlEVvGYggn7ubPQ1i51AA+yhgNcT5T+1OaM
OO0H1W+wUFQSpqONAoYmnK8B8k6macwG1/a+m7wZtGrGiaNpT5jXg80YiSSv3dTrflXuXDLfGfiS
XKAE+TJia8Vf4GnGonreXdIEmmP3732TmciERWzap4Fstim4vc1VnkIji+hV28rVmhVHzbzF+VRF
2OxHImU3JQuv2CAXIm2qrn01Q7ilJmYA6vM60ZhMRvvoCQJRbb5oLFnzf+CznuYlxmGsJo3jX848
RCk4kAXKpalO84VKktMwsW+Q2P7GxNeiauRbCq//KGSaWUmLC5488bbTL1YxEYg8/Eeb4y4D7hCY
8vh5714Ap1V0GkNhkwmutZRvZXOMlx31+3Mnm3xEwrjH8a0c9u92CbyJupmSjWIFV22QJJRj4k0F
7nsjwGl0qKk676y3b1VPSknfKITHK5ZjFQA5NWgH1p8qrJ4iq3a45gWUIuVVbRtQI3Qr9z1ipx68
lHfCEwn4g2zGlt1mjR+wdJdcXIDAwmQ3Vbhb/udrJJ5BfFK57rflbeyha8l1h5376CMpGxh2mXty
wG+iSaGXLPA4m505ng9lX8XjplJN3A531TNy13rNgbLK0E2IeVBoPnc0AIZ/xQ9CH5H2gSCrj1wU
tO0Z1iU8LrbLT0SdAm9ASHOrwoLS0xJLF3iv7aXQGGI3P+Ezou4XcnQI1AHgj3dr+EeYq0TEFhbK
PojpSn4YaxOFbbNhLvmkx9n8KDQB3cx2vDamEh0ZLkamXGHVfNEVk7s30bUupSqpyr7kkDqH+bKc
8SGsw8RRbaURmQbOKKB07xThPp7OdNZQF9z+XVbWYOIquOfG9qe0A5x1Bp/HSP3rxGO8rsvAH51c
osZcgzuM+d2VJkfEF58YCTS3+5oQ+CBX7YmL4NVBJBdpa2bmliX6zOSjnd4ECUtVwzVKxtOxZpd4
RgU2xK83ZmeuP1LKoN2ADeH1B70iG9MY/qiVguDfFYCmLWtPGb94ifbYml6VKz+ftwT7mmIxhg1J
LCplBXXIA2ydgRTiff/0aHL7u1WHpbQnT+5WqBL5SlgLKxqkzZqXUjHYoPpaxj1hunwDVRuwhyig
FRY9LMtSSq0oLNZU3Dr5QZ6cZc6r6cFfcxsTxCHWKa74pnoGsE1E+WLa77hLAXM22Hd7xz+9qedK
Cn143NPHn2zC/acKrzUjxFGVOooe/6X09QcFFSAy4hq4lK0+vD/zeu6caytXmPKr4k/73wPAHw3m
NYjupgqXRo4S70b8wsZD9zHZfmKRs+yRiGa0saPFMKwuc/yvPM3/a0zniuM4eeq4+2DQUf5Val5o
KKVoFLYC6BkxX8JDMkldterkiaCg/YHKUYeaXLI7LhDk8+f9UMIqPP68Xg6LCsff2tu+otuA2mHr
D3KOZVGk+uThIy+OKhjKrn0KAT38xuHSlprpbOKr82+qMzNM/tpW1j8GkW/i9TNlg1l9yNSBI3gU
X0Si3wbZd1zfSNXk5Yl4/JCkGd7M7nZqc+hdlsN6i0lzcMlKF8bsXaj0/5yrS+zBwTHAD5wQSKgZ
Ms2d9N3jLQt8G4h5IE9hm3Yc7I1dbizE2hr97lRa2oxAlWVbA3PnpfmdV9XzEhB55USalhApnLOZ
KiKKxy8DhsRS6SUnzyFPR4r/05qhS3/pHW77Zi86DlEiPC5XZzVc+UQJhjBS6fhhy0uaIHEOr5f2
ZNSbeU4e3th6om1r3lWe6KlPjSqaEmgkEtqcJE5N/ryZQnkfad38QW6Js3gIlHq5ASFX2TYzoLQi
lXhbwMUzSpNJ15MCSn9MyLxYBVASt0WYC9U7mDrBhZYJXpiwCLOKjwVqLOs55EGYuxyHmmhFz/Ud
doIentXbEtXaGHmZfggFIIqD1FbvERDO5sKSlp0GMwXeMXm6OMkg1gEBb8cwi50TgVfNT/RRllMH
pasIG1S0l0dowgWA8iEosAWgbPKyBSLGBHSAPbFlGYY+1vt8XosnOVOaz4EwDDrP/Pr/Wk5/yU2r
nuNdvu7dDGrQvZDekkTdqphGtHPbXd4+IlPH7hKC1Ykr6rVODked6zDC3KJncv+MgpIpUxDjnzSP
+Zp40AU8/NkBsn6vEUpFBwY0+pN4Hc94Qil7dm6lSWYH+qswq05ilojPRVpFWYdtTbRhngCAGij8
oXNsXivjSca6XQArz472W4nyu9Nm2PdWhyZJZMPlgBUhC1O2e50U/URv1subu10i35DQ6O1JNh06
N6C88qkYQnj7nknoTTHLZoU78ORn2CBvgDI6rKQ91WIsyJcWW+Fxu4cs6QywzXB0ZZ6xpTRO6UdW
dkNllSYk+RF1TEr/mJrXTTGqd1kFzMjKN/IgaybNxSi3vJozoRfWdL3t7K8v4+NsZGComXLcL/39
tsk/faur1n0zCBsJJuvLUe3x53xmX/Y1bZ5DrFoWl6+ckX7177jyKsrBet/FXm2EY1032BupiNXE
mhs9/4Fl1EBBzppC3R0uRrZZ6/FQjn17wcBx2rcjPUIza8rtrgIAfLlIxQM+hs5b+E2+J73o91Wz
GkRIxzlHKJ3mIKhYNgk+Gp8ZuEFC8QpH+64YGf8GwNTk62eD5Clkl8uZ2IjBb+n725lyjRFDD9Ye
g5hqtEU8Z12nbFmVutE+ZQDpsmolGzR0nIcXaeAcfPdjT3B7VFqqio0o5aWPwi291JLcvsKm7Z6K
s+jZo//rAdpZbxwICtH4rcFRY/hpRBALIX+L9M8PadFtGC39+e3cz10O8o8baB2MQpzmMXs+HEYu
teP1ass8HBgp08RqP3vTICqscVDIfz3CuITPxDKBPBfz6BrjzojBeKVqY976fQ8L6gcvTh2mIKuu
Tht0jO+McJzqoeMmiqHvnodyzYsc7JNl5BNnyfIh4jx5k9pywpUYEij9+0WBlndKLGbtwmK+YLHl
sEPhlYNKHsb5l81f1Gu40H0bpRFXYJAb3zJTyDOWuMZvIwK0ZlGodtgZDOv16vjfDPV7E7nSlWdb
98jjCSHTXQWUpnul8+7Bb08DQaV4QVWrDvft2MEqyVOsz2viZqPDmt/RChM+yitq4d8BIYwwGMvS
+pFNm/gc9SGBxI4WTGRLJnzXlY2kT1GKAi0ytG2Yq5AqSZKG/iY69Y+TFa+MoSq1+g7RIq+PgpA/
BGRQG2xgOiEeYmYmZjDgFpZVMa4rviob4+eyU4yGD3u6nw8KzttEQkwtRlUexvCkyujRDyP7lk89
a6R1LalmUsCRLzeJ4YMtEMeS6GFBvBW4tcRHgtG9FGPfoyt/Rzg+Y6P32ewhT3ioF4aGGE8hFIE2
ixzWn7seYEsVoO2xIXNrd+dhhpTyiLITsVDGlpfQCDuARGTO9gKNtRRQfp8MfxRLRNzbxrqEdl1h
qfc24iFDsHa0sLhFXXmArgnfSeJ3yfKC7eMSPEGXvE9EVzsNtbfxRq0/DIcDB4Ys23hP3LYDHeNN
LcT/E0FXUYGysZyuhdnhNeI9UgJhEUr92rSUky5w/IgHYFJOxyGG8QUCHtiAtmxR/tjt09co4bMY
2ae5LXtHpt2JN7+LlTHcTBRkGSqxNqCXMZynh6Zb23tMmTpc3h3pImzSa1IZKl8mHAs8ck8UhxtN
8hwVyuz6am6nwdpd+/ksH8TnvPVUc05m7QAC8r53xdG8HmmlgAmiwPyuZcFim2kHGFc73Ee2ZlCv
yqRkskFLnvhCWq1ctgLTRIxqttzQiaTazfA4LJEFYKJM4oVyCpiZvPFea6VnZIy4a4DBbqdZokyQ
ZORhbt9Vp4o+rtd2GVU6offTp9J8zO0AOkesv8GkK4rAmCckaJYpWRmY126U71C7++ghGxQUGWyB
6eUKtZKb/3mLktlyqt3zo/EMkPsD/TZ2rX/NilfsumueG9I0ywlWK/MW1VKK02p9Z9K1CVhDpR6z
WSHiV47267ef1bBOon01RHSnfdifiWRHHsWN/pXw4KsF0iOeuc4xXwJ+q4nSry2wkIF+oTGyHCCk
VgGt3uSGIxwY6XQzXKPy9PlZwzT0q9B9/XN8oB7kNeQMPYsgN1vfe0qbikOOPheg+rWkSbB9yYOC
i0w78XV5ID/tffjRfEEyEdEfA/CszJKtmWz16mMkyr5yDrU9UoJrhyj/N3HZf0Xzu9/m0nKQMB8H
qi4EgVHPxxVnqDlv6AKrBylBQqoSX1jLbXCB6CVBJJU4idURBK4x+g6jcTciJw0Qjh0pGME7+ZbY
32/SGtaDcurAs/3uOnqjBvhKJ85JWH8+TH5p6746xyczP7i25fPZyvf52aJAsWVSWehkHz/PEOEJ
l7U2hOhpR9yUlDMKyavGCdgOOWTX6c1c0XWeqphjHfTm3TwpiNmhmzuqcc43dues6rVdYq1AeRA0
0UihtuPQTY2WB5vg4DbCnAKr2hE4GS+e00gMRB84GTYx9BQZbc9GzYezOuOvcOdXMRr6adqc9Jey
i2Nrchp+2LfHonmnwk+a93oWrAG8j9KEvzH6NPTjAOlzZnfbxzhk42SGtISag7wl1yf2wFNqLzQK
fi6xXdNhHNO+0v9i/YSBXBVhZyPKYLeiCBpsK4XQMtn/wjj1WeBKHjKotMaPMsvOq6U2drbY2jbj
ECCWpf7S0LbXmZkABqLdn30SH4jr4S3z5DYZcOGpZRr2yRQSYuTQcvxF+x/xItScEtPxAfAa+CsO
5RAV3oY2lTk1VQI14qNeUIY+7UbGZ9a0P/X0LaW6DZeU5EPzT6R4zJxGJAnwZMgZxRQoXYsYM4qe
7NDgWwl0Yh45KtYxWTKc88i4++6hP3FwyN2UXHLgMTaUhHFu2K7DytqzMUkUQbvG6PfaktYshUPi
vk/8O97EJ5Z7BuMvlsHUYQdSdDRvOjwr4MmuengMVHBOCVr7L7Xj905Fmm+ZJWONRBy0AIuF9Uey
mo+69/ZOXpOTz9AZcH74WuoiTbjDB2i6BrLAgukZhyiTJ8Rlu9PZTE/RofR+Zjp7N38B1jZ+M5wS
PdWLfj3eCqEHsvzLEyUJbc2USd5xF+tmq1+ASeYDjXGoNZd5ticVq+09DPfFHShvBBGcumllH3Fk
d1f4fQcavZMkDt0xOP4v8PeIpjRuOLdqSllvJHQY2fiwcy9WmKVv8ED2Xym5m3iuW655oPowEfRq
CAcXt09BjCzHveU7yhLX+/dIgQ82oHC9Up6S2KRqVYIT7oMNLe8n49YTncNJYrcn25vZ9VVfzMjc
utc+0hqvAIO20taDIVyuPhLCvGs/yG1lJdC8cabZOhQD8ahXxYlnJeIhQwRTHpg6LxoID2OfShOA
nNirk5dxWdvOtlFdVp9nTI0J6j48L6O1IQSLVBZPOBGUxIlIV/RFsTK5xMXUzzFV3Q40/NKW5Soc
QZfBgtP90rhJP/iBk9/3+xco/n1ehhB7ud7XQBpk2dKyl9qKvJonblNPVmHEPoFEvxdZwAVsHQTZ
fVnAcOgGMh0K1rqK6DEDn4sbmw9842oy0v2LIBD+A6py6RSIcrBvrnKNd330ilBSR8BnWNDuV8fk
IuoXHMFVowyOlaZT8FoCbYugIwMMcnfGKbjpgmC+cSzckogt9QlIZL45m7dqwFVpIrJKiKMtKHXZ
TJ/APpqa+/FPz1izsrKZH0ZcbmFgrJ28ngw2S2OZw2K9GAiavtRNu21hkXYpHR82dEdKYu6vN4Um
LIUtaLH9/zQocVv2w7efSWh1+c2aHZGOP+0I6HArz+YPFIfJL9Bf9oN8G5XwaTSwkb0eg6lCt7fx
YAEBj3sjNH4vBIj4lyt1MSKvoOzW4Brs1v6v+hsHVbS1t6dnUMdL9wQkHkdE/m0kKrDE0LiW3Lks
/bw2AMxBBA9PaFl3BSvtvUHDh41HmqEjC/LrhmIaMiKJ4qZfAs3MHdRIhnRjTwDE6LQROkjBAB6y
476eLOGOzLBQOn25xbB+KWKomQuQOqeM7s1CTCzqk0NbupA0CLDf3+QEKebm5dl6HD/yqecBbEwg
ADocyUUHWqdV1/i8DpnOPeMGOQHWB5OrQuTlDQ0DO95LF2ykAl5ax0hoP852jhG8AWbwXrucC77Z
p0JLguekjJlxEpCxrYmjbKTiYMeBQnAp2jrhnQR12OArLDSwObzRA22UIbfEVcRoFarE5IZw/Wxg
ZScmzaqV1QkrCj6+sO4/xqZVb202hdfSmZMYGGfxgJz+jKYhjvDM96tTffbBz2mLvZomtqbqD8v6
+9j9sOJHzgzChg1HK3VGpj7WgEhHWY6qRGTmtlexT5F/ro6n0M+aOUan6MpJHIoxFIpeAVNZdHNh
A5sRqPXi/j9k/hqT+FTGD38sJSktcwyN2mpDb4mr8SOscYhLy2GgMPs6UHdaJ/jHkJ1IB54dfviY
e6dfSXsuEsA/lyAyPcQDDUWZhnSBP130hNE+R7a4GxWhESSZlNrCFf/0UKdOjlhM2jZjVrDko+MQ
oCduPaH+eVc1B0jwkur8BdvAlTDPZgqUEg43z8pCcsMY2QCttR+XgeJbrGkla04zFgk+KBmykSH5
IGDrCl1MXJhW4s4QzWu5N+fBUMHMtWT14VH4Vgswa3wBx2/xrY8O6Hy/cr9eEuJLq/c6KKLKogqR
o4Rgw5Bpx4G2ljhDtSAkY6rzx4ONJBtoa8D+0U1cjhPMxmnEZ415Zh675VasP0dbRGVd0T98oPkA
BUQD66fnEzMQJtWw8SwNQ7A7/p4A1aMQYr1Hu/E5BbqtJ1SwGMXdyuAzW6h1S3lSXhvXbxha/hoy
FcjWFsssugxp54SMGyIHnnj4BVW7iPr/GDxLLjOPpzytsf5FJ7zSgrY5NwKdO2f/K7O46xm8+0SJ
0wzL6FE5F1yIl3ajbGhDzvHQ5K/tDLmWzaBNWJIPy2HumwZCo62VGqQ7j2zTbTjL2Bv53hKDyaq5
1DHTGtHXDVHwjfxWZdYBGBZt3h0Um6HkAlDW0cahahxnfSC7batmLGqwsmanBXWp00Ks8vlSVXwH
XdN0MgIiEu/zaFDGcfnjJOXrAkeINmflFV8A5NAd3HM4fZCj+BcZ+xavGBiL0KOOPLdtufHknXzw
twMsz7abg0HxP+lm7OYOzT6pGr37K78VWJgBVy/ajNsi27RTCkXNVrA1EdGyoqnzBeNcXY2IP3U+
xUszT7hJbkC0OnEb/jchwgQVdSj4akyLtfidP5pS8xDzdCK+HpYe/tKDa4fevacsyt0g1AcxVJd4
ExJPbIwoKfd8vHf9EyOLnp5AGTwbG0d6yipEGvzaaZbBpAhPiq8K3dOk8ZZALaoWbrRVgbGr8mKd
GSbTlfHGUDzSJnQieuWR73eyGM2aohp0+B15rTLp6GwW0Do//5dL90GvZewirBodvLkd5/bZ1q2x
K0jf/tQzYzQoUaO+SoOKxLRD7aKG+Q+k9k1jSwPeJahwpGouyDzu6DfVzmqWWYthYMj7enhv9h9H
jhT3wMBIhkGUPa9cRqlQpN1J2ZG7JqAf6QEk54n7VkX7Lx0ZN9ezsvZKW+QUYFkwqvSeQSf2LZTI
zrLRtTnx+SYaASHJ0MxQ2pHZgm4Dcs4hBirKm792WRTg7zToW7lKuyuilp1Q6NHjbdSJfbW7lM3/
4D1JVHVoiyCSAOF6qfDOsiamLI6JkkI7r0akg8nAfeYFE2lUvX6iaKr2N6dQd+1Fe80Og64tcfbf
TxioCzZ+kpYLXHZoG0a1h9OBS6fFKK9SgSqnr02DdhuiEhnE3HjzNoCEjg/1DI6TvArscpIDUQM6
j+mm4I9oNmT152B3hX/br9tyFdIxsJSMvBJUsCKlhFugazW7bUiBOvL5Np+rI/VULEovVIHgPBux
+deOrmW9yjBE+xcG7VuocymFkZns3HPixmcSDhPgB/7LrM6ATf8WQbgZMvdDlBRZgjXOFA6yNAcj
AIfmXY+J297dOhItrLRH2FzdncH0/j0RL6r6EHS2KjbSfk04UVIHob/tR2c2LDuhsnUvhpSegi8b
kOtMTZz5vI9iXKxpEBziLmd7UwRZVl/4EXDep+7rVXXxk5W0d8Y7Gg9skdn0VGfC6iQ/G3QAevUT
YUhWXSz3RKRlVKDqwSQBuXFtDXidcHw3O0sSVowzm1bq29MfTR94nDkAjzzGzR3Qnz9lh7Y1rl+6
73rwoxlUBYLG0oxuv2Qi9Otu7ba2m4Q8cg5cHnf3zlg6Mops691yuM0JpesG0dWOo4tbZsErgKR+
RrW6CpEcm1u0uE9rAzi98racaIhcd06TBOfR8sjz5FMPH9npzJGInvpWet/34kSUEF/hKL3Udu2n
RS3v5iHyAr3obtbvfJhGkoINF07NvDoM5ctpKbRob5+oQpRzIYVDbiOeznrmUM7m1Ir1j4UGOuWb
rOSekt0e/oHTn33PU5G4lcGNxjkhevOk3vpLS5022iJUbmpXWYAuRuzigbfys9qse9FCldWuYoRz
BAIqrGMcsSCOKcnhU57fy1nW/Et1f9AiVIPHbkmjDRQn9lfzBmnsRlGNkHT51eVKn/w7XgvmZ97/
+JqMb7oq2ChUuji1zKLasE4QrDe/Lom+ilR4aQnd45YpCTViNcjovxrszKx2DSGA+HeDbM7Y3g9r
DgxTAbT754eSmiti56gu32LihbAcrKEvTxH2waF9ONjcVZofX9Irt6PihUmYtVi8h/Ngx4RRiJuY
g4Lst+BN+b6OIMoGIC9QxBkGKdn8/eoQnlVld5+ROdKvoV+1pMdY0HTI+jwraVswB09iQZM0Xw2f
mudiko3vHyozleJ/nrXfPu/QbpatZI1Rna3U/W1wcNjmHwI831+5u52soLz/mpYHX03rR4easHMr
v019YQ+CILaJzim4AKa6I50w6HTax0ndoM1g2KYJitSTDICZVBE/wYrgeHR7/yyjQF9z9BB7EbW1
E3gOgHElosCEC0GqspdY6/YxmS3l/Kzq3vEJ/SI+1RQc9tAVKnj0KpE1fkGOs6c9MeSz+VH9j7h/
FNu1UoMJZetjzQjSKd6y7N0XcSHgY4DCDhew5jJvgWI79ddyCs8uR+LZWbYkHtfqcZWqJK/PObGL
HrHN4OkzUKODFbNMkYldGXbpFd3ljm8oyx+I2COdtD/y1iapA99XS+aodeu7qm14qBl+CLe1Mams
refwl193w9jLBMCHhOvC4WRHLoq9HW2PV27q/UBcljZuO7Bn/4BSyZhi8f02QqCpD/7AlkTUOzfu
L1aNwDhPIP0OoMC68Qo4fGbj2ALfthikJut3mLPVh7sFzh9v6QPJatXto+/FX3qs0gjaQ1A7uCm4
jplKGSdspSiMUct+VVvFPJVXOR7ykKFPft+EHJGN6vwmEbxKSsbGVq23yNx9SAahBZMNgkaH2jY/
KWeM6eylyqJ+KxWC8rJgM9PrVIPKd6bzbe7Rm/J3o//+3q1u1rugAFPwkANgY8FcSaYEa6wtLQCD
BapUCkV6sWEb8VeOuH1n3vBQh6xKSAjpduD8rRDhCPed99lA0sJC2kLEO+dDKwYbLP/n5yhQQ39O
xiKzg6+iRb2mI2MI8rIdlTMwJrolY911graw69imxzDwhIi2CHcnEKysuqVp8RbEOKKU59gw/Al6
4uDd6NzKYvkmL4oGu/tErkDZRaE7Vvr3jELNvuKDgrORd4hBMgBO2t0WPmKfSZBDmHyP1AwcKQhr
cTcB6mslR/BW10XjtHftxBb4QwY9EZ5B4Av3v4raa93B9FrnqPvSNWkDXTHxK3G6Y5h3Nv2Si5Gi
e9+r2/0/kfdzH1UWbZ2svyuEamlpOV81Ukwxxl2WKg6iHF3NJ4L4zxyvm7VhSTuqdP5SrUNJ/MyQ
C7cNNe4Y9fPTwVP0FxyYGAFVnj8tHAQIfagyy0BV+R84FTZlkFSZhU5fjmQnWr966p1HqDBd33nL
eYs+zYc5hS+IU3ja4OvrR3POnfQOV1PwtHdmFrDwTQGs/lyuF9QhKyE5tXdKFrnTfoxrKK5Lp8jI
h8jayGqGuEL++vEPomB1JDJLcP5mmVmV1h5EsbWoDfarnB4AfD+xrfjLoY6KyeaaqH1DUgM/Pdk8
WuVz3Vi0R82bxu8aKIjnZ6P3L8x9Nk3NEBG8oWnQSxkFIwF3HT89swpWr7NCzMOJeaEYcwd8nHH7
S09QSS6CAhPFyP9c6QQUVhIiXcmhPGFNBGp9UKRa1v+lUkISlUkbBoE860w006AlYdmMv7Xq3RA1
YHtw5SvatUZtamhfUa1xn9a8ExrfM7aPFnyoORzSqGmaZxDFAWYCKGvQMMWH8B95p/BBkF/oFd96
1y/MmAkLtVoW6WaLpSqb+7LNRKjsMP9uxUkLekd7lx/UcKl+LftDbxkoPG7ofFu3y0HFXgZAMyDN
e6EDrCQVEJOeBRNcgpXn0vAqGpwndZtJw8ABEqnSRyUqSzM6ZId+98iCTFOVVXfy+rndPYlCzWpu
lAUJzp/QRKDlCm+/NNcSheU5gSColOz1ad3X9ujzYNzyflchA+e81BHM6xAtfjTu1pjRKXLHyPR9
G82iGCgJ9wweS9QfVJPrWxoejocHddkGy2Y8fWufiaRAoLgCMh3nJYTN7pMmOrKD0gEs6HZITMZG
5HJ9gC9W9vPCwJ4lAqVE6jyqMNk1k4Sb5CZ/lZmnPF5WdLvfP857qsEi5iwbd2rWg1k+xjQ8GZDZ
es2adanS9RJG4d+Ufylcctaw/hkuQGT1BGAyQFmYU3ILEMslcgHSKvXOd1a6ShxBCy1eBYY650yD
xTWPO+iTKJJX4piCYYk1fAJOQ8Y1znb6YHTIaUuXWurKmWMdbn0+K6SbBW0Ign/eR1f1QoAxiR80
kr4ksIySWxDEPKqKFEXPBlHod0pRphe+jEXUNYqnQuub7KBK8Uo4lnmZknBjaOI3+OUdSYy5gDW3
e8ykSTIjkxW4LQUsN/HjYHSxDUOonjqzxb87rXvmwmMYdVQMhDBY8vE93CD4YVCWXbmjluqfr6mu
dfJ/b+1C28QnzyGtqRW0LoNJbyvaOqAdc320DVN6SNuPh1zx/0T1EOWbnkqUWbMYH/MhI+TZXDCw
mjBqdd8IkLvaFUm2RB0i2w3NsV1MpWprq1aKRWfFG9O4+8F1HkXFe8Lc7noKsBqLHIaC+TLiLMZs
4eIns0L/S1pqniX6RWWsZNOerH1wUy5ed2z6y0bYKZygyH3BqIV5ZQcoehfFKlSVGF2JVV/SvSXT
sbhPvG1p5eDsFxWO8m9Zm1mAFVsVgkhkGIy0crMCIbgJ0dLIdvpM7FypoVVniwJkjPgzZlcF+CXM
54efSNa3DAOO/TvSnMdqzd7n947COU8W2N8ZtsnUfzLVEqR6GcTnxqGgWdInjQtd+eTlVyFjbpw4
JpaJeLaMXd9hOO0vPyqrBQ84KlsQzCj64He1ON+AUD4PwvUEKi4zxdvradVF4jnGz+vpCZParnFx
gJZYuXCl0izt7UNLtoyhY5WTucqI/6iWv2CzdHXdYw8JiXXzvZ9UgQJSQdrwJm2CY5GLyQPUUt05
xIGdfSLLxKxJL2NT74jR+g89+5vD1uXV373FAloBsbUPzarZtyu7AQPcfmdPdVDayCNUynw0Crvv
QhXvLg7/2Tk3dUmKHbeGbu4spUgfPkbvy7FfQeGSpZfnf132kp8fofqHz9Kqmfa7fNfUh9ssZgH2
k0coAkCa9Jqr+Kya86XdtDtgRYrzX99x+68hw3ajR/Qvx3Kq6sCb/euwAx8Ry0JUejAbFlMPbK1y
KayNp8ZaQwVyD4083PCviN55Q/loAzKke9zUgoOua3TvuM5MEGyxPV4EwiEQud72oEonxTAlnN90
uCKs2Z/16dXltTceZcSJuCwPssFvPMhFigcaYcDXAjiFh01Nyt1FSgOaOAWsHX2P3Pl1dv14WPgc
pfgiN8S2VUZ4cdfefGHsBuPIGBvq2Ekqmhhtd3K4HJ8J7Dz/G3lzSWIbHYF7/i4S3xr+RHysO47A
/7y+s+gslbSQ4masu2HBrz8R+QpuljLD8QML1/Ct+AjRWEsrmy7YesIUIXzrHEck8JISwOEzZRn2
vIX4HjrlUx/8G2lIC9JiE3pKyHCQ75PGHivDne6868R9+H9wXXHakFf9G/8Ozg5GMgR+8EbOjyKL
LSZXhPRWSe3/R8a1/xTtNiLaPaTSsWObekbuPZKiK81jgU+2uoEBWvP0FuZz5/u1prm9rjE6d/fw
SuG361M7JgDYEly2USkVRvhTWtDDgIEjgg5qG7oR8KnigrhoS9fy7cDBQ8XtZc2/X6RUwETDIRsU
k18HVOnL4S0xIZeQIWyYZ0b29QAJSfkDNGiU16bLrrLCbjsSS0z5gqAak94p2U/tGkrcRIrVc9xV
ECMiExrxY/oJ/PrUmnP0KJaEDLId97BFqMJEWSUnb72QOOhL9yifKkgYyEvPZtAksodLsX39teD6
ye0GZAvl2W0y0VZ/tdWlFrHDqhj5NcWgTQFpHWUgDT46k1JLEXNPPgfHPDYEk9hL3MGkmcT5obCc
R2tSnKa7L2PfIV8l1Tt/PjssGaR4Xxnwp3FGAKT6HwMD2Ypoz8e9DUGGPyaBqgtmyILkdDg/kWkE
a+vysEfnsu+6JlyjDpksT+Z6afm2QPwk6vhVsQQLn8WasgA4NcS8DyRIUiqsytycsUl0xmsX8Mw+
40gkHP2sPNM4mslRpMJm/kd9J77QwgSEK00w2oS/S7q8Hg2WASQlQu5naKppXKtk1tzr4Br4eho4
ErVlYtdjovARsMPkr/FLZ95YnSGY5twAuwprRrWLQef5EB6LD8ynr32tWv3hu54Yw1T30fkT2ZN/
cnEWKywDjBfK5v5NyJvykjQ/hVNps6qOoua70TgABvPZ3OS7p0ISHZ/haeVhap1CgiyKMWxiQpIU
QPIZm7cAzT9+0WiSPlqp6GUj2C+11k7Umx8ca2SBj8fpK2x4W19mJsGf3sxaEbCLoN4GroO5tTs1
p/57v6MQx1+81aDRwvFX0KHa/ntNgZozWtGuXT7qVd7a6U08mf+osLkSsgNCFwSpnitAovF28fV+
sQ2gdJnazlGDu5Q6shcbEU7M/A0OBfenSKDk3pQHtvwiI8Y3f8CiDk2PzFUqFrKqqV/+cy+z0495
dpRQQLFeIVtWmV8Vf/iQafuYN7ffVf/PQFjjDIYcBzQ6ZGGf9oVi9MoCQGB0qTCtnBQpG3Ag/ohg
QN1SHSC7CADE9nt8xg/G9k7+T2vGF5+HAMpTsTVc3f+CBMk855B4HS5DmGeAuOPYOv/gXbfQyisj
5PUk3ZCl4svCeLKMja971J6NxW7Wjm+GC4PihcTFK3/B7Zx+Ovls3neVQQZqqWwiVxnZBZWJRQ6R
bMWjvjoSEew//0tXPX7GV+PP+1v2bzjHuwyVtPefC7hL3b81omOwUR7pP5hN2H/Q5TadQarjz2Ct
tD5jRCiWBiATgh8uwgwKdIqd8DUDmdLV1vdrNOH1dd/WoXFLtn/fU67TbiAVvIkhm0Wf5f2g1BdZ
rrOVfKBM3yDz4cBnokxdumJCu0AXdppS8PnrzvIDmKlJpwK+tTDTtHzjMs2oV7grSGgZHFSWjVXN
ys6LUc0RYm1JWIvFzVrGfqWbY9Y6FO9gEd0jXwpYLrn98QZ+kverprRByFcb3o+5YdwOGd0rHRB+
BS/u1e3c+hskjN02eTKFZHtQ0XI0YAwiv8+2rjuljPW1JAnicRl45ip/sAIQwpfNpUrXjLo3DvFa
pHW3BhO5d6VIsNmS2ajplpBBNwNqxs14TcO0TnmvxqXbYFyPzvThywNvNNk+DGMvVtE7W9yP+bBE
Z58eUFVSujFOkpPxWGL2gCCssbE5zyDTPmnDqcXNo1wboe6aspme9LATgQnmnxz3v+bm9FONIImf
tadhK+r5zNoQ7EizlTehjvNxCoJYxvWnROd7EbQ8Xles5FOYtZivZka03C3Hr4sUDigd45hkIuzD
IBEQT6bb8dTxTdbwx8cQimEKhWUV2MUcLpiJLOChRwk6rLIj/lOR2IgFc8uOrw6/8zVmF4gBI0yN
ZVOI6ulntBYuWLhzIieYAe3SoSZGTly/vnsGRlEWnaG32mzhv5gnuS2rIJ5CTQ5UHM+J6yroEVY8
9N8jqhL4VP7FfRtN2V4pNVNyXVuouwmbLYZ/E/GEHlUt7+yPYoVDXYX35ZNXDcfWiw0dtH7G0Xes
V1Q0JIxRUfjhSVKOU1dQYZ4qx9+MvO+sEP4RlaH5G6WqozJO95D0EUoozdL1F4n9cZeqdCI6qC82
6SvPn59EoTHw3d2bept5b9Nu1Qx/f4quIZJsC+AXQEsFZMyoWCihhr1GekS0xJzHiub0dmxLScSL
xvvNC811cZdmRqujEgvXa8+n0QnSa0RHbRshP8Lq15V8abPcJFbotCJxVaXMeiIUcaDGTaCKcqDd
E3zMLOYccrneV5Beok+yBYE7dBdKzmpFItrgqR48CHPNArb2I4IzVx1zq8vFNzyUwHYXEp5DI2Fu
2Y2ZpMzDDxmTt8dub/GmTeZ+dSTcisckrpKAVGa9oRIOw/vmvR9/chC3PWwscoppaByrrqWfUmRn
KaUfNJVWjNBW4BzRFhFdehgCdCVMw0LFsxr8vQeWjW+m9wdzXOBJ8E4AYzhDegj9Idernm/Af7Ci
+DBv2B0gy5uOrlNmbYRG+QimfxLsWD2OWX+OhenaQ1qoXnJZCwptx5iVhw8NYZbfKRK66ORW7WLR
UaMOpSd4pL8OGk88R812GivtraioMoNpxLvLySHV4qJFYe6JppZ3QnYT/BeapoltcT5+R0/SSgZF
4PMD+mKSzAGHPbQ7sz4jmpkTY9betGmIxkPs1cPMFy/iqudBSfSDGgbQq0v2sDcMQ1JIP4NKdHnc
N5CBv9pUMU1GvvUwudbJNNvd9RxPPJYsyp5CUeNlt85kTucSti2okwJWdkUoQDiZkUDuIFv+24PZ
X8E0twFuMKHoD4EziIYm9R8Lg3WKkNhj/0ezC+3SrLIitJ4IU7eaHQpT6Smy6boQbUYwkCuvqgc4
QA1FgyQgMR7/YhDYBN6vPHujlN1oGKZsJk8c2yNAmKe4hXZs+pGwIVllnEWH2GHH3vTUP74YXD+J
2Iq1lRQww0agwtkb+lcZ0+PMdEkGJg3qdo8fkJQYs2X1/Z35sTWs332L4XCMnKQjg3WgnJR+HzeD
yFpE6Hs2U0zCy9JAQRBSAM1NI/HCpE835w1RIPiZgsVtFZIFtllGqOVaMrS2qSC77V/G9+2NIewJ
HK6r27pIrebwDoBOjpTnXZzVbRQ1++5iEBpjd3RLhKPvEzjl/0xef8L3DBp5zRbJAnFUrNs25B65
Bk3NLaKhQ+tLk7HmM53Vw2TCY3o4ITieGQ2ZsKn5tHYJL9tRAJxfnwySVSpYQJCrsheFDxRVSqVi
SzlfD2IuM1s9Ttr0MuLhE2+X0utME8oIZCAf9omrFlqpvkpOYY8o2XRBSf1ThqZf+wS2B2HAyWHj
4r0TuasfLtUE5GDC6k0vMyj7OF2VSCv9OCYeplXmN3Gt7D91mISM2GnZjJpKc9QtD8Lg9oWWhBsw
DFzvdX+JVj8Npob01Owhoh9k9pP+/l12MdBuZ1V4+03Y4ST0d+HOjiWBNz8+DOGr7nOGRXW6MjzQ
XtlI9EhVgLyNWvIRRkT2toi3C9/WfreYhFgPnqWayVaW/KIOEwx8jFYoKmWomL2PaEFar0Vqi13k
MBdrTwSAohvW6byfE1rkfH4iEcq6nztOMg9CDdllIQ1aT87Tp3TKwyEG4fIjwnOFD5YEXmH9dXbE
KhaG/NSrZ2DTLGwie1Lz+6O6L/p+alKz+3MBSAnYNQUg5Vse35ar4OVwx9+5wDPRkz4DndWvQrq9
/LRQiPITWdG3HkCnF/ZHjHz7+ls3u95ECGG5z/FfbqltcLOnt2vIQMbYyKGpNx2ATTxGY7+loS2f
cUDOL8YBgCuWNADofNLsc3zWjn1NiLrpuoaVnzZWIpKCj5AyVs+uPd3Nc6SpYlUfq2vxB2fGkq2c
SMvhKtYLqr9jsKkmn4YiwfPBuotwEHddUyMkDNyDr3JBkeXv3xZWU5C8OqM5dXFYU5RRVdWCyDkY
s+BJnZIR/RqDisz+B04kU92b8qZU4I51y9jI9BVwNvJlwlgJcjot7RaQ5WoYLKE9n/WQBAJjc3qj
/XTOObsTWIalXWo4VKKeIZjmLTPQA7KqcQkQhhN/dLuhQ0M4bfEU7A3GfviuCo0viVwZIbzKEekm
waDCde1GrUJdbYGWdgv4HgZZ7yXWm1kDHSX0UxMtJOxw4h8aSAuVPEmzV4czEBomCaMq3WjS38Om
OOnulkNh6NO8fb57yuHreWZ8BI41dEa3+lAIyKBiBnp7XtYdTlw0Op4gCDj+nx7Bn74czCdIgx2T
XpdTnD0Ei4c+UoJLvQZCh+swoM63Ysxd7e9BPtSnMdHxOXsdTNQR3Cnsz9BnEKi4T3z/cWg5WzQJ
96j3lQFJ2D6+auSElgD+1uoan1//gSemGD0wpBZUlhhIIzEf3UaTUvlSBaweHpQ90T350IGhSZZA
MQE2fMAfLWI3NV2H0PzEDDZbYa1ph8qSHKi6i8UkBYAOrovU7rYdOJbgmrkDH2g0KHdzdlsdBx2g
AClruCxrdWHq4bi8ZOaQfeOL3qaddaWbUMh/pziH0YrlDr8zFVL4pCLA2nC0unglTpjQd4VHtBrs
MUnxJfHrIlTicrAbRfz6W9xYMIX1sP10vBWHDYcbT8PprnydPVHCzdNJphlj39KMV0wben1kPkpN
cnm6hXMNWMqMqnbax1GBfOEkPAVsSTQX8W9e42rBmct45YcCoeduxK401i8lD6Vb3F45MoBx4AXT
b1C+vSLZJQ/rpulUy27w5Fh6U+W3dWYB4PO/NzAZXy2KFO/T0+TsENHFk6kpXOQZDnZZoZWYoTfY
Nbx2EtvhVizP5xLX/s8qV48LzlbHCbV54KxhkpDA2SG58quabnRzyBc/LrU2Zbkm3+63OvBbi5KF
JxSKONTKi1nWeuTqh/fmjOJJwA/+ZVN5yOehOl/QMkyekGqY2Jt0bhRRDW08NfCZk3t2jJkBhET2
nNV4zbrWzgUBtNLGi3N8lSdAp9Y0YRWdGPXYj+NThu+L1jlpJxz7vO3BCzkikQUYeoo5ToXzH55O
ymxQziBCC8UM1GT2YqzuiACEQ9pOWqA4uoWWEhXRMSSI5a2IeU7sw+EywXfBzh2SFoc4RiqiLoAR
1gRbJN0lIvCmgTahRTK19el3BmyF61zA+qnx3VZnU0d9xKhwcZ8PDz8q/45HIsfrSIXY/TcNtxEn
kJHx0MEvbEfGdd/D/ez9B+PPIwABGxA9wp8ns008x5bsamn1oR6QqJlcfH9/PMyMyHWhntCDgi+1
BudEc3ZjgRkyP8AF/rPGAFXOA9XdWkSIgRjIT6s7k4Ypm/zsjD3X9lWPEgXMiMG6lfmIzhEQbpX8
EYSspdFcNJEtNcrvWBZrOIWZlmSbdtFvb/S/FC1cKOOy+egYJHFtkRi0oQuXnbvkpnH0O5vdetCa
cSepbIJKVPSwoQ00iu7G4Xifq8SIi/mtZCPpKQ05NPCtl5kGLk4dkg+0nDxFjCIP+WGImLlr+AGS
sAtfpujHifm7nhJI7I3hIbj/Ffb+qN24oUhCbXv3TagGCi8HzM3J8nVfyUnuxoRAZL8dt952ftST
aJtF/z1cj7aqOif3q2elqcGkQT2A86TbcEnr222N4mtlMIRcZMDUt5yxNYEEcK61dEzb8vSvPa5e
V8f7pmX+79neDL90fHh+VtP9K0+MWeqhHsNBKVSU8uTRDi2uyHcXlYFB2JLNvhUdX7h95aGIrFUj
c7GY+3m8FclvZ1XPZF/EjEK+GQI3pW68BBalwquN6TupDqbajflHex1DGHFsP19qX+p0xYPV7J6O
O8y0CZMDwCJYOFki9qYU8PHAXAhxdjPm/0+w2b1zue8csgYULih+GhY8/wraIkVusupV1vsXU3DQ
uv+LQ2yQvFJdPQUnoUcA3AqbLgsxVwe01q3A4SIKB8elZExHqjLcre0YLrycKu+W1hvitzqmmcpI
7snJMnbD0FNpjDFTwo7tUTSs6HvfRrp4o6JbYnRb9nf5lttCrd8yMdOq7BOaeTr1G0UDxIM+Ek6f
DfNQ7VPep2Jjy4YmPpc3MBJ0MQaAWeVe9ry/nIFQ0iNSVjoncboRF+wXws6N+FguujyMb/2r/Tms
XblE0piDgn6ZrGxTV+NIlh6xGCKyxuVvUw+V1h7PzzNHDnrPSrYde6BZU7lcVHHkzcxsF0NlBlkC
i9MAX1Y4b9G2uisKYWvMihhO8x/ISS8c+lIPOp6dZLAxHqwFK/UZ7k9QICfF5QcnyHE7xZl76GTU
ykJ1pfnjNEFQb8+pb+278fL8ZP3uvzAJlv1VE2e0B2j50a7/TmCprlhcs9woYkpd7UF1whCGCPpU
jYbWo+VoIyiovGUaZEhakZ9QBqvSbJ/OfWSgW9NRFO1wwS2lz95R24QRIDwUpmMooKmwcQuFYDTB
9HKKqfu8NS1FhFrDvlbMiE9L/eTUEz5LPOriNLdjAGr/hRlyE8UuoZJMvQgRa1paamb9Y72xL93Y
+RmfspP+Rpt6KQYXzZvMmqB09QgAMyvUD1yoyA+np7wrsGqXvMn+aoN45MGGtsi3szDwd1aVxbt5
ImffUmmqPArJkwV28BI7YwJLc/r6Y3OkvdQDIaa7waax53UVI/70RBOR32SexSdkwoguiIxCW9QH
o2LgZzGbIAq1elX4EqVWkL0iJxr7zuZ4VtR5u4aiu1v29akN8E/RfpOTGiCOJmjKRhsSxH3HS70Y
O4LCU5SIoWa0WUzkX8T7jp3nkDKNmtg9ZJugUkKp96mmpL6/YjsPxreBXOdiqzfzcTGNbYOWNyoo
BZVOEGdQDpplfjqbzKA+TH9j0vFjHTIDq/Fck7/+L+ss6RijN3VzIG4qYY0pXJkey9crU0ZoqOMO
6oWJ22HJJ0B0K0iWzyJLtwX9ZDOXPVRwnwxpFsPhDrfO6VfO2JzV28enOZcB/V6TS4fH3Bi9Vz+u
2pOb9EzT9kOeHkiVFKoUPArpHiNIPV+EIFQ53DwYfICM5XY7cixL3qo+Jtd3N83OjtHKK46qQBoq
9mbsLqfxIZu2BdIF59MTi4HvkwkTsXWzS9RQEpubmGhptXPDDJkEAfi9Vw54uGDI9OvcEEGw6l0i
aj/pdv0RPOotQ4wfZ3DVBuUiGSlploM/nDfhTlNZlNazmXHFeC++JcxDi4JUIxEW9h/vtPyeyGPW
PLcRZP20ODg5YxIFUv5wqLqCVU0PU7qIdPGbrdL9V2bgsbVC2Uz4GNdbxEfrtdcoAYe3vGyhyBpq
8LdLKbmh4/wAX9KEyjOJ9M/hInTO/BwgMVDPAJqW7Xdrc3vFv/c3Eaj0+GVjfGlwZIrHg/Ky8Scy
i4s3RU6ux5SNv4aT8p8M16MqRvAjH+5dITKKA+VHalvpb7gHGCLmMppK8C28n0hnGuHRq3GfW+hR
8bG9SHON+4Ixbic+ucoLRYx5oWMbvoEhlwFzhLtB3HMwb8s+LUaFwh7wuRakPxTwTrW3R5YDaE1O
r1rOB9+3sVhmVEOP4WKhfjZYKJe3Dt8ard8HhWNQ4nIjlf6iWw1h/jdVIXmRxySkKacrYttIuPIE
Rkx2Y+ib59Z/qcXKEad9APDpIyjFFl0Oo5dCo5qHCi9mJIhRLSqQ8iKaY5Lz4ArLeD4LhO6EzMqa
hW7Q4sE3XnbSKqP9d8Z0rIxXbrXsQOHIjLom7tdVTyBf/NSwUXwnQlMO2tTPnKYcF4d/9pqjOFXI
JQkx43i3Oah1LThiaWGS99g4ix4Wbicw/4DdqxhWS2/I4tPSLnMBkW+4ZcNav5qXn2dIO7f77ttl
JzYkrcmLdfmpzkV4g+G0eB+i5Z0arHmru22xm3fwIY7oUDwiJ2zM6GtnwgfQFHh3YJtON26qj/zt
+Ypr8VIRWEZAmItikhlXnyBHGbaq+GiJGzEVm6IJLSL+KueOlez3y2JkzuTOCMzfkiiXW7zaWy0V
MPnpt0ckFzGUX1BCe9BGtAMLugsW+HDtaTq9AJCHY4mZZerPtssfnvFQfYBS/ronhiXEHQNDz6eT
Ja+ttsrjJRqhnV8bFwlnQgLjDhsrY+FbxvlgxDdpR8crrOawW6wNj/7Q0tzJU0IWy62lvKIzU+Pt
U8qjIhZ40ta3uHtxS5QTPiJMQqT39z7OixeIWLdWauCPfL3wIQr/4ToM7n7EKPH2FEHYxAOJ584c
ZTkd0aoj0jh77NwsTzWUJqSgJ3Hv42r9oBaF7LjMFYG//ABFE7NjyjRwRC5n4IsGA0VPmj/16TK/
92aF1lfKIJpQANR7yf680z8edMc85iFH+08JXwXr9zK1tBD+ve/RT4XKcVTylQvUxRCwYW3VeBiB
oRohNx+CwKi3QAuIWr6kRl2vT/F2Yk5L2D8JYPcvOk6XmjRHYayjnvZqkGfPH78fbum4fpRmleaP
V7mMLa0JxaIvLGnMjmKCTjOxKdktZBtyzy/7aGNHt72NSn7p1MglpzbEPuG5kGURMG/FPzWMiRGM
wmrF5RyZCcef4+fhOtjRfz7Jmn9yluZLCuoAY3IbSW6F75uX3YhTWfDU1OToCRcLA/E2dR5l59qR
ZsvArGzj/gqpY+5C7Fjx+2a04u3Zzb83KOzfm+OTqINu0+G1fAWT8z7B9C9cx7EIIWzT4Bioe2Yo
TVz300zCSzu6FxcKLE7sExTTHevpE3qXHybjpWA708eZuKsmD7y6be7W2/e3gde0PSITqQpTQO0I
GZyvnuY76Hvk0nLgQckipjipPHyXeIyCnF1BquTIpOy/2MoIZdA/Ia5J/wxWOlLXKaI0ecmaq9K3
CFUoMHa/n6rpgI0x/+waOBKndy35WAD5icuER90eqR8ZA2KJK+bZa3BD0HUSwAvUnvc3x+zM0wya
jbaYii7ly4I9D0HgjzWJlLEVxFDUB5bAIfle+No77SKO8m+fKjFPFn/HMoqysvAjetMlI2XcDxdF
kg3U7KeAoWSf9m64aJaqCswLcZxcPYj0hkNtPxGPsO6sMx0LgOrDBbPoCcYpusUuzRvuy1DSEFns
b7xYNkQirLcPS5xZkUonwn+enYTrwgpPx1/S32l/u1cdW8crYrEW95CQeFSgfPRQ8NC11rI2QRdn
uthC88vb/81RFjQ4k1w0lYMrYHIlvPkygZL7u7c+e7xIKkiBkK6Tj8W2ZDCU61pnHu3mfb0k4n4U
AcvBqI9I/0boZlstZqJsDIbJW/ZgMiNoyXFEVu32l3K4VTm6tJ/W3u7riBkIoP0L3NqW57HJfcIi
lCTlW3rJ1EKAKNkUNha2IKIvGvCmXKUx+C2IMgVuCMvvY0MCtut+VRnprjclkJmTZv3cJ/NzCWUJ
cRRXnjYW+Wgxn2S5qLtqOP8ewzjskcbjl+4dhB4HL3X03v0j7yP6tIAnKEtfUHUsQuaUFNRTHVlM
E7niYZn2ogjNrBQi3nKyAttb2kBlKrMoiHqRoNrDqyrpG9PThkvfIINL8t7HOkj8/fWqClXtfO0Z
NNiKIly2Aq2dYW8h5gmlUnsobL4CN7wlBgLo2auGzdTVd508iXpMZz+gO7CCJ1HQnekk85FSuO2V
QQtDktm0tAyengDFo9YzOqH0QDVZwVOGDIfgy5OIIHyoqO/Cs70mgtjNoLZYFD5T4xPBoQMlPy4j
FuaKzUzaedZbKX0RBvJK9Tj6ax+U8rTEtDF4AXdko3WuO958jFuieNuvIdQzuwT25UJPqSg9Fcj7
FRaUMEbG1LsMhan1K6l2nla4OMaWiyQ8aJhQ/4OYdKBNUWbZ7wlO64O7lXA76vCUXyfqh8lcBzu6
IB2q+RA1BTxnv8JNvkMDJkEwhzi609qSb7Ve7umqbamrK1+wmPmEnWrfcEfDOOTYlgAjO4QLd93O
i8x31USbx22ERUHQoJ3JJUoT3DHQ23GiPxaWd0SYSKVaeSfkymGlBIi3bWn5lTf5nMIC/WAAJd7M
5EO+yHTlcPszAYCpw53+gk92Zsp3+/c1qnC/a5a0Qqnpwm9QBc0LmQLqKnhYkIGV46y5O9wHZK0Z
RXhX5XP6E82mbbOfgSqvF6tHhtXbeh4gGZhwzdo/VqJZtG4/5t7HJf/kRbKTbtBGSTabIHG1BRIj
0ClXTo9GUNiG0glI58pngaYZAA291N0x7lLeq9M6V3RHX4Q1Zu+8B8t8FoGXFjvd3w7+bdI8b34k
WH7g4Iv772JZHzVMspSlUHGwyvkKS45BhedaDN5Z7SHWUfpUI4HMg4cXDqOuVp6aM87ZwKjtHGNl
Pb5ruTxB00rYQWm9sfrFvsCyfKlHigYw9BfIWVb47fMK+qn8flHcJmUgVWnzz3wcMZ/zVq9DbiNb
oaR7ar/XxrjmVmWom/XHsn0tP2BoRF8s8mKv5aDs9PzD+FEY2oBBpgmBiC9/twHcS+y+fPa8K4z4
A0UmpihKu5fPtzcp3s/K3j/tEbYnrh6LPU3DpJ1DrYrOOePm7njzXobuHZfi1gXf7ICXcCM7gfM4
ExqOltgChKVOZJsgSI1HPJjATNYYRe2Gk1uVbSkTlIgRkNAlxismHxbpqZVb3YLZhtir2YMuQUOB
8r5fywqkonHiOK7CmddU9EajnRSoA6/b2RUpe1ZGcagSrLKkk4VrC/3Jj+2b4DFS2GVcTEz/Ah0v
54yrAcwmH5CELH1fiDwn6fFYBFkEa5O8Z+U5E9txl0Rd3r/0EPs/GOmpYe9/PTof+0mBnGC3hAHC
xKGEECG7Fi/4BQ1s/WWLf7+ddLAFmTKhjORHVlXoZo6uecM9VIsSyE7NVEB0KIHI2BM+POQj7FT0
aOz1o3DtReAyt8g5P56yl6wfP2mHjMAvzEuO12YmGdLmwGSHUwYkPnnnzMS6Ex9IVeFjby/mvVY3
fKaiWD+l5tKjULFw9Nzwne4hpxBHAh2nkTMFLAEwmsYCrMQhx0LJS6JkBrcauii1sTe+/EA618bP
qmnhMkvugUgN5HSG5tInH9TzCa8HGkalLffmSDdiIMqLTI/s6V/WMOTbvVdl+Dwrru/aAIiAQdKA
cD/tntOBT80YfVVRz0i2TUR66akf8pIWkoL0Qdx21yRn4t5pIW0TbP6B/nTBkSE+nzMMyNZC1MCa
8Upl9ReWD9bDKpF3I6I46Kgtv+hjuDvVGzsXeE0CSGuGfK1+lHWAirCyawfkqu148unDl+ls3xzY
O1AItk/GPVm36Rnn7T0uKHJMdr9Pib7wsplrdG5J8RwNpMtHRDiMKo53TZVM/W6U3NgUcUMSV4JC
2PmRD5otyWtsbPkji3P0zDM8/sB9dJIxEYxA90V9tGD8EcoFuaJ/rczVOU3IkoUbTM92b526IhOv
lUbQitGRv/B5HH9AwUsvxC1FIFHi5F7yDulS6X3r0oUGRdy6Jd9DyPV1p8Ji3CXQgavyIZ0RLzk7
iYx4P6jmp4B+vpT5lW/8VIdMLT33TS+DMHGg78Qcfb+haQYkQGgZDBu1/49q8zkkBnhtOP9AtTtn
ljK5IeJN8GTZEvYqhrk+6jgBbjbTbXmphjExRooeRClmfe2jAfGEg4BeQH3ufp9MuCT5Vvqyz1wk
561hBrsiZDufnMrKHpOVgjCrKEzu27wVX1b0dmP9W4Muve2uNSIjtu34xciHOko//eLCMYWRJlUI
9KSNMSVZ3yOvNWqr7N2nG2feGoP/nmkhBJS1OKSPeW+DjDwRJz+nejy2inDY36WjmBM29o9Dd7vi
rNBKKke0rUdLgeaSJFISVfd7R3M8aHQPKXNqrHulZPnfAer0P4KK927PEw92nU15AoBU5WgzebGh
UnaIx4Y5VDkS2KL/aV+priabTEFQuQWHluj4r5VYsb0gRHS8xAE6iG+KhF+6PAbLTrBq37l+cm8e
NxsCAXpwmkuZPNRfHyO2LqR1nKdlYMc9R68Y8LRpKaOyOHPqAHRO8Lt6CBRBAUmeiX30dcHZQjge
sYoS4SphKRWXiibvfPGVB7sr7NAes3Hz1Cf1T4T8brAnH/Cl6tB3qhzZfKV1h82ebHVT4EH4CT3/
atZuHa20THYDGYg179VlU/4QkqkF6NPdm+IknztPf7RMTeMqWiAifH8VrQJx5kW0xYt5NtOlX9HS
6oAyAcF/1C2Xn0JV0fJUSi+/Ks7xyBt9yEcASdzJlBpE3CoPaH2reZmIBrk0RVtRVqH2C8u01Xex
WYd59eIBWMDCHCcexFwikgeFXA7i8TQD7mOhSgzlrOfBifU6x8EMe9K/YYctly+FpLBr65ZMdQ9b
EaC7AwDZTRwfeUJB1UQarGiXy+ijHkfjgYWUeTPTuh6SZwndEdk9gE9dhElkJuBYkMRPLXkiIv/K
FQ3xE3xE0Ika8dcTfgF1Zp+eGWoxzRJOZUiMFo1V544sgtvr033DjL6wvcv7Lr3onqQ+RYAQyh9q
gchHLBUBoixwmlp/vhrNfH36E1VvnCn/kGu4L/a2EDiVtF1ZfDN6ib6qciADSyNjXyItEB3VTd4K
EPrHqsr2cALrQ5Fk8ys5Fa5unVtQt8euNIbFAI4N/zqfctPk/41fFep+mb7KiBRGaZ7EFQ0+C7s3
Ao45d7PLHpe16v6Oksoim40nJCMwyA0BlSXS0lc1liwh1+jyEODtzxq7EORrbj+EpZL76HAJvtTm
PVDVG58q6lldsprZdCP7ysFoD4sTqTA0DPn/VyTaH8sS0rs7YX1lxsv6/maWNBp9WXdtRAplrB2B
emmGSoIOeNXYJvnvOMqxYr5SRABcuvGPHAEbnhKmaGAKcV+s7J+Z6qvMNbimmEex1xKtEg6U2gKq
K5HNHBhm8b4A/ynTxdG8114FyD4uUgMy4Ayb4/sSsh9izd/80TZDrIVZAFWginyoMw2YPwGZ+IHl
Wfw4FN549tt8X3HrU/MQkbQ4zjPfUHC/ewaCi+flAJ+lYP0hhgHxEPzZ8whpZjN9ssXjmaOb65x0
bFc2vFqhLA0OVnwuqdphTtaNAs+N+UBPqHbzLU4j5Ad/ha/LMKiB7USb8M4pNN7429g04G0auyLM
q9kZ3LI8NBtbsvAyXmFimu5wAgul4Ei4ObPB6Z6/s/F9CpdsKt1ZCHP8bgSt3UNWkrdYztghXENt
khyyggOLNUft6rILJo2loGPJj9R8Un7Q8VXwjxmkUF3P1Zh6d+BHtvn6oYN5GsGZODx+QPQ8t4BU
W1ZmeFg6fcVo99rkgKs/1iK9oQ6nqsxY6eUy1z6BtLWpQt07sgQEmw+bdqhmTb8+8lA5zWwiScUN
bzEIfmuqT9zSVhVKy7W3Xhd/gSPLVEng4o/jK5nQ9X5ahzLceoVe+aasmG3zg/wA/u7FCjau0+f+
a0FyE5mELdvXkbKwmZRGAro/S/rs6Lcvmfl8NRmLQwtSkWrgEWl8pFSjG7OXxrDQa2vAX9VqOOVC
dwqnn0+kYNfAGwLLgbtq1IAkePKqme5S33vMW7Nt4r+/x5VlOc/rb3md8ylP70fa3pTtF44uVGmF
9dDH1+s4uUTT2sJeHM4faVaylU58Xr0MrV0KXXhU3ZrGDg1nyNv2/gfUgYFdtgqsDvDQZRZDlPfo
ou45ybaXBrjCr2StcEh4wFhcVatnFCqYG6sbN4l4ppJnYyBdTAmanYcQ1kAYnMRQTOJ4cd7Ks9SG
gzdDLe93MRZoLxI9WS0PayKc1uUMTTPSAep5Q9r6yUrWW/+9YolELeS4THawVGl5zekMU7UIPk4R
mEGi6FZ//CKqru5e4dz4ZXtUF0sWw0+zooa5K5W36wati4XAqMLRZpt7CAEKRXx3eu053bA4Zh6g
3kgypigDAWUEErw/tkTPCimEfXxU/gRR1/+7qMpj999HvSN1s/KpIhKD3iVPJ7dsQesn+amHvP7W
ELmiTdiwqOhcNjAGXoq/izmKxEM0fA432z8UIIa9u1/ayXprw9ywXBBDpXbWe6dwbCTbgIxTpitu
SpeHZ0V9OU1beljDDFB5MTG4Zg23eTpoLeazceUhFxBw8ayYHihHXxOZl1jraNo78Ha88bPISM/v
zMmJAmrW89dtQLXAbIO/lkHBDkMQBURDUNAmLTVUcge9HifrYE4KawOImdSPJabuW7W2QGQCdzR9
7d0c8aE2SbynDGfB7JOjiY38ZGL5F9ZLCdwPt36LKM0Da07u16clQ3N0Xh1NQSX9YwG/u3biSMqS
M8E0rKdFO6WBjRMZbhzVkPMvO2HWf2mtYVjBRzLyLj5mmiihRrebNN6aRmZKtNNB/C2zbfS+56gt
fp7ZLG/Pa7HUpL2BQR7uugcjD+ndq7uL4mlv37AmRpsAYDKpourYf7UDK4ts9tgKm2QLgwkIrw3Y
fITDPvJtkuyORiLn0ARvtk9HVASReMRvgqZz8lxldJv1N9KIlpDqB4fLimQGU7oTGgcWMedo3Sy5
t5LVeuRC/3ck9j5IsrqcrOlfelac7vi0XPljh8SCU0ddSPWDkWtbFrIDjSg+9JyDsavtjhsKCnTI
A2LbomUQFixzKX1aOgHCfdXGka1Q0YSolO+oE0b9Hdh55JAI86MuKIKFxK+Kgw15nWyJLHAm+DnQ
siINsA4VvJNbEfWpkf6eDCR6FHDea/S4D2DYwDLbHyatMfc3VuWAgBsHMe0LRjA7k9urtD1Dwmsc
YVSeimBaPf8aiCrGiacAi0WmlfcdcDHXCWqKlpRcb7f/eWcXP+CCHqkfdP1z6HrV+ZiwXBWejXnp
9cL1l9JNf8ELPiaaSbyrhGzhajPXPGvdDi/oDQbrIpL5m4tyw1NcWzXVAEEvZIvOWobYxlaRreWT
aTsUX4+yxa0U13AohyITMqXS3xkY4SLxc1RNlEnIPb/apnW6+yhS6s3HW8eUOlzdfOnUTsctDnw0
wjuZ8YSX8wV2kI8y6gTDX0EHKZ7b57pK67pfUYDYbM1nx2loJBAZCkwPTKpnZACOXbCnb3YL9Vik
3hrsg6rBKSFH4BaIsMqq9n0yvBcLpwRgMGYVfNDBKJ58EP3MT1iDGR/y7IRQ/V7iWsT6j1lmeLGU
sIi54AhncX4CMl8X8iZrNz3kLfQdvjg0NnmdcCnrbXlG+n9GBWoGdKo1Ick3kE/4Oq1YxrQoCMam
Y52I0pe4f82WzC3S5YL1Vg+r4IfQW/kPGNDOaKU+shTIBpKugMlRblsJMzSD1bOEQvdfZ+JsCnCH
kvkUQ0YR2JJFNdZ52vF5WUGkyt0UCWxLDKHpUeIEXE3hsetCQh4mJp0lDxc0l5Q6GfToLwRQU1Mi
AOCovaQTrd3C5x0v7bBw6QlH0pc12gSD/05SKtFDuKXoCE3klYt0u+pwQ+Mf2H6xVYpd7XucrKgA
B+mU7kvehkyK7ShcAyZOZPxKldO1YX28oi6zzvtk13BOMIrF7ObdD1xZuWMkbJHWeNOoSPyixSm2
UTc+th7N66JKyXC8VJzX7/ab+r7AQjfWWIhsaoBl06uW0k3x6kDa4xcNFYPbJ+ycOUIoS8WFnN/3
q3C6IiGDHZuLsVIX3cWvG0Ujz3vIBCQmEBRKIYTqAlPz09o20Zv6GgRQQJ72qzezdvz/l5Ow9YvQ
vPhIjwGL4XN/Rjs4AJj5ua4a5Aw1FADMv0ubizgC+dtSv2YcIyel2/A4cW+4Magc92vfdebAKKZr
B+KEK0ncLeoCt3G/iXS+BNwGPRETJDCpjAO0g7h4DV9f9dCnjJFrDaGriVMsVPp9GBpajTIswpRf
H2kr+Uzwhp1h8PuS0h5d+bffIoHixjxImal0QYBG9zBdJ57tECzYNbFPpuRWAoRpnY+rqUMQ1/u5
S3J+dbt4sHbVCrUC7Oco0CMXk7yI8hSGpt/K6+TqYwAbgQiuXVQMPRyETRVKXiwi8RV+hCiAn8+I
AExkGd020X5+jDVC7qZIFPMs3xBsE9I75z51iun6VJEmlM9G19BcOGRElcFTi/FkImE6/hlWQpWZ
k1QIRq+g3TMQT6xwIsuAp93Ae6OSLohsyS8GaTvH3Mabr+Kyeh4IzmGf9CK7A0ACGs1DF7ce36ky
Hcu8BcX3GlJuJCZWPtRFmwW6e6Jyo8folFZ8fQNFUu4mg57+qUZnCjf7oJjqdkq3IfKWV7VVQ4jB
MPxM7WZQ1524m4UISNPxGa18zSc7MlpnkGxpnmqncyvB7rA8QKDgKaT73+l+P+hvRMPyJlgSl7Db
LIyok/+cBAPGR58kCuUB4yij+WsbrOgvR3uuCGvP4rFBYiMOmM2VHy+8oHWRiiXiPTGRuzd9W9IE
kDjoQNKLmzPQqciIr8xSpehyN/0XcRykajUKOusLgZv6jOw6RBFnSKdlep/gKNiFs1NNLYPmgWI0
cdbzAuEB3xJ1BLaVWZItHg5cJgDrd+pvnE3tR2/dy808Hdmc0BScpnRj/g1ACTK/D/zDq3MmgHKE
tvB4dVd/+xKWUsrq9HcIPWkkhwUGPRfuYbOs+1U9PByCbzafjAPOWgnjC8jrcQBNapEckyzVMPYT
4Nsmrw0aon5ztWochepEjCcxVFVGeaTzRPBF45WX/IQ/lWK6KU90OiI1zp2xKOoVj44vSRXC8j3X
Sso9Jj6+L/31R4gZ5fuzxU5/pf1hqry2kyFPlfAigQ7T3thndlEN24dXS0sT53Ubl7KqJ6cqkFoX
uJRlNQOxqwi5ng9xYYoNkxbMEvs22CmmLWac3untj6tkbeh7/LUkow97aX5sFQMRfrMB7JVDPcCI
ueff+/hR6lwEnhdV3iTLkD+ejZrgXM0YkK2mUY4VB58S3GE4H33Dl7ek/ucuWghOX0nYqMpFicgM
AqhvlxHKW11rgQ7YF2sPNb9Yx/vDP11Kfa5yUrKW9o0tCVWD/TZJsemgnjswut/69PulOFEIMbv2
VGg8MLGscdyNbIiLX2wgj3JjdORQzrHRcW8DXmDFfPWFDe8ufXV/5CiLro/8dWZI1Z57g4IiH5Ss
Hrpgxg03o+vPijgyIJzoV8+4AbLs1mPVN5UuNgw2UQK/4Egk9ICyD4i/MvDFMqNzLqXtdew9ntxk
cp+z2YPrGu5QtDoNVGuFR3ro5t8G5d6zqwnvOSYxqRTZ7uCMT+1MIP6gfCBLK4BoO5tKFTISZ5NA
FE+nlZLbD3nYPn8U+Z73jXhTdT2wVy6s03yNKBy2VuTsrlrhXTDpxAQG6HsGZ0bBVI3gZyejZto2
9PYpLINopmbGXpfrm4ttfrjtfxPbEOmnQ+FI8vku8KKGMJDz/w7TMhpQP+DlolIoWuRuhCNCt6Ed
a/CbNu/vAZC5X4VgdeFh5kOBJJyxq2Wxj1dCc7QI0dzzsgrpkbh09XPiPfQwO1rsUZNzEID/sSlD
q+tyfPIbBO+pIwJhdBPfaqml8lYXQjvObT7cKx/y1oY4FEkxskLp2lU6R+b1m4rSfXrY1kvMFA0C
UiMbWFsz9ZYGbqCvMpe9jegMPGzXVdJf+qp303uIk6ehXbau/vXeXk0Yeq/faZBqPAFy9y9DZm1R
d+VMWbbqArEdId0iVfpXYZB3PPc1va7vr8mEsaRRS+iO1S8F+ieCPWP2NT8/FKPSy2MgkKj8Muff
Qfxny5ictloDgAYUlx5lA0QSiCZAhY3nKdMxxNVBSOt3pbVi2DqDzeT+LG02kQSu5LF64p/rpawT
anL+vZP7S0lXJ1mjCJJguc2C3U78gN5uKkttL5U9n7F/HiapTBy99PmLP0BH6LtR6DzvTXVTh7Oo
kn2KbT9Qa2gab+h8BrinmtvK12ND+neeQve3WR0S4XyL1Igy2rBEHfsancqX3qAeO8wds8OhGe8T
NiR0iSNhGHumjb+CPAKURPzsf9DvjzCYluqHvDkgFlKj/stnfMzBt5a/Zlg00Iyz5rl0RwDac3Bo
FgBZeyfPhCL59UE9HuG+tU9mHSchN4IH0tE6YpJBF3yiSko4za84sVzGN2A1R9PUMFyEuFg1arYN
UcGyrjJdGbkN2zcUz8BossrSDa6BF4mG+YzAXIJkXMKa/ebtaMaE+tFLKU0BT8p5GUdr4VhoRsAZ
Y9IQlOriA2UBIGK1s3qoS9fy6nQivAx4Q3LMxZtIwem1xH37W1aLLU1pXber+e23TlaOUOqrmNlg
KuY8NrCs/T6BPAnOArvuxmbyjyvRF+zoziLImp3g5Z5CPOLn9njo8qA9XCLP8FgPSi9WeKSCyhNl
S50A0S8BATQrts/02NlEYLBGGuxMVtd+0CWpvH2RzPfa7S/xg8NNYVCQoLzY0fXRjWZ2xABP8hqM
B3JDLz3g5U2PEhEwYUV/Z7AatDQ6o/PsO5G1zcyW/i3QICPR1JyRta1rAmvR/16SyUYQAP828OA6
nFaFdukSrKjd/3FtFYLCjse2ATJVDPDQztYs1Ahchqtc0EK9XcGbUeP5UueGqsfWWRZFYKEBLwxy
DJOHczuKwW9vPoMuyU/aE8YULQQj5atvDn0piZu4KQDSOYBTAPtgtcfCjFo6b8IqbT0qemxL4Vw5
DNE9XttPfFc47d3cPPw82AEIbXoXPdaVOq30EZROYRyWncyvB4nCOVTFX+Vs/iw+FzmeiF+fCIL5
x+ooddCFkkrMK8JA5mN7a2IR5UtUIUOoTr3b117QeD1MB2bo9ZeQg0IWMXdP/RtasCiRpO01LHEn
3gYRk2E198G0yf1NWHky3cck5wI2DST3YOlJiCayMPH30GiZK42FtUTCVWCxLpvGW4jnqmxVFEK4
lRCw0IxHpT6OBrK17FIzSRrOenNDt92TKQJf1OT6D89dgLpDKLYRY70fnK/F+qU71SG+azBImTP0
HWPXBVzmSb+OcZnExl6w0aGMiG/anYo7+n4oA2pCetLQuAEQz9Bqa2z96HHcMx2EoRGwSc0NoIP/
qrJaQTF8DSl+UkWL/kIWh11z3IHZGy0xX6Hw4XSW3IOg2LhKybg/dhnTOaDhYJ+KSQnHgmitL+F+
yL/Qww60x7iRgpKvGI4oMT2mI3Ue6Q6eVPTdQrjBEWDNmnycfP6gcsMovgnpXuFAuT8s8Tau/uZ2
LnlXfCDXikiug2i9ZW3sxrGik1kayzmeH+Ya5HQNI080sG2EXuQfjrPdwoBKmx7/yb+Q2hI2VCv6
JiJU2c3WYgNFNh6/1OH6+cqAa698Bpx0c7KskMqu7wSj6kfwLBARyURu+ga070/GDeect1XlvNUk
ypMLEESekXBD74e9PxhuPr4RAOPx90JMD7U5YQPIkEeX/KCdYTEI10oSTHu/vHMRyP2dPr76PVJ2
BRoraTOBWQAbm8ahHmtv+eNUg3OUPQNot8CV5Vnn/1qS0ZB9woI42ahhVffbew56EjgklTz/JrKw
+DMYtoY7tMd21uNSiHJD52iHVrQnSYzOEpZTzXWqg8ntaE3nZM/Qx6AufJNa8TTPX7LxNk+hGOQs
+ouZu8EjkayOXbf+blr8kivri8CDJO+qHNJoRCSQD2ul/uR+bs55WWzn3+D4UUJ22cSEixcGaRZn
aluq0hqMWdUYxF88cFJEsoTB4QLLRyy4eqbOQaTqMaxlL+IJd7VAtcS5Q7SR+fmERHzSegTDNDrb
860eP/BsSJ74xT6qH4q5gUyI1rzhiLdOf2ZI3HjzZjw1adAm483dvTwYHLpUcO9PPf6JT2wba4/8
z0euSI9H4MHcg6HMdtn8wNeZq/dpvWgUef4/U/3M4Hd/uo8tchzGU2Xs4gjUoJlf0LaKgISVJZal
rgEIt2kavT5NjOhijim2ZC0vln36KsOMmtwplj7/aIdkhYArKqaG2jpMQXAvYQSl8GUnWZw1bdtu
7y2R+Mvlig7L+AFOKwRc+kEMEZenh8zP/opJ67rBhjRnfxbELxUW5mBby9y2ITg+p4SFpRWWkW6F
ieZelelV4xU2I7rc1+RKk7SUpuUWkz4OuL8qg4JJqe9rUmX4MYvrJuN1YbVdHYWhJxqgyjYBi5h8
wOM6a9tbvUz/h4E+3mapit2j1mK5MyH5iIPNrnp69W0oQsaX/enNVP1ePlFjSsiZ93VFEOC5BKFz
dINybiidLG2dZ4tTg8VDyHNKlURY2iMJEiVoQKbGNrT8w3Dj8JY0uVFe3PrIUPJTNMKdsRpn0zqo
H2fr+q+Wf7SIYyylYk9aJ4S0/C2m1c3OHsDJHeAxcXLE6nHXo7ENo2Yu2C4aes/Ml5x5U8U1YmAL
I6m2HUNLpFKE/vCHeD8to+ogeNweM7c7dZ/JtntXIRECeHL10UfhS5nDb+Qk1Jv1rxKnOQnDeGGi
eilRF/+WBvOXpl9CAOL6FUnRxQMd7FT7GOmBzYq+tbcS7Q1TxaC4iZcuF9Kgmb4fJmy3gev0wnLI
jAre9Zul3NzeSwI8oAFDPKWnR65vkfe8y5H0WEuP7YHpz0z29106jJlnQ4hXQpaztC/Jt8F47Hn7
CIZbL37GoYceh1AoiL7yoFX2c2YG3It5BfYdfbzpkDSouTb5ft8gXMGGnjQzU7aE8fOWFcS128jz
gh9y9zQmwnQIIhm57anC7WSS5WRLTNPs15qSBThMtlNwL7xBhClPMfSAsEKS+aWNcBtStfKyjyBq
JPFMgMbSiljdw06wtm6UekU2tHagP1vW+YWjWILNMIqFvNpOpIVvYPxsSffB2ScGG6vQD86K3UJU
p9ANonJrWTtifd1pdGi23V7EOnULnVoHKQOpVfDqVKJtnzcvfE6kBy6vJ2VMYXzQpw7bt0eE2MvW
8Pv0B0uP88c5UEyIekqNZCYPoGyLuSNvj4Qi74rlyFFT0PrS5UWp/16xEXVvlmgCa6WQWIzrJfa9
FTDGZ2HTaB/Saas6wG4kkbfuGtMIlmvHcfNN3CR75AV81y9PHIlOVZFSbTOOo7GPy2ULDUEch8br
zm71vQ8qwuRK9p22jSKdTgXL9MO6TgR1eeoUEONcMN/FZeuQSwuI7CrWManAib6bX57FkUnDrmEf
WTZ3fU/qeAS8KUSK6aNAlWvqCD5ckUzj4Ym1YtXtIL9GAcVhh0I9kYgAS5jxbXhVmiqDjCIjJ9AH
JGGqHfmjbIHbJLMVXeiX0haIIeImeyENxsnOTT13wE68twne7yROehPOauPWI00CTkq8pul8bE4X
rjs5QiZ/vV6xphSnJG6+aRSln4Ao1/hjCvsit1L8ZtC3GxqmEnGuy+ZNCdj/U0MVSyZTit+nyjpc
3PbR1d9jMHBlXZH92GgDRJp+hkZtoXaGvBNuQ7wNZvIo0uZqYmkZ2PM9HD0R3oteQHDcQJLs/5xy
mLl8HyGyi5h4am3XxAKvRMqXi8yoZmRD7iLnxkX+8P++z3CxISb1bNTUv8cFU4uBvuwmJhMIiIIS
HJShVziwdZsElreSCPn8ri2v1LDJePQJi3ukWbIxgBU6Cst2XqX6vYNk9dXOdB1XkkH24rb0ZzwZ
EN7pvo/n863Oc9JiesJH3CeLtypI4XpMDjPbpCglHutZTh0UDfW+VU2bqpvCImz9ZYw9P6OUeAYM
Lgdc8mL0QBo+y8x0ogpYCCZGYVaTGOo7dTrDDhNiZMTVCdKFBPgoKAHe4Xp8g1IQdAVoNeeJv+tk
0DHvB740X4E820yhluVooOOzxvoQSsPpL0HIUp+x+oCGKxRwHsRVPRXPrpCpP3/W4Nixyoeb9wJ2
3cfv4jHdFctJ/cMtjcD4DLsXqMj3HlXXIQvBUO0QjFG20RLyvTabOpy0HQe3BXhKxTALLC1ZIo/m
1lZz3e2d6gxZd0nx3F8RiCiVKmOmmPRgGErJABQDwzZcO0v1FPBttENeDKbwi0dlQ1lzkvMDSIAj
KYLZ/S7oGsAA5DJjMyo5WaN6xAQDU3EN56U0QuRXNhaT9kVOkASUUo2RwSSH9BMnHOBAITl9o9sv
F1hGmYjR+Z7dTUNaPrI0pekU12fjuTV7PxIiSp51cmxdL+RGMrCGIuh5k3Mc5IOow8+Qdofj4/BJ
GPWLgKuT7zBOjBd5D/9A8fvGrNbaF+Deay7kgM7Us8dvj4JeL1kz7ZzdcVd1kUYAfwFOqu6vXvl5
uRpKDv/Lqx+w/oYizybjh16HEtECETdo66kuQhccHHhGOeMvKT5qwmDrZ3fV7eH79/97Dn/Z93vn
aaSQVCZ/CRZ1wtnA4xS+c/YGsZ9cA/pXuoB0zYm32hGDHj+G5eCP/xYYf+F3vJA8Ql5XkkhSHkI/
svCUvZTmG0RKV5AayYn0SabbpgZwpM8hKqH5Y82OD0iuDOtXMDg0GkCASVKpHUPh3foi09fgua/Y
k9YnVaiaU3A9C3h6UtU3d8sYMmexfng8EJaYA7IZrJZzd6ww7HBtgiUkij1x5tk2tlXqGKFMKf2M
lZgILQBLhY/NK4oG2OXrYr6v92mXKAwTGKgz/wROn3S2NgEnNvbd67wN+TlN6sZ4oZzIn47ZHM3F
Qpr3gaYtm+8vMJHb3KEsMxn9uRLW4JnYflXDDHs4foaTOTh6e4z6EDF/43ALkZFBY8ywdTyuC8Hh
8q4DsoUA2p9yKRW1GyCf023uFPIE+hEDsvBL9BOD17yzQ1eE72V7644DEDZGpxFbFUyn5L9+lMdi
S06LWAMUprbChIy8pNdfPvL3KL2WGMcmJWPBmCfrFEfvFaXG9WBNIUyFHFscpKFvWQgQJZJKnKna
Z+zmj7Bm8PZrM0wxKAuCgD/WrNbSDV1u6wALQFnFiMl/fbniPya5Bo4/WGa9pBucTXkWp4T+eXNe
Kht4di4B4w3EisazED/9pkY2OHJRnNKRDQQjf9ZMuDtv4sBsiqgz5UoT/F9WFNPAFILyv30nIK9g
np9lawJy5D6dC5aD/5BGwekQWMDs/zT2YwF6CcSDgNYEP7xvsrd1TSGM4Ku+t0u2AMkqxAKOedwe
2ZQsNu6mYApbfwDczZNkzhWlo2TFdmOTsI/uXo4MMkaLZEO7AJ6yW2BFGgmvDfn6t/0Iow6Tcw0D
sXsZ8I5XDipqIvWAKIJtAdY8/SweYaQDgFI+5OfnCU25Np7i93xHh0Ctt82uzuR3ANxbfUIh9V3J
pQ35Vv++JF6NZOZfJtcxsmRuzZpkq2lqQRY0mE1n05uAbDjnYLCBN1q//OsEMo90M+qqSaApZu8X
j/l+AybVESyKMccuwOkIYybvjKuUcCoHo/2jjXNHWq5nCnUI1k7m5HzZcIWVdAD+Gw5a4kj9i8u/
17g+AVQrKuovzUO/WCBlWOP7FW5eXXPhcDhZwyz4YWPA3Y9H3+35ruKImntdtAqMS+dMrY6KQLkH
ph4RjxvFyd50cEisDsdRIYnDSlAFqj1YJtO2WJ8wNvzZpT4/hSPsYuX5pDDbZW9uNpOmdjDF6xto
5LFtI/eCHqMC5/pWTmq8m2kgxG4XBeZZK94UjdjrqJXS0G53D53WHqoM2M+jIPgC70c9H+Gnny2y
x9JOQ/3F2Xs2Qr0l6maI+vTu+0+vCzkcN/lsyQI8KzhSMRqFEKSWYv42U1nIgQ/TEy3ONe29Hi33
ZMsKcx4ocZBzXDrmcBDoVvu7cK4eJ+WrzPmA9vNIrdvkZmthWgwDma0qiyecsJ3lSbrXLA3Of/dk
/WRM5lau7KYpcUhhk9C5j0IttI4opk4IwINEriMRZpnbIGLT61b4CMiekE02VgOAzmwN3ihM38EV
jCkD1Oh7JsjG2ChJLoEcau4glkEsLPg2cuFShu0vnpGsaQUhVE2mPIdUwzBXN8VDUwJenaA4uaD9
6DbRkoDzR/tiUdoxoSrjY6cSKFlSjAN7HacIUOQa/08a9Vz0uE00NO6SYJB2/dNFsRSv+0TpmxtJ
lJ6sUD7LxxGoCIXZlyqL4SDd3jb7cLd6MRS0pJkRXWMgGc4PE+vOb29wtt43e0SvFfwi/vzEbqMk
J4qEsY6QM7YI107/JO9tpGbblZ3L90oJzuN54H3GEAWxzDjMv7Zs8XqhlmlNePdlT1uYkqMhFp3u
wz2G270xbdLC5L4fmmzU/qRirOnL6Vi9xuACZqfq2UxlPLQ2WN1BDWkTbVQplaNd9nnttRE3u0O0
GSLwFgqE3bpRuxB5IgMo5OjewoSM2RMYDvwGZP6R5O2Tu+AQO2WI9wltIhqHEbHWkY0iGhUvdA+x
eBzIvjcfYaxTuE7tBrGntQKxYx1GUng0DS2kdBhKTGF5hBWBQ6KLxF2K9Q60ARwGPBaC4NWo3gsT
DzEufwhFMLFzwkAR6nlwL++eUnWtPXy/ykYEXjg4G0W3iXdfRJKptg2du4OWmRyciVHokHv63yQk
alBU+f9dH/S0SRBavIoqHQ82ZDjKbwl/WQNqnkUPT0pwoEpuj7AkLZkLNuB2wKmpKQdLQq30qXvm
QnWhzfbEg5I/CPxolrxvrcNrZfiPRnd+zymu3E5Szt0JuuT+RlG7kItvm66v/pMXPkHQqxyukNCQ
PDTF68W2HHLh6FHyn8bBkMinJpeGBA3lyje2hEnlKhpM4DkFLbX4sGTYI6UzF1shnr2Pl/3UsRtO
9yZrTIUGE97FMU0QFQbMlOaF9syCBVNv0SRQ3yTNWVkXRRsS1TE7mu/OrHczoM3FszcoBmz2QLz7
V9rZ4htf8sO0rt8WWvPOXSP98zkddu7t7Kjjj++20BBLyPSS/dNR/na4OU3FPiY92R5jUz0spQjq
ldxZ0Dm+IQCMscH69R8I0UosnJ0uMBqTXaM8RQ5T6OCwNobox25QPVlSh8pZq/54GZeEXlCkJURx
/cYVrkSFyDsr+T74nUczMfegKbuc4Mr1r+jqva/Aq0e33yD+yQtJMWC1P33BGp+z3uu86V2IjzQK
JqADs8BSt0lWDL24/M+hbv0XDdDY6RpNEO02qtStKKG2+dvreyo2JkSvjI81BwObZl3gBl54X9Lm
hgtfr61dR/XNW8NOsi5/FkKFSGRHLUWyBmjFIPF+Xk77pQZxAWjz3uncBa9aZwL4T4Q9D7/Lmhj/
+M2bTRJL91YEYjJg7I9VzUHCg5RXTQlanWnVjMgb7FUfj2Bh9Mp5xVVY5kJB2/+cEj0zm5tv7ouJ
rd5buDlA0yVmG3dEWZJZ/0ADpTFsGNWpcAkZR2JPm7QH9h/xtMc9CHWiW++gZrYSzqAtlysB1Dac
qQAK2/AnXkyxHH7UNih9Vl9mvw/d173fsCa9oLptPvem3Mje4cJUFC0laqY3Z8vc/tYy7rlNl3XV
mepIMij9TgQ4xcPKcmg7aArhWEBHCF4BMMlpambw3EbQHZkugLroRWd7MZhyrKw65s+aUrb+dz02
RCwaSxI4jWRl/EAizYRSHHKfSaKdNN0xu2qH6xxFUjjRo7bzGO6uwJr9f3grmh6yN/HgbPoHDUTU
et34md0Ib5CCcTNf0E+FfkfGfI/Zg0tSXEWFw/9s43pZ+9uEku4DT5LWrM0skzsglp6HgzlL2sz6
UtwJJWDouyadZvrQTDuG3J5e8udiBYqRNll552IATajZMaBxHTuyoEvGdeMj9/kYN9R0La+F60i2
y+HfwgT2yBaOtn1YdG+mFiD3WRnsULT4GWadelNNvxhEW72bqoVQoWADfWMKCq0bZgDcHxetTW3U
goTTDDFLD3P7BFWWIVUIZWo+nLzncoRNGF8/GLjX9EeOuzjoo/yqe8AVsoEPtHEQS3vDjq+k/iF/
aDIRktcoVNJHQiFHVbdZZxK+POvpwhi6M3Tt1sQDy39BkD3D5/wv0kiwu6hL3nySPLckrjz6CJrh
NOie7cnT9rCKd9oijrDK7IXYDxldV42v2ntWajneqh2rFhMLKBRc2vDF5MH0zFIvdMBj/DM1K6HN
glYLpPOaWLWHqQszs6MWjNvO2qqyG49GsOoE9fPFUguHTzalAx/PMs1bCwlrgfC3PF4/DrVuxAJI
B3vctP9m37i2rXxFdVCOTrk3SeSELpkqLTHxQgEMioYvNkpJrGPtAtN6+juED3PXAM78bs7XWTAY
4Wz043XKSWzAifgM1Ae8CqozFE8cpw/81fNHcvXEin1s/r0A6y16XOiD1pUclqkh/2QaCaxr264G
Sz3yaX8UP6+tjIxl4HXlkzARgwBPk0CNJsq+7Q1++dSiA2jQpLZSFQgY6YkgYb5O4N6ApVadKUuD
36+WSvZNuRDVecSVPaPX26a/2pnDSh/YKRNnN0nLUUlyWcdBl+8MqP+63OtViQZfazvAoZ7lSh3g
qzY/va5Dm1aGqeHukJiZqcQuIdulAgvHKGIp5T4myZlL64ngnCSOqIxGh6p5fz85wr/BT6uuzpLy
ogPoFOkcm6J44D6wds4C84DyfGhsHF7+8K5CMduYhjOKmJnlDv874tPK6ZcTcs/NCoYufEala/0a
7xmt2hRKFQVAMnFJOEqVL7X5HS6pfu6wpAD3w56SKkheH0tYMtKjbnTJaUVf6dtu2Z549SFS5a7O
eERDLbd4plmXLkNeJVU37JrKtiWPMmtQ0dpWgnywYHQYbQtLxC4tlub2zY+z5WdiGZVY5GQ9FU+B
CuejKw6RqRhTD8g0TGpP6pMUzgtBmEgO9cT6Z6dYc6y58PTUlYgzaKil1MaBM9F/p1EBay/RCN7T
/rkxdHPCy9ZBcZlvyTpHcZFfwMZPxPgbjaybVVgRCevm8AJGvljs2tkjNZb0fHOKv9BPLr9S7QL6
khgR9mvzq7MeyJjgxljihdif9kDs1GkEfVi3llGHkHwFvVNueOauZoJ5+1PDvCTorHEn61L2j+jG
WjQcMdC0cE3IsRCtY6Erbi59iucDNZYt2yD0COQvuN21JdhMEF15suExWUnMJIG3k/m5NnInmFwq
RUNfi/MlRAavwF8pJIBLHYpwApeT1KTcImkox7YH2Di/laDuuQuOJWT27LKKrz4ABsqlajdq5IvJ
prX6366tZMntsn7znmMPEl+QrD3uhpv1FY9fwE0wMGXJU8vmFWdPCIzpI8W73qHFiZzC+MzWb1dD
1Osh/ry6dLAwO/ocvXN1SNlru8via/B7o0Xffm+7XorjglZcb3bWxskmkcCLgdEldnfdITSyTx1O
4JZPMwnND0XAaqrdQZPOOmZH0uIR/Q0ZmOm3CV8+VMuWvmkbz6B7xT17poMDcDzV96RopmT+4yC4
7dKEKgpwl5gUn8YS1B52kA0+S2lAFTGhYaoO0q7WGm2l2cPryt7Mvi2AMhmxoNjBk/YiR0XDUWNp
EyvzBgKDgsfeDtQd19lOMlPkVZYxpw3u2KmYpXEjxGNeIwB11hTVSo3oIGxHuZcD1tLi82EG+0az
fdEksPudW/RaPB5LbM4vdx4XlaCb33hqKfAdIKN60Dbs0gYL2C44UFMPztREmx7Ssr+vQI+NyzOw
aRmRMszYDE1uDmTbLWUYLrgTwWDcKdhWR7/ZG4ZQ0EhkI/GyosVb7/zXs6kdxU7Y3OTSv9SuX6Q6
4UyDvdtTcFqka5DDp8MAizmiy8YNMOcx9YGZ5xr6SWU09XNB7Cb3MaoIdk928yytgWpOdlzskwkk
Xqk5zK7DZlzsRpoWrnSlqqYHkDDn9PebWQRTubYEqP9G1jmlQhh+yaWTsURhdpjimNk+SXu2QaCz
vO3f8XDYl27tcV1G9Omk+Mexi7uJMqE8PMCaiFGQ3xls0VEK51VduWyUAXEhZH75GeoliBiK6VL7
phZNWfMpDjqdaH38qVjnjU6zk34LPmPVWTta9NgNY2DAoUwk/m7PC+lnDcSKqAO+TwBE+axej1yd
IqlDf/W0wd0y4jZXGNsXewUYRsnllGwHRfAlf83L1CN4riEOb6w6uvFKPpPyWujKFYUNndzhoiSy
6JDyN6ugEmq0DOshK1M3AZdzwpkSMH2UNX1EpoGvxWdUkJV4eOkHtBBw91x1CjWVFowPASeekOXs
gKwq+8a64PIZg2mI/ASxCToIOvyMPfcgSz7WVEgikLX+xzOUl04Raf5WvN+7r0UvAj1zpme6AHGy
ZZZ70gvlW8V31DEbgybqLLO4TqDUH3qleBQzvbKMpmJK7Uj115TgsK1smX4KlwT024FbwuGXIlpM
z44/PGCBB6oB+kILBDVTFkY64BWE5yZwgcNQaGiaBK68kEkAqHayK5M7o5GaA6M7nu/CzCro/jo9
l0ES0NAGFac3w/kXvpbfxgaiLc0qpQHmGmKR4vG1gonJ4DQToP2l/eJZmR5mLP+n0V4ydqsbr5/J
T3zUBQTwhGfns1YP+tEzkts6kAdxqFoP8PF8FqpNc/2DG/tFWcmH6oo1dQSQr99IxwhbmlxDnZei
d4r+5N2A+r3paj/QBBxWJeVXAWHIamxjOR9Wi0EE0qgqduuLK6yuk1rLJry1JwvwlT1QylZCWlks
YxTILzDD5EJltvl9LQDh56pr3P40Xa51dsWiZvrgllNdrET3lSy3qaMnFPsllziKHIFjq52qbTnk
bhBZjI1AkZT8QuK3xxgmYm0qBZaQYCOj5n/hGnF6tmsBMB5F1Ztyo64NqKn0hS2biNszFq+c5B38
wQeKtmavllP1XQiQDt2/bHt+D8bj6lvy6AQ1wGM2VLyddj4/r//uIVpWdlat7wfTtoKKPjAts8zJ
ECp51BV/pwc6QvdPVNJCON3Mb/+7U1c2QMpLUECgqm6WcE/7q+7qEiziMYLI5qYxnBfgDZJaAbK9
O4FPIhAsA0kT9OWVIyIhjVFfRuTv56ZY1evV/gcXvHHS1nrgmXFbyLyrWRYGkUfvyzde2qeWleJn
QSS18GBwCzKS2cp8TkRq2QWog6czNguYvqBfJPcYnUUuo34ZUtxwUnZseQDsa1w8obElzxgpKcD4
2IdeMNnc6IVxxY5Ku946gf+a2dz46f3JVAX9gB1+pzMdIDyYc5FqgqaCJGDOFxeuHFAEFEY0Kp7X
soIqkUkeDuVxQR5WV9WdcNBWG0TG49RTmTJyf95koI6TleB8Z5+LE4gUV74FmzkEEvEO9okLWCsI
VZuSPRjEgAkBZzHyQEvBBcjQroB1lYSsPKXIPv+pmus5MdPqCuNA3MmfMZiQAjbEKMufGFy5E/Nw
6bIGUonnPjFE7RUrrZRdJToTvby9674SA734S2XgAB8CpCkxrnBF3LyZzUEa/D2Nh5siImyihFbT
0NhUEID26QqPMGWXCcNJodc5BKtt3OLwYO7qevVm33uowurM3FMdQHEaL6hiqeNLd0Ki8q0R9nI8
6SctbaTKplAXjDrqvpo4LPppVl3OHZIcJ1oTqVJjeezPa6OlQd5x0tLE4yoC5/Jis0ecofCPVAVo
vLkjDcPQn7SAEjDgn+IpG9em0lFQSdKW/HaRrbeLaDXg3szS0wB5JpbWj6V7GlZ96hj3amhCSigg
JABtj1iUn1EiNMUWB1z9O0GAd6GW/vd7s71fv+Y0v3fAW4cQDKAPpI/4fxIIuBpt6A9pegtD0BU6
8kJN/PQl0MpDK04nwNKkG4PjbrPkDybaRdf6el3tie3aemrOTXs35z1p4DC6zFnvfV7VizmVCDH3
C+GZxVVgX7Qi+5bdEfQJRFk0mKxjCOHRALKNJ6xkRwOY4U0VdUUk9fHIjzanoY0fFtHpdO4uh7qs
+kKOwXmneHmt6nKbZ0S4avG1pZiBJE6z5rOKfD3TbrMEC0iiyghHjApNRVVIDu8bVWP+/kFvFpEf
3xTRp2c5W/ec3iTQy+exhSyybzsmi5pLqSdSlmdoY36/iLfRejq2xKSt1zD+I82OHSo6frXj/VH2
F2M5dFI9M7k5LkYbKuAPG1fdwBi4dQY4Gx0E9r9+g8B0jc0AIO/O1qGSiEjc7LwhBp7Nho/4qHmb
s++RdA3vMiwazBQLiEEYeX/2MNv8n04TlWTkSAhENfUlZVSqqgfXBPxHnxZ8MpcACbQ0YSKzmnxA
HuxYl2HA9CkDVf0zxw7OVzi13owawRzR94on6XdQMUcI7K+R9Oxw0LQWldo0ExdwGBr3PX3Dfu8/
1cDrhvfokxvxRGbwTvEyMN+ewFy//XMt1YCZY4TeqBQd9h+mqfkwiPMx3OfIrn7SRtdk9SWNubuU
2xHpnlOM5DSWMIsGAylRPqf7MyFt60/ijJq5JbuzLIn4ti3EfhM+i7DSgcLjlQoKVFe+2NcQo8bR
EFUkpoHPI9jvTU9jTisH3HEO/D7XWyuebWZj4EqMp1Y6aVoCIFbGqcoFicWnnnAcNHZjnsjDQESo
2lbIAd+pSQD4LL3kHCob7mCHbqvxHLHWXtD27TSCvE/8fJdMp2cEu6pIYnz0FqtjJs99WCeWx+3P
qZUtOTi1iKvIJUUwpQ24skJ3SI2qlGnNGoeubBPrkAfBdMauhoPqQKDUdtNfr8z6n3UA6zOp6UXd
kGsHVA7T3My44ot/4Ro2bed4iSvrVRz/cU17MmN/Elq8fwDMrZ6oLBUaI77KTKssGWZp1F2kkWZC
yOeY0nbeimj+OAqclO+8mwM5+aiZWXhyty7tCYVstdlOIOqC9g0cIpZpcxSY+Ri950AnLy+AnYsA
Ng5WZfi5GnmdAvMJYPf9qGUeCZ3a4rPFm9ORATSmFGshWwyvPN/v8VbdqVNcTjFPHN9GSbC1aGHS
rskXey4hnl5CRfkjUhC9VwXrQhoy7WK1TZ8nOMFyAUYci8Xke6/P4W/O8LdrW6J+UFCb9iiEUe7D
PU0YLpM4Syopfj1B+HuG6fS3b+5OvTKQ2QrDuAZaucrpV0LqN2JK6OPkdsemc6uPPSc2duGVWX/n
XiULE/3/+fSPRUROOO+GSnv76JCHSPZ36EasBiuZzYLZCqm9nwgXKu7PX03Qoc3T+/qq763+7NYE
ZKxikRojfNAT/qqv50fOcJK4aPDgj90p1tZdBY9t3UJ97FsbCQHcDS/i7utV7b+cYc2wJSDV2fzE
dHYIkzD4SKm4OsNfBzVNMK3nRYhSm3/mCjGnk/BGfkaF+eL+NfW4xPadvqaMiS7DTfred2MbOxum
AOPOW7EVsVZm5gPgnUh2qzgzMP7ebSxp3a8VEO63UIufZc26j+7PF5QF8y3Qg5FjV236EAW2sXo8
cEEcfHeMr0rzfHznKG8V17mnc3snr3EnZKK8+1XIN5D6gSowoUSWKHAIStNGDOFjmfadW9J6cjsE
yjatzPuYrqcr0IqGrdd6QsiC6z8QjMP2h5gU1H7Gnvw4/EThHkCUFMg1Mm/AJiBpWs6clURyWs1h
ypLWJ05nEmyhlO9HDAeviqnqL0jtZ2NrSaoDucXStRejzvnuipdMLFYSwoKVXQkkiTXcEuO4uUc6
Ysub9CFaYdbh4a+k5Z+gSnvIwz+mdyGu2phKobquWLNozv1I37O28AIJTl3mu0LznUUGYT2r4RYA
dRkc3U0yRt6Kud53GFwYJiL4MzKwenRCB9D4nF00x45KF4Ebhy6wgAInhGCBZFveuTEHlP/TOHgW
D4HjJDdYxRGLW5KkwlGInmCJvV1XLw4LcoZBeNVdmlym5OBNsr8X33iIMt5/zoZ3p36cUW09VAox
5rmG6hTpRnzlHlqq++A83impbGu4iQe0Wazdb7uORP7QzC4+ZYT5cgCYb3X6zKlABuD4kaBY74XZ
Xd210GpG+bvzS3L9E1VUfFgMP2NXpwq6kGA/8AYcKy/nmRHsxliSKMOwJm09P/edYPrZzyz5owvW
GjlJcjigfu2ZAriTiPdAPOl/NweNJXmmyBWv0Wfvhof+QGhc1hjsjNmfES6g32+3f3eDAiVKN6me
fC/tpEzKJtXcza+7tVQ6ej+chslGVOTxpshy2c4WEulncP89USbZ9FxUSDY7lwfMuJIry3C1L19x
2iGWnqOHNwcMHLhzP1AmXVWoEUP9oWb0yxaw/8rdh2aqr4C7qkoRP//hpM3EbsUweWWQ5bGJRObj
Q9E4JyASNc/snf34739uT7cWNWnuOCrxJpDLkwuEqtN7YjzERM2o5CxXxJTRbJWoMLvEDhTohHVh
DsXYLsUft3GNjCOM7OP8BQ52rgo07Pbg/8/mlaPLOwDC/MU8augGSKPbdbFZPZZRifXs33kzMGY/
Uasd8+BZazuMcFEvy79QFgOg0cOCJxW5BN6GJ8y3psrHY8edDBUUTRupLk0pEo2VmHJJktbZj5A2
vVLlzNIdLwU+f8B2AgZmdZ20N5JH4LdbIpouCm7X37kpr9xPFN0GI9JLlBkjgvqG/zxT6R/Oc6rS
ENohgbpx+9qmJ/oRrwKMb0w/QctAfhm7I4f8O6rfPK2C2gZgOHLfvWRs3iNZomjC/rNr/7Rtxsc1
6pI76NR9d73oyKaCMUJFFGrlp2IBVrakhjfKV21pS88nFgTmIsQEGQYEGtYjSJ8CJ1juWUF6hjYK
J96jhUnOtCyk5yrnr8jR2ZVS3S3R6hkdvV9irxJbXo3IN88xOLIJp4Z274Adb3I40QFntR7taz+H
o3MSrf1oDvrQX+PeK8TXNOSE37NcvT18CFiqFdBXTLFlDT0tB786vBv+CUugsn3nIEI2bs3HUuR2
98YEjec95nHnLLDVp+TxNkczZJEgMnijPrKzvexT5NEKwRX0bDD6/RAc7eFMUAMZpBcBoaeJxXk5
g+akj1TVnJs6Stf8Fj1bahmoOqoJUs5L0fr29a8dq87mn25MOpbayni/KShiDByLPU7Q8vt9Y/4D
nS+ICYOkfWgr2Kk7zTn4eGi42FsNcIiS8kon3O06HEE5rm6B+JHSAbeEva2juViC4dS4TzsCGhNS
YZQ1XxxPhbQkpBCsnZ87WtuiCY9DC3SjFd/x96MkiqF8iBADyVwFqAVItQPLVBdb/Rdl01KEaCB1
jBvx2ZNVdyRKyA7xaiID0R+F2NLvHvp9HHHlOv4bcUGPxbodqLk164VDFyfXij5GPzBQ3DjCTT6z
GGM2PWDg5atTA/AcDhOou2aUkHdlN/iZGFu84wZBuL4vQLwipFvjOegYrh1kNl4uQUMv/oONSOJf
xs1xfzGILP8kH/N4peswGCQ/lZO+/PGT48IITxhYKY4udHwm14RKPQJxPg7Ud64LWCNArXZ+xWET
QpstuByal+0bLZ+lrXzQcF8ub0FFHzWsVizAcN+BTwM9xgUq4lFFkxuehfMUn9U6+XTnWm/RK75e
veSKd6Yf5HN56h94B1fKc7PgWGdd7Usqb6kV+JqPgS+uUsg/uWS8FAeJxeKK70uoNi34dfg+GQXk
ShZ17KEPH+RxrypucaooeM9IjEUIYsuB3+ORsBx1t5CJxjDHHU+l4GlX+ZeUXy1cFyoypjDd+lme
FVEbB2lJZtvzijwNaeDW4XQPVfwtEuFcH7coxsH2+fGHZgiZkUD0mRZc3BoZqr5sHgA6YOcnTNeT
Yb0wzUXQBiT6mrsaJ4TPikPEUPzbwvMOsICPC/yNAmTFKCM0IrVmkVxmuBX6Xpfgk3RHrskRwkTg
Y+4S3CytzPI5e2s9mT1328OcRt0tGU4kwrJEndr3S4HvNwLcxc4wXWLLtpqqNgpmG2PmTfWAgaBK
YyayxoL558Yk5sdgoc9pKhsHRepABLAx3uAggWokMKIgAf4YDAZyqqlAD7KR1s7DKOHPyueA5ay3
U4+IDImKTgoQwHYSo4BEsi8yxcAeKraM36V0o4z+8p5q74BbrHEvIehpuYDjhMGRQWShYdS+eefS
JvWbUZj88UGXyL2Fyph4rUtrd/4UJC5cwf2jzhJg2HSlj2geCBc9rE+1MfvUvBgq3WkgzLXDrsDd
vXjejQR3SRugtMe6ijVqcFg+JUVKxtmA9Tz5eDz8Tl/9cfIDrcXo4guDross2zQGkR/TRFZzl0gt
xKJo5aNltFPyml3do44cPmDdizWX1a12YZLSIhNVeFp0nZ+trYHEE0ZKNXGXAEOrzw0o5gzzuWYz
kQU2LXzxCJU80+NvU9aq69JwDTkI/6v8ZR5GJcaO1wxFc8z+gkG1l2X87ljY/A6xrIo1RwjqmCvG
RGpVYB7GBCgfupGGxskNzWGsFMcLePDvvZEV/rW1rqseu9CAg5ucRFlATkKjuYDSqTpEOjgXICmF
rPr+zwVqYBE9gam2uZB1ltHYUVn9TjNIL/ZX5psr9QVRUsh1I5A0Jf8YPmBJMdYYfDYZTQkl0w2O
K8CjDGrUXPXGnw1W+8iYEpYt52PApBrud8GLz0yDBA3x+w7mDZsEzS5SOasVmOt199xarZ1USOOO
bQLEUvmwZXvQbR3gUdX2/zO/WLOX4wukiDVOCHN/x+U1S62N0P0EVR3veu/SjRnv95rso1lHO2DK
tEwq0yDWZ85PpIDS49Bj479ypl12I88fHhfBFhbSITq0w6ETKPaibDwvrcLKpubmtxpkWZKPClzN
1jqBnA35Xj8omO9GZwkkRGvI4Lk0+IUbDJbtH8S7Ib5QcSuFgQTWOHw06LKaZ5UKBGy2XdC6FA5z
CSjH5frMM6JOdGEZxYsT7vK3AJ/rJB6qgVN2gmE0nz8R73wkhT9VapYaFZ9YYmJxtbimdXB0he1M
oJWn//OP4Yj8pBETJnPSOUL+v1ctAv5bxdZn5Zc/BQYXqoCQVkiHXOZzINqXJdsd008fuLPb2NGQ
srFGk+yCYLnVVkgeL614DCCkp5mqW9plgkcD5g2e+qntaEyKt2mEXbwxutsyr+PRi7pqXaktaNms
fHznFX2OCl3ls23PxGWYHd1cngZIvn9/7XwTiC3kn9dn1tASNuVe+mSWxcRAqSMINXN0beUBZnYc
frt8TmHkqocmKFDIGSxAFlLa266MskRDDZChAaYkJjUE/1Y1bn0Fdi/ut/Y8kMm4I7cz4ccOucGj
eW9fCM72hU6VXc5wpMHr2H4vVLg3rm5s5l7itvCUb3Fahv+nQKAqk81T+n6essg27xSYZ9BfgT1V
tLqrBp5cL9iM/8XsSsvap8z+XByMpqs7bFMqIBLgDwnq9VnoXwnztKpSD5mWAGeBfAwT5kRQGtNV
rAVdjdYYiqTi1WacxbBtHCF3nlxXq2CRZXDpxihJDisQ1Pth1is5UmXpVm2su/CGz5JKcPAU7Fho
J9BiPTp8XQ3OVrmo2rj9Sq6AvuVmOJn5uFF9UsCvTmRrJMGo4UAInixYMEY3q4CB2bTzH6F/aJyG
z0MoRaYB4jioS+ECIYYNpnjUSfXYKoe5Qg73e1eI+gLx2sFT0Wr82PeVoC/aASmCLz7DYas5qfzQ
ut5TvCCOcMrTQ4f59KaXpZS4oq2m0T8Wok8SgQkYIIjWKxKNIr61L97Ngge2lDCIdgDkzAtdoefb
+Pe/bISPKYOQUG3B2cxvs5sU6Ki4GwxsQAxMoviZWSq8F1w99JoIt7K7MqCvek4HVdhvnpUbAhLW
20Jsm4HmMgXkaPP5oCE7g6WxT0da4DL6cEo9Sx61QqFCxuneEF0P46PbIFlhs55eKIYNO+equgfV
5nx/VRPwQiS+pcEauXwowxehKDnqgRMJpN4kCT1oY68QsY1IqQEVDIkRdkqVtlQqcRlnKTiAPpYI
bepSwWZrah6RGaqy4Mh7ms1G7DLTgKJB5IGeRRNNtpDaM/ZYegMDuxtYZDlQGsJ1i5Q6LwlxmuFA
fD860lIRsGBnpvzdNx5UWPP1BGjKpfYUw0HbPiUsqGif3pUWchDwk7WwumNEEl7IdioFQnCr7kzn
Mf19+ORDOYAUmgWGRZOLrHmYXgzYc32nAhwwca9mxn0lZMTLz8gDl08IRgm1hsseirw26EDXtGJU
GzhkX5GSgHT02AXrXict0U+WtXxBB4OqXQwaPGp4MyqNXCR5O9G/pHisJ/N64Kwy5tmsKJrw/cPC
aoVWZPf5a+4ms9tyvbxyQLRpDS2XXDw8jrZICTNItm3YSNLu8HHuDgOallDuPMXKq8j1s8DScVoO
rcSTsu+UvSE3aVCQnAmYwp+4JtRaNseH4SxnRChbq4GZmTXtaeuyGPvepNAk93O7/RqeZwjUf/Os
aM9JuVyjPmbIvNLTXvb4/kXNGSycVhwIsaRR9FEu+SlH14N8U9bZtXMHuYaVr5ARBoc0XENptAY1
eIE0p2PayxsxWlKQDhWW1Fi7Kq2ixcvTotV931HIbd1XJDN1zO80cTwZwtoZIMPBZFnZNncVBmIc
mUpp7cb9sodKeIeyTm+XGh9h5KGWfzofv3CXuVYSuVulSSjRuoj+dEKDmKlzzPkxYhi3pj9KGUUA
upRZYtZLoM84ch0Hm0UP+ITYwmPom4BpmzTDyyy1NxVod/vsdWzEVa6mMGgngkp0oiRU/e7p0Ip6
jFvQPZacwGtlYPu6PR8R3lHbxtqMdGuge+RfBg7INEV/rT0SG2cFKXm62X7nuNDUsvK0WbyF1QaQ
R+nd4TIlisR+YJBLSGWMpczn3+5zCLKjTTMp1z1nik0FA6xdoXEDm2CGvmbrUkRtvFjuhnFYl/ca
Gv3VWHBYvorI3EeJlL2v5utY1OAOpZkbnAa1Mx9E6DAN2B7VZ5RxwIhzhimtaT04i5hWonbmdwfn
5oO7KOGWKyv9eqCiHgUkb2Jso+4e4dkaHkyxKZeNdjNiytx04dQVNP1UzG3F1rfSdLvG1EB7QKfJ
bJljvexFVPKPV53QlfpWROGSs/M4qIW0OqhVFo4yw1aX7248LQhBW23htIctkQyTv7nfDEysJwuF
+A8kmrcoxnrlNNE67lzHsrqMJ99NSk+Ku7eR7BKDfAt21YxfMm6QBj0Zva/8v/vi4psAgqSWG3GE
1S0OhqDozQ4otCbKJrLLyr+3QkXvE/0DcgJMzGR2l5+jKMXRzZkiDMEKDHmXNKSjnR1eNR8fChkj
1XdK/U6TcGUH5EbaUdpqa2iLhTDV8Ohp4LJF2NTIPaZxdwS0IctTynYjN/Ymr5f51ZiddW6gZz6W
S/p6KxtuJA0NOLiD8YA/C76iyG9VOPjVgfFhuHrRaLBCbMZnAZwwE2Hvhjg1mopkqoVFqpQILSGe
/Ad1SoVdqMwXqjnlVmcpfvBvlprBbv2akPzodTH8fWd2YEn+c2AEWrWHsC5x7n0TEgc54zpT5w3/
kd58tAmOF7Tw2V5Rrea9Xd9zdxtDvpzUgMPb0bBibidjoNOss1UjT2LFhWx4W9t7hZzsSeKwDbjq
9W8B3tW9xGzZiJe3A6SYavYyzCeA6S+4bIYustGm9GeiSWnDzGVHzkoAmglEHq/mrrTamKO2n80r
pPPfBwv6HILTl4GsFMB8yLnmv7GA7zzyuJvGI44ZMATMBTNjIpRUXN0F8flWAwQGHgBJb4q0A6xq
ReUpWiMVffKJigapV4K1Xfmt7FmzT8IpZlIgbBigWvmnnbViO1SPcvcX/Htz5d4HReUUbE7110Km
JVNT+8SM1D9RON3aapGLaTlShdGSNmFtfESVdq+imIPlxMp/b49dMYm5/caJBky1io1cxcwhN6aQ
sBK1E+23uL7JLlyHuSevQewQJrh4coOxBRmCYu8ww/E8JUMAcApLD2umABONQV+1LW8xqPju9Q34
vUZNfXNeE5Q0tcPPHyXta3KByyWr9CXGCFqTqdCt4zz6FO0cvxfbsvVyb7DhL45Jsdb8LFNgNsIe
iLyztHlAoCmkwIMIlVyEv8E7JTRUDwbM+MHftarCUH3JqY1YtYGjjZLzPQMTq9otIBDSxXN9aaEC
pPuhSAzpITZpRR/9odXis915tP8VY+Mg8Aaw4pgShb5cyZAl+AE+Hwf+q801OfFzmLmmPLByb2ye
LuxyDmwWi/bmTLsLZpNc9PVcOT9KgSWnMSJwS9P5KxAOLgqVjnVLNHCbG6l7XIcALawg//NjvbyL
5TkVgVlJ3zjXk/wSIFXUO4B9oXZs441Gg5bEtMSdJt76R+e0nUS8PrlYKf5LJzEIbj1qhEtAnJ+L
4ifJ2sOjhNIsOQzUyYjlAQak8B/Pm4r9m1CUXQois1Utp8LeluGtjJGCqMnIITK/HvnFdAUHvM1S
36Pjd59jY8JGYXDxcqLBDb8GjebKmw+jPeKAzHvGpFOaVcX6A9gwXdPL9wE5YzwyDGpit0/gX4JW
CSWjb6Ayoi/G/UfnUTkU+EwiWtG7dOC0tlGil69QDqMPN40U8fQK1iIj6W4I1wWZNOL0EB03BwnX
4M9guSMc8PN2X8L2iXx6hz+13TtCHWL15RUKeWtc7+S26US3yPiamNl1y4Sp8ClqEHRMSp3PRDfl
Wqx8EDHh7AXHktMtwoApjWR3LZNXyUz6dWvWQxAOYU0l4MwJQdWKcFFcvYDSsFRDr2ovY6JKbvQY
A/M16u/RnmC90NbrUSmlRzedsNVW+/6Trtc19L6Gwe0JWmmMU81144rQUmqT8YFdBOd6SFY9pFYF
PgdxPtxsRTSSP+HBHf1NLyEJwyv80DZ1XCP5VEquk5v2JGBwL9XfbJy61bHRxcUGHiiSmzQsBYs+
dGeW70GtIzaOYWI9aEFc4ktu63eZpnS3q59vxjgQYKSy8Q2lf4Dqq/Kf6Rk9qWoFg8UAmDDkbhUK
Nkr6pczYJCiUB1xmuVpJKtldPz9AgHJ3SyqaiSvvJnrpTigcMsxyiO00Vtzso6kt6CTpJiRyj6cy
ZN0OpMNnqlRNVkMsuIe9kood4vP4eMbO19stj0RDVVRwQCmMaiBjU2aZuMTq8PaiHJNqQyOFwFru
IGWf5uQCRjeZxxjPIy/yYDv4/1gDE14qf5luiytHUaAwBzJcpI3A8tuIVYQLRUProEwQde/texQy
Tqtm/xKmdXGoVyK0llkfFmxp+tkV3gNVpUZdmxShxKqNAbwbf/km/WjeWAZ4
`protect end_protected




`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
U3sDNM5d7jYJEIZQTnFuo64E51C+8gq0PfGADcNjuAMCEE266ZL06hQGQBM0R+DrGmrgQrq0Wrge
uPAkNN5G+g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EY+X3Lbne3q/n8WMTQaQXRPOg34ay2XurtUPGUclFnWfBmzqnpUa8B9ymki0aidTUQYQEm2sh4CN
XOEOFCD0dbL2NgHaa05x3mCcSGq5dNxdn2t2PxrhLN9Qix/dsXnx8Dx+tcL5bK98qHkWv5TlPw9F
mQlgxUunse/mkLNp8o0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qejm1NMrPCpKtCQM6KmlkujDwbNyPltQGSiXBml/xklqOs6mwCS/d6S4AZdUpLLD3IR4u5jDDWVS
tBHBVK/11sIMg2yoMUaMj3nQivHXak00Ja3ku85yUxdiQBAhgZxAUSIYncV/h1DeR6eez1FtmUiW
k2R5zoT4kmn1ReKvyHBVXzIontFMNGOVHWDd0aaVAg2L15OVyS1Ff2rAUNHwsIDpfbkawwiEWuBY
HzkvTYgTqO3EjjRG7NHalOWEUrsKOiTJz+TKrcCeI26X/hw0q7lqif+Pw1fW7NKExvU0pb5zxe+g
dasyo7ekd1eAMBAc2D2qxnWrV/xT+mEZ2RjJIQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aEJMsL6nIvSfDKkxRVE9/86hi8XegqbQQaRNO+NCeWjYCvqPygToNaA+KX5cbTCa2ZJDNbNP0LqZ
Nf/ztarS6+Kd+yLfIhz+p4i18KkAcbPbJDi06aJfDKPZPGwgcfdAZCe9NmwjCDsNRUxF84DUxnan
NNczASRvUbnjFxV5LSeJc7fgS0ON8ZzZwIxYYN4UBE95NRZiEnndErsrJF1EiHhWW2etDqHUak7M
uJPvDNPgWyPWgFZiZqs1RYHjZsPF/LkSjAqW/s9C2dc+h1j65xJ/pXdhlNc0rO0z+LAHVHsTq/xf
4rNNAVJQPqr18LJzZvqQRta/I+LZd6EjMl3I/g==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
opiMI9un1L5qqubBM3bYmRo7L3zSLSE74WOKnJdA2zsZxyl95nt1F01km6bhA8+lOnRZr95jKUno
BVqVLm18ciDKeyCqB1ZqieL/IRXh35qDwHXUpEYaR9qYetWe96Rfmlgcs6mtV7gOqeNSetRrCEQD
RhAk8Xq9TPOwAaBY0GGCiWgPzhrabcl/GNYXx2aBQMmW0J9rLQ38Hixht17xBx15Ai50jBhhmsR0
lQD8BTlJMMD6fMBR2PAXv2wncn8avzwlLh19fU9rAxcZyfLMW/X8q1Js/JKQFdm5L0zIKmMh+rTG
91V6Q9ApkyFQcPKOXaUBzTBYujWOxjb6150fdQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
V5+XqY6/KmzZKYOyYVBUe+3bN870OFCeVmp/kcSjztpDExtHlsM7vQjvaeLLq7LgsTUWchr91fDm
BcWUyxISQ6O0ukpTvBtXqh3k6jhpMYK6WWG0AxglmJ+Vrcm2v1qCLAeC6t4vatuW4PHgc4HBloHX
SA62p45b7fezLVMI/OI=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OgVTbizwEz1D5fIn9QVCVHRE9bQ/skAgyhfFYkAxhK01ppsQIEw/6DODTHQQRJeXHNFg19LWL6hn
Ruy/2+40tEWd6FxiqzXIe9DOhxqxnB9lxu1o7DXWYZWCOhfKkVKMsMlTDbTvFpYyLOkwA8aFzy19
5qWihLZMNVvFPKjEJdocORPlHzJ0Y9x0/Tlhoya7V6F7b6n9qN9zK43VZ755OaAWnh+gfIIqyyof
8C1umBq362Yld3QbRDyVlrkdxHQGPeCBFNzdyydAoDQJoNbJ9LdU5xTQJaXbQTMbdc4nayvWBA9x
Bp2aZX50ImADwqnWUo43b23foc8li+MluopNZQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 71360)
`protect data_block
wj/+h6gd6HK34A8makK2ITvIR3YqbSW06ZtQsLgb6kmch0bn4LM6uwKufbjte7dcwr7rpC3wagvl
YWmkni1XCZBK6fOv4cmXqHoYYzV13j0LkDVBrbt+AwsrJtI3ZMI1ai/Rj5w11aEFYF9BOkkv91B5
sNYggApG5G4weiDWZmqsUmZKETliM5M311eeeAm3Ux9UA7Y4mAjgdpMlhhj2L13RXa+GWZtLELE6
8nIID7+cU2oVvS7TlXrmHsScG/Rd4mEfGi92KNT6MIVu9Pp1rdPyobmdi6+SeSFTdULkZ6+8WfD0
iB3323PnBTpEvBC9ipIN0WiEOgCn5aHdbF82VHWelpuwq9s/uySlcBde8jXQ/wXqm5rY4Z2DA5T9
wD/IjbVu8VwlhmXJM+u9Fhi0o+iDb1noHjDMcEHa6M1W5eqaMqAnf1SAh9geOAqTT34HJ72UZGVJ
wxtiNEv2+oTsAQRrbUlTzJtMVuSkHnQ25OJk6Q7C5Q5jWQ+nVtdfXi4tslLQsEW6rqgg/ugc79SV
94Eb+9AtemZbReRJSt7VPjitMdcIr4sLbSWt8hv2Ar1zJo6uhV2GUivmpH8jzo3w9lYelqXu7Nqy
cwIExdpqPUTdNGIL3IRog5LUwmQcvoQDiFb5vpUAC7q09i0AhnK9S7UYqeYdut2Biw6PEAfesIt5
RclveyGm4Ko+FK5rfl95Q5zO2KYEOUJiu8WUwaShcHKx18HjjUW8IIphp6EHbC+NHMW5OeEqv90y
76lWcQOVt6LAQay8eB3zRX7NafEL+1Qg2WrUW/eeV+WKSq/CtIt6dTDJn9qQUU9azXdKdzUGY8H4
ln9ANKVPfqNGynpwjN5sTupQnsstEOzm/MJrWaL9FBQY/9L2grg13b0fQrRyxaq/p6pfA82mR39Y
cdC1q+g1wnVPrsZtY3/m9/qZPVqc2lJIsfN1fkrk78MmOWrPh83DYNTllUj0P+XHJl3HHuW/ysgY
9bh1MWmyuSaEeFq4bnaEf4M33VYUb9YhGYkYEOZHfYmXeZ4Ql5WzoMgR7eXrLK8mXT1uowham51x
i4jnSL4PKF/2KkQEQZinYSW/f7BwduA7DhuftTaz0Oj/tLKpCKA6oh+0tRrxxXuS2YLoeWYB8uR+
BtWLPhI9jsF0V+ScpC4xs62Lw/vtqO+Dlq4AkX2Dtw62JH8rLbjuS+EJYh3Js6YOGlgCD85scg6I
LArfIVd+jBPrlPo7wViPvaJZUBA+NQGpwuMJjrPQWnTbJPz1CivXHg1bRcm4jZhyXICD/vE03Jz5
9G+q3R4I+1a99tK5atCIRn9Wo/PBX8z5400aUGFSDAuBxgxUjLE8GOXd+3I+zJsU3jRu4wVhDoM4
PeL7inNjgAsrsQcaF3UxixHpvLKHEX9vhvdmCIYWneS1cHOGHCFTwUuE3dNlpMtjXclUQVqE/w3a
fb1dQYtml+2ts0ZjorkqY4L6XnzTvE51ZEznrDORbm/FUeIXUj8dE21LZEkfy2ih4rlZMSAWuf0X
y95iZZcmItcBRCT9oxE73zQCt8vcM6meqpWX40dSriiGSNzGcteMZGxNuH/1VkyAYdSrdxPZYQwo
iKMwIb5t3gJURp0PhXYZ+O0155u9G0krcMbmeoq8tlvSkVQBp/INuOvqiw0XInhCJS2/6MuslsoB
UdJwQJghSkcSygGOOHPe4LErIlOxMvmWs5hbKjgen/QookWf7R2gMAbungOXFwNjKIf/nqNZzuzr
aZPxuG2ylu2fIUVZicSG8hHlg22GrtzCaG4G4KmSBpmpwGycdONd5d3SAW7SSXG2YmNvhX6CgCzY
86iIpGXAvYdNvmm3Lybn0aYqfMeOxdvhFvuyKBycgW9lS7W9DKsF+JZXoxt0tcxkyQlwEXxizvEb
DudXpobeEuB0/SyVnK92kA9rODMXkuM8SEz5QRei1z6Wnc291l2kh4pWjMJ7Fs5nfOoZ4bI8J65k
kXH9V8fg2z+TGJKQlhj5rjMp97msGZADLfKOUBCKCPGavY5NR2vpxSSUU6zf5HP4IDsJZudnqwru
hwL0Sy4s8te5kF9AG9HTas6CEmEc2ByOrYTTYgAoT0W/LcNKvZQtkj/zahfQfbCEuPd2RrapI9ce
ItVtjduWyjmwJFe5/oZJSyYFwPMnxApnLZLij2Y9bD+LkEJSX2a9P9Wi0ceOOJxSWARHCwTXypYP
4x9Elh81Au0JfGNOm3bpq7FGaa0uyoHpfukrUT4gDGq9PPmPQVAs14Cols1Ec6HE3rNtcsXKYVg4
Ez6szJuq1K1SXiovVnujFP8MSbe0HoVrr8ljUdVelDoDvfJnHYGAVojF/2uWzOfyzSZqZgUbs6u0
8NcAJ+Fr9d7Fws+um/qc6bkzawIfm+3sv6l4SwbvQ4GsiDDvu8kN53RRiWWj2fqERW+kx0bf/n7J
dImRIc+4y84QfDvOaJJslRtS7dQHdJn34R91c1uenL7dTMQIRBKPih9gd9wkY3EqqyiWxt+qXL4G
G3WzcxOYxa+vIClEbwQcbT1dd/RdzyGZw1NRBBicI2o6eJw4QZAW1IOOHlCl+C5sTpdB/rgv3M8e
9xayoOQ8hIUqKCi8TRwWCLZRRhBH4cLT3jvWtOn9ADAl6+IMFKqThAJq5oh4h6vGNbkoWEnN6HKV
459E+25xKMh791zZtMz50I76VF1UTlXIVym9qLdBu3mzU5By6nlDO9uQmnYdMa5mjo4f9IrJ29lt
eS8DtHz7erelgur7bQAb+gAD56pWDG8KaOgRuwODbT7Vf6ygO7mHJfOQ7/1fT2iCALDDfO77/U8Z
7MKprb2nlJpjpy+JX8UOadCUIdpS5iQxriIWAPI33neMFIZt9hUpEtmjRcxBoPULRPkTQgak/SbY
3e9AyzeuETgp4L2Qb3pqa/D2ehXr/D8cA98pE4pwuIvNK6v7kGDZreTXrfFp0dRFMSAsEjK29xXh
8prAW27AzdZgdj80Z1iTVeIr6puhkOX+UwEnRcBAq7yEhW+5PIPmsmffXjKUTBidathnqGMwJsS6
B9Mwyr+8cIpY5ec7UveI+t5n28+HT7IdkjNca+3j7b8BMceOj4VLjBETpphkgv1Vmv04Z+LY89hA
BOi3qFe1C/yE6Pa+tKSh7gZR9p9gbvhBIp+jC8VKlmsQb5HroAuSRaXtc5nsnxox6Qy0iM3p9ita
yjKsgwCx8nyxbntKiIA0diXrDSbD98fdwALUWIZDoIOKPHcNRYJnDW/40VIbd/UCxFNGcLckZWSV
DxvLhIt8lM7ceNf092p6sj8isH6O+oDoX3qLRC6gFeIidOR6mmN1BFFa0uM+wiaD58bzE0Ts6eWC
1cfIyAYd0dOjlkQe+6HXGlnad7OD6YxcjU3dogsMftMkNuM9fvDcUe5ljnrCAbRbgYuWhMnXqG96
l9niYyhqEbqOAZFxIcO4Sab4aVA2kUvciwBLmKaXybfax3OF2sI3jG9lay+Nn8N6vYzN/tHxm1Nd
XNwxvNu3XAoQrl/7xekJ9UvdCMo8OqNbGuLL8ClrRRwQSIqKG6dSeHDjfadD64h8e+yCyjGXIuhz
B324nW8CqKO4NhHXdt6HfXzbuoGs0msoVmoYRd79g2vSNBc55oqAg7fjmRc2WKkk/YFJ5IRhhiWf
RbGsB/Kmr3HtZg9U17gVOcQCIv2U7AG5Ge4WZQbd/kbydEM6tkwyGpmI8zwbvxld8jKwujeiZ8Tp
vgT5n1S9ZJdfLZGWW+LwRXVUmZUAd9fgnk9v0dYin1N94Binu8V4rlro9A9vaIfeRB98KQzik+5m
MPR7xpFWIf5TFkD92TOXN8qW378sD2C2JOM6UldMbe0yDPNYX+Sv8w2WJ1mh3g8UbXkMWGUi9NIh
vN9x9e3UM+t+hlJ+f468CGU8fazVa+EfPuzvDq69GWOSQzzzuQRUFrVVLMPdBvpORWGQJ8NmizR8
oerrGRgVYC0TEn0E0X0LXxLyFnCaxQegot55MxFKbW8LtquccdstAWswUDTsXdesnzDJzYGYNPhA
qeOnNzevea1XmY2MjOGasl/gkuAQZH3GVZwuxKpCEOxGaDN1fvIxN/Q3PYT5s/KswmCBr58wfRXi
K3+WjEyxT5TPssvOhZnc3lahhNEhcvvGNEnNWXOsj6sEXxPxWU6Z4+FTRZEpadgMAsqbfzM+7BLP
sCh8neo/Hezb+YYUE6A/RJwq6hsmk30CocvTAem8PaJrxO/LplFZ/Dm4aocu+6SMe7FnbrIcGYVV
9sknlFZe6DUkgxfvRIGpioa41Tll5qhCeMCipvRZwJ4Np5JmpI2YF6mpuCvRJwpnMST+nWqPGEHd
PRG6StB1nw6gEVnzPubimxduVb7ADit9g2+kr6dP4Dr/mptZmmv1ixTQJnmq4/c6FexILTJM3sKl
a+qpgCIczGF4Bdx+uH4Hn8kX4JnfbMtzq3WE0J/bmEePaKchbBqmxU8TCJ8iboxEkaEnl/HPPY37
UGqerg9bFoo/iVOKenr4lB+SiY+IUtE4pt7XR0S1ZfHXt60H+k3hOtsTQLWJe5hOHFBtxHAZFwmm
0bS6htx46pQgBA1KLPbZxktPPs6Cgq1nNlSulE226YLHkjVrbd1FVchGZ10KVWBi5vGuz/hI9OFC
usk7NtaWPHZ+9m6fBvIAseH5bsdOzNK1HaJ+Jh1rNvTTQhKWIAz56ypnKd3LzrWx87iZPVqqKu4f
pOVpERp3IbWXn+3LujXsEYuz2GVGzHBHtk+/ZKMTPbx5DkWp5bUvtqS1r61jU+tkMScD00/xYYvx
uEnm7ccCT+qj8VNGIk6nHEK26GhqiMJdy0WHbDNT5aXJIBdxURFSP1MP1hCUclfEirGTofPbTnR7
RK3jOOONSI+MTttbCvIV7Ut6k5KvNCVSDrLEumoB+pRaZbEW0DEX+43xo4DdrgO20SsjXxpYVFXj
+GPzHkF0ahZ8mzvOSVlKf2BQ6KB2Lj7OJAPAA7w72NtMLndge7LyLXohLG0smHHnwhDWlGG5IOBp
wRjaS9vtTbvx7CD3AKl5JM80Kl+iR3PFuaHm1qLUp22x11fX1HucF4ByKnI8S8TSQngxEMiYUJcI
l+w1sqbWMhQD6oCuXog+d0N3WvwZuKZ0r1393FUSPcs2Ph6TDwECuj4tEYo1J4mpWBKtCoSf+ynB
mAmlAkihw3hphIyOXlZislS5/cRIOWoLuEBJBtGmbKKpKPr4MkJtrpm7aVd10Wzzzl9EZCv0DQAN
nkUvoSQDmmJzd2GNQQppRiMitDnfCZk6oqXIa6rdxlPH7CVrhHrUym8FJXYWrpdoLSCqvZ2pGIuO
hXDnlDsTZv4ZpSfINxiv06oeoq7ZPuzl94E5vV/iR7peaDSRLTYnagI7Fu2VyUfMzkJ6IO0iAyGJ
SExUNcY3Ps2JtVVf+zCnHI5TjI59KHXEMvfVB1HKsDhq0MQ/Xa3MpNo25DGyufAQT7UZDl86SyeM
6gtuccW3U0OBa+klkNqdnkaXCQSx/qZFBwkmGN43qBSJ6+f11KV5EwFW1lbUWlicBs+s4YFYIVYh
f7N/8MjqsO60GRFuDZgZZ1v/jB3NLBsyZwTuulRni/b1+hqif5r1sE9KEzVt5eqG+VZ/12FqR4zs
vk9XVoWgm1nMmaN7m9LSmNzpSKkPFETEGxPFwgKMneBolwNM6f630WqnN3+KkEebzOfQL9bzqLY3
pU6XQTIVgXm10aPFtuCAK4B15+zfia2M2LGBQtdAEW7c1ZYTarDYRQzrIbU8Or10tVUM1XCL4MqK
Lc/o7xcHDAKrbKc7vJetDMnrza3Rw7PYpiOtZYdYRBA+52EEeYKdxhXrmWabrHBB5s/+RbtaSIWn
oM6Hz4o4dc6KRZ5mZwEA2DmYVQAXXKW6YtroCFCeihthcTzEhyLzZXsih87lZ/NG7/nZcRLolJli
eO9FIrG+xMKxKNoJnNLE/Bd9jMH60LN02z1at16hz7P47mJg+mlKZIclOkeolk2zLNNx5tqLwZi0
FS4/h/G2AGuYslsyuYHcIoN2M+a8LJxMJUwLTIQ1QUpeh2Ppn+j9rh9wlndTxTse0Xh33nhCw06S
moUAQsoSrjSmhid86nmyjKw49D3J8P+gICeTl8i9HSZ3+hwPCD0AcR8zzNB9TK4hfMyWf8XNxrSY
hHydVvvE9HQ85LEb3HWoAxE8HXFo+aejF1XBplNtKVr+4j4U+oiLJGXFhNNQ+QGe+o2FMEEpdThu
0hwDQCYA7s12etYDqxmq8zVzTvcpgZJu+BJ+KHXr1WxkQNgE7A/a/6FoBwRqwFqOPWjKYsf5+1rR
60vJnFyhxpa1g6vUQ1suKZqpv9M8pZ3c6t7OzoXRE7kNcMQkia1BF89XCJ8fMsv3Wjm6HPajZkjI
bAaIZu9DSfkpEYAc9eRTpPgv9dOvwBrYixROkItI/RoRtq70r+93O0Kxgi74UxOrWemQCe7TYXyJ
e9sp46VRJWl5lOT9VkkK9PzPz0g6kZ4IeyY3qAG1UQJRWVBKpX3mZBhmaDMXw5An0/J3I8P5QmmM
wtyiY2i2qXenmtbQsIPefcK1n+vtGrEsBqCy2jTs74kuGArgkrZE1mTpUrO2HSK41Z/A1D26u2S9
TAf/XvmSBe8aw7eiB3S03UQe4Yss44GiSXrpDs5r60XWiOKXM2482KkUtHe/z+EMz29kdwuNxr0f
mIdQrzKWwrZac4v1tpL9Z46Tj4F64S02uARU13JBqNz+B4Zh7QPky/4bFmBUjKrCoDkynd33VDAL
VxgCasB5ZN/EV7c6EeE/gVptPJpEDa7mj1nmR6KJWq9uSJ+4qL5VHxDRI88tuykCnsSsIuL4jCuV
ONuDwwnexYJTE8II87M1yQTNe2y7UaCjraus8T4W6C3jaTlDpRmm7szw1iOv/KUm11+ElE5ofTlz
i0XeE3ZmQ1ClhKJij5gJrFgwfsVgMChbacvsJRxxLWXt1wQHRFeyCw6Mxc6p7Mzvvbkd0WlatZDl
bidkix/sE5OqlrWus18h5nfEaYQzGSDtJREWwzRsXY3XF3KlE9IF7XTJ/+4q7oUd9Bc0ltd/90/6
QVLkOqSFRyHKYrAQ6n/JxwLSnLDIbHZ8SvEMjfTONJ8ASlaw6vCwDBGu1iRAQCxUVkHQPAHTkp3j
fbobRmobVfpBga/QNCkOAVJpFi/Jtkj5vfecK7vJKyo0qa/jpliac7ZzjqzIpQB0a9H3S7BI01wv
Mji+6G9WSmEzI5b7DsNPD+54ZxbcdetOc3btHVzdYtsg0Tu6sEAvJ1OOim7nO/4EeX1QuzPoRKma
QYiEf3WZ6g1xNfuVvY6JC18Vg25LY0ei8oPiYAT916NWv5i7iXE8KMo97NaJfABRbde7IXqZDFs3
h7rBtLgT8n4Nh6xAgk04iWUaI7RzbV4Xwx7Up/GwCqdOjShWiFQuqGe+uX1jGlxEvLiem6f66VgR
RxVhzrRcSO8zp28PWBLKF9+B3MGbEaQCL5qEoz24UKoCnteu1rvGj+pU1jSmGH7z6UPEWbs7p+C/
LuFJa4O0j1sdJ2Z3ig9z1QXSZnXBR+BDTygPJfa6zgdDI6ejX/GIW3GvDekI3nyNcLSgUayGrpvt
LIaEQta30ErgAzX/UI4c9IfARQtbYf2I+idGEZHC5v9gasV/HRTB/bFqxggCJpoEb7MeXf9DZE7z
4bwm6V8JpSWRT5Cj2WtTOD+et0aEqhTIG/ZAP41/jhv/q4HLIpYO5n46jjAKjZMmOaJ/e0H4mi8S
5BRn0T1wbKpVPrAB9d/4eY3dSzJDQ5bP4ynL8FlFyiKAEjA6kmd1NzBRPE0PpMM4iT9OTmDreKVg
cW/4F+8RR9SNfWRyqKdOjzu8qR1NmBx7rzz5Z5dIF2B3tnTkj870xRU6cbkUG2ZidYuDIVmr3rSn
pR5TYEYh6xLv6hT2o/G0LAxUZzlevC5DPS6myN/MoV7hts99yn9qpdnib4prQJ7OCuekb09oPXWQ
0AufP+9pN0DMvN1xDHhPnmywmWBieu9nAYkGlkjNYrbXzD997c0uzX6VNMph2m4+MtiFFZLXTOlS
MRioDPl/cyUq52qUsxLbMQx9mjz+W90UUoKiTl3XoSIjUBMPd2Qt1vzOEMtE0YWW/5wd7KbkChg5
DaRtNC3vRnPSBkz6pmzg2HVFtf/BejGITacNNYt9adw5pwwk1QQfyZsylL4oc8JBay4a786xkQ7T
DRklwOzxOvvN2PLhvz1g9HdkprRVxfe6vssV0GMJ32Mg4sOciBXkxi17E/tHPNyfZS8ttFpBvuMx
oJvX+UszfN6lHZ3Jk8Vuc+Qup4gPczoyr1tSZVbxudIlBiHrJXCI6qpQChOGe50NsWppkFVoavAI
+tNHWgkxw7p4+SbiCu/A7Jcpaf05BwMGSPKaEqDAYp1CROPWH8XvYTcelS1YUqbgygCcNnFqphEt
XPXvll2GajTKBBimmfN267L4QhMu4X3tkWk7biKsgGoK+/Gty5XngamcuJBHi2GkH4la0FHpeNHC
03NvnRwFVJAOlXmIsrDpGEGvEkSabs1XnQ+9IHz4Dwp5oAcUgVmopc0dAdyKW4sxurV0CmFgVJq3
+YcP7Tn6vaA20o87MNaGwrWVuugAl9Zq479d4EepQ4KpggPYNHTxRIFBg1+OYYdTdrfL4TRGhthH
HR+i6smTHzYqSZCsjijDWFg8NIfl4ywiE154TmQbAk2hhaH+kTeH6APSEdzTPkOof8XVvSrCLXvr
aOtwOJkxw2fjpvMn8gUoonkuqg+MlRAzimJHxADEbZbL65hvr7ClhmsnPZ9IfigtEdeSFAydJyre
nIZqfuUM2WDBXTOllZFyL88wEl+ZbN9lKM1RRCx0kU5u0Ya+SevKHPNm2c0dQygF7I4puzJHVUg8
5VuEmL+k/zRPk60nDbgd+wPofnRCwgJUkpYZCwXRt39jXZ97lqTSXejkx1ZqZRAU/JYBBx8r2iiv
4v3x1y3Ypxvha+X+axlEpvFB8u2FFTzefsuTOOcVB4wyTkhJUlaG4XskAiWTd6jm/li8icNR238I
mIKxwNN9rPRlaUd4Bl9tm+4jTDxyHV2JQSh8lcyhn9ownNm1dYqwWnfavLSMHeevhh2Szr/SlNT/
IV9HnhQ1uby2SwfurZ6zR1G/IChuHstlcl5dvM0MGhNq7KjRglkmvE1IhzNf2hzsu9L2CX+YNt59
QNFp4X6K9wNeM1W6wt73OWhknht/MdrmPiLCZGelV6xuNo5rOFLAvHDmvEQOXYPXW+mkcjb2H7ZE
jyTO90yJ8yIycbcLsvGhMZ6C6IZ+I2EU2X9Te6kRHUpsi0LeFKoLF26efY5+kmRZz1C1Qn4yD7Ie
MQbsStd1A0T1gdXHrI6FtPfnspLSJ5SKGSHAMkyafuY0dvVzAiDmqexvtbNbMON625zxubhKfAxA
6wSKFlUEeMo/+zwlWlvsVzYG2nORhbjYqsx31RWI7AAZ4VABdmYWnNiIoL3MBLRhvTUzNnVPCopw
r1b30nXjQK2t1Whn9L/zEgaj9QxturZLEQ5MgNv8ylGcLNjyJqu8Bs6r6HPfwXrbLUH4S+apvvgI
cTk80+KVUL+evuV27xOn6Nau5nI2GCy1bcXu6Bl8F/ThVbfIafIhAvIfwn2y5kuc43+qmuHQa6vA
h68/EZCae2EU1HkVt7hx1PHo8RLQdinVv25InGuvFBSrNv9Xeam42k8zj1bnJVoU4J88DiHIQAIh
s+sYNK1YtDqabNDtMYuewPzFTWRWSADJueDLfMMSxsHK1HoXndw1nBXlkZ9k6H0EbqTfvUoRBS9Q
ibUttFpUXCJwte85w+EHFv8G0v6kTdH3L8WUQQjhUuq5rusllnRaIBr3XyM5D563POwkmQSxUQvy
Z9QrAkTrqvKKc7z87GNMPiMT9GlX7d2Wl57Of5rn9o80XmUhRJvmL7OHLLy2eaN3mFEuLFwhLe4L
QCr+Nq1+ZbYc92PEC2ocIH372sSAbqxb4QbJ7C7UBSDepiqnvuOvUvdeDEStzDnycD38aWdmc2Tx
RKey9G+/IxJaByQ+fVqRUIMT+HW1DAEMjjs7uQYgHsZZRFUTtS0gKdVAi9D0I9UDMSor1fcZMk4X
npyo3930FCvXqcYH8jL8tj0U2X2Eqg3IZ1WkcoQyuDpdDsaUFvf2XXSSINJz6DmFy4y0ci+hVEnB
cwNekmSmhAzauViKqBuhJUhxtKmXRuZBmg2LhBwi1YDucFVAqIvpmhl6C/efYWXvYgq65eSEKsFb
GkIhmK6LvYhK7Uf9KKs+FZ1Ejd4+iZ7fCicB3lsCqPI6EgpZkqmRUnPm1X1pZr9e4aAqmv1BQaTC
xHECNx8d+w13MdsYq9FMUsEbyETRE3L90teAto3vx2KA77U6BMG/BUFZRYQm/CQE0/KFjYIA3zGm
6j5YFt3XN2Zvk1qQGPcS2w55AnsXDJ+GZBu02I2heSlDy5GP8iKkkfY4bvNDzz8vXZ2+n53FUGht
9a9eSZPHT1Nc1aDOUmDYCJDPWwzDZqJHMWZgQZlP9bOHGDstYeZIdx9p4PVBI99LEGORqIi6UO9N
gF6JnL5ppXldmuhol8cutcTTRAaHCNyBYtig6h3F8LoOTa8zg+OndQ3QzN0i5AtKVsnxAR8nGm4y
a/XisQKxjPTFpaVLkIKJg+IJIz/ZHMfeGcszF2cDN6GR4trCFur2m6GNKCV6NU4uw9JNv3sbxw+P
t6pSiWVHOeQQPHNonEuKwipK81OfdtTcsId1LvarD60aGlgFK0gUwZy8bPEFQM29yupo25wLqvdk
d3i2K6ma3yxrgeSNdiIdSac/22jMcEpk2CJP8WlSehNzt4TKWo0/H25+OYjrGLZsqNxE9XPmZDXV
Z1bVS2+EKLKF3ZCIntMD7Od3deto1mL+WwEkWvzcriNtsjCDHRPdggtYutGEZVMocyZF3RM9zpZ3
GB4RRlC+Ip6zXcRt8nZ2otF8UBBt586RqoviAg6RqUjjA+QsjZgGZ9CivMER0MT3sWh9gHPOhOcR
0p6rWEnsoYv9BQX/PVl3jvPXEyXqBt8z6UM4vzuspRwQgMHTeyWQhKpHOc1aiss7dqQr6jl9Dxe1
0S1TaLJN2QlmG73DKn8LCO/silTg+VquQVj+CLwojogZjZdkPrnBh4MWDoTQwphLpAI2q6biUEAh
/RH2moSNWdUAIn8tkb7jrwAyyO5879GczEoGkbbQi+875Hqz+dNlv0f7TPmqCL4VIuuGlRaK89zl
npvKgnTqH4jeTkAoINgP3bWQQvaQCCUxJ0DD1RpfgigzdTl2g0+usNhMegPnp77scozHPGrecBdk
5xsEwfxe7T+zZXp6fOBdvVZkICqE06XGOU6fB62vbKIUY9iRGcXZvxe4SUE1AAIhem3hFg6hT6rJ
icapj3yndIsHbNOL+tJqeVJmb8ejjelVIfKtpwLZOl2AhajTAQrVX8Ae+3fqCe/KJpAGaWUMZTy+
cstwBfr5eNerr3zw3bvQ09Oh8beWvqWssFn8nKdcIfJHf+PJE8xzHqU4Uz24RGiVMVLWo/VWpDAH
xi/NMcaH5s6mjeoCKLGlYdT40ikGnHoZsqrVFDgK9a7/lrEgwhnnRcymc223wgor+xHZPi6u8Cov
kmvl0yp3uo9/j1M1BgbtAmcMyAblfCJwW2gs5FT6T1jbtG7oRoq7LXm+dZcVKeAn9A8cx0CvLOpD
2eNFACTtcihsBDZCAuZTCwsYfSS1YcrPuAZfUyf4pGyv6eTYYhgW4HIUFotL6nafGrpbntotOJZJ
sL5ZS4ZSZqfuVD86zS5c8PW15m89xB5QVvrQqo/e4UD4HZ9d62mTqHXjdaOlKm8UvSAoghOyyo0t
01thW2wMugTZjQQM8DygkcW1w2RPS1di0j772V6JzSeLBRMj74U/t/f4MCrf9rblPdWSug9u66jF
QJ62/T5jDY8XAU4NTW6bZ/0R83rTHSJrwLTS2N8XeEVuqYCZ8SGo3Bf2jqhCdT5uoF3ewqE9kXd8
MQdZbjGBsHhvinYjyFfDjhkG5ijLYp4wi+S0pNko+3q4tQfmOmhuF8HP72IQRfNgg+gx0aBOQGob
qRNE5pRg8uqxnAkekPko5jm8UAhZNVOhYbUIy0PZUybUw/PS5lxkBZZ8Ret6Ap/WULIUXdPpgWnF
7oIaLSx5oqQABC65JmXbHUrGjjCFSjMZtmIYUfZut4dMoBC8H+7RELN467th47HjlzuCKcBRyDV+
KoNt/z+bx7tDDUhL/l0ExrHckNj1SJT/nYEIhCp+qD8kMNKtxGmqrBf8XA18sRlifYgEdF++xSiR
0/USzQYG/fK6CsXsiOPtgr06cJ5p9KGdnpDRLSmXVNVa4C1JLrPnw/sfRLVBAQFXysRV0juGmuhd
W5oRwp3Ndj+wi5vW97xX5/vUFiuLtDqYslvQU+g16uFZXRAMcqcaWm82Hv0LfZaZ3JNMYGSVdEXa
vdSrY6xDvA/9Q657evxxSztWzdjZDvsTo/15k3D9iRa9eSJwm0fwaF+wKi9JESTVcsHJcuVWc8cI
/uVvViFVC/EYh13RcLRZ5cHIZjSw/BZM2uprACWqscJrCiGDlYmla8FdCQuWL3sf1i4PxRrC9RNX
xJLwsk9DLzcEEK0Z/1umkUM3wJ1MBrMK3XTXL41gwgqVlKGvNL7oa6txskDh2Mw7ZNJ4mBu75tmb
ZDvjD8qyHPoQchYF8PFuQJ3pxPqIwzJaRyUm/5gHweGP4n7/RjYVjmO1QJsU0XIAOubLWVJfHKWM
hb6ETm7NpTOnMmxKz+IW/8FiNkt5RFO5MzW05gIhvY31CkkYFhVua8kQYXuComiFaQVumMRn+3xr
INu8eBzP72XPhDkafh45eKGMQ0JsxcHmI2RZUgMifS9TPkxRfP3InGRZ/ZioZWz9EAhiBvV/tX8o
DvbzJzxt1f67UqvWtwi000qe4l2Z5+ARh6sL17EjPkCOtvM/hltR19swts7V71BeeS6ODMawz29x
lmd4JA5AVYWcNloNuE2EW80nnaxDPYScpyjvDIn2YMOw6UDDFwsR2ItqMCZBr0d5wv9dKXwBTO/Q
IeFCh7ky+YwI3y9YdYKKiAIODPTNF0vyv26aI4jwBTRoJglSzkc0mtSfG71O6kZ37y3yRr0zvpy0
wh+ZR2KvUpC25tgzl8e/QTTMuV6GCGL4zPV+abde/7Fr3TryHdsVwlno9/FyejoOmZHFFPTUeg86
HTCW/gYHztHcdFY8ziT1XFs8QFCrEi8sxCkRZO26Ws2d+vmhR7W13JykJKKKy44xZIz9rij3Ym9r
B543i6uxts+8gPknhciQuUra8kto+uuTv/D3m9ZaJN5OWCwPiRtqRILZN0qNOygyAppfBmGQUU41
p+BJl9+ceXBhR9USh/QJigLxazzZ37jmoTfi/gsigWLAMEE4WLfsqntB8ntLnoIkHMehEOsUucsq
6TzLv6+G5SmQvBSJXhV/biPA1IlbOMHqluHBhcIXn3Z176yodUwlmVlorLR5asQERYi5otiEnekC
BvDJBQB1WVKh/hWNrFkZxCLVDmZO1i32Kh1K4JdiNwSJP5vbrj6INHImxn5PRkcFxQ/qOwT607y8
LUGYUvz4N7Hvzkueu2Tj1mUDiswPUH1ArbRfN4IBQWPuMgcRz5hoAdqQPsvmn/SRNAYIV/OcKQvp
FYDUN5gc2/Q358wHPxAKBJSkIZ0TYdVMFfhdhgGt/8pecyPG/5LVqesN2z0wlR2M87pn94eyIc22
NuKv9byHYjJuog1AjNtZD31xA+lUUj+kUKdrSNoCgjkRkRFdxW7w/qmzZ6Gi/p6qotP0+zZFi+hn
8vLMxCMH6K7MDvbIvmas1GqhB8HnRFy20MX48zOzxmiDADdzu86JWFHGgPWPolwQv6DKDBRPZtSp
T+enydgBQgg+3lI0JlAXfycF8zHQsFdS3td/bqIAJCHr3wHGGWXDyf3USmbYvhvOtU9bd8PbhGPt
C2ZN70b5bJtw49XRwpQA+TcVDQ7JfwjqYSnYOcLg39lJaDj6voLAkFMm65U2wTti/o4gmCBTFBZw
dzv2CJPWX5JDt7XD63Ff+RyuGdnkMMF6TO+Z003ut+IUdgk5hwUCBliJlHgTzzNHhy5s3DV0iIF6
P4jN8j6saH32+uSlTrMSwygHDlrYNw7PGi38HNDurZEcCkYuZMzZOZVSdkah0VYPTYrj9J0f6z5X
JQdkNJzNZO77RTpPfZxfbSmjFQ55xOa5hy6vWbxbCFoqFBl/IF2W+fIiY+A/cWG1pgNR0duu7rL8
QBSJedpHfE8FeUfDkcv71ljnB/JOW3grG32RC9qZZtL+NtO63flxUcqc2NOXDQleKmuquKwS9QP+
NPyEyl4vf/xTyXAKOgNP6eWYPmCJOUoA9QWhm0lmJMfiUL7IXn89HZ67yEUSOfPrvqiDLpZrTLpY
Ue3/PYbb2FxDZwVsmXOtRU3/C+oFECP2049qXbrd4UtcUO36CAYBBIfBUOZlLG70eqH/qXHvxBaa
pXOsa4UCOs1E2C0x6QE/hxv59MJSVTn/h7ZVVqp706N7vl0Pe+yu8GCptLd5oPw2VlIHjxV9yPOY
6+rLmp2kautpSX5708tRy9PO7+jY30OElP0imcvBBahksa8ymaffAGYhXvmxVJQKtHHW91XWJHfm
KCvcSNSpzllebKpyYUtK7wthTEKf0JoZbPm1rLudP64qTonKpryIzS9qfMgbyntkmSG2oejs7qxZ
JRngVtZTihywXFg3vqWp7MUFk63KSgBVBI7jusGDfF+96TNKD+3WDLBfRC7pF+1JtV1d459YMKHV
8jX/Ko9SFpCcKco9wcN2TCsW+j9+eILvE4zhWC4cGkPDdWedvxHdwjXUocNdvnXRJ2tT+ke4q2m/
auvFOtHP9HCeRsbYMOOeR69UTP95epoPy+m7cFQfJRIiOP1GOabug1tyuwCOLK50DCC1oeBoPpD2
4FjY8JDVqbeEUWdrQYZOT26roitmXXDf0I39xjetjGkpNlGA6Xvk7Qwy8C/CIo+gvUVo+dFnDIbr
7PcNiyxYN0+RvIgD/n++9QV4P3t+tueeFWyE2/MjC07kxdhYVb/IDBoHAVdWAtoIC8zcpekYE5u2
XnAH9+ucc4pEi0C6Z2DaTsHEUQ547BcDtG93yT+Q/l/1kvZy0+47VopOr2WvpwWRwDn/lfrCxFM/
dJ5o82D2y08M8bHJuUVUrY8Pyg1Po/1sPM4uJEhCFS7hJoDbTIXjKMbBUUMDRu5zVWNeuzbQG5uX
AfZdakU1H8rjZ5ZdfM7casZ3Oj0fRdphHi4jAcaS21+yoYTiPMIAwXf6VzAiuzwEuEmgZCJEXav5
nkI0TkZm0oWbXXO1ibBnx849WEQk/DppnJLtkg3vZMkZjVUOaZxdHrEoGg8N6YZvZQhmGIDcTXOk
LxoYz4T6AgWTAS4LMRQs82UbKMbwmGOC3rmLetilX6XmN3KRyJthRl3HDmwkX8RRruxFg6C7/pDy
KcxScHSw9cuPUNc1xNYW4WO8yU80kYMinf8r17k1cNrGpsPf0vdUQdYw1avchCCXTprVdJXDaWXe
U0Xeq3w4h7MZndhQWZxHql5ffIYaROOIiA5PBp7mqXLsEan+BuRFeQ+JawChb4TAqTKZJV6WZW0z
au7jHGBYXe0VBGPZdltihJDs9+LYJiSiud/2P79c82LQi6zSv5L+GQBkHKHexkJm5DTacLoPI5En
9BHEBkjN7Pspxg0DG7086m+JrBe0WGojJ0ol2NOZWUtN1tBsp8CU0ckVGkuYX3t4qwoT4mCdInI+
RrAj1YSdZajBIUO7LRC4B/f3AtZkcGj5tdLiVM7f6KnhsP4xNg+I0yJ0wBSpug9KEu9GNLBDBO8r
E0MO0Lhw9znlFTBSJeC/mwhe1GHbb31k2Y16AjRgNWZLKr9UDUdibheTnyk91fu0mufzIweq1L19
pqY4aCBkmFNFqkAWRGdHosnrD+85/B1Wae0Hs3r/Voe2fgcRq5LfrztnjXPbsZvc+fItFtkxoelN
hRHcd1/W61RTbALcZZKOFkvcgVAq5FYVWGa+VszdCh6U1+uucP8SJGNx0znDLQKeQp30KPTd+krh
PvwvQHHaFz06uD3ea9fQCErJJVHN+qfuL+b+CTvaKO9F+hCP2gUFGoLpb7twG59iVX3rOZ5aTjjn
mEsxQdZws98neZCUSMJ7SEFmTmXF/WQ9vw/AM12Y9qvcGk0hjSzRw4B8G6tRHQlB+iXiAoArImaK
5x+ZpA96Xdf8O+oi390kKC77kUoFbGXjdGNvUyXewgf+JgeAn/bv2u0/GzYz1q1/KKY54D5Epang
KTQh3gKebcHLZU6g3P2SaR4+rT3FcrRb7DWTm4QaHER0SAoXxeD/w5wdNQEVd1d9yrsUXgy7zUR0
rhSVw1Lhn1HLNVmlm9SFDr7TEZZcn/k7dMdTSloXfteWYzSp8d1/KlDNsV6s3kooWnqPp2tz0nMw
sgQHg+15O/UQ1nd6EfIVrP/+biEMiZNxW2Thw/6bjW5wBoWMz7J9te9V5cyvHpaWNfCC9rS1d91p
4GlX08DiLa5sV4SWUnwSi6ijAGUdAPjhjLJ9syQHAExhaztozQDZ772UyiDL7UNfftqJuUwOEzsp
XZa8EHwCCgJe2WXcCKJe5oJQUunL27CQFMKMe9RX14PJNZLwmbVdUo9+7iqxF6mN3bkNbv/N1yhH
fB5O401ank02Mf2AlOiuNJYlLMUy6nTBcThwWJ58+AbPPS1pjt8ONMYOkscmK9SUW39ldd6wkf4A
qv0i4hYjFPebcpNt00xRhrHm+kg5nT+ULk1TFaOD5s1KXDfnqOWA+KX2bV/M4lLlhXI7CsjEYsYN
oRV02IN6s1ogaT5pUFwjCWd44xV6xXP8In1O+g8heOLKS4Mea1BAbgUForO3QqsghuTPVuY4u7vd
EcfatEX1avIiEk2tzCk4fmTQ6Tl5Sbba25i0A81u8ZnNycv+5hGVFHB7zOvXq1xUnp4Lu+XLa0Dz
EdxnRpufLp2G4nMsAH21lhp2/d9A6MwDUXCT2PY6Dh+eBT9bcwOcnNtWRam978vogJBux7Ah1iLH
GNfRz1Kaz/1wCFjOMfv3RbtA5LMHkzyOv9nHDuY+sCWW4V1vFC41pdxX8UsP+7lus4ZaZy0qlHCj
WMHrotqby2QkKVOvZ8dFppb1g/SrItJadFNPTmOeTk5BwLFA1KrGtwsNUJw4a4sHL9ebNcCx+ZHo
1REtGA6IGBh6SytWja6xjY9vD5hwSIyqqNPjjXGDwGOkdHq72KcT3GjwIHBx7sJuO15Qhy6KSHQC
YBE05t1HGjTo6hPyFOruvTcI+DA1lxSaaN7UAv9MMG23h5wufVFFlwaWAcYThMUueq1DPNx5h9s1
OrrNfj4SeNBKF2HrDKq5P66J4csJaNJaqms/fn6HtOjAPs+a86KA0aGfAQZgUu3NZO4+S+As9b3g
mF9v9gah0Hq8i+40e964u0lLrr1qlYjJSva9Jk6uPWB8cDeBZe89VlSDwMgRm7CNS/CPrMVddhg/
OEd0KGUsjxWoYBMtVlJvTJkI8sra8vmk7HA0xD7d+27lwIrYJX0ir318QhSeexcCnBt1JRh2QRDE
Knr+lrpfYC61EbwpVrfPtDkOhgrN8jNrKUeP3a6vSKD69pITL44bJRfaYOgPHMj+SE3Zz5oppQs1
BlhnAJPvCEwhPPXTeqMKaAOnVnIYdSNvT3Z/gD1kXwAyPpnVQMN5SNVvJJo36HaqRTSlof6ZfeMb
ebXjhLy5JzyiMZGFYLT1GNfp6oVhQ1IQmTg4gX9If644JhAoDhPk0lPiLHf8dsLDLl0rO8TjVxBg
U9GV1Q+HCl4s9GlDk9rTEimYiya5FTBhO/W2Arzk6VqiDY5zuUcL5xoiOJ0o2qFGw/uG8Wepuv/P
guk9Jy5lHu/vO6RxO0ivR2qmk4OHYCg8x6LaKkfo23szkBgStaq3jBER2571cv0yjmN8kURN3tv5
0GlCSik1uyxq6dgugzcPJzZJMsjAiXyJqermjCfQg/p65D4AvwHkLTIW8r2aBW6KCYQayL9untpZ
1oBu/bCM1ETUnqKrRXXIPrM+24aoOkW9rh9mVKpce9QZPh3Vw0DQ8LELR1tGn5ZzHVQRSGj4CI9a
Kx70o+qCXawSq/7jYTLcOMIRXwq/euxgr8/C+gi5ADHr+IQDy4BXpR8eo21uu6CIgiRsXpaJitEH
YqSMMawk2U1k7DXWkfrGkrWSXSTCoCzY+Vd608BLOPuyjhfJ7/NqlCYLgd0gSQKSSHnAOaRgSUrc
eH+PhrkgQ8kRQGdI9hSlX7bMBCWTCFSZTeFRPZd7UoLtYha7erHi1jxFFddpBF3lKISBbycOV2tP
zei8dPmhf1AUB0LmcaBeHkviucvIgB7fwahKG/PYNPpPPH3CzhGBKs4Dk0FsPA0tVGgHMQxYBt06
LoXUUX+m8SKorrzeKTxS1K6okjgFGx6PWnTC4SqK9XYoC4HXf9vRwXuwe1XIaGD8FwNbjaHwBVXR
puk17QaAz2fLvuwmeF0DrKrcr+pn3qaFy0GLiVgAniQ9rkzIp9Sml/kQmSZnB1JWEKNTdwFRjB+1
7fvi9BuWaAUIn1E/JQpAwbie6kWGyG6WSXfl5E6+ankkhf/vr+iBS8jcbHhKsSMeDXaQhEZDQXW2
7yjYMPYEDknJlR6KnvBPdqwUEYFECWLqlfEex3ot3+/vMymMq/K62xxsY/JHmqjqsxRFHjbGapE1
OmtvzTS9L8P+07F/dY3LlgYeMHyKvimLLZP4nfE+T7UUsqiqUD5tEpMBig6NGXPhfGlB/lZjjGN8
LOmnIB56SwETChf87XMNPcwrJg1CLV43kCbSBcZAtbZR/BBzyhkYLhLp6otuIKKvJG+fRcFzaeYv
iXAmt6p+yYhVx7jUPxrk8BC53Ek/DWZxsqBg8sz+Vhiz6YpEL5bMy/rSIeL0H/X8iirbEG7wUHIQ
N+uMpAVIS1GyE475eL2kgXv6aLs2g3c7ij2S4DCBAeRARF3MgdyaMYBUpxWuDchd7e+okek1d7Q1
3M8DcKVH+qaJP2YMzbp+7Va8Jm148uAoKD5b78rMBIMpnxjEomAo/+G2W0DhugeMsHOeVs+JZttm
h86OXv3rZSuQd32bDP2hUUiTefufrqd1U8/GnQ/hBMjkES31D8S2N4RgkrIpuKTEO45gI/PSm3/0
nUpFM7Tkt0qADo07fVOZGLuLIVB+SrxFBxpbRxsPwBsTFssO6cy2duW4P3DyIBlq3Lzx0+3sVmRm
3vxf3WT4x1ixqtsyTzuRtg1r+SjAEK88lRZfjt95LCzsU0YIOQTe0mXzrNd/snajtayVT+xZXOSc
ioEOYsd2oxCw3meVk5eFGUJ3DaDBu753mD7uwIGvrhW+AjuuXi8HZJa6YXGQO83zJpeuArfYAJ65
1CXMd1nO/mwxK+v9wpI3Pd8lQoUbTOumi6VGc6HF2KnKC6qdgd68QIl7aty+LDGwfQ2FCUUto4Br
Dgbz2o9B3QJbmcs0j6Xi66bQUJSgvuoAtkeeuDdLgcPTWxrcJuBYWcboyNqqx3bKHVwZgm5cqef2
aQfYL9RtHDxW9WX5bb/6hHHTf4Ab4VuhqU+G6SztCv5shjBkb0WwQHtGbeMp0tCvOXfTOF9f8Q70
alSHQSsGFja8j9siF2m20Br+WhgdbLttA+2pivQVusWFOuAasK8YuiShH0v/bYlWIgAMBOW0DEMN
xUAf5HL3RW1llZHjTAZiq4TxEza164LUMboXxP6xGcuZCOZyKffVYAsC9ChyMEeB7khFAjp6rJfW
WXIAhfRPl0Y97PzqaViZiToCH3Z1XJ1zQB0A31KnxA0BA97HEuCvsE+Vsan15ru4+vAfCbjoXZ9L
4IzqdLs5wb+Tyb0m5QCHLlg7mieiog37it8stH2FihXgUvmBbLyq+ZtDHKgZ//aI3TzWJquTv/JC
cUFpV//IZ2ReavAmLjd8sVhmA9+RypsmdDMYSAYXuV9Z/u8sKGQ0Se6UH8zsOBak0WT4eTxoFw58
wa3RJGBVnP7B2KvDC1iQvuuu9O6RUXgVJcpThxX4WOX8WgezozBfN/OS5Ux2EYO3WHo9rL7XJJth
kJXSctdP2TlY1g4vOkTLEwtJAnnpghOdx3RgrzSRWojZnt5/+SAuAAtMvv84g/1ceRMMVTIdhhFn
jyzHzNWde9hPiSdOTNhf1mohOc7XEn3PuiMn/80XUWUExB3Y/nSkxIZ/BrO2wN4c+p9FBhDUfZKf
6zR1RbNPTCIcDEvpVtGF5Gefo9DvXfAyA3OZetsF+eigGqYhj504LG5m3awcdkGlLccj0X+gvjRm
wElSSvNkUVMxkLhlPpCnTgXZfg0EpW+mx2xAMb5f1evx0PYLfEXXMLWcAf+a/p9IF4TsIflS/l9D
YyOZLVCS/Oj/eNsAFNV9nvIQ7/4YZjt9RQCz/a05+v/T/6WFHOCaroa9l0peirJCf0lJq/Fatnw6
Ck0vepTRx1WTGq2K0E6riztpLJaPrICARs7wmoFFhe22WUOm43OFPu63p9TurIKrrhosyQwMARfQ
UwWcIdN4qwoCQ/NAwnHe5Ts8+yDTF3O4PnhuLHzVrgbOOseCLJSJ0TOiuNY1MdfaQIXxniPWf1MZ
12C1qpMeIvrvvvbTfrbQQ2M42JWr/la4yQW4f6e3lb8l49TJIlcXiFknSfjR2zb2cY9TY5MmaHDo
abO+3McZWHQDa3uup7yPmtILMjBSiH+aGkitCIxUoMhGkHRrPSM2ifEoY2+7mWtgHW0owXxLUsea
lGgIhjEjvpLRCJOshCt0wP64iNh9r+uxzwbTYbMxRy5YJFQs5vfbgCi/ip1sChVap0h1D5PC4Qia
VaFIPqL2WZwito+ENaLJKkqLa4ZKs7lP7H3OFwqlobqQJ8I5Hvhm0ZK6VdBs6UcAjL7dsCyZtBUI
H1Q3YsZuuH1EK9iXh30v9a8qK0Hlm6SQtY3No6DWJIZz3OvZX3L7yHlKnFsdFr88SI/1Q2cj7Rum
9EpQfpt5/cPXwDo218IfcogqLQJF1Sy/5CHllZDcb8gdqXL+Ya2sEtUOThl26Hhi6qTJS+JHWHK9
92MR3apIlTOdQPbrAyUhfqOgtW5xdJTEjlhwHhPn6X43dFTHmGvulwADwmA+Y3QDGXGNS1TPQ2k6
GWRNcUQjLUSuW/dYkAr3Lb5X+R37SPxpuJG/n+YwN6B0GEln7RKeSCT/VAbM99/FLm7ytT65nMYc
vNgcwY6jp3Qg57hNqOIxVqL5ClHtMGC/w2RL9OHLotGLheMk092RpnsVhKWyfuH5NTu6c5umtvmv
kgMvrC+v5Q7ADOVKshnc0m1/RHxysdF//5R9LFfGCuK4YDB0pelNqqfWrj75zfGSV+8pxwPDn30a
ff/eDVbXZODi0u/kYQAkrf839orCxUvSMqvNa3Wtf/ol0s3ecDVU9/RNN5tXxLqm793dMHiBLVTl
ItTRRON64Q+ooLUAE74xHIB8KkzBn3IM21IIX66iVZU42fazA7OsDOo8GB9m2jSk4sdj+yEzD4rp
dzQRooy6Gk9Zfu3PZ7tus1CN9po40UgHvGHnpMDBH8LUS6KXkM/K+GyQuoNFAODXb+i/mY7Bg6Br
byb/fd9qg3iNZtKCah3ABQSz9Uopd2p7ntsoFg1Bmq85dk3TxPW+QT+IfboTlk5Q34ujySbUxU7u
sVC3hROb1vNArBUfVJxs59wZZgcHArL1miJeVvkDgvYY3HjyrYCYWzQxSXEllflKVdsSKZIMp4FE
JkUilmiwHrj8tSkw2WbOvojeptsc8GcIgZRxmaimEFJ4K0tFb68vFVCn5q/zsW424r3+aQVygg8/
D4VM18ZAQKID4HI4K71DWWVG2d2hv2ZEQ3JzsFegoK/C/n9pGR9VarxnpaG4aWcwjYKiyy9HduVM
0mHOOCpy3wNVVU2nxSXEj7Ma8YtWu0YtDTAgGfIxR8UwObsirl3+cF53d0mD/q1cSF/yG9ac1UgV
YR6SP93kwwuzajjPZrB740fjz8239ZdcDCywiOmYR6vLH1HfV7dPQK/LIvuggYNJ1MfbqqUzbk2W
OhWAHgvDpWdAmVw+QDlJv1jJ9s4hZKSmUipyex9sxtkC7ZIlqhuizX2bnEBItQYt3yd2EK3mxhcm
CXE5p3lVL/5ka5pfhmpycHnJRsLVGDoKNJ3BH/d7Qik8r04GfI867a9zpOQFUNil0a6E0rZksLle
lxiBSQRj7X3OVHkCPY+hNWPzACKc+ksJpCkxxhMX/uLlq84LoS4JCBNIr7JSs1VB8kh0tRch8KVa
Vk4UlMv+JM0oMCNV/I1giMV50JUcY0mUXqjBe16IAGmmGpR09EPcBt1eASvCpE1z7AJwO7kO/F06
AxW3Zd5tbRUVBGf+Ti8eHlHHQopZPqYLx4/Fzs6NLSP7TpsCylcUm1mQADYyai/Qq6sOG5jMURAk
W7ty5UvrDnDeHgz3eiptNL0ofFJSkX0VKDww9wdv01AN1DsFW7zEOIuvlyVSZZkhuTJ/iDXoynwQ
Fb537jJovumryhzMOlh8BC498eGU87lpApRU1A7MvQb+Hv0a/Bkq2QWWyWXf6psTvqleSxz4MlWg
2wnBJGn4oWwWK7EAtU7pzZGwCBHHm8mGSUGS2qWIlOKCEJJMtc63+n8AAN7FHZ0MtPsh90jhaJ0R
5BC58LLG941JD0+8p63sUi8CnLGFXfBZil3HvzYRRBz/cToGL4bJoO1w3tjq+HY4WHKpn1VsVHxr
su6F0Uwam16i4vMnAtxHvPTZdq3trvJRpPeU8X6j+W86niUOfEY2nSGwbqxYG470n1CUl4+Ei31Z
efH0mjzaORICqq/AD9hnYnDJJ67saq3L/wmpJCrQlg0HfQD54h3OiWyt19paj5IeYN3AXs41GD3I
VDWZGKyjNaKeNvIBQQU8h6i7wSVhp8G71v7XlWTIgPOuDEyzSjxZ2j9gEiNKSa4jcRiHrugUKDzV
GTAzYRHkgu5pOwjprhXA8DnokE4cBD3ugIi8V9MwyV31dOoCsQ76A7iCJPZ8qoZ0pl0afkHorlth
NDXREQIW37zrS8UF9p6T4Y1YYYrnUmtmgvKwQv/RczI+29fJMEy02CDpg/AFU5fWj+/7ZFkBXW1t
Y3EOymuAYS6+H+NOf+ksiQHlKbn6pluBC3R+R5kkpAM3s67t3l1ABAg5mX+EJfsx2tikRbsSPdeZ
BX7IVcHfJucbqoaflnpoKwIbrxpo14NH+GHg/peYjYUiVJ/vq0b2EDIJvBnhiS57zDRbVASpQPii
Owrft6FPs3XHOwAnu09plcckw4hgTq81hYp+O9kt5tM3PYYJfKcYYsX32oXv/UXEgaKiB7YECVDc
uhRbpe6fC755dtcbw3fopYZN7ydPAZavCUB+D2+oFWaa7grNFG2pfffxhcKP9w9TevHi8Y3h94L7
TLIowLK3ojC2AwhR0LzEQNU9b+151o+fTjkVlp0CGoimG+4uZ0twkcVk0jXHaorjWovsoAghTIkG
wSNmXu/8HDPizA8WyapfdotHo2yiDjBCTl7BIcWUFCoRCLtolYkdl4KAEEwad9HfxvYLi8jqvgeE
IWGB8yGvqU56yD78VbJjxDE9JLP8+bcs6b7AiYwPZbP5p79n+z5ojMFVDrE+gwpi4HZkIloYwGVd
XFd6DiKJtU1hhim7Wfj1h2gTRMHWm17pjMgwMgurixqCmnPenAVSgvIfJ7+XdJX1V7PNpOUKQq8e
3jPLB05blHMmJu6F7R3DcffSWgeEkG/oUl8//KC8a0YKfKftKoyqqKg8j3gw3fic72h1DVLwpenB
KSEKwaGKAU5zeihDggTNaIfkMPebpKHJqPsOpEaz27vdNpkOLxtV5v/LpFnJoFSfos+Nu9RhiUCx
z6Tbeq9vi2XuxbnQS1rQ+PVEYgEETY4CMZY+SURCfxMDAtfZ1Cxm3+081Gte3D77V9eLJ5kznO4j
nNkJZFDla3jwxprzDcumsuIRzbkkzlynHa8U038rFGD/f1A343QMVUnGTCyCyFdAhtz5hrHE6zzS
BAUoKEHdJ4GphFVFJn72vapXin6gQXcHVR/PzgoCumqFfAIUwQbk5zo3WeK+d2nijHii0pgoFBBL
wSLtMH5VwMnfEy6Ebqz/H+/QWqSTfC/XVeDmIsnyUJ1Q+DZOTlk8JoEM/nH+VKgxe3PU28X8YR/q
Kc8Ie6HODDncir/Grme2mD5QKxkv+ToEXAnRIHYqKTK9vBPX85M/8YDnatrsy2VaPtAKwpEYCTF0
AVOO6BaCnWmaLhptbYQ9IeYbe2APpW5k9P9kakUY62dZh71MCV6d/jm3DtFYvh1X2T37qfEnTsv4
bGyD5+tA/ewtReB/7RTxMqXMPS3DDqRQDi6il1l3q/UiNPsvFfLcByk0NZD01yDN7da9wBAtpq2O
Yh2QpeF4oas9fU2qaOV1D3YFPjLPo2s/41K06GihwtegIrGdQU/81lr/G3tguS4tI35Jzl16iNWW
51S0Yai0KyS2arFWLB0xdIjQeHPFaKnKK8CybwTIMSKLwspMkmFTx1AvRkqaLovnAYP99bra8SS1
IqcUk001qgh6FEpHDMqGwtQcc+ctUrndZGqEXDn3WtWAAC1bSTQ9PcmuGXxpkxXeQcaMPE93dHbj
TIoJ7R9eJskl5yPm/JPi+bNOUz1E0KN80NY6Gd1v3b0RMwFkoZB8VIR2vazziSwZg6EQF3dk/H+P
T0XU/EnaMCYnRSw8Fr6/MHhmyEBOJbv5RWvbQrfsggcQvsCuQmTfpzzPUZMSoi78IjRQ189llZqb
onK82KEQKaakS9NlUQBPbo5jrsiQ5rdoRhoNqb8/o5EzwL7WFsyq3S5sabFxSwqw9L87pgnmX7RV
vSgv/b1hlxqHZRkSLOh9L3V+yFPdW3lxVLkCTGcV6aqRdIJ1IPwnsi9w4uWDqjsO5uPdYSbK+H+x
hCpjCrAtcaE5ZRXfp/lR1wThk7xvGUt+/i1yyKwb2eTmeF8g+ZkfVyPaG52tUNr+b/M6uQjhBwUn
ddtz9OnXJeK370SyjHHErA/dSCHCWk4kYhFnambPUajvHTTIaQdLMdPkfQeC3DknZDrSyKLH6Mf3
IE9gxgQ/GNpX6ySjnaAeOjLjsfPD3vMqQxC6KCHqA/EungEV/Xnq9TJYPBe0zK1shP5iWbSTy/q5
of1Ky2p50z3dxbL9M/91yfDKe6C+hrg3RaGBS8K8xLLIjxSTZzXVOifWwJpOccAsfk4z48uInbrC
C57Gi42Z1MO6bX2zJgx1vJA7jfqdYWdaTjsiQ1hOPF9MDyc1Rk9boG8quhZ8orT+uTPvT4R5CXow
B4tzEM9VAP9iCdvosceZ/it/eRCVvd8Dg9wMgrh2f9I06SqE9Db6lkEBEbW8EMkv3U6bREYudxXx
yY0uyHtTKE8H0qKl/nO4B4eCg9v7xD78AYbtu5LY39JRh+bEW/SRjfMny/1SKlOBRd9V8eXqjB8G
wE6NN2BpfOHVTXrZoGd0LX5qiKPXV5Dfr37sfJw/yD7f84G4h//e9J+e4RLI3cjZ88gMs1HlGDII
+wOvq1/ofmosYcFqmdqXeuyREnuaiRjnAlxn95MjkvTv/KezCa1/6FKFmX41vUzhD+3gFJtaJous
7dgoMw1Z8MJ2Xyf9g6DkWZKBHwGUsoY8lTZYLXLi/E/ZY55ZpXJ+ggRGN/X0czmg60z/X5Zuy73c
fFLSuOnyEK35LLWlmBj+Au9XdDsORRqoZRpGWBT4IUbqZrtu9o3sQ7yEDB4D1fo1Le8nwIA7TEHO
8UAX1E4Pvnu37hW+FSnrPOfB4c+6UAMTd7sjKNAq08OP0AJ2yztAvEwNWONynnVRtqBfTavtUbAI
MCDmSNSb6XzI56+k9CUlrUmyTWyy+E3rKLQ5EqHYKqW9fXCaiLGdW7WZ46JIKt/3tVPaGm9VaWF3
C3yzUzkHQ7ElnB5SEHnuHis0WUlHnzJso0VuqKe6cqfZY5a/dxNimrcZTS2vT0ZSryUQwtvu9+ub
Xm7s3YTYMXRFr0osp7YaoKaQFqpSNW+bIHOtt/cs9Kh0I0f8ufFHKYfqQtsMSE2k75lvGgT71eSF
hg4+hnOQsXmdn3jWJ6XFijl/L0y7/2b0RqKflpJzMN+HODv0IybY1ceOJ9vhQBBc6/vQEf0XtWKS
937LItoqgMeOcksXJnsLVfFr/ge4yH+ITjMq0BggpSJIGR8rtGYomtia+qIgvqtlg61t8gWSTvEI
X7ui7gDie/c9iQBstxAD7GQYFV4FHCL1kdizblU8clPPoObOqx9i9LddAdkR/q83L8eRj+R/4FoM
emK+sdXWitizWweUcW3jikvJwR9ZlEMQsz14fhkB4lWXjCyB1JZliPRcVU48AlFP6jVIMwlHeUo4
8i4Q5v2VAMI/Uh0tW6/OSWwnoWC8efeVynVFwRjLmSCjaFgeZcofI8xBBtC9UaDWLMHV62VKLkVw
kpklb/xHCXHCfZOQV281aSW0nhNwDS0j1IthAgvzmfDnVaRd0/2IFP9+UeSxm1djm1YRJ5DO/ptp
DiE8/s2yKtfFxFWl0M5mqG4PMHZ2X5IKIX3JtTBc0RBUgwfzxxTf7jmsH5i/qXTz3nkhVTcnwno3
9Ze27x+BzWHcK7URTjsSFTyjLkdgSFDGMISAwmYEwRt3hOmUilaQgWhafRat+PkD6uKYxaxbWfSV
/Nz5WGLiuSShNxVCH/aNddwSJLsss1b8VTAy5OWiAF24cKfDXfTpYD9UI4nvBzisEFIyYEY5xuw2
Ojf8CvkYg4a7Ikj7KHCGSvlaMtcpRcgz2vq8tA/lcvvW4AOlg+M9I2fRkvZuXqU0W0I1xXTzaoxc
20UeWAX1hIVyLyHQStk+omozc6uLknftzPzV4EV5xkYsX31x2/eKS/uQ3IPoNj1UHUAQqIMcM6m8
fCwojvOiQZV1jN6L+px9/XMP0N4dYX/EYyeKNFGwl1bxzJh9Iq6EGNp3mjT9RVWGsOpp5Zz2eNaC
WfOT2KjvPIt+489cSX8V1pCCz2Tp0NCz/sK4GHauGIKLpQUlMAk9aXu4E57Eje+CZw7NQH4bkxtz
dTtvqNeY5lzT7XZ3TQaJHpjayTgUxnlH63JfBUMMdwRkSijEM7WQC7+JdVq4kAA0qyvuQAWAN6gr
QLtT0Qn4PibY/2qL1NuzSah7zeO9CKuzPkvquELQ9HwpwOUJ7PrjdNmNgyhJdoY9AZ01nbRJ+G+0
9r+o9F8nqaeIHjvqodlyQrX0D8VSYXm6hjzYgjpNyYXjj9UYQFjgvoUoDkU7J1W/GWTYD7lwskY6
o1a9cBPWh6bpHtCBTPqN90Y6KbExbXi4vHFBxW3+kuwJ6qfJo7WMcLslJFRdikT6weI+ombtB4C1
fVv0EDQKaHOhIyAmihX1ESf/pldgPKYtKTi9a1xcc/qkzjFGyZf0zwYIsRh/02C29GEknjymNI8T
9AsJ7iBKxDJO/2efKHsgn3gT7zLHzaaz66sTgh7DuxWbIP/bfUD1a8tDPneXXjFIpbqVu3uyalEI
s/0S1Fi2yY+41KZxx+Qa0UG31BQgJgNFSKO5Psm6j99+qoIFWVcXV9uob4VXjtDKqv26UU/dra2s
dbrKhgAgkYYVR9u/zNcxV2MGoTofMC0SRK/bLOZrNznpUZn7SAdtRJr6N9psw6zl485N1Lw3NNvj
ilzQw4b6lrHkGMtQE9l65cohc5FYe9db/g01270yraIqcfNaqJJCX2TjPq58T3DU7htVOZiCbOXw
/JyfIi79TPfma4t0PLgQX6A4yvISdZbcrn2YehJ6OWjDgdzu3wVG5liq9t3fc6BarMnXruuw+b4H
WUFvpNfc3mK44mqpyjSUUsK2U0Q99eBen5m/5LWIHfnFPF3b3idQSwwVMQ31SWlBoV0TsN2oCs4u
JZOG0UEoJJ1gbfx5eiB2lhYa/gqdJYiUTvx0UZcwWysZQNCMr9h+C81w2b3rxnOCdqkeemwLnwk0
gU8yYcNr8HiZz0/O9BPGyJ13amZ0/K0Mp8mgLLx9Q68rXKd/4DbJf4NMj5FTNq+DyYwg4MIWLAKQ
Tn1kCn72rCywR4zQ54X6KCY0H/JCv9Iy2PE02XkWYFB8/GKd/g0VURYcgBh2CvRVYS0gzgeSh1Xx
kjkSKZMTpn/7c0Voj8+gIv6IAkBWgNZ0lWjPtoDsASiuWS1rfSzma6tpSq+/PM5BwSvxUIHN+9iD
6knk4GT1x2IjXywZtPrzjcOYQlLFK9pHvgLfaKnxNkOf/A3KCR5KvmAz59xKw8WTtun+F5cHIyPF
Zcdy+We9rmf65CNgSG/fjAH+OhZ957HpsNJD3DqvICyDXGi1Uz+uPRlgMNko0R0mtdcHR570292C
jr4DP4CFuBr53cYXlRnmEYO2fIHjl2qE7nkA5J28tVxiahV1KwpbJs1H61MXE69dJO0gDJx+uuUu
EOS8zuwSm/Hud90ZEH74j/4CEiDspLKQwKirZhTOAn55EqnJWCfuWEoUN69pes6yGj0vDMO09t/Y
4A+OvA5vYU5m5tAoQ/oEoP9IvtyTfA3EE3359cB+enY28P6NEu74rMK6hcU2vcMULNyh3erh6U5+
rnOXRSchChg7lcfNhdJMGbvCnYM0NmlMVTOmvSKEjvRh4gzjYuRTqF4fqrGKE0CezqEfLadw9vyP
5etdpV16dGpl5azBa7/5kEQHmEsBqmuUe1yxlxnxaSYvN/gL1oTYX9Zf6vF2D7v2n3M0S6fLIFJJ
zxV4xGAn0w8AzdH8S0u2oXirptNHnV5ULej5/S6NSIOL9kaqurcmrDMCeTlVvaa8x2FIwsdAT7Tm
r8TjDDXdE4n+rh5hQ8mayHotwQfnFLPUIW2pHFlfTVocRe3o7JpwcqZ4hk58OOVD7cDzWqe0N9yy
KGLR/b8PkjpafeY8vYF1UP9ND5wfvfkQpyLyaBchR0IBdXIB2SBgCwj3kMFoIPOTR4yyWmH4m/7V
6crGrVCPYDzu1YJc2RFUrOGtkt8vzWNSqCE+YzA5xcAf5pe6nz3nwA7dcAavbn9LvHlJtbAjvL1G
TxHWCy1cd7rtS45i9XiXjTFRCtqOdBRTVX3mZwgDYqZbGSl2P+2MFj/V17krMv+JRhENGU4e0590
cx0SVRiGks96KHTgmiXrzM+GTMPyx9XdSE2MsMv2kkpozJUnv93OtUUfSsAqaDJ05loS6ZkVKr6a
lldf6bqcx3pbIhTIEcb4ZLevkMf+NUIlMDYo0eDAPvS45qpwuoK0WnMItov+Op16UozCt4H738Wf
Ndghuo2umQio4UBRroJBnyxwL1IqAwGSHxMmFW2b1k8CmorX7N+ThEpJ7R+ajH+UfZ/AizCYtBay
4hbvJlviCz9qUpco/PVy9V++XKldl6Rwq1WOVb8JbywVHlkJf4Uonv4yoaiZVFnscst5SNXcn9yz
1SNUDzukyu+j0qUs7wAQ0GfWk8pRKpQwkbcfKbKJzQacPdhEngMcO3mLtbdvamq9SqFoylA3oNc6
htq0nmdIHaJCrGbTdjVw33K0HYPWQOCT2Jk7whX3wJWzJLhjyNf0rwQfWJHk5WP9Kw9y0Kj49i2I
2cMfLs7Lgz4WCsE9e1EMKFN7EOBX1mo/DxGGY7/k1FokdwJokcfPy37OwsVHrGrr+6YXZueeoOtB
lHWBzw3JM0nuJh131PapXPBMTY63PM/UCR7nkoiZVblJV3t4d2RskYFs2Fgwaat6s8eREDH6YSuo
lAMvL7wx15Z2kChBQWY1a57xm9buXFqWFGzhErWRmrYQqX2bivGMynAMz/awK1GbIa7iwfu7641Y
yH/iRE9dFt/gWzU4k8VPqhufJ5M8MPgDTIq7Sbgt5zPl6HQSJa5nfGKHWFZ4ukr9S3WltOl/277O
twJufCVIxeF3YWcOm8KwmCmSy9Heq6oWmkYmsocoZLtvS8WyDtoWhNalLSCLwN03zghwyhq2RLRb
9neskZ6BmjefHa64YVGCWPqy2VJchY4/iVjkiZo9inhmi8qvzUppEbJbZbGPUbzgfsd6jhQ28cp9
yzTirN5TBArTynz22+McT3dsReYQIdp708gNtxf0YbTuZa3rLTHePWPduPd8WeoFFDIUgJxtzOIP
ZsngQ4qViLuhpeSgduoDWhzU2wCk5XbqEKMWVYEvVoIJABesp/eJGvY7lQr4j9C9FSQk2R5NqYMp
4MijClpsn9B+0+nJXJV3PHWbc5kcsopFzvd7ZsESpeUW23pVK8F9whuKevWo1tvKyxz/+xddu70V
LIjn3qYC0BBy4tw9qpx+0/Y8A4U9Tnx0lXFDHWk0LTrf+tDNLm37BKEph/swyUC74TI96hO8tFRf
vhwYWAuvAZeoXyizRDeQG35PTVL41w4dUmjvHdTL3t/hisoei6jswhbRrtleSZqvx3NuCr6fBDA2
dkqBUrCKMKy/T3YbGO/BOw51+i1iSAG/1m4Lkhrrav/DSLaQyaeLhhnk2s4Ri55xjHjDcTnUwfje
mHPrRFlYCTBQ55+fBpU9eJS8Pi7OT9Ovh+go+VWqTXtXBPO0gbfiedK9PIKr4xUTxFv4GpnnbLkU
hxIQmU7v/W4po6ndc9YiDWGjxSYdp6vvg6otpVUpRaiFMXm2lxY3EwiNmP7LCFAXp3K+P2wOMhio
jNYkj27HvhZUnvp7BoJOmueQrLSjQvV/GbX8E+l1x9hU5EVErdhYuaEgWz6pdNtDr78xpJq+oXas
il9a/+y6oqtjx83m0goXPg3RgBuoWBv9mNS0oGcynuT2j0YTQzFSXYuLUc8UtvfDoLK3nVGnSDVZ
d1YNvHXBjA7ShF1sOljz3zRmoUW+aJZ7wTSU8BW1XuPB29pnf+TrwCuBBddajXx/2RWuf4qGm02C
1M1K2upE6VU7MD8C6sZ2sgSaWiCj8ABR7hYgWyBdf5/2wZZRvKJ68AxdeVqJS6D1jiOH1zqmWBca
03QxS+VvPKWwnLmZaZS1Jho2eJrLUfqXcAXC5mVauSI1LdgPXFReV2+tvu7Yyl+cfPDyH7d6MRUF
9rw8THLW4AVK3GbvOhtjlNBxDpufZeoO83r/nZRHmevc2Z/EkbhdOoaCpOyvfgo4MSwdHGOtcXOh
TWy1pzYP1ITUNnf22XMIYlscHpB8QCMW6sA9kgto+5SKm0sJ91oIwKucoNqZVZ9NkwsV+lngO+5u
1mUJwPcuowNPpbz/q1WlBIvddh+TEaapIyUZ90sz8GT/m7rNqWjvAxuY8PKgmYK1JXf2VOoKRBWZ
FCE6aueEVv7494oJRFe6sV1+5qpxpjiamFDJogj0jFHfFN8c1nJL7z9KIyygVhBNYN+gxpAcjZOR
4FiOyj0m82pQMHToiaBEGkvSaFWdpjVdfd6cjAvrcHRgBBM4VeQKpOtoDj2Q9bKUbNH4LYo8seFK
MhS93RN9gwWxPBFvPjcvTCMksPYksO/yx7QS32oujwN7KOGpac45mhwXLnKfY1yF4iBzjTm2Ni1k
klWUT6wpxWljTIKhTubO3T0I42Riz9NONmpIv6n4MbHMC5GMy2vfBHe3MXiTIX76yTUWVm/HpPRl
rbXiuWCiTL7Hj4Tr1wtbeLHf2MlXM4DBdVQ2QlRdj57aXfSbT0TWAsAg+wDMJ7BLrRr79RUfLnx8
q364UcnQY6bApOt2t8zGLNFSbBqQ5gvbx7Ifx8YNosGce1mUtzRC4ywhCBaG/mdzt+8nWTnhH/bo
R1oRlEmECVa5o8yRWD3ym7S75QR9bI1ZjCz8LFn394V0+8yDFCEbRfsv/GlTsdXZLyjS9I+VRJy/
zYXsJFOQMpf7cO8AZMVbXIXHlVg4I27YSIGOeJ/RBTmIRdddiHKFKhATHW+wCtVDLsjk5mJe3PTs
zIYSQ3MnzERneXD8qFxDq2bGSP6k/pe1EUj3iUXCsLgB4Q+hI4MceYrYHBYlnePMvJi6NzRgOBQR
YfXefwHoH/AMLqpqv2LOAnkSUMIbZT9C9D6yz/Wzz7XVzLjsIBKfTtHeH6kIO3vbUbLRGk0wXa1p
6fvSBpPDCzM6Wixj9b+nqtWczG3OTsgwsmUyFxkReNibgq5NTGWLc7g8kVS5bEl9jkcuwpssod4A
LeErDV54fHbdBWZ/HGlxTQesVKM6VcYDbhBdbCq1KasP7siu//iRjXp3lhLBV87Icm2gHGuR/k2h
wRbz9Ab/8x2RzshdDGYlL9fRAf8AYQchpdsmG6fMQgzXUqsJYgxVeXU6tGXmV5zCCQsbpdOQCSr6
ptZ5OYWB7TgkXtE0uOvX/nMHmveX+nt+sx40CvGXBak7OwXLe/eNUKuSLwN810X1tVUclC+XzrGZ
FANj3W4hGGlEV3oQeJYfTR8sUKwyuS56VP9WduqiNcGc13omV42Blgaa75RsA/5qufZ0Xhy7AqxW
bZzNIORAqdhVywtWCjQ9O+wzhygUZSQerLuDafUSmjjZdeVrrf50hxlaMaK2yM3+EM1ByoObYwh0
DiYnXR6bINOinB1kyvAKDUbTXZTNDXdHciamfTjp/PbSQJZVuRD1UYZnTGPUWTJXSKVJMu+dWLA4
ajgwH7PduaUomXIF496xFmkWRW3PbThDxV6L5/gMPCFzq33qx3xUKeNaWRAB1OenWdTvQ+zGV0HR
pRrX8ftccWveEWYuGHZxCX10PYMVEVzMbze/ahGLMoUi/jOKaAbeqOTs3ivrScYRoeTXd8Lvzfp9
5PR4fodqFYAnttMXOVgSb2oANruNFSO2Yb29PvNWrqtrIEh9x5zZMDBLqgso3BQaELxl0nECsgB0
Dci6bKOqlKEjbNF4R9jf3Xq351VzTzX2l280/WTZEQSRLEtjhyXZUlblFkNWfxXh3Dp3AEitvaco
P7PKRvvTj5PudgxLkjr/2ZMvB2PkAdfdSutvcHYI38B3U2jmJ7hVPUVNMxqAOkrIsTae2ExnQzV2
/g6J6kOptJIy05Lg28RMPIUTfHufUC5/PbEpIn/Z87XI6ZA75IiwktaD0U5kP1GBjlwpBR6oP8cW
UAjJU4kd29E7+LrdKsimFWNlUUWzxE5bNFBJeMxt6KXO3DIY0D0dnkTKsWTbcqTnKCTbM/IUEDMG
ntjB1+zAi7ZLfcC/s72708cLhxhKafzp/BVJbVk8/rLe6Kez0k3ip15c6sHxbf4iYMPlU6pjpVgC
6O+EOLCCTFMcKF1AfUWmfJ1MioY/8Z117JIEkCrh6fTh1qXf+v6Ltq/h+7vIoAUy4nLimBpX3hxo
9B4Ox9vZBFvxXwXRIsSzDIaGCnaRzIIi2Qabua5Y6IW9HzHPssuG8j+Ce4H2q4XXmlbCIWCvYZVs
ZR76L+Uvl5OcAeWD3n8TGlQHW+QqUYwE3dnvrlgYH/w6GTyDDU5EDKFRcw/U4ICe5A9dSOmCP+Kv
Td+kZaqa0L+6e9CWTjrISR3DStRb5/uRci4Ujsvl2EaSDL5E3SNw33dImRsCGTzp8YCqAy2GbHjI
rU/yq0ZTXEnHI5zCuuDgKBPf4aDlo8xHvM3N2NxHm6m4tRDxEy/wCEZk3a2VMlCwalyHfNUvBtNh
8YxFKnNL5s74apeFkwK8lHDHl8iccmYiGoQnZwZCnEUVo8hjoY1twMtnEEvt18Ut4ZikQIQ/Ugdw
ZMg/N214jrTTpF5AwdrGODt33wPCKlAQMTD16+jAf2ZDZit/B4h6Zmxopv2Gwc03zQJU/GgXIYeJ
z5ba4g7Q7xdTjUiP2KGOIyfZ0A3sS2dT/lgofhREZEY/ytSiVhjXiyze5gO7cGKKH6SAytJP3SAE
b/Pw8NsRyBdbdh0z+Iiym7DL3JwgniNsOQtWtDaRJsupzLT7GcLcG7R4cgF6gbmU3yPhCxHus0Jv
mBVVNsz7JIz6CX806UCyHR0SYR0JtuDpe76R+fjlkUC3FNLsKvuHQqLazYvuULf6ChFQSXwmjaC8
ANyb4Dlg7bjgCJnaZpvMsj8UBaoo/R4qugI4YJN9TfqMpGXz4i3EKaXg5S/UESppTtZ2bplt9Lac
7xpmmqeM+1BOlXdAJYxGOIOAadC9P5YMmQN6i5YpL5cGFePbHCQgJUjrqdYgdFkOfhSVWomOvIT4
wBEgBmflCvvcwdIE6OmtCobNw1/m61bbf3IeFde2fbgaBLKoimwId5/EBpcCNxszt37fwUKLa7Kx
+0RV9WybPBC5qypmNf1Jt0XDqBA2FF9cn6V3J2NQ1n0L1cR3+/HfWmmu/BM7b+Ka3t7k96OanmKB
p+cgXSjoK/7P762I6zwnFZuapUZwvZImyRtd3CH/WjmPPstOt2S1uzaV7Vr9AhHWJF8v0qK/T74M
MXkth0xjVE6Ke8q3tFt7ZRQtREH+9AZr2jXS/5LBQ4mofcwiUD5n70BrM+UePJOkcZRlvgaikr/2
joEysYtNR4Dqg0JGk5fxjShuyizeCwfSj043HxivqUhI34uu3sqyUMY8D1eUjiwBoD1tGGJcYkLN
7wcxHtZYdl8F8BO8CQTent565KmNebHdSPnuw04hYWBs8Ou9gDtNpvmg8UW6dwfw/nVi3ou22OQP
Qji3OhuE3tBPZsvWA+DbJ/hAoN0A2T8mjDi7w8yPdac2wP4btTLV562NCmwvMrpLf1YSiyd1Scrj
e+av/t4KjTT0YVHEHf1Wm5fsTDwGYZGy33g5Hy2++S9hypFpXLGv69kpSo3NNplZNGzV/QvykWdM
6u58btp/WBXARcyKVqBeloXSanZzb1pFbBtV6n+zyyDQKl7JM5RqQAaFsx0bs1W03jcd8rheNm6y
EkRA8MJbD8aDRI4dvLYUY2kaEXusszhO/K9hh0MAzIqqiQ7gedrLowtxA5h+C6nwmULKldJMn4pI
uq2Soai0xTWn/fpqjAZSyu9TfsdKPk8e23+7ZRgk6Ilao1xmzvX0/UFayo/Ov7ov/dUs8QyqrwKj
8tXFboxymHbM/7J7Z6LMOBHpOe9HxFLHAbwmsD07z2xq0LakoquM2IgGOb+P9sD/fx75NC5/qGb0
ZWoJyeWyzyNR2XUsqpB/DdripYK6LSYXA/ndZFEIQsxUYW1t51fLO91VhWzWofGxm4OOkibCzzAm
tAugkhJZS8q+3N6tZaoSdfcOhbNrxNoXC4EX4ag4PcH8ejiOLMO59axwJ03ogiartQ950kYxDED8
hDav1Tv/cG+Ph6Ncxkw70xQJ+L8P1FEe7wf1et5Vt1lFT79qCUMVH3xYs+cX/uP0jVW+Sx9uP2du
eCmuhjpMBksmJTz27zgH8g43Si7vYD1lYoRuzUvzNxfmybA6wjLdGnXrAm2/cVr1RZdaE1GfxuBa
pkOF5LOJnOcE1SmYKZK8ucoNLqbsmtkS1/WCm1tCLY4m2K0OLZleRzoZ0S6Ci+obDDgewTKL6VA+
r9GBcdJ4NgiekjUwN/bFKm5TmrjvbhvhL6l0RlYVxlTKgw31DVxvLFRxQBboxIFaJ0YyrZYiCR4j
JAH5FCg+BOi0pq3XgUsfapgXhWy6MA1F82UUgBzsjVcouYNjaH4mOyYvkb33n12OiPQNr7X/KKav
guykdxVA1OlhDU1zFUZmymgrVToZkzOFQheuhsLR2beqr/p7dBWdeKV2XvpCyMHsp++axwyWJotg
od1KVESOd+Rn6JoZ08p/7yGhh8XePZbJTk23eM6f4Vdh++unvMralmXenPRCILmy1snSFquON4Gd
VfcGXokrZ3mmXlhITBiHSOa/M2gQDBFThePAA9YdIhi5+pRTiFZ27iH1U3vsU7mNqr4agns0V8Qm
m/26W9eXtT87nSEa9yoLYfeLPrEDcGrO/bF8/4REjPVrVvKWXeWZHwn0Zd+p6adwFYaGhHM7iT3h
xy1AKOgQ1cYDQWu2XX9syv6EJFD9A62k35nte9kDC0YLTxGTSi6XHcEBwNtp1ZUHdTXPtXQsgANm
d/Z+l4KMtohYyxghI5Muav+JgFjYfczEdw8l2WbLrSDFtKA3PW375273FNz8Jsakcjph0hog4ito
h7a3mV7rmLIqc1eypMy9oeW4AYvfdzvhU8jZogSbNDGddhB2BubYu/759gGGw8B8kvBoiXs4emKI
sf4XsK+QLULyG9VzykKBJvRlGUPZoxCC9dWfFvPhk1LJtM6ztHTy7fdKe17DCGO6STO/JXOd+z+b
ptmKIyeswQugh6xIacwSpVZmPMp4rs0Rtt7MMBQuiHUTdLo8rKrSh04PfwUUKtitQfDdcoI1Z+gg
qSCESAYBKKTAWpw4gh4bs0ulGFiv0VDgFiYZMfR66me87jBiF6BepANTQ57Wd8bvS69cNVYUFlKa
rkwQgnstsUq0owrB1JF5aTVOy4UFR/1i2Dew8HNdM+ULmFaFNL3AEUPDPIcJm9LE5XRvTpi3j6oI
404Az2cAlaSErYs6GHKR30G5AMXsNZcVdIIlbOW1c60pLI1XQsqU024KE61Sx0b91h2MpESb+w8I
F9u785aulqMcSixt10SKvd9bjDN6K7xbl6X8r1AUYC7m3VALDQPvLIvrtF54zDti+Bl2EMMlDkxn
RE+995BM4D3n+tqDAANr+aCTc2nkWPZeFOtzeVOvtO+oigq47wdUc74Sdyz3j2dXOSTCu7LSRDHi
dSzCZrhLSVJVzHMNSIdhdyofXE83sOXNNpCtbR3fdxzHLdQ3LJPG+DmrngVMHtae91Ju05qrv0RX
Cel5ABpl18iJud8KxV8WNs69ogToRIHT0fO33AAyjjl40HKw6QMpqXP5jtAA7u5sg60z2/wKb6Wv
1YLayJBvpZ9ctb1TZSTHbNOqa8O/uXosiEa3pvRcvLbcxt5SNkdAiiIxOwXsA2wV/HJ93AsY7+Mf
3fIZcZmZx6mdhDMrmbxbptoh7epPl/DesL+tOqVNYhlmeheFcs6HNvlpX2a6GHbGWw6lqWrBCOkg
ufM9tTigP4AX0cPJNAeXfAzmwxKh3cjGuhe+7HqKf9MzPUyFfpCNNjx1BoC47f+NOHOuUeS4K9Uh
2PtTBSOEw2+IlslnGCbYN/lieCqknhIRc9gY5aSCygEMyMid3jU0SlPfXOPluAr0aiWASp+mAKGX
fKB5RqN018ZFQGBxDjJubrDPX95knP5hQGF5eubSAG8Xt6Dw8leWzAoKegZE8jFh2z1ODzf++qq+
xzRNTjNSaMwb19R9mbSL3H19QfvL/zRgKiTB1qhoMn5ZHpi02hArTje+7cg3zCpWS8LUvvxEH30F
gQaDOERXtyvO2XWSAtWHV5EPGSu/VrrbMMIpaUArLowXg2vsUYNJArxc/sAvl8YjortdeIDbMT0M
ZGAk+osEv+yeEvcrxBf7GLM1s9dKvsuR/+c8ygutDSZMtOFWhr7MSBxQyR5uJ19mubzs180UXkAB
mVrIn1OMmn6olRwa7mRoLNTZem1DrEsWLYKPu7NES0yuSiEB8aQ9xgRxq3F3EBBMLRaLujfLqnOj
ACJCyTeZz6CBkiDiSdStpNbKrcH2y8lpj+JA9zLQWBqPgWoK7cnv2WvW/1HpzbYQPQQn9eIiQucD
PpIMAmvtViXwz2BigamaKNYC49RbNYk9psbg6Fz4RIAnfncFmtmtIK8g9rRlOFqHz3rjdJfacwbk
WlvGKoWWnFz7rNTSnXHrtpjHxw1tCDAqxEUuzcgqpuxOuHJ1RcE+2QDZZAJ/6p0yixIwPQKKMWxQ
6g2JH1i0NEqe3F0GUO4W1xpc9j4Y4Hn/Aass23Wmdc5SFWfQsaEF3ILzvgj63yzllKtnHBAtvFct
jzA12zjC9eVv+S9k+EgOrTSMPMWGIOChGGqZEQPcHbeS81nNqoI9jfi8TH1wOMlTCac/KNccaged
+5W1rbEOnxF1NohkZw6ETB0aFqOihuteGUjwhzLdMsPbiws15QB/Yo4v1aofkcHQY2rfnKdZtWiS
Bh1dXRbetZrfjcsVYL/RnBfFBaIiQYoQU1gBuYjfM5jL/HN4Ecp+ETHhoMghsFbPD/I6KShV3vTh
vg3t2H7qhXsCiF/hYSNsD8n1uwHaYm8LU+lDcjZUfYBvzcq5g4dMLgzAPYeuEef/3h0KchtReaQ7
wafxEOc4RCYSJ/4dRAzbWIscc3PrGE8VHek35TGTQYAzbCvALLA93weMJdtaAi+V/oL4d8+Qq1/n
snNnYH8GnRHfh1Qr3ChHHGtMpJycJI9C2y6YFs5VF+TXBXU2UyLmPuCnHwBLXnaWhch5+b3PS1CW
1gfGO2o46/DzO4PkIQS3eMWvPUQ3mqkTmJrzmGS/6KtoR1dpLeExw4PL8VH1eZrQjzyhB/8060io
O7BieouDvlletyuJ2T5rXKcOxfqYeRePlo+fPTxk9eBIrmw04kg0z7gZhFXHp+oC4jJQgznYrzuc
drSLM3+dWba51L7ADyUrTyx/UlLdR9yjvOde+C8GKIOxmltc9tcNcnL+JVmilKLmIZckxHp9A35k
HD7yOQSr6gGj5HICy3U60+GdZBXxI93VIRLsPWEb+ZTW72DgudNgYI27stIG+KkHIb0OAvfsgopu
NiRuGJYtl9hjkRko1OpaavqHVOkBGQrQ9n8Wgt5wKlClzeXYOt5HQ7XKv5YJGuOurX2y8gwNI81y
55bT01HOXStO7SW78AQDRkXbseA1jPEyTf3LgZDOwf7b/vsz11yx45PN005wpWMjtRZQWI2/NdWX
DRJQTISSt0Cj1nuZVkQqLBWDXV+CJ+xgnw02gwJ60rHhJixeIf57LsLNpnp3B1nnlhd84uPmbO+y
mErm0RmmlEfqMRP5WPRpMowJmnReFMzojR5/V1l1RMhxQ4f/97cDZzRlMHbw+fR02A85mFD94b8T
rnBpBM9HLqihyMlSTBiG4IEcdeFbfYUOd9ZhWc3ZTLZPiQAJ48QTvKN3VtIqrjCR7Ce+MELWaDaV
6deu4b2nJmP6ZCsDBAQitd+T8cWJmOZ8KNJdp+aSYfx2LtqyUKmq+28WY/dxRo5ONYtxIfp1Leyi
EtO3dBAcn9ntmfYjCF/achTIns7V23h1kOCSW4JlRjDNQ477ATs2W1auv8CVnUht4Kh5xSt7mOeL
hzEztLGCmA6V7x3Du5ok2GCC+ciQCQUCuZrw0w0QIAr04rmeFwshyXTm9QKWv9cczwMOa/HxUiO7
iRlRm+amUkSDYgjLneAV52OD9Wp5sDAAtlahbrICJcpDz68nr3SI5no1Z+dP3UwKTjTZFLStFRZT
E+RFHf8ElklZTMztkXZWGN9/bxpY428uq8YOmg7wav67dft8A41QgCw/W7HsnKirv1DE90SU7u6w
ieZMgk7XEjAyI8/zrtsm5CJGKTbwbLPjllLwCZYEdozWBg+Bv8pMwBT2HgrRpJWkHZ0QGlQWtgqk
0XrRLQG6R5i4B4slR8ZNlDSpufRh72eavj4ff/X0aYC5FK+AaICBBRYdMLmCNf7T2gSea/clvHmb
ms65d9t/2X/4KKAjWCcDrJQx52ax4E/z87YSUX8WAjv6GUvk2CwJjGXkgGU4sb9HkzpUniCfDoo/
Eun2en0wZTYjFY6aC9f9FoSxzssU08xW/xr4PUyYVfjCf57iarx703HT63lOP/AxSlENzDcCuCTm
9osA2OtRgNMfWp5FRZPz3ndU1Z9Bgm0EwOf8NHaZia6qXKUxB+GeihWA6tiZ4soj4E/hYUjPIaqq
Or7Iv9VOg6LR/WHaLb4/dhrGGuebcxYPcmZ6yDnGqHudTdIkfl3XPrFFiPg5bJmewonWfHC0u4Rm
L97sur9vAj1Xp30juLTRAcQjTe8J/OomDOE+uqJAdzhYOTCHLpf7L6pD0Mg0atlYPqcgY0ug4OEz
mN7VVkPsPQkjsYNZGJho913P0najkaKxACcKZ30ZoYPll+Q/zJbd9OI4e42rcDXxCkQHHUzhq60F
YwoOBgGkU9FL9b4mTN9Y9crgnyoO4qsee/4LEhnL/GUkjnQF/4MuERsfsnnZKvZtMljyJEVlXGr4
5NRzxFJQjIeidoLCYeqBTeuCZsuMb/Ac8oplR4pCAUgl0YTKymLLwTEK+eZGwqXQqr9Amk6BJu0x
escddN5OKgw0v6ye04ghGGhmfgIFsly1nnomIPtZG+O7AhkCwlEqS4sBoqr0/iPpo/ubMfEyUR35
OCpAGbPcQN9AVs5REjsVKIjvzXxMjcZaMrF223t/Ts3ZWlz3+SHXf9ae9nbQIE44a6g08CHKFMPT
hGiBMl8cN/Lg3qEttAUaIpMStwDZvb9a1AnnkgfLhlAwY6blscoRsdl0c/eWp3isFtdRAuiBoIX2
V/UBY3RrkTI8iC785S1bpBwS/nujS/QCHb3lU45c8n2+4jwzjEsrm4YIwrxbq4BFJJ0TPcp1D32L
SK7G+j/qzRM8lxsC+f4+2BSs5he2jm1rwsELNgIuEHogQ4ZHxZ7ufAjSTchdR1yk7/3Wg+g+a3fg
9jD/JSutb9eAnvToAl9mHTmV59bTDVCHhELd9zFGBIXdsquIVIWFHSQyaG5GdzeeM1QTbcKFB25j
aBWUc1KLZa0AvIXxkwHUGddMqbMn1MGr+u3e6g3b7HjoUu61T7oFzCKPQp9MNapsZLVca8MhhIdL
1EGaLhk7ptxXtWQ/MPJfLztWWoyIvttcoRGHJggZacAgoAiAonxxvVTcmpAbUftv5cQdabPGej8W
Mslb79ziBV6MuorNv+Xvwn94+HsDrSuBULbTRoC6Q8lB6BOZ6M8hwL1mwJYNKtdllISyAPIfTlt8
L+OFtSGu7rLAYW4oE36OsH0oqdAGE09ijdXv63e2+Vu/Xk0lAou4v+4dM7Q3dbQ7KqJvkNd0qWK2
eTxg+rh1kQ8Ln0dOjpQFQCTVpyLPox10BYJoVwa73OhS5jGA3RU5lzNoHp3NFnXCEZijoOSX2NR1
7cBue1r+PONSJX8KEZwf+BQoy2Alhb5XddLko3YDl1+8ywtF4C5YKkm+2eUwOD8jG+obWVn6E06h
V9TfRgwN/TZnuoMPVRicLgZ0NQht/YnyOl9TfQRK141Zs7OFhytC5J/fdYxdjhZNssUQf15XqcDb
KVgUHMCwe73hz/Iizgoi6dL3eaq37/8/J0PBNLUsgrIe4isBjyhY4W+Boa3Z1DIFpTjo3Sv5uPLu
FFzs0LrRh9hyVRN9EVQnL5Wb+xBzuRP1iD/xen1eavEztJ3WdprnMV2LlcCpiPAKUwIHa4NiufLQ
XPAhuMdtJUFLiT60xzfVKR2+MEbm6rvoNLWT4HQKeSzgn3tltjgGCeeTj+DtmYs7Ce+o9qUCH7Rg
hDXzJTH/vFe1vEUCKGPJKZgQG53kOfy8tpy9OM+emeP1v3HcAm86usPRWRNzFiemz1Ux985f0ybT
CdUZ70VEnJFnK6G87oXX3WBhkRw2VZRspeKfC/XlU+zrpLxp7jF7zEMoV/ZL2rsJVkSlZebeXmiH
4oAbJLpHmJtIEy92r5g2lZKGmPq66ZNZb74Ym5lhChRY/bTDb9lRQireP64LfEPVVjKpVgrQgzWk
V67xc7TmnEuRp2Mr7dq5A1AaD9X9iIKAMu/6jgp2YDCvC5n6IDCsq9IPiepHh/4+iaC9DJhAev9q
Fl3hfmy6FVP94ZmW1dlvUFMGvl0HNdi55jPmYPomSa7uFIZgasDHTmno3/1LLD8lsG+x6Rv8ss54
e5r8TWMt/TiYJEvkrwBxWJv+KSGcFQpmlnNtaPN3omVJGhZ8wfZQMnJeyy1JSbsjwi2n77VbGFct
qqlIKjymMSURMa//pgPdcC4sl1wPgvcYXeFJL6oKyeXaol0LES/wDWw/2DQPn9fUbVVF43Gff/rS
JcIaJ4lhWP8vsbjzo6/vAPRLZo+fXdx5woStBLHYWU4L0IuE8PKEVNKiIPRYDTvMHBf50GZVcLI6
ulrx+pVO1GHNBpTAYjSJ2mZvLjzy2IgQ6APaN6sKguaYXn89ukZv4lqZXmnyjNTu+B9oZvIuEHZw
lUwO+nq6W6J20n4xegd8/eQoTcmrAI0DnV684s9eqKwklr+6zbevAmZ5nQH/yFCjlgXsfuUORBeB
TLiai0TBvvdzzKSF6eokuNhDau76PGQ2B0pgYKOuGckOTTfIlYq5z59l5yHiKLFVSFYY9SQI2OZR
zmnYrSITOJ8z2aNsg5E3bf+VKhJ/gVVJMV2jsEE7pQwLY6nhjFmsI+TpL/UterpagZxTxs0I14+F
nvGUfzbLCPHQK9nByfzR9F+Lu3bdntFHmCVdtd6OfNeMO1IzV+9CEVvL8uq2bdx/OkpPQLzzmzw4
rankpyxV15Dhjp6LrwZxMY2050OzOmWEevIGrfLf7JFBhPEjTLr9DrWFEcjNqfjv7nXQGAzALwkk
j18NW0EWAL4KG09ZSKUAiG7QaOv5NNEusvnRHtHWCjoRE41ZBWlMAnRhrHJD7pnUH44vyhF/U61t
IBO/lek6fi0bh0I2MfSEEyGfZZ0ueyp20WpIcwHZBwJaHpV+DC/eNTdlvilEW8C/Ol50IesHtgHM
9WCcVM+7qDJhsJGft0UGvVJeh9ZLOIYAhjL1agUrWxuz/1acpSKLpQueDQLBOowdo3Pu8kPNI6Bn
/7Qpmd479+AJpxl/yv8GbL9A8t2H6sx1WyVUk9fVOv08Yezv49SxSyeSgT9xNdi5MNXSUjU68EJs
JJDGndNKXo+e6Lsu5xGWaYv/DEn5w9e82YsD5oWcSiFNSyhkb0YY7JEeQz45MoVXn3Ku7W3IVvza
xZ3HEbSgDxYjftUflAlUJxjqlgmwe66iMi5pkKhYZQ8AhWAj34CBHBWhH8Np+0nXG57t9fVWK9L5
meDPD7Rbvj2utxnnzireS1Ae2a8qo8XpvA40pk6y9ETf4Q6bB4jsA84rv0FTEt4ti0G32EYsaJFM
QjhOc0j1T46Y8HtcC9AHZeD8rnXDcMi+O384ukIr7nGohw8UlarJfHue4VGmprT0IehmwCVX69iO
b3zbviHkQqj3BuZ0+eu7aUNwoZOrnAKGZ+lRCLsvUXrCWQySw7snw9gZ+24y59BzEdxQEr+44vDD
hFM+NY6qVeN92q/9KwDsx5hoDKgLADx/yC0mD3yRLasKyV5zJhPdOG405G8+pBMrUAyZKMXFa3Ka
Rz5nIqMIP3aOiT4Sb8bjcjc5ISpUJbnudz4EuSs8ZlpkEoUTC/ge7f+eejn5JvZhceiWWwv6tTCH
PkmEubze9ENPOomkXxc7Er6c65KlHJ1+bwTxQvELhSMJy/lciIW6BQFbetlOT5Hjw3u4ORVEui26
XIzRhx0wuO7CQSDhDLoFGmMlsAlTRWiX0fsL+6sFBLygVJLMU9WFNijYXjn7M8YB4GIZyVKHv85q
ZoV5kJ18lc1MnHCK6fS6LZd/j9uuvWi/ANrawa21FKXovZysv6cJjnpS4qG2GWM3uTEYDcV9Sfaw
FA1c2VFpvbA06RZesvKPWJQXWwiTiwv4dxtcppuVhPUDu5hr1MYJzWZRnZ9FNA2Y1j6smZHZVNqY
rYwCvwq+M2SfN5DJ32zECpHnDo7n6mNkM0yA1N0cMjMuw/F9qZZ8Yb5oRoqdH6Tr20/8ugw1l3nU
Tg9s6fuTX0/6Jn3Q/v3FwMecOHfkVw0bCyp0gRUAuG+hNhmMMD7pMjX5m8cW+fXZ3ep9gNNNVGOz
72FBBJ5dT/cTA2N5csVmJqta1odOq2xxrhG8WlSj8ExQSPWQcbW9RkJK5F7mJyhp0W4MrJko5KPG
LewRyEE+EVFO/qinkzFJrFdoR4ta5hRaWqFRQ1/7u450iXXUNApWwA1YAFHi3bNfCUzwBm+DVYp7
VkcAgroTslruTQQ8uq+8Fm7xUt6DkssnyO/aZSW/i5NI9vcLrP02aj3tsmyxRE0DY9Qh2YcXwI/X
RPYtt/Di0pto3Xe8utxsKB++DYT05dHJyi35FpuGFxUPHh8a5epmn/SPT5uSnfs0w5SRAuD2CnNh
q/FnNTkqnGm3UVwU66HfYzcq86gUEftcJjGeU61vf0Poz/OEPaLMvjEls/MTpVhlUB6VziijfTy8
4+NzYcYDQkVe65gZeaMxK6pkF7GpBpVxZ3tanW8mQsd4z3IfGgeYVyuFl3b2Cjfdq8SDJHuctN51
KrHZG1+/l6HSUUYNSwIGGGHX0q3+4uBxpHFXOmJ2ocxS0w6HsPyvR8YpVD35XsckNC6CNsczCpQn
kPrRGiOJ8x2UCa5Rjss9MCbEtMhoKYl/GrI6ZNsS7Rwi4zaDQHNr23Jm+cgJVw3ZaOWxQdOY8IlM
FeVxXSIlNOAxUp7HO8XQk59p0euP09B5SbuMJuVmqFh+2aHwY7Bs8liHRKFU3eMaILmoG10NutCn
b8teqNUtHJLfM/8ocqcBKxPgDCyGulNUbqMljJBGS3v7HoBIa/jGhCVEhqooEXnncsk+6Q/CClkZ
8zu7yjEtLzAqiSSvYi9FNMNF5L02XQH/ERvDxFYYtqWd9smG45pYafNQ5yYQDSUoJMb3VXzmfsn0
2JcC6fNJRZBJCo5ZZ7Q/uImSfkzc1Z6sfcGvReCPOKCV6o5Lnn8BDv2Ta10fJSzm5BVRPElLDKjA
bmK5bPJv4EqeWFxnmzxqxcKUa4/XUwONTqQhXKp+xTYmVN/TkfNge+tNO69Orp36zY6o/PkDDidX
OaCGHrS4sYVkqWtS3MeOeB2DwhiZN48cks6pw2laQCqiQMSjN7h4xiANQuo+/hYR+q0lZbgW9sBQ
a3tZG7Xp3Ne2sLiplWaYDGxXBodLi1ZcTRuIuFfo2A6yyyNIUyxeEiBRCjGt16EZONvBXF3pP7R5
9ta1N90bvl2y4miSAG4kzUZCw5kZJ1RyyP1sKhz+EJYZcI1ipo11z+K0UqpSsPL+giqb13uGQzyu
nhPUnPW0bY7UCt+uId4JS+MubdBKgXbajvM8ePy0dKBeDE5l+I+mNlcNAuK+7rgaoOmieoqYOhbZ
m+Qoy9tHqXsns46dB4mHglCsL0648tn9hmWC1E5I/Al+2cQsSuxBqYxKIk4zNAPciOg9veMyk362
N8z7VE0CvogNX9pt/r0I8mcTs2q+Hqe3pTfs26hV+557nE/EEzID68tqpLYSLlHd6dQYhGsm896c
W7AOuJauJ2woSErAApkj0lhZ8lDrbddJUSxXLEwbf7dAiFWBJWSTj952R6uipjnXYd2G6Qfz0dv+
PvcFQkWWn9nhxuu8koSEe+mCh5glZF9nMoHoH8uRWaGu+hhSnVrCcjxOzyGaMQpiB4wiYfwDjTGB
TmoboiIUCMbpazHn/0U6060lXKqyAEalTkJI5++CKhbnNdsYjn2dDYA5+3xnJIBoDST4K490LOU/
1rBUt1KV9j79jrgLxdxC11XVrGQ7ov4pw0egSKvganTQZw4aV451SDs3sNWs1+JOk2kyHDDjF7Xg
kv6CPldlsHehVY7/us3GccO2G2Ea+/2hiDoob+cjgJWIXe2/6pY7F4C8BaUVU8uz1/30LT8l89hM
4SBRD5wsHZezKqnePNPVkvzzdTiAhtgV5gld5sUcia8sbWgW5RJSa354P36aikGA/ioWSbBwkoTi
u2tqfo8rWIHvBZJODHJcwEbH6NSMWe/4KEOn6OX1UmIn9ToXv8xSlFlNUGF4wOBf0EITMn808tTH
bBicXdy6zHcoZjsA2rHPdFvjg8kuahfzUWhQoMeFaoyTg7qY6lFMX4IovgbyoI2RmcXGwWOuukLM
pBBpmmk3H3hIs/LR/I8xRnc2ommpcKrt5Uw/b+ThjGQ7NkdZGgv8Qtk5s8hb561+UNIRGA/OPnEf
tfaIlBM7tFK0lDTsA9p+yXPRQlIKufnQ0E8q3c6+pD58Wimf5cZAXN0BA1aCOF5amcdckDzh13/F
CGh9mHlph09p36KKj7h55PjK0/KUtzp2S9uMnqqWclHGHvRZe8FdupxcMomEIYrrYLFHsKeg5BQc
mwT4oYN+7Cq0LNfbBc9tz7kJbdO6HwYL1qumnicX+CGXvp1pYXHgMl+STAVr3kK0xIRSlEhFhZPg
vVWvqzgueMFJmiUyg8g9X8/d1BDOx+IaNTRyjp32YWK4ksdpUKs7K06RX9/9IsXmDmOX3DZyfLKs
I3TbXYkob2dyUpyBg7ilRrlk8r/o7yri4pZiN+gRdydv217B3VdWaKbYr1OkW0aEmim7or45kPVl
+OHSinoqqJCVoU8btSsUphBaEASRouxSVJA/E4Xxq9XJ97Wsb30vsp11a9vtusmhc4zb9KVIt0s5
3PLuZUr+k5XODPdSepCkzU/uq9bBIF5vcREHS4QzohY40pxXTfLhVDUcclM0jcm2ey219gOc3Jh3
byEHXNuo1cmkLDCFtELc2V+j+/zFe+CmefvNBKd7xl/Gw55sLmWs6Sydl5vMwnyKrM5Z7yAZttgs
eTzcQVdrccI3BV7GKyZL3W5mcNGltkNIHKgx46KkPbQKTB/m9YbLamBwmdcvYXTZY2GXsfKdvTLa
jh8flprTd7pzrvyFY14y+FxzJQoxvw2VUTWhtnJo5Q1izRlj2ZKTp7pQcUfhi8NO9T4kJwm2TCNh
nSI8nRBzAO/ZTSA2YSwX85/NVOaxfsJ7q2ICrkHKXLE9/sxwTD/Yc6gNaV1KG4FUiFhecwZLR5k0
qKz46Ggrj3xDHRZwCsyKYFJGirKIk4/QiTvGr6IS8XdzFCxg/125ABVoz452zuykj9uBNVJ17deU
mX+t1tgAKGNTk5EVQRwu6QgmmWqB7HHqVROFwClV6MxGJIN+JcNsm77fCR3fzICe46zTqz51Mm6H
VyYsLaOUVVBHcuKwOG4AUVl9qk32Q/u5/szNGREC6OWdxPdSU50FcJ74Xwbf88SzCY4OvpfvRtMb
3AyUhriIkwQM9HCTIoA5b6FUWFyBml5MlZUOHhggNyEg44L6d03PE2ADTQ8heeSJNIFTxTibE4KU
NeLp9Qjazes/mUZ5jsAKe0fLdDVJFpDGi+EW/G8lQwia3jYWqeYfTbDgX/VygJcvypWgq+3nENMk
PvqSmVSlX3xkV+ViVthnujpo6aD9vFzzmyXcgJ1INxdloZeWrfRsSnIW4pldt22eAA+u27vkfHWZ
Ao/NksJWsllyJ44zlEBYpwkLp1gC0vLcqUU/WsoI+YXAbMaphW6rqpExPY3FBKkyX/rzJuisFysQ
hbngaSXdvYrPoIMiUevmEGUWLHr4+z0VG8GRRRRPi53Ay7y0HQ6oNKHzV2mFEKGK1hSAx54CVk9w
hQzbIIhqGOSxWq9qA2havfaL8sLODIyeO6n7AG751U5NODBXIfN5imaxXYgNsZ4ADHott2Q5WlM0
GfKOOw2sgCEdteHw/cGBUVDtDIDyVV2XrVuGdOHJPzLRQTaQbw4j+mSv8nHjwKPUC5fIuMZetYb0
eGpDJ/m1RaJji8eGuzkJwosY3qUl0266QCwVOJ4TB/4SHUjDFMl+OaG7aRm/RmAAjoSrCgzL/FTX
pRWWQX0HyQF9yKvocAvI8k1FAHhpGfmqit5zJPqtAjB/wLq2eQdGQtvMEuEFE3s1gUImUCV00mxW
O5aGC4LgQM68T+H+NDNqhP/X7SV10LI77kvt1CkdhMl5o2zh/gf1sCLYKjcv5ufE4u0OGymZxEPU
I9NWF7kIhzja1ki05hd8Dg8PVbN7bz4bs240zdnFxlusl8TvjiwkrwJHPU/jdaoeP1a/5ykAriu0
PcN3P/U5ihid39QzL1a4wlhXKI8jRnQyrkdupm7/yk3UVzWWcni1QZJmyNw4YiIPe7wO3ZKjruIH
IYWKAWxO+jiADMHps1hayaQ5ryPE8vA3LEVHyHJx9kXxXjSb6ZxkEF/jHoKkRuOspJXkJg/2ZArU
HdG9LMJ5YYgLueCPOM4YtSXgOmV/2h7p+SyUcSuyzt/zZPQIWpquKGxqbBzNtUMBlDsvNZzC7RF4
p/WxcCPzhtpSLJpfpFKpL1JbvVfp7ROOOLEpFg9/MbPETnfvXn7GC51aGMGpkZlkgrJzgFGaNJWw
HM8Ly0M814um1ZkkfRpTmQi6Em0U8aBnGos6pQg3DElNxnjNL517EWrX8Hk7Zyztf7nW3yRauewB
lH08pa+ZXkjZ6/rMQNAunePKli1VTw7SF0TE/aVXIYB+J9xKZKFgl/qYrZGX/DYyXHCO6GI9GLRw
P+GM7p8GW3wF8FIn6y9CTW9nLpD06Am9chsmj6EiO1nalfFWbl0pM+tsDCszs2EUaPZsErBdopiZ
P/hafMt/8kf/5Lc/Q8h3EmcBlfvoSCTchsoVVb+B4PKZoSWvaiXor4MssJNmMLlEMr4krs1GRUEI
0TiLo4zQHgVbVlNMgaZn6O7hYG9m90uKG6XlLl2tRxrYQKbL5TYL+aoy2YQu4DTL9iRZ+DV/bS3s
UzCo2wyrSCXrD11oDKmlUP1o94l1USe3ZqySUeRbPtTiP1AgMO/kAIFyqq8z0OFhyDvt2zh+jweo
cfn74LQqawYgqDo3v2WRehxvUGvw6CNDJ7N+YK8NJ/uY6SoTxWP9unuJqEbYf0WUkTbLDRkmRfN6
kX9x/GUScs0X0O4nHFMucKSgtXE6A+AQ5KBZMh7mXrZJjXGHX30nkL2EXKOX6z5ohUDkeHl3RQYH
k8VhfrqIzidMJflrO6PQ3Jun1HbnBk6hdnLHHth6ta6NCjAbnu9ypD9/bDIpm0aDtb1gul9ZHZlY
edM7uNQ7UDx1MDGzsPHKhligjCLQ4gENS58mxHWzHUiNGjnUTLJc7N1dydGG/FHSGz9ty2Cj3kIw
rlPAfSgJswgUTZxlhZgeiftPIxsavuZD4bHVrsw1JbX6QHvU2B0TIWbmd+TOxXZ9PGV/pB1hWeqf
5/AIgyTNjenl5tlfg1fItpbReYnMGwrrDObwtSr9OYoMuh60+c49kcmYYVpXjS7qebbLhfhxFh1+
KwiBokIr+jR9GQQttUsYUL/47DWkD0pNpeIa6LuIHGQvB2snT26RfZJetulwvZ7dtI8M/AvI5Cyl
s798aG89PqzdbjyODAQ+L5JLNy41ElOzLKwHD1+EMGFfPINQBMIu3ByjgJqvIBgTsXbiDMNZXz/f
abmICv3dtG+36dPqSDS0RjasR1H8b4ITQ8V4V4/5VKdpqKaVy+dAXCgGrjhEWxvdF6usr8o6c5Zl
q2f+/6o7ptTY/OkUrwehoVD3P7o+Ywc0mUQ5VoVWZBwGK1dwdkTJ8YfZKhx5RxVuDYrspQ7CcTJV
HX32ScdGWr7amof80mj97mvS/dcSxyCM3kZmAgI5E82p9vqQsTa9goizSkdAYErIK8+5ncsvRCLo
tVZbrNwbrWf+4ONd1RPzXofeSdIgq/dKUG/jGSD/71qA4cavj9OQeStpvmEwRNoYUi9ZJql0hxwZ
Rz2O4d+EQWDo1g03hJmEcYemEmgFBLGgZy4dQf/qGroIaqpxLG9mHrnKP8xALalMsmvevVohQenE
/pOsmDws1ditRqPgqVcJtl+B8xsBk7ZkN6YuJurwaD2k1oCP44hRvOTxRUFkuvwdfYUwFbbPzqnf
1jbGz9CTEbwAfK6qzbUkG2+Y+YToC7e5CMo+1Sb13LUZ3/1isZ+2Xvab9jOeWBx24bicme2uW2AE
wWY/rIlDH4Loqg41NATr6K4BLnSH4sVXpboo0Vof61eF2N03QSyOn7uqTNkXRmi1cAvqdRi/+5Lr
lPnpeYuYGFRCrxYkWwfRJN1tvCp19P6A2lC0dMONfeQ2WTwkVJJFT9dezTHB+x8fXMbhwUHH9Dbc
i0C2FgmW+jz7Vf7H9EvI7OlyOVhstrz220zW28AnGeS/uG5Le1SUaBO5KmVLiI6Tu7ePq4w5SzZL
X4I4H3Q1r9BIhL972kX4qHJs4a4eIQTNcTDr4V3VEzGHC3f6Y1aJnN42gC6bSFG1BkPFtGaNhODS
e8sdVbfj2HgGPI9Wq57I3wHJIQlETsN51nTYU8tehIibxmWf/2mscj1K9R9jar1xT4fJmVENJf98
3BwbItYOR8+oO2Trq2deniyIktW56ggJAmKjRxGLzVYYIRMpnjWWB+/FR2JEQA1Lu5LIDN44WM8r
G6NRRSCtKVxsG1lUKM8YWf2ZxnmxH1oFp/MgYsszw0jAxJmEOaWAPiSeaZsHFEp2Bbqesl8IILbk
gjjWDHgBLC85gbePv3DWyNnDlXNT8PWl7g3RiwMs96Uf/y7HPUW4QNXMwcZ5jk34u8Gls3aNuvE/
0+T3gea7dpDu8e4hJ8ue7n1mqfjYumnsu11Ndvo+w/rhlEeKXw8L+j1erNPaD2CpsuFeQz0ImAhK
dVAPF1ty0RJkuPi1UXiYLhaP8lPMoCtdZ/LRGoocqc67NRZ2jsA/ku7xQ+kmiUqMKoJ+1Yehqt9m
xhHdCmOJ2lV14cOap0dVs2mG4RA8W++5gRNFNsHuqjeUwalMZNesdnFbnW6SkaktbgZYcEvM/MRR
c3wjG2YXqOJbI+zEaLA65jbEOd5ipLRRWgDH0HFPPgtkNQycl1y62sLKTjENTSQb28Wn+0exT+FC
DFBDD78aIvn3hN53c90/CrGabo2P5KsS79giDFodkDuOpEzTASvQriDKnkdvcABqP0dz+X0pzGnl
Ax9j5365e9gend2TzTWvkVTQJncBf4t7QjvUuhswEey7SgtI3yPskBycK63v6NMTAgTrDwDEJo25
Yzv14H97D2tFK/Mfy0xbHv32lghqmd2rvUpbpy5UUmofDQOsEGHajSob2VVsK5O1NTndtJrbEEJs
II69nk1ltoYj4LgUI+6HyUxFWJmrnvXbAMCGdkdjmtZMHT34LnZ+s/F+6g73od806BwwJuHrR/W5
JhPKc0llwr6g154BhWySRLPTUFmSWITYhQRftQ5a0fX5/ixse3qCXa53q1ZtlOS7SdOpQyogP3wW
A2V6taBGkg2RZ46S74hlLzN/6vh3lc+J5slqR7XiGBhDJbB6pXcCZjt/VEgVUVX6nIH3ECiygYqK
2F+XWbSCtejC0IGo0yeSjjHYKJ98f4qtW3OE/M2DMHdhgBylyRnBUJlB5BTFJm++aGZvf4vw7Fw4
g0Hfsig07dKSJNmgcKdr5IzD3MP5qNgSzD/iJRGuw8FXo7oiO/6N7AZy/AL76SAuE06phmiqeaBW
1nRqPzBjlg7ZtsJWMkJ4GXq0j3T6wWw7QS157iaKVHpQ4XMszOKAUyfpqpB09ccXJCaDRFahOFHx
7YHH7TIGnAchaSPLWXKVNj/UICrym7CQon3+RMwwFEMuKuGDvXhPqPVtZIAqVXvq1KzvilYi2WEP
k2R0z0NXJUr9MEvuPijFvn/W0l4CKzy0buKyjfLTKcGW2bd4yAKLCGQjPOisbAyDWe0Yv8uyGOL5
Z5T+gOyrSs3Sb93+27YSczobdujicYZVcULmabJ/mq35gZOs7ewpPObLh/F17WUbpStYsyOrlHGn
n5Z2dWrg0O4nMoSjsCF88FwHIT4URbCaqdc1UDhJKqrsf/Lhp6xuFLoWo3v9Yj+iZvdOZQR9hGOb
X38RKMr25pyUmrA+OE5uAsgnUZO6KUntzJnMoQO5vhv/6ab7r3CFz+flva2OFTgxmSCQOvtBMbI9
ZiSNfQrdBWsoBn2EUSRO2f9XAa9CiF+tkTeDJeDw6ZjFqyGb75YG7ltNzSEs5euHfe0/Auu4fTFK
HMAG8JSVbxkWLYVELnPNODAagOfDL2l8kjQ6y9yhaUn5PnltDlLnlu8FEzHL1dtzkMHqGQcPsoad
X6KvpgE+UDEtTIF5ZCJ3KeTBDXsLKXOOLIlwuMCQ8KyMC6bxioYZNA69tf68OiGWJXOsTpl/EWVB
Boexn5Zy7qfJA9+VW1G9Jp55EKiH3KHVGFssbyFogMWpHhG13a7r/tvYvzH8bAZ64d/6LQwOVv1C
W+TBdN7h7DPuhe86XA1iyVGWXH31T5tyCB41e1NO9poVO6TjEn40Jbdn9U/UNAV4Luvy7esRm9Wv
htgD0Zm60/6QEaoyy+6S5Hetg62Y7hPzCvN1eTsjXBSKRC2BRrq2v0xYNAs1rB239bRv1+POZyK4
aaClrRD4Qv3Jw3uvDvQr9UNGlk/FBa7L8FtmrsmhFGQdByFOyO2cULxy9LZkNU3HdXZyRqlTikHv
EDmyjIbjaiIV23T2Pq/LQbbKp4jsdB0YqOcAWf0Xd9eu7E4pc0wxTb1ET7daC0fEW/YCXOBH5Cad
P7x2D4shElptz1QPFhfeMsvsXUqiZDKwSj3/nBHqPOmG03U4ui6e6gRSjanreGLYBIg4/YB6EzFH
RhQcVgwh1clrPwhIFusTicV4jcEycKHEMQP31ZGDWUu0JGJ798/ypf+35oOegeXdp6CeOm/VXvlR
RyT0JrfmSY9oah8h7PidDJDqm36Fz+iz3qAbEENYDt1xyTfeAgaWXTux/Bz0fV8pgVQkcwzoNGhC
M718RYEK8MbyXqS3RebXdx1R3kbgzXMkr9sCTho6JRXdVzLAOAtABsVb+OQQTHqrRdnCiL/9QpkI
bxqj+UTqnuDM7bO1VDQ2EZMV2kcKPNVHiU73PIhTshmKNaPzjoYCkLMn4pnUVjLsw/TsCLaM8Z/k
m0cIJ8HNwieui9KPkH/gSjAYiyQlD2r9ZZv/MeqObkiuUeRW89LRWvntMC4Ews+atJo+wig/7iYg
SPS4Bwy4nzV284nHdpho2B2RrDTqSsmf77CDwinp0QEUxCuwAXAdPvCA4I5bM0JZLoS4hFIF1M0r
xBMJYG0uuzQQgJAqWMIaE7cLSgezMPeDjyiya8SFrJaz7/1E7MwDl+MLVPNHXDzT43lhjvNC5ZkO
oV/EvVTOCx10ziSvaFHoYQx0cLDYuIegVgxUbhtZqaBf7/XHdrCNEaCD/Xv839T0qvR5B6ol0r6u
ipEgnK9+iVJZKiFFk0LRUHv1SKF5za3guF5ghiplPXsPure33zPPkoixIktLLmE/bX6YobOalaxf
scdKWpVPC5Xt5OKFpdp833IVZV9xtiDEn5Jk3nsIoKJ7hSjQlo5wBtxiH6/R6QycYZQ8BjN3Df6+
D/xYgOhHa/t/20++M4bJGMD/Qp8mK+1HsLL8cDjx0wW3ORmVdk1+tQWFf0AFGgN/onWf6Zp8cNpz
VRYYg/IJDBvog82mh7wyaRAiIyHXi5N/okxb58WMtJxcUwva69q3DWVmcUcaamoY39tciz9Yl87D
C5G+TpR9KBiY2MmK/w3Hb2aRNB1iOLy462wrJkocDDYzuwqlc+oQ/WcgkTwCZxSi7MZd2UG4PyOb
TBArg08e0d86jrUSxvXMabzOLAvo0Yulwl6z/FMku/ShdgRpPwKl4VYFhecMW//QRVC0jOq5cOij
7i8Jg4bsTD5f+iVYu/0CB27xVjuwqYK6JZqQvgJPk/R+Vl6C93WWs6oBDxRONmwLa98PokVVcTzo
ycZxHxXEB/B0Q+ddx6TKGfGY1OF9MQE0jFck0aPS3zJ+qi75GPFPeegiI5hqv47fju9e88IKIHxb
YPZw2U4Xj59/vgXbS5C47TZcS0cSYDTWtBvskjP7rdOS+wmSJYofnVFo6uLE5lfR1FDZQuOVTteZ
sABwo3hIAHoJg1X9z6XGVf23tz4gIipclnZcj0TAQn/uHe5u8lktarJ+WDQnhtJE0I8Vhmhl79F3
vpr7qIQhXxkVl70RUmxapt4lAtBXDi0fFnm3EhLXVUuGgSo8H6d1cjqyBXl6Syt5RxPcE4BVkWkY
h6SAJod2W2b5f5/4Aem/ZKzKagsQtuCVZnR3V6wM6WCisOGQHpMhZKOMCWRAzQxWwp57r79lP0SF
UEQJlnYC+oFl7OzGmgz+uBpXi9KGP8BjhVBMQswPg6+hLwhdwSgWGBSgfKCKAwiFPw7EmFAy5IME
/jRoLjFLe6h3yFSpCM5xNTnjyGnh7XicbQx+jOaneeAtgKv+m8H5VDeb6OQ5MavjWZ5pVJCdL/w4
ZP2Ny+ed319k537t1wgq8CZ68zK275ySzPYcuB7P9XKbvInuylXKy0WF5EsN5K1ctsLqnComjGCK
BHBl7uoZJgb0d8hn3MTW+7ADQKncULABMBTHL55nMLZnIH1GDPZ5d17O2G4OrMCcr6jcETnk2LbE
HxyzyjDOgoWBSAmaTsDTQ09vF+sYvK5WU3HCgMnGMcg0HNWcJ8tIX4BgH2eI49vUR0TV0mr6nCTN
jmGdvFv7lZDRzO4TiOfoxFtiQtI7XR1numcdHQOx8YVLcWp6zc155YQkMcnxO3nbeWW2aRWwjmlS
EiS5JBg69e132DudRJ0mvOqCZImdQCgjt5FmK1WmRxuUJeHO07ZR7o9RV5HQWziKpPKXD5C5rdWh
ARL/pl2fbQXDcRJfFeg9Mh/2lby1lp0HH/66Jjhs5o/oW2PUnkrVdI9yDZrEWdUM4u0ReR3CihEX
YHTzAYWd5xZiL59znCxzfxXwpFyRJp/PfZi3W/AP9sJ7E/NIH3tYluJPQao05vonDlSWhLYn1n3k
0XpPKLhp/yQWIkngEGvTpdDqhv9sFkFBcOmL4oW+g641lRRgJWuq7i3DPWwVOm5xUV5l0t05UoPp
jpZOXL4GmfJDm2nwyAUWAHw8G+ljoqBgUKq37eibmYnANpL72+xwk4qXSbEHGtS3Rw31byIpm439
kRLY8ELXgt/zClDheTlvap4CKPwsPAewL1vHpG1j5IpXRk6WKSSPokrKsA1eZXvvxDTXBfw2T//m
tE+4aq6ZLTnHdiyyUtkBzYPjqTo1cEJtkd2FMXst+KX1jw50esNLZt0bSQ+x+T5YSjdf+DVLyUU6
WH8a20F0eonvA0ZyieFsRQhHmuvZCZ3bcq2+w9oOKAHsxeTgZcxDt9mbazRz6orQTdKcTyTu8L8e
7gp438XNta3DIVkkrLg+EBLjaUgZ+NUI3vq/+fyRIcWeiSQ36D3G/G2judBKoRiOE7WylrVLoSfi
nkQzOZ5Qld8/kJNjYd6hkE6+N+xJ1uVity2EYQcQbE+FDTwBwRmPqSxW/2PNPUBOpmQSLdLNA5yO
IwGnY5SF7yKWwHtOMxfD42j+0Yf/Rh8tLCrx0UxRKXbQe2VKJSqnAQQIq73ZLCUmMSi4tWakhlvK
qRo7anvf/oGCW+apb6+uKr4UPBxO8TVdrc6OwI+29J0M7c9JZU1F+JR1uNMKDMgqQEve8iQ7SFOJ
IRkFLvkhIfMvKszwx4oT8bWP1ZTywsIRHvrZQCQpgTNOibhVcQKAtm0V14xI2zyp1Rnh3Yc9760F
tr+hf7UBtUYWJAKQ7Zc9278ySsQDqBbpoe6L02p3elXShiA89R4sdBDpB1qtPGmvcSKmGHSFimcC
Voggkm/BzZ/IVCSstm75P0iI3XesjWOZwP2lhwFGvR290bR8X8SB/+wzovCxUTUrSwxZyvkdW3Lq
XMVfUyL082nv9VmWGv3Jxpo/r+Hz/tAGJqQbEH94aYdknq7aDaM5kP5Q5LTlv9wthnZsm66AIE63
81oTKDnUwWR7niXgAbNFpg6k305cJqVujmB6wxBfimX6Az+FYUFAi/dTlvpNRMyEPlaH9wHlNShZ
1acx4JXSA90X1vow1Mdn8QW4wcI5RHJmUSXzhy00XfnRZ65mwj4fAjZPBuUcyHIsBQdw8L5J8LD+
hKC/5FozwIdbpILsRNGMUgFV/LI9Y6dXG+d7iRwPE9OD+uVG91WtA2RWSl4LmGvOEHYheo3BiemA
m8kB18/PNj/Qc3iaj4ecAXSFmf0IkyT/4HgJ/DxUV1hW5MO5MkZlwA1TOwU6vJ2X/rxsF/WYIzRj
ks6nCVucf0AX/SKH3DCFJHDzpf16WffybtDvpYUaQz3f2hq92l2zbjZTgRhLAfUl8y8HmL5JUkb8
KaRMvhMO2cDVSn5kjOkOrLSwljgwF4ZdXOJMAqaNEy7elSz7psyOctvoC6UkCiIk8AzokIokUc4h
VG/SRjw019o3DS6XT72JFmd9ql3YV8BHl5FYtsf9ULNSr3I0xdzOHjPZuEE/BMoe1Hu9JYtfvzaJ
j7QLtI0eck2mMl8fxTOzUQAkcJIjBP5rroNLgAa89+i7AuqFdzqxlhfkac+5cr71A8XCOj1EMV3l
1VhtkbH1/xk2sqKL1GH7mPMpAWkxfDpq6KQXvCClRgKE6VD+ZRawXHVg6ImoZ/1IuYC5AwAf6778
GVgE+ph1cQbzYN4BtdEF/jclt7kNg/hilZcRp2BIECafZIvFvibStvvOgWtoCgyuINZI19iUAGcP
m4gdRTp/fNYPzWWIevg2U+JgJEo9g02PsYs4p2U9toQW6CLgQXWnGIdif/yGR9vlIjsKv1OgSIGA
QU1G4Bg2Tb2soMMWEcakMFFEIA8w9TOPD8MlSvcKPbRq0uecrAgCKOPEPJ4v2RrpIPKfuVmO9Bwv
2VkgfHUQCFR0ldPF2H6VewKDgXAh3spO1v7JKm+Zm8QT0JVokaJI3qffJQrJsX7DWhjKscVliUZn
hZBDXdOXm76xWqQqIPoOtdMULzRujkDd2KMgqeffTUwpKgb6ft3N9ZrBbbmmJgWFdgdOwckD/Gcu
gRAqfXeRMShD99m0t53yNBpM4+Yqr+uamCd4SsiBg1DQSjb7IHjJj6VXdnImo2IYAF3d8R5we2ko
plchz0KpiX5XmIDZyWKo8hMocNyI0cU0FaCgXeCF/XCht/YiOpJRMSH3z7xc1ZIHlDOzVbZmPqET
CMWYzNKWBi+c1NLNu6P3+JJiQejxw0hI0PGpvp+Ukz2ziP6IBtqUw2CiFthsou8gZaGXQGvcA12M
KFK2ZrlXcGnyYW8cOgnFAAgQVl5XXpGnQQq10dfzuKaOCcHoDlkcA0zWIQroTAD1D/+DsuOTZiz8
DCokNLbTF2/oSlWs/uhJ2f0qy8PiJvdqEGRjWJfFHs9mEW0GWtcxnp84IqAlU6peSLsUAlM/Wr6K
N14GdaB0gDZAg0/jLFxIwrBInjriNJGBWJUbEIEboyOIR4n6C1kYZ129fkfRghah/EE0Ho1SXxaz
wm/fuf+L8tLw6sDgkV6wfi9YFI9LDbp15CGyNy1EaO8IhgmHKL4w9Rt9l7A25ZAwtzkOpnviqLJl
9xXWnVSTHyXMCXZHIZCK3NmtjibNrgqQKl5Osl0ZZAAMOZjKvCV3co7grKKod9uEn/uopADDoYsn
0WHIblKFqEAqQZmAhEFygbjDdv90t6poM7UxLFeMyk6JqA6uP2GzVs9IezSCf44ipmITumWC5a3p
RGbkIOpPMOJKn6VP/uF6jDJhT1W1hvwsyIqjxEZnjN2psod1S0OpzPyBbKDjegMVfi+ZDUGtSbkC
Fr52NoUn2nWoz+E/J702UNl/VgWX1+3vQY/1ZlqLfy5G4rvomTNURXHX5pc3i95ChOdlIoZxMX+T
ncm/anN1kIf9EbxIIWXBoV4q9RugaIR0ktUAwnD8VFZjum96pYu61i8+jkTdj+TefmR4/eo0UW9p
Iq3EGhfDXMJ/nn+AyIcCEG1ievwuqEdFv5vwA1gLoiPLYBALWsHBLD6CEIfPPV9LfyQPryz15naA
IpLuC0uxwxyAxEf8eNSayhStWYCyqeaqc65nVwzVteUIoT0aLOhjEuSqwU1d2wldkv3crvhqnLzt
epKjRO+zS16U7Vxh/vvTfIwvQvuVanRhjvheLDErrWGvvGuk4m6oOaGA+OEF604Qg1Y27S5DnqwM
N+7opKYIcPLTNUmCC6YL0JkIHIT5dPwCspofKBP3wTzzZvoSbByNd0k68A75twXe6nUunoDVla8M
TIC9yDgLF/fLZTzm28jhM19ugDnI/A3qKCwQJtt8varnHZc9T5LluG6VWF6YdgbW7mKL8WVVpoSO
1EibARFYraYHJP5zedKLKTxZFMq6JkdgJ6CG9V8o3z2XasehWZMYt4/ApKGzzGGe88djPEnaG7Ss
YLTle0xasoIRwo45Ev3A4WOQyzZdMU4yVU7qev245digqtmRD1nkpdvlnSmRvZi8whtghK4z+DHh
vGVsg1fgxrxHsx+DiI5Lak9C3C+4hSI2podrpH5HIu5XE7qAgHWbfUjjWhVfV8c2T7zAm/aYuTAC
v6muRvXlmrtEAfYTD4OpQkmwE/PMJNRQPrK7zKf/F6J4DTaY2EQ3sF6oowSBcQabHxoURe4I+OCU
MpZaq8iXHOZkYJTk1AafTNAv0WB9CxzoDkj6fbWAF32JJhRarTeiR2iqWEDqNG0yZFueYHH6/rWF
pcxcaHxCFGHA4ipZpy2wr9tGwzBya3unX/b0AEaNECQwARzW+OhXMUbICnnjy5I2MV/TD95sFnxk
bQCA95LwSnc6C22Ib0nF/A1SXJJbulLyNHZCZedkrbSlLsPm/OlerwqjYfO3XVXmdzG4Zf7jqf/I
M+hJPQO5BkyGX31HI1ntymoHcyxj3vDqjcFkuj8CwOfho8reOswHJz0lyW/1SGnHY4fJT0LKh2xR
uepA7FQdaELdsoKzXxMtz4N2J3j7OZqEXRnY7kVHr5I40znMGe3u2XDP5ytBRQPKGD3P/EJYhp/0
bOmLdIcIbu1huaCODihWp8k/fVv1Ce0IHej6umxkaRteBfy1ZpYuVCS7ds38RDz5BQo88luwxyEA
YkCeGzK7EbRymoTwN7d2oMzr/a/o8/r3Gv8qNSg62nWGheveJy9rCvhmpbjx7eUdXEiwaDz7+uyC
EVl2m5kyuFhzqGKRtDjkWvMxlBdAbcJ0tWMBjJ0k3pCo8jZf4yIF+GF1y2PkAkZ3t/ZtbFlRxN48
rdY3iVd2JbeOymB4oXHpgXi3f3uou67++HhSMPhGvNsvD+4UE0n4F+bNcQ/SF2W3Se0XiBVEuRh/
ekv51IUTXhm+IEq97EIrUvR+dkcBm61yj7ssk91OqKe4yMQm1IvAV9gRpdb2I0IkuOm1bbvO/K6Z
U0SVwD9RnT2Pw2gABJyxlqWTxZn22NfKDikntRhGEEmGtnqD56bZW70/PaUU8ImwXqyxV1JX1ylg
FNumtUWDvb6kwquQDNMK3mJGkthcRdcg9a2f3Ne/6zQ9d1wgoxuMJ9JijRelWGZ7W8GH+kiUvFgI
hU6sHUsvIu87Jp7o2wi+tRYGQYo71t8e3x+FhklsL8iaDWSF2q4XQE0yC7loaDoHsB0gvu6Cyi8q
352HNY81yWFrmbvdjhr1WL9VNHnZml9NkZcRngvhXRZWk5U58QNDLLgwR4LPgD2twWOnN3/pqBTo
TJX7stEnyvN08TLpIMYrebvHhYLVO8lO4jCEgBBkY2AEeldcbYBD0klzuZyaOfFs99cP//NSnEaR
YZUf6mwqwkg0x/TZMMU2kiqP6Gk/dlwIvxcOvk+k7emvL40OytYmVLBnfjG+H7CSJTB0wekptXnA
5R1veo7V1jUw75HD+s+/R4iWKl4MmNAIZbifZHDfzkGcpWSQOog8zfkUkOJ7ro99Pq2adRtxFH05
2XucTCOiRjG7D0cPO57qSY4Tk16bgl1Kkrf6E3+BGbDzNZwpr1/K6KCTKRqTOST/hQpBZw5iT1tb
8Dy35BTlsyjM0oHHpK9NmC3Xw/D6eOIaO+hi5OtLIIpKURw9mNg+flCE/vGs0NR3DGi52jmNjHDS
aq27griA2EBnHc5wyUDyFaxahxTvGHxKnvLN1pK9OoWzNTaPLLocypp1OyTW4tQe/6+Nfa+pAbQK
2AROy4yzHvHO/ZzVHyJIDG0Yo0P16RwUqVcE/0gpuNUuiFKTaImHXSuSxwlpDJ44lAJUe8HoytW8
h1MNC036ygQGXX21oC09IrAhy336zJVlMwn3PW61CCK9tbd8Sn3+BoDOZorHTTlBJ5yvaL8tppPW
tz3CiuaDZVDjM5BZcRsCUP6C1RdfN204T60cIsyKH71X1hQh5Z/UwFJpVtDOEmCyLjwIoACIFK59
ohaiNLGSFiVOEAeo9umbMIs9Ak83D1Tjt3DhOTBJcAbLUuEUz0iYSPs0oCbS098l3xj5L/NLf1OO
LYvj4VaQlUPCqhBgu1OKf4YD2mA93Bt+DanTH7TSNwKYSLkAmBXQPmypAlh2/YDkoYNuZNPPoNY2
pOxTRrnxrzbOmnjOaP1rxG8M65Kh6A57h9eFZCIDi9RzhsZuDruP1XoPdxEL/Fd4I/Ctj5r9Uqof
p5Ia+NzpLCqUskX7cIhpk58ORwoXBvV8XNVHzWbIY5Zn1dFZ7MjlXft93PfWnhjFutm60mYJEE90
XSnW6QG0oNWT4kRACCk7gvLtOAQ2UHvHVEhDogittI4xrd3QTcpoi1tMUt6q4pBfv8S265VRQt6h
Sqy1ej95GvmuLPTffw4fSkzqSyYPXF+do0mozb8X52P/xMumzApmPf535idh2EfWJMe8LPlcE129
SfS5dNEq3u+2ur+2mhYSU5ydShT2uF8s6XlLRLMZgRWDh+FHOOfH3H3M6lla0cB+0zgfhHRAGuZM
42Ei7uF3EJuT6/sZTVpwkPZTYUBPhHw+9k32I3qTSduW8oYCt/j+jnCNIB1HLC5C1//MENmtaop/
UzplWrU65JkPAIRp5WzHpwGNdb5lil0gO8EdiZXO51HnGOB89yrxSCtXT1al7aJnVScWjF94uc6W
Zxvi9K1UtqnYSYq7IdlXnlA/ZbzrR218aBl/RaaRNFMeejy/fPeupp7WapLkFMzZ0WldZun3A3MN
Z7OW/jGmGtr5r6jdQEhMdrDGG8oce/eh/c5yNXRvEAGgNT+zkdeQLA+bBpxt65sCkxpPx6odF1Ws
kN5mUIb360CboxFNcgvd4KHomdlus1+A33Rz8yAiki39O3JlWBrdJ6D2z1+8HvDIcxOulEk1Ii08
J+CWllCAQTie09OslT4TiAqirLw/sDEumoycGSjGdVvWn9AmVfvp1cugzdtuG2PDLCOSg8SlSq/U
DmWVtgH45MY/AuvUUWh174gsiXeVlupuPkP4mMPGapfwQG7/Sw5NQze1hB4ezQuecGUFMv0aECkM
a7NCmvbcmR9CzXMFNm7njQMjekttCpv27giG7rW07WaDvJqDxfzEit2NZg+5WB0rtQiCLSJOz30o
iGBvGvMHkGPqSvR+o949mPUV6WLKGvfwXkiuiDFERMFD5ROeBhYOzHDcKIZCPcuWOoBL5Gybrezs
Jsh8dAZnm1nN2ZDDgoNZSkEHuIy5jOySkAtucC9d5MvNrfPPfF3HMEggyTrjL878yrs1ZAqTyzFz
NH40YxkELPfO/fYXwXvcqkW6K6HVt/jXq00ws9CusnowoLsX6jSL+Q4ZhoiNZoZbq9ZHBBAi23wZ
Pp5fm1iQFFftP1E64whnSZJ51ZNeasHRo4JWjRRmIVw+0TC+cdZHzDBIypcGJU5Szf66KRFq/YC3
W0qrGpNeIj/kP58h7eRDgAYMPOlV0jUQM5s2iySNqESLRwBOyG/65Gti6ZKbO2Ry8nJC9rfT70Ef
RnZ7zvw2zGcv1nJ4MFgaexUB7xhuOdE5QYCAY0GsNGBSumBt93tkSoSwyAw2mNvzSyvnoNxZimoc
p/FA13cuUHoN7j6tKqZVYND/AF18+ltli7DYr+NSZdBEWZhbY1SRV69lsSvrxCMHmsOYXvzYrfKm
AE121KCXaL9SL9415ctJuINu3e7yefkCfXnCJWKrs53NKFeab0cuCaP5fLHy7O0ZLqRoyyrOn3WV
SAIaaaxnXd9NyVj8DJWb3mIfCXgJ9higXftcDrJbQ3gW2J0NAhh/bAqUutnYbtCGe6zO0Tulk1Gt
HvrLQQaxwJOKorByjCc34gPLLZDq+17zftq9LwYldDjbCBnoteKaslD9qH07eaHuKXHvqzySut/r
e3sZndAkHlfp04RrylscDXvrYFKKBdWhVVlJMIF+4WsNBosBIAfN2NRSyEHD0/D1HytSORGEpQVh
OshSqRgTnvzPRurcYIMoXHanupstc/3BGhyCmm83yuPyHWao3Ftr4iSY+nLX+/pd2FG3dHoxMU69
JGCMxrFqm1igLWWIbhqjKuhslOsJ7nLDbpZOsRETcqgt4D8nwYnfdcEgRYVtbn9odbalPhcsDQzk
+Xeu/M6DFXoCFPZGAw/Yvj8eLKlUp1pC1L22RCq79BsfNEB1D1Maqm31aY1ZiPzfzCkvA5Dvire2
9vu/xajLY7YfFAbOfnkMeIICes8SQmteQ8s1YKfk0FbpKrC0VRVB0xdf2hM/1Dje1aTDnsRi6Ryw
oh6+uV9iEZO2svxX/2KPugAcWLrBiYkZd435H9FbD82VkX5G7ECQnCAf8w+xAODIxBSe19Vmy22Y
Mk173Lybqb2xLStoj42NPHCmYj7IsnEKb1aSAO/wKofBRBraRhNP+cSwNBxmQVEtJR0oUzOO+IKY
1nJNkItJsNDXwmPtXiLli2I2jDf+Rcod0mVd5s7EDoh+fREa5tpe7dXzF25mET2OARHeq/0pStXk
KCqpuAidkEElL3Lm/qX6s1I/FIY8yXxWIsDr+8mUS4b1Xp5meaHBQF61wSryKg8wK6zby8BiWPT3
ChBkSkTiY/iU6Zg0qo263/FkEvV0FNk3K8/XHOxvzutfAwaDSheqje4YBxIt2Zz3MPa314J75/Qc
zibOZgEBBCKcd0vshPnkM47/2ZD0spra4qYR66QGOcrmZAen0kCHEDYq+K430uyfqllMQMLxEwHd
CCYJzrbQeZIz5tPJdKSpYBAHyh6RpqFjOIgJju0qi6iDuBTFUB8lf5htP05WLJpQbUuSqY8S2jMI
17nefDKxjMdEcLexmJ3vvInlL008NL/znIg1gpFnotXHoSYVkEUL9/g6Dl9XFTrPRW50hYjtRwO7
8yBIj9l0PFm7//MFS1zvR3+YA3jrNDztfgo4zd0DFwNszv3kvZYNQuJbYFms3YLjtpL+KAt4TF6d
90iqxYo6sSdjv1aEeqZF5jdcod2jwjrmPjLBaDGG5izNNQiZTAuFUxYh413eVl8EqUqJTFan5N0m
QgM294wtu0XAxbyB3nkLTbH4ldF8x/YNerHb0WUN0JQ0EhgpcB9sqoeb2nM2aHJfq/hIs/OxVg19
ThPPwdzxihN6k72fbk45xDoANeQCuhFABbRQZaDgPVJoptrvlYrqk/a3GLS6PYqI9TWgPvvKvUX4
MBsGOxoGyXDpM4e7Rj6nYayW7Kg6lCz1g27eM0capRwZwhq18CE9y3yS7IHYRL7fdjkQfk3PQT/H
r5W2ywtxaLQqUsxom0UotOHXrj/BMCzSuR/Xoo1RWOZVg/1m0EIymiLMgMiwv7QtqRYh1EBx5I9m
NaAJXi7UN7eEE5Wp9qM8dV1TKTju5opBvhzyup3JB3g2CGnWpqujtv9ORRN72dFlmtrO2cbazUu7
VWqIYtxHtEDDS2UNq3ZDXZXb2b5QyKrQ7h4Rbp5Hpr/4KiMivmblzb9f8vdKgjk+fVkrsXizespN
deMO7Fwo38/RelLN8QOlaRcPzZddqsYXix3ckDrFJ0YhgE6KjuzFq7Erg/XissseOeUCE5n7aPGZ
T9clS0W2+FmJB3Wg+UblxQVMFMaUiGV6OEXsSSh2Tx/t2AV+ZMhQ3P5cyMZM+e6znEfNizq96c/C
/0zxdkJoNIGyvJyN9WvXgu9Hr8UHL4fwkCwhaeIhzkxaLjPl9Jh+CYM1TwF8V+CDmCA5G8b1vrwz
jP689K5at0FWdCPt4WNCZrkqnLFymFwFbpHVyacmPQ+cUThCwZSNdL3gidWIZ8k0NnxT2+iInEun
dlbk5dZHmvRfyp9fF4KpW4KWz4gc7shyIedBfC1Fof7S0qD+WDjaSrBNWFRHaUrUglAup5sTPydE
LYxGwCgy+tSUdu9s7h9MkE7q/5xFq+RZpgRWSXE9PvDhh6Zhdp6tfmMpNG8RR9DchIRoj+4As9WS
EBH6YTfZ20w7DRPMGywqLggXuy3EsFTrufawhgg5mFRFU96OHm6cHu3eJxCQioQuxygYGeJD4xES
bvuoQa9CBMLHZBCQ3rIU5rbzvjknBVhJE5Rldv+9Qxh7eO2Jz+ie2Iw3dpHeDyEndg8hp8rTDnIP
/v32HQUGmFeIjL4Bvb3s+KI5UMptWDSE44k5tQJ7oU+cRwF+qG+FYOGpqem2CWv/rE4xIvaYGZTw
z+tX3kTFQTd4XvHb1QcKsg4lD8ajIJpSJhHkyHCO7MauJSXkwwbkMPq8h3MiX5wReYCJ8MeJw0pg
2Gz58YSRAIeJ/DQ4JxFYMY3KpAVplVhI07j1RXRcpts8ylAn5Izo97UMsWOQmIDECk9xnRmhSkTe
0/b9XLDfAFf49HQjFSYqqady37aqNXwxTWPZsNCCtbc560j19/rD/wO+cx+2fFblzlhFdKs6fKQu
oDaMevKa6Ey//w8geo9EOZCva0fumhklGwP3CnwdDkfBtiNZsu20U/DkZbj+B3LQCEYZUuOt5YtC
1dxZX4+NOTVLZob19cI9rU+DroOSt6M5c7aacWn9Giy6o8dc5PlSkHlLu+WhTT3T5Tsx9T4qTip3
iVqlyzzxL0p+VnXHJTBG2TUHlT+dlCRDKUxerpSeVsJRqhG47ByZJTbqUqyjJzotJBrQKCYJ0BxG
SAkaa5q8aiPUOPmax21PR4E8PX0dV5+YnkGoGcZTxKSbyXQO+gv7VvsURmCyjPZUCE/TWfY+eJyl
m2JpO0uM8a+Dt6TN/Cd3kk0+j2NHa+fDBv7fPc3WXzYuxFb5wEFRd3qoO3uCU7xafG8yxZMWy14W
c799f3Z9E0/TIAe94t72a2V3/TnaK2etRJRVSycpH0Sklpixy00gZNPsG6zU+KafoFsjg/58dhZd
GFcpp837uLYr6xYVifFG0bYhGtH2Hjh1FHXhyLe34jHRrOkQ9kra+Q+2C46Bo0t0Xp/QYvx3d7d9
/4TKxopmNhZp++YCb3w8PIMaCF3oxOT/FbZz0e4gjT2B5DdK+p0R6yYTcX/OTLlm2pDviCX33U/m
nKj/ojwZyppANLlySWfdjPe0li7ichPzZWcbAJ+fxeXCdjLqhTPVv94Kq2kYtbjTIyUu5w6Hp2jL
h+LOZLTiIh+MTwzSfsKPcGhxUPXB8sRr5Mz877/cuC2iq8pMXl2NenuX8uUs+GQvZ/WYmSKvoDRe
oioQlu5xuwUonf9Gj6s08sd52eqfjRJDdAVSCvSQZ7AmTPnARE3oxYrGi47Iq1Hp5tun7gFry8pN
EIAzDQmKtaRZ1f5hVqxud8wgcm9QzibMvQ4kzPTc5nwEg1bKfxCKVLl8tqBrW/pmkDIul4Fxz8fE
5vpgTExRqjT2SgGHfT5swix3uqFqeHBaFiWPBdTYPMU3OGEc5o4m8QMLEOAJ603jVaMlcYfKQJHz
/26F0MjCxa+D0crc28zbeh9/ioxIFPgw2U66nownSh0CjfF24wocVfGY6H3SHW2aasKQTQyGteQf
0Ue2kuzrVXchX2SpqTTiPpz9GrUqOD/KxuJbH80fXjqUreXkG8FP4emm2YDDqORoRUQjK0rFjqAx
B/L5KKmx+i5L6gaf/YtAEwL5vHmQab8bD34y6HMnLHDJm23hGsyYG+hZPsrw17UBh1oOeE3Mw+iH
bc26h8pFA7UNdKShlNKVATVPhEi1/nkAYSSH76MEJh8TBuRp3QI+1bkQRgwqrJHy0wKPWQK3LGzo
xuhme7kfK8w/FeWcoVW6dxHJFjVw+TyJcnFNXA+3lg6vhEk8s1bhE3HOVzZx73vdrnmT/+6MXVRu
chU8tbxsRsWjNrjM2gqRSilPigHG03lf9l1MpNneVXDOFwNDu6bL7AIHk1bxc9kUqgkyNtsq4yi2
XLJ47XEcUSwzEkZv2zVTmaKHrkAZWNcmuL+n1HWFxilW/J0yBeSKNVmkdzMEK2kscMWwx1gJg8j5
Wq3kTp60FJkqxPNyw3JYb17RBNBF5wKR4M7I1gM3tb3AKKVeQKnYV5pSAsX+INsrR9F1gydCZyQ/
83nv3Cq0Mmvy+qJsaVzOVLDMJi5RuBr+3KD5ZYmr0XjHC4SRxx2CeHLYYk+FuBeWHhCPnerL8qhI
DFIsOvgFjUe/0o9xNPSWKKBBz/gcuYwp+WTyMhe200V72q4rQD37+hxpngzmOpAJVd2doIGLRhW5
sFY3bdsFTdGFR9m3P4/FI2buK5AIhc4Ey+ag01N8h3FNYEWIOQ8yrRqpmhi0ffCzRQ4oJ/VKRuLf
VWUUatrCePqHsKGM2ymiBE+cAFpdkMsuCrTGkLHXZr1TrMvxJtbyfhelX0Gc8SsEC9gP5uYHN18O
4ox3EH5v4FU1OVoRAY0S+SYLTRqHW92X1dY+6tEMGgNATEg7m1+PH6AkiPCTETuP08xP5ZooG6Iw
h7Az+WDLNr8xUgybREF77neS8Nizxg+DXOHtA6xfQ6FpxsTnKihQqTGazo04iXnJK9pXO1c/q2zF
Equ7SP2w9jJWLk8d/kUjouE0Dr0DUderG7RSdBw/HYOa5N361pbxYBigMsfJh/mYTWmdWPLRLmmr
KFRc30hwuFqQTF3SLC10TshE2bdWhiNeqgSThjLkiRjgVDTgn60JMWbi57yA/NCYhGEGlL7ZAN+O
NlfUn9Yv6f62y/lvJwiVACu4DUbZX8fOgxdf61H7cWpR6rvJerYpvqS+hOg6ZrYZ4ER5mhxfMmFY
/jH7glQYRlC0deoCfG8q7hkeoJ6hlVAUc1xjTEwZ69GYT1d8Fa3PoHrDxGM2kAC1IxEWLthuYkRq
HWEDehFp/ynHIEL8G73DU18L2Ad6dZ4UPPH8ULmbrtZpFPGQ8fczGjQYBmZ6J1/ihbciKx6uV0WY
Gz5kXucFdRSpSb73BBHM1zMao4sATP4rKLemnfT+VNm9fmxkNa8I/y7saUCYrswqqqcxmDSICIou
Q1LtBjj9V45i33DdzxpcssHEvAIxEBp+wA6irRZLPyBVpczx1xa7TafuEeuxGy1hR+MlTRrWJupe
rvdUJyFQ+HtN18n0dQkNGMzM0A25Oy8x8dwPZxXnk7rOYjyoVloqheq4WITygW++FX3IRgPT6ycO
cRLUrqG5JjMBup8LLKEC9OmgM8GYzFINvzaoHRYAb5GxgwCuE8ldccjEL9ar+5s8opVqjIp3r+Mu
5ZiRd3pE7VggnG/Wnh5/wIa5OoBQS34z2O07G5/fIJgNtVjhqEJfBxJmB6RRHgPnDQZbquHKprit
f1nL4SeyMoWa8ksTF/I2XITH0pHtEst62Qd/0swJquVer5vPWpCYn0ra53igunsulFTae3nd30Xq
lkq0CmyUarjegZBiyrum5n4Lbb07giP07hw1hn6ILPj+jBDPTwUkgiLtRptGR7B8+PkryJvPNpzp
UCSv1JibsVS0FQhs9cPW8Vm7JESb5xCXgkOlShnArci0fNcLLtp4kPOCdCp30xpDF1EtYUSyiTS2
ySsn7pEueMnfp+FpgK0MZwL6SQ2TyybgRcKg6mlM0PlXyGxBPKr4Me3m/ixhBbQCGdUuiV08prEw
fgwW3BX0pRPoyfpsXN2Q2BeGu2I0tcr8gCEZgPhJMfMoJuX07AOPCli8u/HogSquSd8VQTWquJ/K
SL1zzoAYLm3+K7DXkVZXcABHjdpsdkWSBihpCPqk283j1Tt/Q+DFHVME9HiVSqjBG3WL21cDAfpx
xEnEN9VahV3rK13en/LeehJNM9ROU1DvMRmnLZ93bSX6iGQIXkjbo+YF967IFV/DOrvGHfXZanG1
lbtmze2/uIbBcz0lxP4vZ9TAgVLC6ZvoLoCDtrXcexbAzhJ3z4IsjU3YfqipfZQ4rLie+vyIk6T7
VPjbP+46a0/tkBTEUV5m+igvB5jyfxznwaRJOMQlYavmYxvp6/TDKCyioek+bjemXea5GMBR0SLc
AmECMOfWS6KXZOqle9KCCQJAI+nXIcGSKcbiJkNqdnodjYRLMgufB78kIFPhNm4s2IwNcd2hw+u0
7PoO/s3OTqSG29akJ0GPNIZdaMRw/QK6dcV9YNNYA8+nksC2Ic8GOZiHukcz5QnMwetN1pxEd39U
IOfaxkXc+fvTYRn4vMr9MtWRLEW4nKzU+hDH2ip6HFfxHVlq+S4pQdpHkQIuGqmwGLJIOUECFVdz
2vuP6s6YzpevQ+Tmx+QC+eUmWIz2GsFTKdRDRxHkD5sCjj32dUFArvWexVYKeF628CHHngpTmKt/
9eFu9XXnyAVekPQqk7iEhP2S0AIX+hCqLsAKB5SOsnDwNWQzA8zSaC+GEAKcljD+FCDUdr6U8UeI
NcN9B/Q+gxD3nuljEFet68Dq3K5Y4gjiRgAxeZeGeGgEiprplmLCJe4AE3EhQ6XZ++I72mwADTmo
GdhY741KQsIEfO3kOxS7o7Mry1JQl5Koiia2dJn4C6eTInrMuGa7pcTQQ15XyeTZNqTD2XLloq1I
mynFCogsmmsRmgKz0lV91qEC6VrtOLwpcr/YEckcqUjxOh/0TGuFE5EDLLUMtcWcAHcaOuiTmjn6
2eoOZGQWO5j/KbukHE/GGQ0ZpywYAriaSZuQyWFicAOesaXFcIWH9o8e2pabmjJPiDk0dVgRQ25B
buoaJlxwYlW5DVCOxApjgY4aEp0J0vDKoGCrgZxGa07nRMEU+t59obJuN/PyfDLDMxaxKbQ+ypWT
+6/oohYlw0GTErt680b6/KZsE/VkrNgbc1UP48MT1sKFqcanjLrySwCmm2D1I6Smr23duG3skaPG
4hq+23KquX2DWUG5BQP2l0XUPQ6EURuansMhm37zFVs8Bd7cImUVz911hxcJKf9n9/05rDXwNXBm
jKGWHXZdw8nGwPH2gpuQtdI/BdYuFSCi/bySPL0n8yK4I/U7g0Ar+Mly1WOn7TeGPSLXGkyQUng8
BkdCoDVMK+RK3/G360DJl/P/0lQvL6M9rsaZ/Sb8GYAl1QHgcReYGr1u6lwhjyMmMLoxkLgdqLrI
Gjlj7EFlfnCXlTRHU4F9sxhXlfaKpCq9v3tsiIbV4THVWovjIA+wOKBbjQJD826Sh6mKb80EEWZ+
jDZq9qGJN8SqAQbH9lR0aoSdxyqA/UM6fRlURFA2RnPqulBsLvttVtSlUPJ2newx2lFgFa/5MTuv
3V/FuLhno89DNWajeZ72h38d69GQK1ayDNswQ+oBQrFuXrUgQ3ulQdGp1fDVWZvj97hxH67apuSv
1meaDySc4LPsv+hJ6cg2IEtdF09daQOK631O7wiek+oZ0MlA51kINcT46+nvRzl/kqOtmX+i5dFz
pqK4JAvsuJOT+SVhmXu7zTnOfsKeU7qelJVW8tZ172fytYFBSinRkSfHzEVO7F63FIJSLyyxXWJq
pX6Y08p8P2xesO11BA92+7wm5l5NFk3BzKt3wyUrb2pWTzKpMmFvUK0VWyAlqTojCzCibGRfobym
cmEOyPZIdFXmb/RlsIMdnFHIpVh2PfrSpMkBRGC5Ft9b7cbUWpLmTpwMp5+gLevjAmB93miichmz
3tUrN9Xf3lzBefSLH/z8HoqzhERCKShltfMKwes1wdTW++jq/1MzmD7Ugx+w/wnol8oFVYqXWPSN
1UjTMvKveOefslBdPa3tdLLSZmI1KIPOUjviTZJWwKIPzRmYcH8VekwECvQ3wWHVEbocAPlqVFq+
GInijiakXN84y0riDewKFv9hADLkpMjC2mDtxo8EL8d7EGd8N8qmY6YHKOTZtxLJdZAab5fOad1a
/xi61+6xZ4Kf16LFsfccJpdLcUOJxzhYcUHFoNUQuvOJkNXlrrNvmIcRWcIWcavQIFwBdPF/Whue
lZTmnsG8VGFdGFH6z+OTi7tIan4djOFcYU0wkbJxLaQ0Nm7ziG7uUdLF5oF1NjM0Xkl4jSKvehLz
saFs6dB8Jtjtu26u2ywWYQ0OHY2MzFeRETPyGzUeyPQ+BaexdekncDmi76+n/FBFDN0yloTbKTsV
wwCdASZYARl+pAMgjARpzEsleQ/OdvperwuwWdYTela8434UBSlyIGafIwoQM0G0lnBR0FpzdZ3v
dXlVCH0xFt0fFQKgRXtlLgZCDKYNv8AWlJc5i6sHyeGOXy6n8BOFtqQnA7d5RTOuE/qbOlLcaN9j
K8h1Zcp2aZaCa/Ze8Bp6cZqy2ysUNWm0UGW6rzpd4RBX9pTX6EYgYC5GWX4SG3pTKYUgtq8ZIjZy
1wKmV1ioDn7LeiOhS5rFNyJmpp/YlaB8JOprOYyjrsjz1o2GH9iKFwqnyTjUk396qRB/86A4aTzU
ZHLrOLCaLU6mrFdSTmV0txXJQSNhqG7Y+BoPftwGGfJzAtWynSyAwWWbJ898VlNTSIZNrfbl5ti3
TWTvuYpkqup/7wze+tJzr5vHESC1gPyAjBqQOpH5lJ8yhTiAioEcPzSjlTNocD9Q42WDNxMRECoY
IaFGIDSEi5nYe+D7PWaoLz/+IUGqgJTnW8kTIfg/Bc3WDncfm5C6ZHlyhFQ1jfFXzORGvVaxPays
mtiejA6GZxUQbTLJgZ+dvX7QvstPMeT/h0zKyKt5NlJ1NrX5m4cTzavaOudc5nlCyk7kkEu+cY71
hcHXAe9YF4DKhCQogh5IjprNY+o+8Y6P+o7KbrOSsyx55KnPkcMEZOZqsli2h3YGTVNbm+K3g67G
MiHBtQSWB6/ocvU4wq8XVls7oLIRhJDQdeQFh8fzCAy77dxHiyfTL3zKkA6goSzBT30kgUEot5sD
EOr1qz295BOp0y69LvC9RcNoopWhq/YDtHQTIqbLhhWE2WafEc9PGsa+wrO7PyB78Zi8b7jB3d2j
PIArG/xh0+9VOvF65EjesJSdK8GWvy38mBu+MY7CDi55pJPFvDm70EMhlQiE06bDLCusg9YQv7w2
+hpuxP/Xs5G+gP0lY0w4VD/rxXDvDkz+pv1er9cYjBTh+LL0sEDMbl3nNQfvh+a/XbYNWSsm2g0y
Ho+tnJP5ZWNxLui9qGN9WODkUyxa6NyaXwUklqaip7btwXrf+P6PjROUUM6bw+ze64kiwUBZL+03
zZZ0nFVM2L44VvbSiMT0uu4azkPW+Hs/xBDn9517XHaDABEgE3PNAA5uBpyuy/+q9Czfun7pBOT/
zuaTTDpHGbwCCtzZvABu/r+NI0qjFX42TV+nzTCqlxILQGsYhhAUS9PVLVh86nRaRkbEpa06ck96
U2lfbVaeFmQbkpiye/c4l1l+gknI01ZnDXctdzZ0U03VQxJUZblBUruT0JN9XswrOFLU6kDJFBQK
0vfAIUdIBisjsp2VejCEcAwXFL05i/eMYVytaT51aSvhn7aUbD1Ww5HvfIffH7ZaKmQ1vqqijVsD
XbothUhZTLMHSCdN2Fjd9BuRblyuPRSM1IFmcTbgjXBIjrDIukYXjsJR5RP+VrAjUDw4HYwDqXt/
W5HMCNdJOfXLBiHkrYclBF54cFSxQaVqvOnXzrHAytMM+qwvYiNHL5HI99LKcFX5bc4rkzpV2HpM
IEkfcOyTyZ1IBZTFFcsdY5gWZe5BiATxld8yHRFUTYKowK1VrGFb9IVIMqvcVAGeWWuefJcXvRhD
ERdgWW5Nd9gyCSCRH52A7FBxllKnqG9hJOe8mI/MoaLv6GgiR6cDx164/q2gJR609qeEYWWRHHHm
O/5q8B79UMF6CczkdWtBymjUIxhd4xuCPykmRR6F8pzhjj5XlMHc2olqsZPdX8N95rFiUGJUISL7
n941Fefj9GRuuhDAeqPLX1C+c6QxAXA3WK+ejwLgCzF/IieH9+O2Onr5MNK0JRsMrs1o5RqUbQwc
9Kooe26ozcjfaSSGO8mxgbSe/dZD5my7aoTTB+bqmd0ZZX8Yzo5XEYzrEp3df7FNrz5+bnc/nAMO
VR81P6yM2/64LWOuoHiNscCLVs69ugC9PXulVmYX93Fk+QYKdoVTr/q4llkq6wSonnnvWFSqJ+SY
DLN2QLMvrzcY2L6pkfxrPAkAc2XEJOXvXcrSLrNmrf66Miu90pCbrbvNfD4ygEKvmX8gpjVz2fku
yT2XFBN115pfhFTIlYZzAjxFyBlXuiOAtmE7pzI8ktRL3a6o5RjKT5c7Ue+Q/BRBkOSt4U0byLMA
S2F90kUNIdh3eYsWPu8BgLbTLdXDPvwetxGNCShM+7Ctxm7l6AMRfjhL6wfieWtVvfCeJu4jj3UJ
xPJUIEtwrarcLkyvzYF7wPHLf6KnTYEITnC7KeWdXhHOwQse96B4wqnEve0qrfwd1T31koWx/ScJ
EPtWFOEhxQaV+QdRAtlZ0wuqfpavNttQStm3sEUedACxIGLMj4pU7aoFPP3Vn6kGsSYKyfoqdceH
sSYzKDby0l4DbKzOKMH0MxtkCEwIyhzN2DbYC5LiUj5u5aGgX0avVg27JRYai1groSsd6Vf/x+1f
SeEXEd+79QPoesR867VEOIZ6skSQ9WYMK5/ootD4i0F+9NeK4RQTd4LaqdaL0rH52zVfNta7GCUy
gr707qGZ41nAV1Tv0mcAWUwD5cRFAF5UyG/u9TxLPafTs9eTbFuUt2yHttV1kUzuwzoRM3qYIx2D
2QM6H5LXmMts6xsdWvwjpJCF6Tna/De5hSkqfCqpDvT6z+zK+q5DFHFaPCyiS7TFppc9e3TxQZ84
mswnGXb+gLAg4X877uLXjHIrbvMhL6JJKNNwly4toZaC7YRu0dLPGJ0wL5dhV+Rb4COQpAe4efmo
iBj4vXBPiQVFA/Ii8w9s5Xt0Xk7a9OdkQ/AqudMeS7h+fKYBoSCopkFn3ApU/v8GVt733t6CtXkX
WmQxxoJ3VLlxPLxzNa9xPlhEoN+hyJUlofYY5tyo2WtEs9s0d996v2WOk6jxI+UyDk0zSi24XvHR
MNK3Kk6j2C/oYlRnzp8F2LXLbLD2Jv53+yeg4z5UBGodMjPEVRtTTxKdXUEalEd6mAxVsPLnnTpM
PhvSeG7orKkbc87dmsHCYIDHE+Jq/JpkMoOlil2JZJ4CfAvX0163a1LSYufvlXZh4AN4u6S2ePBm
cUZ2Q2vC9DIvS2daun/AhafIQA2miq1a7EHKYkL8EhEfc4eRtJ+1lEDuj75TKdbCUSqCMGPN7Hfw
EepsOyP3EwdMz1OntzVewVaYlhtLMekjyZFIxoK3PyLn/VincGPV0+ZPWMT9hcKIwls0nQnGiF20
lCKaK8kqak+UshrU33Z5kAqmCrU2Dw9Jmr8UE7PplguC/524SgXcDqLZzPTO/ZaDoLn1u+bdH4O4
X9uoVLLFD3DzEiN7BBiukJD0Q71uEoWlW5RRIMcxXk57IyrcvMD9cD/GU+LGdLQhOqjXEfOODLC+
yrpTy5oPXVwhj7xiQR+0FZz/6NEi1UZdo6jgbIOoWdXbNiG0Ff+9CsTJkr7FtOipuwRHbkKnnKJL
DSQ9n3+pM7uesJhBYCRk2A0m01rrchyLBZNFQPfTNRTLx+n0GV3PTrvZpvSr4XuzvgZltcpCfLkF
Ia3DNge1fZvmNP3z0Gz4DQZZI7jbfVeF4NUiVHQYprQt16nNTqCNdDspPfdZ0/kVFNCtKyOITgV/
mV8UoeFuCipKu7rzj4N5PQQTcm7CC/tM4oa4gWFsbiQa0pCCEhzjLaTGHgpVHPiLFqWJ4Td1R2mb
UwfD8Xn18EIGmir5Ty0j93CwsS4k7WV0IEX9a87I0fYjZgK87PId3YAlEmyuXEVghVORG3YDoy5Z
shTM7DHKNjPNAzstRTKfbUDalv7KlrgWhLtdHUpe5Xac6Mh6O+U/4NQ40kP+JlyZ66DBMQOi4eXF
UsJDsmL3MSiiSrpEE+AFHucsTFNwQA9HSE9B6boDbSVNIL+P+P+YaUL/qLfK5N3x+9SoaeIhEJM8
qHRfYnkeyiO04scVHliMcAc943jrQMPX8fsmrSUhEpvZ9MgJZ1oiJbRVwT0s7dmjG7mgBqDcDUdT
EuIdXPvdsfUCrfFIh+S96AZg+F8xFVGcuXrWzQre1lttQ6TXFA3JOMx1EQsZJy5Qbqhe03MsnDhE
CT7VnNdq8707ZuuV1kvh1FEkIb4BDNp2a1KzSS3LO7BKUCl3w1QvW2Fr1s0hfS5/6bBVNzkbftDH
ghRQE/HSua/Mon8NUYVdfKdiKpdxhuC3azgH4FUAA6jbmYAR8NmGm+JCOzXK+8ko72IX9F6x11Hl
Tnf4ms9BQpfICNqTOiELqOyIO8cKXyXkGnIJwRucnYVlO7ef17ix6Hu4cZw97EeJlGF5GgIRmoF1
Nnq0VNau1MdCHP4HRMzR/bLqpyKaST1TT/ONvTnwVQXSpE9yoMrpz7bHv9p6017pRognUpBPJwDO
+LqXIBqYQ1IxBjWUFX4HrLIxp5c5j19YOkIxQHWvw2GhnierZ0jRGR1WsMNnwxpNR8ndn6Xo1RD/
+1KWhAJNLekll3wIr4dk5/OLSZv0aJ71/pxio53AgUSvCrQvF7uVFKYBj0Oihu0DC94zSz55e4gC
dhJzDnh77PkjBwryPRgpkgM4yzTi7tvNNBtmE8fB1Dwzj1cSx8rqfIYwjlVNObvfDXlZDAhmI5zZ
x7koJa01vKdR97b5CbH/cBUvuS8rslxqiUbvoiWxmDsItkn01xY67KK82ZF7q3rW2+fiB6CsiA0g
zsED4N19q478FSX+umZR4WyXZhw0gcrBjis9R5iCkypRyc8d3O1N5SqWNAEjjQLmrgByvpWIa0ev
sNzKdSyC/DTB+VEhlPYVM8TavnRYKD7j8mhcg7O38Yj165ymTYzlgdOCP29+Afle0/a6SrVtC0ry
zzl8ytsjBM3vXmYiE+xHvnBzKxD6E9OP7n26kYt3SVyGqWtktPAfjb6PbXlNzkthhj4JzaIKbFeX
/Zh0zv3pN1XRoVL30g1Y3vbgfP5rtU9TJQdJFgS2yzi+jYV9JRTD0HfKZAcWOzvddjhD8DuTRKgP
rOr8HUm/EjIILoYOSZ6CENQgMaHOKFzN9MotboA1U8stu34eO0h3Z8qvFLqfnesnVgJS2LZv7iL+
uYBsBbdCPmcQ2nIhy1VOvWzBzTcfEgYOWR0O1M8HxX1SJLHcoNpcQFR/596SmdqO/X5JZxbE3irF
HYnJoz3erzGnpRo6/8ytskpYRl3y8SWZ8wrxTcYHt8xzV0aZSivcblO15wxc1xPXnrBlZwgC4SoS
lCe0XEZ6+AP2SS7hgp7HtvMS84fR6nxwus5r564KKqOTN+bssvOcwKRyjXhw44fdc68IHSJkpUSt
MPrpep76yriauYSAm01w+i6OPmbDaIzi8HKy1NuDo2LHjf9F9ywIvGEwZAy/3gsepd21F36mQhYr
UIc/GHjiXuDou6DrSPEQgfXTTDiXoLErdwkXJ0vyWa2f7FBn0gbzk6DYelLlLa+/tXUkWHP2V6LO
zS/FyN64DjyzMdnyFMEPOCSYXnfrFGZl9PMp5Zb1QwbMnXgjhYnpNAifOftgdoG2Mvtp7J+QBSS6
6ehBrVfCxJIxLoO5QELv7k1fU13J9j41LtLijeodRW1HzMfpDQGygiNUOF431K8nwmV2opA1Fect
u1v21IZmZ4LbR1KvUHeAMFMslm5yiQCYRr1vLY9xPa4tMhhB0KCHSpmEF4gTyc7ZRr1dD4QxCln0
x6ywzukJwf6llW+ZemibDpjqHrs+wJQ+Sw1AF+GlHgy01KsaJYo2ktqv0ce9+aEYEMFjz+FbPlBN
Xt61wP7KEbfUgP/WICptIIn7nYNq5QHUz+EURqSlr2Rw0kpdozKPbjnQoQBF3JZenmyej/i538lA
KqBryYcmL/7q/gB0bhmN11qZVoCqnJLw/sPzNWXNsWTudV0W+aP1mQGMSjCS2BmItvL5B1jRY2bI
Yge2Tm9G3qyJlysZ/VwXJEdBsUHXQ3xKBJNi/iViJT+mcq+MrZJAC+OXJCKOS5jX7mtVG9ca0TYA
CLONVb78oYXJRLbSr2VzvC4cfQ7UhmWSZpAsTIQPIADofNjJ470aH6Z8ttUnnBkVoE+sa4JinBAc
glnpHvzp9w2+d7Dp795Rwu6ajBUnwMMJUA6ts+C62MeTREQlURNKs/0L3borokIjPGw31jS3rPuw
UTuQW7rcvUpPb2PFulkpFvDEfLBM5EKlkFUDNar2tas38JuWce2LPqwBiX2XLSUXT2A+S8kfDkfR
PHvHcLRro2v2QP2v/WNvUJU99AKP3E1F68id1mZpNmbajwLCi8AFV7FHISRhylL5saQuD5ZMcytg
5X9QQpgFTqmKwJ6iEjJKngQcZKud2Op9hIy19UAFmkjZ1NwNz/g07MBtM3ygH2ur6kp7JY+jICWM
WCMfwQbPFhkHLyJX91Fua/YZmNCLY2JunO0ghLv2DMLXi3M25qF5u4age7yX4Sd1rV+eoDN0OFzv
YZR75cGzn7CSyKmekQbFtU4UTmExIATl03DaXGxYOdOYycax95UiAWJdZwNBhjM6rM8Gr1yJfWrw
C8sD1Y8GxAQ826IRqaI4xkgVQ/GpK9ra5XjELe0Np29onxBknCJf0ZWfGGLS6xWCZ5mbHQ/K2iuE
a8BAYQ4Qu0P4kD0D+uD6jTa2cBuu9I2rE+7Nt/oupc5d+V1pP3tPn51CUFHVjidSKxW3p58Vpwf2
7ynaf32l/QuPwjlDU34ApD9GM/c3qCyxeVxUizZ1IVdQawsmxRxNrTLeV2EcPJMC0O5aCR3JAvOR
7UmtG9oJC277mnWQO2yTh/AI1ShFh56D8tp1nOuQgewQdTwtkUDOWL0fAN58+CCwniiz0drd2pqY
blCIUTI+VYM1tsOcV1BXRwh8hvsPlBICkjEZli2wJuqmbqQaXRfg4zGhQfZDnqUKPfb+xdd8eANQ
OGZ09jr2V6fMHkdc2pyYrlUt5H1nXb/T5WNEqzqK5rBRlK1dEKsISNRFG7F1YOuO7MVaZDHB7+7i
HBGRzBaMc+h7jvGpIT/xy+XIMpC7WzLhZO7sdDyr1TtmiRH4MGWzarYzMYgQxXnOQO7e1vcZGTAg
hS7Azl5EKOdrnTiKjLPUdE2GYpOutIJQP/uh4oQiJTWgswKKfWcGKcsAHL2RhuNZy4Y1Hl6IxmE5
uxQPLyqpowvxOucCjWQK3iP/TOHoc+gWhiimt3pD5TO9q+j+NeftOxD0/MZIHR9D2eyNxTDPgqzV
vjEFgK1EwP8hKt5QZCTaRhv6GQWyHNLHxViUEq7j/RSh/PBzKArUGRQyY2WnmU12oymav6//bUpx
ouJEP/vAq+oEMwZr/Hlg0FayMuBm+tBNgyLUmxYf0otwidk+MAHa+GwX7zLftLV0QrLLVwzvdIt2
SeH1CZzGU7iUgtB8Rcp6bij5Y0ck8WZl85xtXDLonoXqk8zQaea/AWKoIEzpwrTXaqleVhL9oo4K
sXbdGTVReAmYi2Y1QgyCtPSkFThhLrmF8s/qQcv2BBZi3KCmVqSFn5Yqq4d19M/tbiQIgXP6Wuk2
OXzgU4X8tZfTDaGJ4pNW7ULwGHC1VIu6hu6Q5bA+UwSZrMLbC8Ae4+XjtG/BwrcEd1FrsgtHSKMb
PPCtKwuXxJ4Y+9ScRz7+dd0jkGo5U+g4tWWswO6E47J9qpGcOAk3/F3ecvV518ydgi/bJNMYv5vT
UXbITIKytCsyOez0wl/3SDtxMu4M6ZzA6iN96Qq8NEIdQyE1OET+4aS7A/xSlRnONTW4jiR+VeLm
jz/sGQv+mO95lWvlowYCk24Y8W46uOLh5qk9SgW8al6yoiAkFeJH/bsXjXILtszLf1TvGxFWPvg9
oyXnLwY04L5o0cbdOgFRVS8uaQ43nGk95DYPXsMm+PSXwVevcteo38DWY97o/rsZvuRKJ4CFuwMj
OT4LRaRmLtpiPXoVhrS64zra+GnhAwKivPzYr5NQMfwTkTEiTn+1W7tTDppWZxcDQF4ujymBKkHP
OQehq/RIu0D1A5Aere1BdtLAgkIX5CZmYa/+90zCiiWzlVhdHVlUtOrVVpwaqKvl6qIm0eV9e+ix
LYWFl5Rb46uKgNd5X9XYwijEuupftV6LkNuaa0oHvgJoIz6g4fF5+syyRFxV3zkWy953hfu067lR
sS/6iTeF0G/DBcQ1LdvlbDzejd2CpprNmNLSF63R7geC9BiLz0kEiPTDQTBiZpRLNKl40rgz760P
PpxwGL7M+BeA8RA2MY2qfbnAPV0zEwzapC2eaK5qF+fvt70ltc+cta2QKAVGGFPXnaybMN4pNis5
9PdoMDitiOAcJffEP82Ob2qz6+w+0xltBcoo6ZZm+UIdQUW0wQ6JiTbsj14HlBOdioA7HNmU28cZ
rqjakojqBfeB8gjdzRsYs5YmTPToYgbuDOcPUNVGgPktSsEju6Kc9hYfkiqh6pv9CTitRlurZOis
rTQ+dKBaLekapzALwJ1z45Pzc/EM2V/3SAEWjjwAkpi9EJwH+57cFQ2ZneTMdBeSUJkpmvpLQcsP
Hj+/DlVybXeZmmvBeJHt/pS1G39h9NhoVWSUviW+fWIPVF7imfJp2zDkCVgRlDDCA12r8/N8p53u
gESTgw8C3OaRQ1wd33tk1jQzP3DOGFJ9O3fR5mA5IbyZv5zFpzQ71X/d3nGW9eCPhcp/3e1M75Kh
kiY5FDNpglxm8MycEgyPFYhSfmj3odzkIEAUQ+NU4zGpd07bl37Nz7IlY6aZKItaH2eydVBbk83i
yECalRXx/URT/6svhscHJCD4IXaXDY0a3ilXyK4JlrRLGEfnwycXMsaUXa4yCXPdxOL+oaRf4ac+
b3UsjXLmK0ydOTJTGDuX9vGou5rN4x2Wt6AxmWKZDvDtpo1i0YwS6UsdsuAztCa/Ogb5ZsK9OrvJ
7iu20VrhT0i65DayV/ETJ7wBOv2HHCa87bBlfy+nM64B7pQ2//Srr1YBcvDl4LWQIsZeEItXgvpV
dgDr6KeGYbS9uFXrVqOGiO5C5LUkB25niX4jftaERNOP9Xq/qDYOx7NgX8TMj1svxvFqgcP2QyX2
o94PUBYNAoGvKb11xAJX0fm7SUvGLnlF6k8+2GOPH+7+Np9DpLzEtwpI1eeDDixMOnivyDyGP1g+
W6kw5Fat87aV581zBhm4eWmn/QDB/bQJ0BUcOK38w1SZj/qNC1531If7ceiQaoh60m+RgIxw+P+2
l6aXtwYNHAYQjGWE9yJ+uZNcLYvQc8jFM5IrS6DWOao/XGku8DR1yGoBCLCHQ2qO9JiH+7Vx+yLL
bsY67pv+Rr5FO5tUHGqJ3rwaYzb4m2bXvGk4XnOqaOShCWEPtqh90VhJrdc9rDjLEt/tqWio/w8P
f1UbdDyRDjOhs7A53VY91veTjH5dlYt88x6tzQSgCPx6WJZ2icQ+VwQJc5/n44EOtuMAUuwE4Nz9
SUVKlLzUotGk/5dzjPsR9W1Hzhzqn96Y2Pwn48YZ5fN9H1aUWNO125uepv1aQ+yG8Jf3EdgonU9k
bPOj7mBGZC2K24QuZqEVNUA+TCBJTpLMz7/3dsvJI4dJ8pQyqI5iEkZlDVjRrskucr+/wfQMwZ01
QGPK248mm5vWVsH3VetOP0kaU1Y6K+l7wmBmlaj0ynnEE2GkyPYIEK796V4dUMCUGX0luxC3zbvg
0cagNAhPbifWnh9DoYv1ohePWxhXDO87EJDWkmvEfB+R7Y+10/K6vsR2c73A7GYN302KyQlc5Gyv
0XuhYZV/fyKYRIJq3AOuhant7A8twr+EOr3ejFYl8G9oyyMD6CaPHdhu+dH00+lbE6UCift2zo53
iq3fY5a2Az2oJmbCadGWh9UPekq97q6JLV7UtmJ3uYtqeMcbP8/zviX0euLLHzsFg8kF5kYoBWh2
p9mluWi72j3ldRfG6jpgpTQkK466vSY3h9NdCNhXpWvvcb36cPMT+8JRe/Cd19JnQpwT1ytPyq2N
bvr8mxlAK1aEM9ZDYzVLtcufzDCoDk6I8oCwHxmCB7cxcfLWOupevP43EYRwwEnIOIHmznf18S/h
RoG9I3ANYEVPmfdLStkAFjAoBC7b5/uyybJnvTJOZk351BCIgSbQ5I1YRZwDMO+3Hb1CLW98SK66
xClDSg2Blxk2o/6apIEGM8T8xLTGao6WSO5hjGLfw61bbi+nwkC+S3y8OXu269bdLTEWtnNpStFK
xIRX6F49lfFW0j3LGJFhXMH1xfXjOzV0XG0dv4tfTECwMsYn0IczRRE5i2o1Jqw0WYplrcNXXcfN
U3ALNW/Vn2vLHeGe8GgLnpdOavX577mnIv/6A4AcscibUkqY1Mr43KaL/AeM5YtFwvM2B99fsF73
IkcyjYjXQgSJSgAOzmdYX/hYPSjVbZ065sTerqwI2pLKfiQXhFMxOgWaJ8dgnB+cD1XWDgqjUC6r
gw+8tuTFGsV+4XCMy3W+VtdGk+tnnKDx6UVD4WK98Xt6+GYSiyHb9hzFFL9fmhOjtgTZ1wgsETNe
RX/hc3u1Ada9pkDOiu82I/S2SX6BVBIeukqSLAvXJ3t+3nQNLpTWB8zVn8lIo8xN1nM6wXMy9JKu
IODIf2/6DnZU+HAiNGLnYyHdiBYCVD68o52la03IxtLTwOOVYTqEyayQiH4ad8dZ4ethdEiEfDea
pOfBHyKKk4Bi4g0I8FQSPuZpL8bU/v+djIuydi7F/ZPVWhX0GMzMMhRxm2Rglma92PwOHOBaIzd+
ROVaFBYMbamXoJpXIVP8fmfvg18ehnFftIhYF61EDBkvQrTDbLTp/k6BV+vmHZ5ikUrI8b/jn0p4
p47rKmZgrwQJriRC0O0xeyAvu6WEf2GppCttBw/khuPcUHU1DW/7i5GJ0OKJF/TBFXqlBjhUDHqe
9k5MXMAujLoDFMCYbBsftkrLQeG2WASUshZuW4taqn4OtWoSE8gRl0oG5RCLgGEWeZYoAlS+F3c/
Y8PLtK+yxodYW+ia5pgWhCB6On2K4gscQLm6YC1XsN+0HlCkL1KN8/JLPgQRnwdVIWPu5AWLD52U
JObQxc5wS8j2FYw2uy3k/iXKkO2eKc7vzmuCVhSamQeMDxF8TYjaMaa0bQfIu8uPhXUG8SSVA69b
DPpwUxncAth67YjsnJjGt2tUe2rfouW2AnOEMvJ59ZWDVkLE4punJT7atGTnhsBD6GIYOjvT4EkZ
tB4Qwu3l4Fw11laRxyBBWtaBR99aqWckUWk1WFNJKCmszdwCKCrvLeAy5FAyxMTAQ6vm/83uGHp1
C7CH41mcIEK+VebQE0qZSObUq/OpitS2riKhOVlRTdmyCQO01Aav8KynIgagrc0mvpqKabpQYTNC
M2jxC2eoQMOdKiNGLa8hCGo+HnwGHmnXiHrStRwxZyXa4rgQiuQB6XlTaPan3AE3BSHuplk8esmo
PO7VQDf7eoG66Gze9dsyQeDE0f1ERgFGwchmkMpmJ/B/GDtl+m7TTzjtstssnaeO6H5UUqfgZw9t
N8Jh2m0hYV3SL9BjF94xaq0l/ZEz25Vqt3DBD1iTQSP/YEM6/m1cgfCErPo1xehNXpOi7WY24WPd
g+YxOe+kLuEb5CwRZSLG1bkgI+KNNlRtNl9xyA6BgwQ1qhTHm5QH451U2x/tHAi5tLwbNgltyYjo
5KOCiE150zg7NyFNcAP0SAUWGwC7Qo5wOHsOCHhj94Y2NCb/erTpVrgvC//e0eVwu/AH5yxymK2t
jBZCrpVVAKgD5PbebO4wVT2wMkFxo+R4eAAAm3yf/DNK1KN/ItN8QOQx6bVgDHvNdL5jWofEbdQE
XT+o/wFtmn+h++hDM0uQ3UdNtEaBE5G8Z9jd22OCO6QAAQiKI+ZnXu3noyRyIyPCWzcg+1Ck1CZs
y+Udqon0Fmrm5zJSQSxCrENHnRfTAmbHstpyZicLYrXiqyKgAVKlHT/7KjXBFsvvpVxHspipK6ZA
fczkhOz0hFuCzeNG8wl6lEDupkUNwQo6tBeWEdlrGEoCipbd9CToSI/C4kWiuaGa55XdQnpFBsEU
lwIeV1c7BmJCTB45o6S3fxfICwPWMNQOujpNZIR9qcTsPb5LUjzynm4EIjxECrEkibUsMWxDUxC+
6wyn8a85ENHOR616XC0mL/qRg6nKEk4r9QPJXEcnBLzjq0u87Z92JSUVLk9/6LjEbXlYCIMvnr6J
tsnyVbxzxNFvHAIMCxymbLbczZTKlQyGXs50w5oDgeKxE1Wk/9GwDhYufNbaUZz/8qF3xOzkxTpT
LJfxJuD1ii7oLiAKBVG9qwpvNetLYXIiAI28veohbKgapgG4zG8UjP5VL66CRutSbHIx30ZoD9er
TBI1Vq4UMwT6WwFD01G6YZDwbbrHd/zu9eWZVJwLn5+oBAjdgb8irWHkqXck30WyVccTPQhGmQ9C
AoA5eZ2GZtmzaR+90szsmE3WIeQu8JLKZkuA6CNquqjwjNcjXxlr/+9Rv4CvmmBHZKdN1w0eHi+W
ee0r8Lj/y4r0M66JhmCTUVzgF3Z1/G6nzj0USVWkH6Q9wRoh9D13r/RNFqiB/JErUmYPIzxeYTxI
tQKaWdHFSjrA1Pe9k2yghS70svX6JogfJoAn3ZFRks0j6i9YrKa5nVaSTZ5qC/ixpFcWhHaLEI4F
LdBD5yPdqyDveRppV4GlExd/YfDDv9fQMQ0Apq8SC7WLwUTLp2j0uZ3WH2IUW3up+pw4y+rfVBew
lA3HNiGdPVuW8RNT9DkMTZNpb0duq5bY74jx6rtdRhlaHdagKteZRnB0KFCO2jj9CnSGuOd5ioFZ
2V314XqFCwJ9+3MMKoVhYWCglxtLbSoYPiTw8M/6PSlKF8DUg1ZUh1bLh9KGmnTgnsBcAEBgG06o
pvFRk2EIsTOV7h5COVy9c8F4cp5Lt/X55WC7VQ69/3kt7ebuIE2vFO024WgpbhCmxWd2n/FMvJ89
2tvdCcQA+6wJTUum2OP+CnOgY/Xi9DFjVgqVxsTZfmlqQVvcq4SXtqe/pngH8Fig8Nhv5rWKG/ZA
YZcZh2ez8BCQKQ1LhjWcKuB+Yx7MySzIJFQ9+FcCYV9Craaw2r89jRxaAkFyM2M+LU/BcL7m8+db
CXOybSFT9vAZ8qOjKh4P2tB6yerWAGP7B9G4W1x/y+0ZbPKzOP8MyYMNdgnT5b2Lj91icV4OKavA
z2bpF8l33kWG/Gf22waTgm7+Oy5QZ6L2B/7iTpMxnd2qP5wM6RvCslPnUXNuc6akTtbM/gtKhM0I
FXUwMe2ut5mkEyn3MCjk6Dt11v7TasOCrYcvHUyWN9T+Gv3ae24in+xVT92L4paThhrWACyjK9TL
nkTm5s/7FZJ2yazBxFRp6nJFV+j4jukkz+qvf2v8b8mJVcLgW7lNHBrMvnjO9Ip7xeiRM6TRpFRO
g1v3JGmPtJCl146bVsawcc5nIpK/Y2cSbCHFvsYFcY4DS+okutRcZnqBdhlBR+zbno2k6LLD9f8e
5vmLZwIQmSunHszYoz8NC6sgjt+uKkLA+OTw/ExdAdcJ063qrtEzO6WAntxmqIM1CTXzow3avgAE
GiXO1oISvBXFGT1tCdEX+eak84hsBCaM2kU3qhJsw9U+En6JtEWiJvFxEzyWC7qOVdNowDDcrXUT
XDYrQflqRpYXpFcfbFrQAeR9JmiQEiqI3nomg3fcLzM08UFGnhBB1ci8ObZoWqfyXAoZUMTg83HB
l1lKtP1WiwC18P4E/jG1iub5gM1gk43YTT1QB+6i7G890Xk9Pcl2Xp1b7/KVTq1o3gL6HgKTSEi5
I24vDGa4ZlR8tBPHLxzYVzonaH3IBZ2q/uG3PnWSNKdJOUAP0XhENvrFC55idLpv0p/IJ65bvD1u
pCRZh7NTGGvkc4IkLhwjUkHtHVUGkgnlP8GbekPtug/0NbtOhYASopiFfCnYvgAbmMBjd0aVTcsX
MNeloIZ9uiCBP+HCwxjmQgbZ61ktpzpp3Iiu9oWI/J3ZkxgapcSVGhT5PSEPX3IdU7otI1HjeMQ+
t9LoPHZdoXksheuNOGWLauxnxDUuwOih1WfmWC9m/EXwnJ3N9Sd6iqTZlvmnhWoJ6uFzuRbM+roJ
StIXrGYEsBDboSFS8mtWhEgtFBvb1LtqNFRisv9yK1NPVZdAShI1fXzE4w2rgeCKhv+XXH7kWs+y
B5VT2iSLx3v7FXH3vqFJw6MyHU5M61MXUYb3mn8GM31Ps+vtNZ1X3ySj0v0/G8jZKdkENgBHdAaD
T2g/Xl7rFTH70Szlbn4l20fb4CLlV3tQlWL/6+W6ajBV6b7k+UL3TahdK7I8C3agC7gHAOpEMwIw
4DN0QaeAnxMQvcfMvaw+heZvHgDX6wdD3Ae2g7CYvxsqr70FGmwSY4jx/720vknqJXAIBrtU7Rlr
l2BPHZI6+/LjrVI3CmfPdzJCXmzYIC/aE16F/elTkxIs/SXhIqod+VOaNXSk27aPbtXbpDULI57R
wvc9tbsUIkDKsZQgoQZm9zxcTH2vhH09K8jkkZwP/PJM4JmCPH7TdpNxGkMUQPWhmuB60Q2ZNfiT
GC8TzNgx8skhFrb0gSRAiJ9Lhwe8weA85cBwIoWOpIRrPtkF+iI0hajWcOnriD3RpG1yrx8h0wbF
yB5AqkcCnZ5mZrj5C4pO7KH7AghzRRoB46h11/gHmjrmRcDjgC1ePqoQBpntt7qWEFKPZdJxG1nK
q/gj8rmm9Lw8Tixc9iaZBcHo4olE4AfSC0SdjDOTKUzKQ97XE0k4FtapyOw/lhGB4nGpgl81GLXT
L/9pPON9i+dPhDXFrHa4fcZLvL6HVCe1bDtV17KaQd5VcxNNzN4ENp+dN5GS6BqlJUCEAnweBP/N
c1trACD8hkhbF6yR55u4Y4qBcJHwo0i3K6XmNC/RZQFNL7RFdClWsCieYlk8Rh98VkLYmuUhT09B
KO/BiWzgjarfTv4J4RQR8DwY89NaljKqaRzQbTcrbxgvOmUgYao/K1oiHk5HlC2I4poSVGD/4Ioc
2icM6sNZVDTUPeD6miPhnbJCikBkOuLq9O6PIto0qBmwm8a6KXN9ZghhH6L6T6JzOpNur+Onj+MT
Ybo5tiE+8eA87dZ2108chB7Ok1WT88fEmIC3qMbxipU5H66Z0MUxPuFCjn6mClQ388p+XPw9sLbE
4FvoWwMF8JEjaz8bmgQcHSC2noSGrDGLgtu8svuQuyz0SHde2Tgc3V9MImc7+3660HHduAInCi3J
JC2gs23VNvfX43cX9J6/xjrdzFh3SvD7KTZcZ6lKBtb9PSG/cHfNk3ZUjaTJbbixI1l+GN5Z+gSO
NboNA9ugP4F4O/T3X88sC9mlhkrm0Twn3NBHGIS0+c1eULgS2IjE/qZe3aLMX9XPUPMLpXVuhxzX
ZoDBJjwgK6q7p+BWsltcw68Ru0qgzBqQNM/m6J4YUhlVYDcdMuBDA8+GDDqAMWHomVy0A0UcOxm9
EdK70n+W0v0h3Np9gcBBDYYja9x2HUZuFqtlaBxTvI9nvcpfgxiBUgvUw0gk6SjV/zASCP5Ghe1m
LH5qzROloObw0vS0muV+jBhrTRDFdklyflfa8lpUfnNKEKPhVQu02liWvUIEXmtSWcUa7y43Rit+
KUNnaUxfHx1dxaT50kIrkDJmqAm0Mb7XuzTfyjqn8eJBhMh++cnmNCXm0fUn5ml8+s6mv43sxRd3
I6/4uAqXJFiyf481FvFhzzuvYguCeDWU558sIvUpYCDeJCHPfSeOO09I6ADfUSKtbuxJSe5gN5l8
q2eIjpZhJ0n2DHc6pxn0L4gk85g0B9+URlC1tEBn0TNhPsKrUNotzVHx5SbqaWxlqOjLVMydjQuX
QE++4eDhpCSX9xhaL7Gs5tRiFZ3gQFIUDbYlAXAlj+oK8gyyOneq4tdGe7O14ESxtpoLQRvLCM5Q
2JpAmMWLXj79LzKalQ3YxwkVTihaH7hqd0mGa+9zd5sUw1XLaYsNNJI8VCgTAKG4da69mQva+z8C
UMuQLQ072uOr1Y1ZGurUxCtmxneE+88w2xvmt0Bg6pfBnM6Jqv2MLxVlysKRn138xloz9UCT3Swg
iUUpBy7fDyBeOOoXsUHv37pqAs1+j/feWWtiyUQEUB1g2IygjCQGSJ1mIuyHolHWM8dWYb0Ec+wh
wGac0DUcyF1/RVJG10ya6VZ+4Kmlz0EeM/FRPpSTRTKAd8lM3E7idGc/tpGUGpGVqzQFNf/WK7Ho
9OzvbK2/vOIEEDOT+LgWYTyBIgACUqTlEDaQUupEIyP9UANA3FDVZCjBwnp0mNz5qnRQ66vAQ0o3
bB9CYewTnfiPc5dZiNQUGtQBEtnHdnwe5ODOoIZFuCzYZ0bsX1NgUMVsNrtpsSKABQPX4ONc2rrB
vtFY9msKM4IjEvAoVCLu3LNzZVp1HMoQI7KSjNV0skRTK5WYNQWnsmjbV5F2qg+YJUqmiGiARF6D
+Mf8o1Ty3M0q696J8Tv7+IEex5sJxMJ2jKfMhk9k2AUHfwxz6p8l5+4ZREp8xut99ejsXayfgw8o
UiAmdpxL4IVxZKjBGjcbncMtH3vj/OzqLj7b2paKP4wtnhBUeR8AtOPXIvqbykMRgmw7ER3GQ7Bo
sCRwsuIyzc2PQmIv/yLurCwBMvxAnIqCQFXuqRYqyAhkJ9RGFQWH/6diebeYNBaTRevvM8P+WpbA
vTPspVenvfd1/u7HurtuvBiwl9Xs1ATtdDClPEvLve7Ehu0IiLTM+BKPzJCABvI+dnnFwoBkPRe+
LsIjGfJE+KMLwSnxrji8jHTnVq3GdXBtae1yNEUVewWVMYsGgsj9Xvh1LKbeOJxl1P2w5KfFxv2e
ji5ymt2L64Zo8kviX4/xPIlT31Tr6ps19e1hBhRQCtbCfW5VOZQ/f5GC4zyC+C+2BVTDw3Qbmde+
MKWshvf4NpgM9Wf8QdQ3vO4wGAWiiZIgSNeR5aqc/pbnsuLAKuOvhoQC9lFEtFzHigy7dPWdHL4l
B5IHUd3aZPutOOIqtNPrDQwFIPrypy2YxmuPqNDiW2DJ1BgLZaqZYkjzVQWrz/mfsEq+rjliBD7w
aJcQWdn0xbzQnlJWQss6UeDB34EtVU+PhyIecHV4V7a9vbHAEvMOrM9dNgZuj/aou9cnhS++ckxE
HSSjIplSClgZj9B3cK8xVf8O/P+hrB0M1HsS4osd6/5HhauB1Auh6n/cMUz49oXorCXGNkqxgIcK
NdoEuA5pJNgi3KC70OaWWnrS7SusIDOp90DTDWlTthjSqJdJnSOPECuQ8I/UoLmaaMIXVqfrFy7u
Xq0oeYACZ3kbLB4rfl7LWYR0BpEEgIv5pcExgecG8so7C4ugH7IKK8lv85n3XlC6o2b4q65Z0OIH
i2IBRwo5qpRGEmAoqX+8OgUzAit4vROb3wcsnIWd249VkV0bdx/dmWpp5pmh8sp7/mISAQekx6NF
+vp9I7GNXDQA+rC7erSFsVIVk3A8gf5SlphUioC7Lk7NNmtPsTbzBfenslDrkUBo7YDbiYJQDwn1
klX9LklA/SgbotEOPoXhYYEYcyub8/kSnewvGSXwNJP41rnMObezaK6RvOqWkGD4STrsa7fWSzjH
emuAsCx6EfGasNbeL86emV9Kz+FO4qlHCyWjYK6lRzJhu2X+T0VN5ei44TffVMB2ZxbxVtZShLFY
eGz0WHaGoMI/ST4/CtofIE20XngOX+oXG9B/SGIHq2h8GJdr6rkxvr65hIy+7PdRgZ4F07HYu6Kz
u+6r5V+wPqTWrXdzNJdN92udqmBqBmfFgIU8KDrRX5fWxVJEtC+Jjel2PXuAJuxDFo3bvelAllSR
3pSwlwJEeZLhRRnenkJox5tU8YOMcrQEMZhIyAsKOJ1e3tnYbcezjKLjth66MS90RJCV4v7NORfz
036thQjOspaNgeFErp91peuRX3R0jp/pC3I6ViWKyeHhHV7JMppXxdiXSfVSQYMJcFQBFP2SpokY
kWFDVh9+xowgXMqSQ3GciQYKw5ESBuWkGzcrMF3doD89Gvubd1cbDY9/8YAA3/Nvery7GcEsj5qV
+8EZTTAZdhur2Syd4jOY/hoTG4v8fQBG2hFpoZ5VneseQE4af2NAzxXVA2bpNPMqcpLP6rp0h15W
lx0+CQ0hjy3sz8Fc124XMv/2W6zxBpUIEcdgRUYMvcL20jmvMhbvotec3bCjI4IYLWvSk2NLtZJK
0wKmpvSuiSpzPAVARLThMMuPs7iKNwPUXMcm02P1So9sVRLJzvUhSkTs4hYve5GWzS/hlBRVFZ/c
xEfuJLYwuUKCFtOSEcPH1t3HnUoTefP5PEZtsAmJJPWNvAxHhJxOLsLCIRXpNdV5Kb+5z4eh8Dr+
8AA8rm/dx6D+wd1uDBmpUtRhKokwwILcX677gXrr6P3zm32o2Q1Vob1/5MQe8xeCZBlTmKnk+i8o
UUBJCWzeZsbbTpDN+ZzHB7RC566ZZ4HwOghLh7XxMUFP/aTCOKqYLTsmdW2EkAIt1m044hVC3knO
/pABYLmxfd5OdcvQRuzOboJ2djdeSl+QJZf358e8cWJSL/KoGavGTejcM29Y4wQ75YtRaNmNcJ86
ys592clBacD7MlnruMIeV5BCsU0kH1k897JTv/a8MJ2/MePPUOff67tU+ETNT8WkhxHd+xdXOzqU
e/bRKmTwonhIrhBCIYBtmZ5LlH6CjeUyaaH75eWSD75Ae4/UBe/9q2bhj90hCdnQjjL8sopAEmUN
EpR63bwT07BpAGdEw12j8TfejD9TDHunK8kUErCSC/IGhM3Y64fl2ihuEV56Te6WTXFDqrhVpO0L
0VfOM1rA2WCaBqgY1VFQasZ6UHyipXV/e9co9BzS+UVuXtjpj/qXL0CSuxJL+ocYoRB/mRC/a5z4
7PLkvLVpPEjl6X9E3YlpSzsK4BvK23pWPTVv+EiM7vyTGI4YkI8PtBkDIjH2ngoV0kT6o+KlFjEA
v2WlLBft2g/SxxW3ASH0n7YU5oCgAcoJQkN4TLjBRqtSqWz5wbg1Rpl2LOt2DOhUHVSHzajiYcvA
5/aybok46E2lobProNo7pV4V4plhgBoJMx4TIA5f3n3MyObmTWt/nkPrIe28aaVQ/ApSq0bgNWfK
qsjtx7hOcQl99mkkCa83obz1JOf5obdLj8PQdZIpAyV9oQaI+QE7NQspKzBw35HV4xLQGTzNOWZs
54PisrRascpqeV8xo+ccZ/u4q3nHagXcPooxwniPLCj2Si8a+MuDyDi+/B1IeotljAIqKnGavjV/
i7T+KrhWVfHgKPQQu4ZOychbeDvyWFPCFbn6DbEWD3d+UQm2fA8EEwxwWTVtfHPB2YbAH9G+UxHc
lbQ5Bxw1LrmgcYO26srn3CH6KhVz84074ZOjETEBtJUuq3yqKXHrKWQQjPh1RzljJYVDCLBmhmty
DgUn+Tj/1auJIHq/W+w+f4VtN/zTPfwW+g+f8cZiNFUdt4OvNuuRzPCnyuVd7zdh+UBt785mFS8m
6HjU7H/BkRkMK0MxEhgtwm3iayN2uy0DtVv8y9s6rDkIrM88QJXijz/kiszPSG4jLUDyttOizA3n
75fahey2S1a0NjcXoCOk59TB/NRIAGiXpNm3WRgqpS3WV9Pq6Gyx82WChex8W4q6ukecXO7tYIhS
JYsnzAr6Ix0159pV6VNujl1xyM7q1ef8tGjZ/KE5xOiBjdY5l7eYpLWsvAioux9JQjaAHEmUhj+f
fQeqJu9atqQqD/39ckEeYUa2IV/beTR0Af9DcFUlKIrHax8oQyv8es+dQaUe7Fvo8sofBbll/ByO
0e0gH3SDexVdE3PlK8dhH9Wz2BnKM9jtkyx4KMg+41tX2jouJih35f3nR6bSRt8rZ30EuMSJstL2
U/y8qGX3O1kWFavAKtZXNEkQYMCRkNayxfjXqPAz80mHa5HcIBOC33xIJjgZW9hzjCGB1caqG5+o
hKNJvr96bnzwAlEw3AyM78kf/XfbvVMFsCUBBjKTAdNccXLMzfKdx0y0kPUwsj/rMjZVwm3sjNBF
cVFuGTB8OkHUsZ4k/g4y4GT4WVS5sPlkWFRbRYkYksojmhy2JElDLAmYPZGc89aom2SNlOfknUxC
/x0z93kYLp/txbQG8usj74VNOY4aC76eGTidzhb1N9vc1PNefsWtGJ7xTwNa/ORrvOneoT8ekx+s
IBgbySUum2Nfc30fFMICRxn9oCjM8WoDSIA0E76WGOSJ1EVZ5ZYwEcZThsu4OKmPZ5VP8ukd9ooJ
TayAcPHfhl2Aw6lugtduG8Jy4DAvV6Nn8Zmegf2DIkTYU86iB8yD96qusDfWqV4gi5Iiify7y9T3
wvfZ8fm3N6jZBY1zy6ISrNUOiVIKSGP83iETldqkMJb1b7fQ3m43wfPxnH0+IQDrxwpZoqNl6A/9
SCcVUzcjRIIdJIjoAYLDfH9QzX7kBv4N897Vj/h1eeZAByFWO7g9w93gNVsSi7N1hQDb5jfNVCEN
vS7PRx92Om8LfaFzJhLW39yodIKDyHAdCgCWvPxyPBM0rM+4ZGYc+Dm72LiPdDVvdqfquswxQesw
YIier8dGl2FAncFrHQ+45SzImQHRnqBsCowVCtdhDRZ4n+l5N03mz/uozRxeG2WXeIZyh+PjpJOx
j+PNVS/YAalE1awbnHlfSEnPJgWvsNiRLpIgF99LPZJtGNpu+ZtfMyvp7a7zFW22NmgZ4aexOsnb
I63YrxlkWOzQEuvOioPBAocI5UuuXxAggxdswF1bRGcg6TA3K26qnqfCr0KG3rzUdFTWRoSaZ7B8
u7fAKMWWD0MRsFDG6JQA8r5QuvNc+lEWw7NjBaGKUiBANyGS4FYYojToBuO1j/QO+M8QtFpz6FIN
5LEtMunN2mk1pArCUEs3bsLK/JfNHG6Fk/M5Cfy0I6jvyCsiWaKNLPwGRuxgj+J5LCPdiMF3IsYW
EFW60Uu61oezEeev7FVdA/xjTgFkVblr53rmPUB6OjF8jTx/RUt6nxJZT9uVQGZ0Eeyth7QW+344
FRS7RA5aDM7GqchIaFdjIDbDRnrB1cGBLzDhSoTeuOsMes80yedm1sMEK1jWuewMOkIb5Bjx+kWl
3cGEtTyCizoEuwOxiqeFrE4RIWI+Db2XT1R0m2bIfyJby6fWH2WLxpZ2H0I3imwLOiN8eUyPWoG7
QkiMNj/jYJNo/TmHuguW7nWeSzhz6MtbQO1ES7x9MfW3fOQGURJKZ9Hp6k4Kb7PEgMY14ojIgCy1
s3mq7jN8R4qcFvZcfNJP7A0i5DJ1Y55JgW0zq8ogGdHEpx5IubVHojdnLA0p1HNqNayic+Dinj5/
0efiPXTxnW2Qty3FJbYUgbG5z3xo6tZjz0Tqy3bB5VD+GLQnJCFL+cRvXBenDPbaECp6hc7mxTk4
eJE7w+NpiI16tJIspfD9nbPBPuP2K/s6XQ/zfh1bmAVmzDsIYA1M1TsL74dAIUV3q3j/+nt2PLgi
PWaWD++gpfGvRhoXGjLSbuZroPQjKTXYtNEj7KroIlYy+SOMv0sxtR9qgEw/9pDj/uJ+nlQR1Mcg
kO0LDzCMYncxxVv8URgRjwr6TbI79QugMdsIbRL+3UPvQJCi2Wy5PlWCII6MyZdXe9JmzWyzYcRL
ll3pZmgU8NSNltJ1BSlSmzNqmIL8QZnBavEpIozTZeCnXJc8s0nZwd/QowwA0V+/bHVm1Tq8R+ee
bwmzh8/r0LHZWQGEozA56QHqixL2XvyYU9bcxn5/x5MMzcshV4Euv0fpmgUICX4XxQXoFX+eMlx2
LGJ0puIWGIFtVyuyi628nc2AmbvDBxNFng//1jaelNUniMy126XDoRa+ymftUzWfPVoQRv38RQGW
rWdbpXfio/xbVOERsFpSWYsusPHIQNGh2Th9aR4gglwCMHxvJMxNii1AR1PxkL4WPTy1A8AI5SNZ
pbginz6u9UPzmdUyrB1JVdXk0wUR+VsH/h1XLtagwhS5fjRyUVTFIPT8vDzcava4hC82DtRbMGMG
ylL8QQe3hRmjdAMhHr+4ca8urKBtsDmt5p/5PbyZT9v/Vtvv2Tnf52kB3quViPkWTqQRlJh3rhXB
37lS8hUbeWXbSVPOc0eB8OGNeljISgWaT1uCHjhxYKLrTHmFIhmWhv8Qvexyo3Jxx97AdCim6M2N
bEZAiGVQ9WYjVBNNbmaOSuYnvjlKrCggY//5dQwjPJpVznW3Tl4bUECeKufFTRMFYYw2Vd2G+hFF
fmsnk846wFMIW4Lb0EcwJ+1PlKEqFFqbbac95qa31Z+TKwWja3W4d2D1kbCG8AhpgWFpcBC66NIx
Sh+e5XnT7/usRBMF2E+imO9HKUN0uGhngNLenYfE/SMGCMRaQsNSVo0IizytsPIPmwOhBdONssDZ
r1bPUDmNLCvEBrCbo957eYT6qrIIZRx8OyB2qIyOWRnQq5w74Qklxf984UsUF9EQhFoFxtVz73ZI
MKWLo6Ww9qWTbs8tA3wXjIkamBC5yjZXZVDOtF/Yg8HZypbJoXMOe9KBVIUaZZtsbVYGlI/61h07
XXnSbvdpbC+WiG0GozjTWx79dCXyYvaOMB50kQmnKp46RVyraz3PJtwuTIHQ3QxiXg4qPaJLUmPe
t6NlfEF9BOwyt1H9XYJSYabfhWP+o6ieTsghjt7jB4H1DQ8OUmdqAgRT59BKIYjLsPFULV9JLRvr
fRIPxoO5utjCrUkV/mVf3SW2JhQVlIDKGOs1bxaBYSndFTMHnXom5XTbQLlWdsiuPyuF+jjmNTLW
sBXf7AffeqAhf5q4XU1QvGgy6peWjLyWm4LT5peaSxkL3VQiwaTOHy2l4mMISo7LSBtkEbc59RkW
XoPrKRvk7OpoG/WEe8+wbm/Gq8TC087j49vQyJ8NcGmuwK+NyiGtou/3zOKVJ3jmF9IfAyZ/T46p
UGWz/xSBW3WsCLqo8EfwcGQeEvPAHgr+TmYu/HytG3qPCW7q0k3Wpi1tqgrO7LTRIIZ8t3VaqM6V
u4dqwxTbY0LRQMdgLV99AI2XJXTrup6nMQNOMF7ycxmnVLgU+q5oyTf7/bVvngsq4ZBnEjBEXbZN
NHc68nxkjqEkBzGqGMDpaZ8ySB/SowcNt6CONAnSMKpKKr1zuqXfgkWhzt0NF4v2D9Js9U56VcUQ
j+zsSuEj8i7N9rmtLOKBp/O1RqwndHhk5dAWVNsNpMEu5aYhx5teFsycbSrKhfYw4PWtPEMpptTY
WhL+IK+pTN7Gs/IciHjqNhgo2JLPo5+pFa2LzP8bkJmlBxA9pBHkIUf3y8/YxIhnXLLgNM8nJawz
yaw0J5yB9SJxqwdQxUHbb8NqeWIHj58eTDwvMKrk37OGNsFhUFQDNvnxTy0Q10E4tm1SF9g8I3L6
EcPKOqNqeSSnEyHoGmM+UNzXAyI+oq1ELeM6SN9csONDK4Sopdfyd2vI5/xaTlLfdTuMMzOFqUfL
7E+i7c2lcjLhl36gFky8jKJsrSEr06ltL4f9MVObjYkOxA9C/Whu5saezPnZTXaA9pRqPU/2K3Hi
c3r/qymof4cPtE39sWp87upvn9YxHpp/RePWs5eZBP0vGQhAjIr9Adr/xQGvDYlZrobBYB5u8XQ0
X1pcTCVbDcgCVxflw1V3alFSUk47d145LAbmzmWJmo38wtp8NihCIoUFCRczKGGnAVQzxfP3ak/K
N1P2Gj3PdZemXf9tLq4CHqwaP8+IsoOjKT3Ek480HZjBHDW7394vxUXlGfo7wN6omgpYn95C8+FF
TxYZhdB0mHrGWD74Fic0eibHRevAVvn+dYV255FWoFFPoumNi3OktmpZrMIhhnXj4m3yTByMFybZ
CLBFQ09qufazuQjHYn2EZ5s04XfEVToxa9Z9A6YoRazizfVH8XcBfV4vQeQHUGrHxeQlPWtJw8Ox
zJHfwYhS05SmBcdrUnEO+sna+LV87/IQ/SyzYy7Z5tjlJbsTTU/lJHMOyPCAqd9D0XLoNNedxQey
7SYuOOmpSXLLsx01Prc/y0HWRfG4x3GIOTOugq+31KPyiF7BTTC5yyrJy363wr0ZTD5rJdvsJF/+
3/XkhwF8lBndg07yCzfq3FrE2hcG77UUetDLnQJBIeWias+z13KrpcDQHc4lCSNRCXFjAFo2GO8K
la+jANSVoZ92HJoMoILS78M9/rQrr7wAPI7VwNh2u0ZOp0NV3yfrCS+cKM7OFA00dpcQcvMwqRuD
k6qR5qSGXmwCstYx3Ui6gaSoJbhlgRgz//kD7qQO68lN1gVeNZu0kpegqA5rfOskA7B7zrWNER7h
dN3YZCSrbHAdFDphaZ2KPgMHsF0SxTUUpQk6Auaumf0L+ZgnHfmidvxZ98F9s5A2lHVyaNIVkHvf
sv+r/8woX+dO+Pi5kQeXhFLy5usq8D/ppjiouLgSeLJTaYaUrQwoMx7vvUgnh1N41tFJLYqYZfLj
+RB4hOXHcBN0mRnQouTI7T+HYSSwrQB5hOzyC/qS8ttMxz1V2WmFLZCkxIePsaqLeQTKwytGz2mL
9DNZ/S5WdWCdldE6OYzbgA8H3hx8qMxohPhm6GIBjsZl/QsC8SxdkCQo1dYXVYOdkBkCqNOnXW7e
MnpAJdiO1MsrB1hl59WJ/V/ERO1XtlotmStditwIHgiJai0rQCfcD47wvnI2h+FP4ZBpmPAutVWK
5L2E5Xqoh1aF40ZOjFM6NddPB3H1QwcPObIdq54NCErUn0grBoepX2bHsFsh3EMBLRz5KTjstjVq
fU9dix+FpfTl8jKv1EX2rq/73cwoCtP+VK7obZG4hnaggibIufHJLMevzGlcWSibQvmhSar+Ptt1
E8FORTD3U1BJlloEaIY57DdzXBApTE+wlprbDZqafy+muXcsVlVWPqc/2qQdvyf0VXpDHOLzpaTI
UFaBj4UNBsEOxB9voh5P1yAsmX69JrdT24Og0E7lYYzNlGjxX+msYALrox62Xn+4iZ69eunwN4HK
hCitk3g795pR95SKICrUWZfxtsCdbxWst2dDiMzX/mKZE9RjFJC0eocgZ87v5wo0rhoRQDRoW2ub
7sjLCwy7420Ni1ut8iqhzFrNBLxUZ7l80sWYpeveks6Bk5qK66PF5z3ZRUHon8bTXAOBaspN0N0J
xjrcYP6/8uQUtDI94Jpg/GG6Zv52RUMbfamC39nEz6hRnojolJQTsyoQVN1Fbs3rtYt8pNRAFxyb
I4OI/4RVaABx4ZPPW/m5LwqKWHx/WQ/z55hzDLrUVeBovUHMNLFJb6C3L7JXkzsE3zCHd3sXSZbm
xuHqFCppkKrd6eAoJlQC+pfgRRWHfHcAmf7dMaLu+BeMEUzTFsAE/yIsPd3EwpVMLBBHwEMVSs5t
I/BHyucog14SwX9HW67FWpMCAeDarlMTV4SjxAeOcDkmGUUbup/7uDRH6/cJaVK0RBH5HIlJdPxP
HnDfVPtZovL2Y+RgK2W7FZ8sXsc2Inf5QfAR3WUSosdgN2AGbArPBIp21TlIDQN17b+WUjw=
`protect end_protected




`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
aEP1OILvWGtKjWJ9kixzmYvznJOBoMdsa8poNaZ43LOZ18QUTdSaI7tVqsqcSdJld/hZgwGX4vpc
YiGuAlIHJw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
l/rNhyeB1JGJCJUXztcuDL31yIHLYQxo17fhqeGJoNYFcZSiqjWmAySwcUG4zBHR1APtJLo7G051
9tdb3KT4WE3AR7LpCDGJjX+Gi5hG8PN+tQ5wjzPqgJIxozJukRyxPojoDUQadWN4/DERq2EWtnIx
xHj3TPeYzEGZlAux8II=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y+mQpaUDSo/EGeBgIWxq+cVimSy+RL7rNbMmL0BU1Zq2lhWTk5wgam2BivaxUvfowRudDeVs+dCd
qw6MeX+4q5e7qffB3svTMsK6GtIkPBwvjmKTFY1i72y+naD4Fk1uYBnWG1mM7jYHcMohOeM7z/hr
BsnQazEVU+OOBMTu9+O9ywsfiSoZ4PsG0b8tam1zWRo2nR6yADyI2B7JGt6k1EP/JNbi471aWmM3
aRxvYNFMk5xHQYc0qI1w/eTgn6jAQlBKpLstyMY079LjabjqsWdifMFtakC+Q87oh57fCPTzl1jx
mEw+2Uacq86XtFrt6AOYoeHKQzUr9KFn+6iRfw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IeWYh46T7vsV4MQeHH+N/qUkzU3GPD2WBJS5Sie4GbhvDCG9lnuCHO3bU9Wlsj8Bkp9jmmQpStY9
rdYuZ3Ssy+QDQAlnKxUcLuB8jYp9bvph2TJB8XYuGY1prxOwSKcCK7k8RbLiJUhmU0kwTF5Y4zMy
9dW8rr5aM4IbhIXRV5b2MyLHZJIChC84aGTCHP8ucL89nD2AEJi1yHhrA8HkTOPGBiBKWV2ztfpz
9H9agxhf+JI0tkbQ5N4bolXAgvBL5oJHFCiwdG7fUET9Kz0CFeTKOuLHzhfGB+xIochUCVf6Plum
S8jP35WRpKAqqVjWgdORvW7ym+Hl6+nSeV23bg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ght2+y+7TMk3O4nLiLJq7JUA1YBYAlvbqxbHDYHaNX8rOMa/arDbgd6lQhD5mvqR4p9aAUJg1i0W
s3Dz7yoFoXEXY4TuUjvMoreYKuit98q0sVfbZwYLS1ihBD1HMnop6tSMg8RlAfN1a/PnubxMhHfR
UMz2zbJ0ZLGAbyR6L9oShCNaqhoODAx/xkWaLb5rT/2aOsDm47V45IVQje6IHECQXmq4WcQ7lQVF
llBmS9dYmANwlYHGZak3fDrPYLCrF+h+L76zJCqYYmwNCGCekdLRZR0im2YfleqY79zXa/mEl4t0
fx9lhozwLYO+4X4vIOAks9EmHR9LZR/G8543iQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fOIP5LVhSnIiAUKRajU9KKldDIkEdBJ5Q/VjqlwPh65gKGK5zGwP2dKNLPHncvMlMlnbvvU36JQk
0gygl0E0B0348s6QYqAsUCO9tT93O19EpOI/OmEzyx2K2QLZ8syV44XQ1EmkqYauWFL0HFyOq343
c52uDO0x0AyXGERtSM8=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FuSzyNx+2Hsv0fyn00O9RmHA6pWNoNGZAruOHqbTsgvQeIuh0JebjUxD9OJ6clTtyTZkN5PkCvyE
2gG5qutMcl5G+yyxNrXz427jLlRZu9yiyTlPCRnBkV4/3BFq0ulJBTPKWBy65xChNDtEreBuTvqt
vRnkzh2HsVnpGByv+bFVl2IxrXA4osRmx0Z7cXAgshZh+g13Z4D84oSdRxd+BW9L97T1B8zFuG0A
szqpsscbv/XzJH7bkrGIfgNnCrpMvaVvnp7dF+7f357WM5cLHjnVv74aK9pSQyXT6koPyFYgC6Gf
/4qFq7FKgOtsor5LxlyOcpGj78lednoa7XfZAA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74064)
`protect data_block
oZWAsaYK9AHYWDZafGFokEbeEafo9xYEDooDKUBan/GgfYyHHxtnM67EKYoCu2cC9lNsxb/pp20P
jQrOIzruL0/vGimYjTiGSfRDbG6joOEKGmbX1dFKLdHs1jLXwS5NjqlI36Y0jZJ89jQV+HfAUdR9
ov2swayBilE8TEUXCBT81k31SbUG/ut712tP1ZNGE3jU3GBgJXKK78oTfDRmeTt22W7HRTxSzZSz
WmwIj4yobKzpzN7C2fvlVdanQQZtgWhuft7jGLsWyB6Is0IoUJGlRuA49P1sRoXbh2h5HteQf7jX
RhIx/LCix4Q5/LP75NFWfUSJYD1+6tHeU0kSsnp1ca4RgZ5ws3ABKlDtx4e3q/9vvy6jJ30+JwDr
pND205Y5tgw1bHBs1atr/TOxZ4wh1l/2Lhvfm3dl7qIoI3MMe+st2LlStqXkr8HwCm3j7A6UlbTO
Tm7taFS+bm/fN/xLIZkJhZhcTbCIHG4VSPKsrgFjoYIpj9/WLrIpRfqBuSa4U6/xElRGM5aC4LnW
KpfwvT/DmWSoD66K35yUdtpMiVEzspMqSc+7i0aVO/QdNp1NrpRxj15xrfRC5xmJaQPblqa4z7r/
b8UPCtHKe5+bC7oQK+WQ7X8zLsFwkZraDfoePzSFwvGPlpUjGBDYiGS41FNA0gw54Ksa3M1aLl1V
rRKJbCKeEZjIVQD81LooOjv0+pXyZLiNjhgyf0Dp+GBWmCvX391QTHqD0FOB7kKVPgniPLsBWhQB
b4d8ByOISaphigQoFAzxFY7gBXScrE7pCgw8uvND8GsqyvEgLxqiJ9Fnsqpsj+BkfzyMubXkiNgW
pkAsrBDS28I59Ni4K+T4DCBB/1BjXdueddQKi5ezW8H1dtei8J5Gy/yKgDRaGpuX7Vl9aqN2bL5b
iwFI9blye0sRUinNdigMYqB4zf6AzoOobm44XtaYQd6utkuvBfSwiLRNyiOMsTbme24X1BKsS+S9
LbGPdBpytPJoTA9E1vrJguMvBo1TJ/MEz+fdyHlqU+EVSwfMkxW/vZKCSzIbrEQP+ZSUKDarxuGh
ikRl0DWYqlHjjR5HhC2pLB+8v+Kl+a2AOgN4FaSWlr4L9QynSSjGp7feP1864QFj2nq3l5WvcDdw
qXOQN9taSogW0Eb8Ftgtv4mnqXyQanShhakGAnBRh6fBGA8SDXbHiH/44DbK/yMt+WZgJ35MlwyO
ucASNv3SnrkbvqpLFr0G8Q+HVwgozKpb7OS28+fUfcsr/8o/1OHfwpIGB4ve093ZwMf17xAkDOSj
GxaYdcnZyg+vcknp2/dx0mcCrT+IP0TRsX4EWrCjJA+KST39cXEZP71z4zQ5JIe6EtmkPln1lwXK
cInpYipLmpV+lwUkIYHML6PBWI/mR/P2ta1FwZUUGHGRDaCJKp3qf0pk8JS3ev0Q2tCgY/qWjp0L
Mr7GLuMKmDT22+r8kZFZktlK+nq1K0QzaIWsEEC2Mxmh0SFxM/0Qsv3PbEDWs/deq+ByrRcjdVN9
Esqs5ijxgOnpsDOTrUN3mYxqxMoyjQ9C4T3O9CgyrDznv1E6U1XgEcoEoGlg9BP5D/H0nYWbKD7o
/K8gFPMeT9S7HeYJ1lwODPOwROC4ygfg+gyN9qc+cdPenpjc8n+bajzxvmov+IA7VeB2HAsYRzpy
4OTcCwuMhpZz3WcdudhKtiSf0njqHSU0h/YnIlZgk8wQFW5dzS5W5wyjAKnoKWJG/0vQUIX9PEjM
e9o78FvNwLyqEgoKrGIyTjcNPtwrZjxxPbpb8Jbup65ris8gSeKJS+Z9KkNhUJgao3DyCZuHI/ix
aP62FUayQtVeTLj9jUeb9kOlDV8H1lMa9ZwgMZ9QgJ4M9KIitcORkKbffN9iYjcQ+BDSex/By7lG
xs1ZcehP2NENcv+AKzJmoBE7u1huDAjzilMDoF+/jXtCk35dVUZ5h+kaDC3oTtFGj/VmTvJVyp5n
NKyR0wGe7PdlJriE2rIapAN7nqUf4ULoo5Vb70drhqmhtr+sngKzOGgQwrrL++MRjTpIZ87LAbzt
e04X9zlCR9/PmMuIZVuLiSeir6TNyxW2qKo6Ut2pr3ZNfwPAQ1IRn5/4wlpvbSADtZW2kJSHJHBr
PF21uTHuwwHEqvAPyD3FyASb94kga7LOfw3xfRNkgfu6QmqmaY7Cke0aakTjBn/e/zkD73cTDXyj
jR9HbK+c7t9wwBBJIinaUeJE/QHaTjbD9vb1sQfiofwWREh8Pv+ixGSgPQQnQV5j3+QGTdKnm5x3
Sb8TlSlnS9CZO21JsfsyHbABSCDEa4KtJSy6xZ9LTGnSCDh1X8lmrRX0IJXCrFR1maKpKBaQsjPd
6o+LhFrnsRRUNpgWIF6ArRt/cF5mLXbUG+isMCeHzs+r6nKluVlj8baBzIz0AVhYYDt/KrYvLj+g
lPlB5Ez3PKgib5E0+RTWRYR0UUlDod5dCC02GGejTJXij8d6UN27HYaeX4z7wOvyx+btokoNlz/o
eemGNlVjFc/lamoT7kdh6goDl3cNQLfDHwPCFiwFp73qeFD/10jVoYHbsCQDW3zkwz0Xhmj9SK2o
Tduj2Dui489XxaGTx+NQqxKYxLlz1cDIR2d47EYJiX7eLXi19Xr5EAfn3vA0PpRM1cUx7Migex6L
YUyl8PEnAxnb2tlKBwW4fblEI3xDhcI0zr3WlRVP3ZXUIoEtd4RQYk7f89dzUSxqV16ygAmMmVxK
QRVWTuGJAR8B8dExJMXchNvDsZKqfUFmnRnURyKDsztWByieV0//oZdkMLk7P2zp/CJGTRjZAoeu
M78IocxXnOTw/p0fOovF1NUSJ6aTvQBPko3YS5l9YeQ2hyeL7b/ZmhF3YJWQmuFqJlZaRHCGUIWY
ndL5rCgviGJ+CPXGTdxrNMVQhdzq4ObQh04Xi0/2QCgzSzUIShWTRsE1A+L7W2wT2WgTHHAhzi/p
8tE/ARtfCjOmt1MaX2TNuCaMKF0H6fBaF/ogZl1HpUQ2KbRR5/+dNk244vsG+RvJv+yvTVk/o0pr
xUFq6kjWEnOf5ku3CrW4TnZnwWdtgllDeyoVEGecBeqiqiXcfQkhNsIg1lkwDppUfkJfgeTcT4wW
dFSJby1ZysqpJyRhKUza1mrgh2jli3v8g77L6B/8QRS2lNP8O1PehyMs3K7n/rEDNl8Em/lhP5X2
PcQ0/XbmmCQbcKsYS/lc9/mAZ/hq/27ZOSVS5BljOzZelfWeTJsCiize9FglfEZtQoyOSjuIURgX
9GiwePDsxJ1FI0gJFxlXmBiYUWJv+ehR8pF4T6KehG7wuVR3C2lqYDRP3whg7tRVWHteW/D8U/aU
2nQ2mwM5+nXZ3r+vyA1raQRYbZvsvD1AvmCosOGuRacU7EgS8iatlQTHL2MFEy+rYOOphQVspJly
oCJaxiXxTola9dWg6jDqIcanwyohM1nbfkmiXkog/NLUC0az080j8uYCsIvF8LV/bitJ+VFLtVE/
NT3WkEJD6EBhg5/KQPSczz5+wK7MqwE5I8eYCav+e8VEQ5n7MMhcu4lbN+WO+Feqs2vfiWrSjPsI
+FW/ITZpzTuFt3ZeR4snHwNq4k0GYOy52FNc78jWc35++LePwu7GY2PO2jQMqcZi2K8S1W2sTun/
o4o4MllR8VuICqylT+Khnt+2l7I1VsiGxO8RPPpTYUIru+RW7W4lv/rKl1Nd2YPCOI5FVFHG4Aov
Wr/LnPs6fvpMPk7lye2AqbjrV2gkjlR4pXPMbgj5IXl1uVwX0tDDvd+JZFbgVz8P6pqH2Walvxen
0GmF+cIkCafQgtL9NHsWIFpC3O6IJ0NbdpVKyah2Y9aTNarE8bhsCH5r1iumWGuCYvhBZo/LAXAt
G+fqaDHQXgwq9kEI4djThfSTiFv/UOVsDJ0Vwba/XHCNlmkBA2uWIwGCXXLvgUcpVDJgNEHRdcYq
8OrsK8QTXNWtgrnjX5wpCyhg5cvO0wneAGj5s6KjsqVPQML5tnjZT9mXdpY5DcKd31rZSxuejhcJ
Stn+d1OwrWeIF34f2Mmcx8I8zh9P46uDdMK8tRR4BJQag37gsJ82XzJ02gKxu9AWGLbEXC9zMdTl
e3Xw6t5LMzMzz51BX4x+OjgxMpGGFqPUxvgr+5FZQAjOQ2dydlU7aQl5Njn8l4RoOF17naRI6tLu
ioe9YjwnO4k9K7f8CDsYtTW7gt/izAwb9yqhmtmj6UD9YOeYkt7h0XDPQLAjbk2tSEMiBlFvbctz
I9GJ9Bpvf8YhlYM1fu5IVI4SMxmAtazuqdQWMbnSIer3uliKxJPbW5nOJvw+sh32d9TSjyLldEAk
8SVUpEsa2j54Jrw6W+lnn/W8wRc/7cq6xnuaT6cvKValZ6IM4JulvKZbsvGdrHgH1phrcP/GpVBN
Sggy3TTBLWKHI83CDTMxVt/iZBj89zEU5Jr8NdjFxbVRrBwnRPwaW9ISD+ZOnxjNYA3Fi6WTXsDK
aguuYd95MtUK/JGa3k4VoQFSSJshyRnCnvfk1uvzm7b4ShgXpg9UCtK/Sn2M1wpVpk7b+IDkv2FX
vQCVAQ9h2CStJUft87KLzJ2PPspN38+zoVqi46hqdpItJFRsOIRKjlMAZ+xMZUVwqhoUv2DkPTBZ
BffTVeTunGfQ/qX5rHd7OWXJzUkjRz03+5itqlm07vTolrXQ2UALhFjj2se1gKhyTgSEm3azwyVP
9f1ZVnOOpaklMtWEBGX77fA0tfotA/2nKFDusBiILNfwRGwuEUKD7Wc7aWaJtNoUgQGDKlsNMBnK
/Unrnm2zC6/3HUlXP4Ix1FGMz10FOaKXG5NVOg0x3cA9pr96/awqBDFHX9go9l18teRGEvU2AA4w
i9APX6b3xIdtjdYsTrEcgqtGiwpw8xYwKw+11CLFpm22F+iMIffOl+DitMYEdU4HXcJVsR/78qlq
LPTx6UgFbEmtPtu/akfr6CORud0emWoQgkglVEKOvBweKBjLiTeQayf/W86B9ebtm99t4g8xpEe2
fCV9l4frxV4IY2uzE97U/k0WBpD5oJHC6ZqpIJ7wWn05AQIm8vcpFMdtSakKVPd6p+i3B22OIfml
Ryq1eqoooMGJO+O1qmQpPpPfOUm2lmXlBpdyyPDRU3FYKBex+tabcEol9bPRfYC57hCLn/LufuvW
Jq5F2nd+BMQZWsYCWu6IYGAVHqHpgKjT7lnYM9P7tMmALyN6gr1ZtfVhkPLCtJAl5SdE54VUR5dt
06we0tHY5C7Kgo+8iaO/mOR5+QjzwL4f6OF4rslehOlvrPbpdpQ1YaKY8Fwabu5LVPmqHPqcRWBu
MAVwZCnpmGqRGA+3JbYhvsptz0FauK3xM4877CK/bmftb5ZKetXKYqvIv1VnCAZh74fdeP4WaK3/
vrQkT71RWud+q+YWDOAnJ5gk7xxCfs3hd7ZuX9w4iG2v7hHCl2uqqeastz08HR9Rm/4Suwd93Sv0
4HtX31vc0KoP5nPK7RY0tEOHop1JkoU7lFIFeQ8DtBuh876MweYIfGXPSQOU3eVdYkcyf/DPBis/
bX6X1WeHpSUnreL7Z3/TeE6dNXcazEKv4q6jV/VgAJkS5yU+aBKxWUNrPrIWe4YV1ASMsufiI4Nk
Yn/Ow+rIwn8EXinhpwSYh58tdFMZWEv1fRBD422SHDfikK27daysJ2U3jvUVTZ+SIowMRxdcFYr5
IN25j8hOEm9uo4LQWidBJNTwIKIC+T5EEcUJbm+4pmYHGBU4fux/aBE3y9M1OP+1fdKUTD4lly1U
BLUlLKRJu7FCKu21rZBB9+skEIirMgMITHr1rA3nHv+GGbmTCcqQdYIqRrt+RogEvpaczBBddBhK
+L3XT5JD1XdLH/1S1RteQiRnOhuODvBzkQXLRUqoYOFlCZZbC2POpS06slBFeUPeGEUqm6FVVLIw
vA/sX84Kj0TLQMFr2sWZnZOHkchPa56Qh/NbeBixJ1+ClTItlSayYCcsKTYipBF8lcnKBbucP652
pj9C00QT/bZomspBEa9Ml3lSKokfR6IjtpuFxt193EbI8nIXGHZSMYwY2dZ3YHZOXspk9bX6dKym
RyU4OPeTp9t6FHCZ5kwSF8Nix+Hx4VRd6FEbhf/OVWXYpJyyMm3X7pMW9mpq5kGRf5Md5bmENoC8
NN/COw1Pui24Q1hn/K4K7F4H4wVyGW0B7f3uZ5c07o+atMJt42kLc4kidyrB1fzfaUKV87TZOvyx
9LpEMtG6QaEQsaoSQSAZ8hZmEDmqJIqNzDpWQqTh8gDkP4QRvVi8b2V8rlYsaglhhoX0nMBMcvZG
DaxcFUdRRXS6ulpOpwJ0SPNQuZaifMBkMN53gXb0piq6JrboJ/FgNxyXrkbZTOdno0lajlTc1xty
XufN4hp6Q5koPajP0EPR5FBzRVgqVTesSEMZ3pJB71Nmlp7fHSZt9yazVvIzB2Qld40hpUmCKfrT
MBXydA8tGpd6JbMqgEgruqBUnDndyrTl+ksXAMwXa2zZiuiDuMOTNC3fdA1VAbqAd30UqjhRmd4y
z7I+ucsLHKPc9c3DOF7ayv2OO+jilf7eWifcGAyoU1ldBHE91dmgDU0x2opuSs6HrauJqTPka6wb
eKVLr0vlem48QZsC8EKe8zdGAO1CC5RAjNFfzcgbgcvxnecEnhgB/ZNSLoZX7tOC9iUftxWM7JNc
49haEOfK+miSSVrqMixinfUovta00XZKTQqUYra4tqhNDDcg/IDnPGde8zssMr+7rhpOMC8UcUMZ
1MwfiIyrjhKeizcBn5ke3lidnCn7qrYtX6W1k9nxJNvt28Hrsy2dBgtBDOvWpQzHYG3wHnARTWmS
lr3Wx6QzEkrrsYtOA7U5DWrVVSkUdnWEg7RvejYaecWRq5KV0gKayjnPu/PF6lmJUr49z/gqKNo5
ew2jwFy7U0Ku2ciX9niSZom6QzZwmkN4QFIArix6ivby84GWgdBs5fIUbEETZ1sf/+wZ2VFMbcnp
my7I1dq/Mlo0r53gP752xBBmx0Dvkv+Wpa/Jr5IMdEGJrKFfciznx/N7qrph0zEiq49b/FGNEbaW
EpzKqihWs3ig/ZeRoyvKEb8TEiU8FtiIGSOTIYE/16aahJJFPQ2ZcX7JsjDrhOvnvmna/caEQXpt
Sz2aBshvgFG42Z7Kfrt7tRT72G4bqRMQ+pRw4dDYYCj6yKnufyKGMazApDzMMAmqx0V2IjVXlWPA
PkaE4h7f0Ta8b5vmKo0JLD0oFc9yFgNKdxbZJsDCjC63H3bCzWeiL1rQR6KAlF+36NWxymlIqYno
eeUc48zAeqFrkDsdjq3xf/DWqgIywQZpvafJAk+W2ZFmKaUQnugazhsuWDsRute9NtEt6RGeKRVk
yxHxqoktLSvKlx15KuVBrh7K53K+Yy3YUZ5m1mUKyOwKdTzW4DBMPAxP7HSxWuR74Izj1EOkGBG2
ntSijz0kzss0NaVYSoFXDFo55UFf9oDzsBBiUYMSIlFsJqvVt3/Fk16/lUObMKavwhXMp/faxJ2f
WKygEkkzeFTsbaWw86QGz25Vdyd44E1obJWsFK1l0JlGL7Lfs7tGpLDK2N4YUkECpZobje7uuOcB
Dlvsr6pEZ8bTvZ+braBQFgl23qrh+vNEj0vsA/hh059CX2IS0AtFhUK/VI/j/E3JpptgbEs2BODs
Mquz0DX/c0dRtZWGOIZnSgIQmR7N2AV1sY+pG1vzmn2m7amTY3HvHblh0nNXbtt24BRt09rz5vSk
P8fhNlm1vVHRYn1ATEy1JrZDHE/utzisQbeCEycahFi/LD2JQ+Ei/GuGacmleS6blhk3aghIabck
5FaMWxp5IERDLjramvh5ZEyjm8cByIZoym/TmS5w3CgArU5SJ28qzEGCdFx4zv/sYK0lpKAbHMpd
W3ksG1JuczEiwz9MXtziEA4/2gFrUN/xmlpTBOOzuDLutzCKg3cwGGhw030Krdin+cNVjlrTIvvY
rLI1E5EvgAEn9mbs6g8SpUbBU+0XYo4W2Td0YQiyZjffygqIt36o9o8vTXKL9hRYXyrcGDM14YN3
kskoRZs5jxrbIno3zafNRk+r/p5jPOheI9LtoXZ1TYvMxkuy7qK5WMVl7D4xRgLREabx67+UUHIi
JZTImmDS7kLWMkSxH7zMjaZNLNaI6r//D8P7vlczaNInF6hmz04ixH0oUh4HYcGtikPuodu+pTRe
TWMuC5uN9FUezv7bV5LF+pk3PF24LkGU+fTk1HP487LlaphAickrPhHddQ6CO+OVBJSjcfukBmCf
/dedrTi4Q5mX54z1F2UhK8HHqq7L8bGfA2zZ3zm5ykfukb4hrBgGJT3pxByTHTeMfS6pTVFxBjJI
QdC9bUyuR/owdtB6ae+XxU5QCfVUZ2uQv8bP2Dud5rm8o/rTBobGdFRjIqrUvTFp+Pp5IIG15rJh
gpIoURWV2pdoqrCfqGJ6XANngz7dHl1v8Z0LLubmquo3UdrWeO3hlHMmAAlNwgyKseuKjf3o0Y0A
6ICGZxGN6I5lzN5vq3oY+D9KLeCefb0Der+VYPKpWtHRXH1y/OQLLT8m66AjLEy4ESBuGwAfZ8t6
WPzpO5Q+peZDQxrE9nTpkyBjV9TP5wERMXmG03w+RO8qkppKOB/HA9PPmLiin1RzDwEGoXcIoS8l
7lSskeRYXm76Ct4qVdDrbCwfMBEBvszoj/Uhaq1Mg1hRnyDnpqTkKxksK/5M+J2c7cTx2c8Nh1fe
NCe+2HelT+5wZ4qRgxy9c2r+WNw+DhZe1ArTdLfBF+wVzNPpbxPp7TrmF/vamPe1et0IuWhGNne0
4Kem/DbKeEANBx4p8o1Bd8ZI7HsDj+h/cQ6vsCr+STNCNXXhMoQ4VhFTqQ60Of7yK/6ezWik7gt8
+eWmIOM/r/XNqI2o+fQOBnP2X266iuCJ3JmcN77ZcLEGz21CV/QQMPG7LLxVXlSY5gSk+LA/p6jB
R8fNXd9Rx8cLXFFD5RcnTF5Iy/FCsWvqeX6K2ZyjJgkir2wS//IO26Mk8SRwo74nvbqrMgVRknyi
eexTgmiEcAnT0UiTUvd4RRxGQuk9c+6FfQlRPii5mdL9Fo80oZSNMD0yUkdq5vlAIAOY7LWn2vuL
6hg2av5Hnx+fk27Hjoso5zD6aCWXnuTg+0+oMDIMox6rO6tMPe3eWgnw/4MZ25s+qelZIA7Xkula
Cmo4ugVdCSimVzREG+gl2OShQZzkgZzwAs/kTueAI4MPuuM//6Vk7J4EMYVKQdCUBm3ZGex6Diq7
CShr9DI+xfPnO3g5vFsY73Yz0p7WKVwbPGO1wXTjHgiecyoEWqUh5DJ4gdK4b7IBR/h68RryssUr
eOBFnVyatygp9er5ALH3jEyroM40jhd2bH8oLPAONndUzGqa4dqCplhNDZVH4viVukAgGWVaPhpk
/Jol1E6uJq7AtohFHYNlsMXjTkmOdns3pUqkJ7vZwFKLDvxNOTAHXFFBirLOv0RHmBMs19j0gIgJ
ASu/+5ZaeXKjzxMrIxpk7yQdjkIdAbtBM9flv5MvsOKaXuI0+p/sN4UvRKj46S6m3NYzFHuRRMg7
EvdimwXMXJXolmVjy8OL9wMqtkgEJ2qNp8egRpPgQsDv7V0/88gs7y+fCbm9WpVbO40D+6iX454A
H/w9hD+yNvoK2HpRHnucbBo/PWQVLs3Me+BNtm9MtrXUNqx1nHrYvk1Yl87pdV7dVcUMe5M0zgsj
xOeJL5BprDTHwbsviUBfqYVEqX+MRBmkDsN11bw8PvBXMLStybuATEp8CcjYc6ciiqhN4khZ1614
ck1bpkL+Yuzfl3fKCohsb+abF2G/ba2czRV0A5h0VE9Qvd8F9qODhgDCVRIQjfspepgqJ0JF1jwQ
ARxy/GiVGtJxPy7x8fGbkAEtbFvryQXJ0eVHzUTpbN2n4DllofVBiZNU2LM9HCpQOtKCOHuZSf19
s0DKa+8MnpaddSDPb/GZ1luD22dGrLaPPWem/synVRrwEYelT54LW+6Jhvvyps8k5ixKGD3LpH0+
Sh9DbCabxF2LvdwmlQM3Mx506ddw6lA0Qdwu8cV0/Ch79LrJyZqXcjBYKL5jArUtoRpM2vQbR4KY
k8CalGZ2VAQDLvan9649cd8PipPS7WtM3qMF1fzbxjUtsObaa5KwpJVyfDw0jTQkZ6hqWNhS2SlU
l1Ngy66yJUnDWwYRSf6iMSRkus32HvGSm6c0zfESmTUugEk2FM5CBvAVCqpcu5yYPVKbFVai2Gqc
/CgjtUrizqp0EueBJM+DwGagSdicEYJAk6O/CblrthDLxnL0xKKl10HAEyZ7tWrE8NrAP6TbBP0x
Vg2a6z6lg+KvSN/WGeFlNiYDmcTBF/DW+Ro2SyzfL0FUAQfSwg/7HHawP5eGFVPCEZPKZF9luyEb
gzrTd4p5y5XR4NnC0PKiyxvKlT0QDgPpikXpCeyJbZC5vZlhdKq5ZffXFueGaEYeN+Rdh1Z8yxYx
LSWhnE5CmPaS5oc3KpOR2EyIAZMkyD9lH50UPf623P8qvURJi5kuId9tJyNL0HKsOjpKkznN+QfR
/jkyP4XVYxHMbnF0xy7GQpi4bUSaYkv7VSDTgCa49iQM6JxD/o3rlDzwrjyTdBFi2Q2cLbS4vJnR
/5DQWK29mNvN2zsu7Kw2QMdHfc9xdboC5pLgDyJX1n3/KK/zczH1ghsCZIGns2qXE6OnTSCSkIhD
1GOnX52sNCZA8mbkvC/dmm3K/liRd8xT23D75eWr7btcIuwaVZBcNEW88yFFAZ1q8RQpkamPP9jO
dBLURNr/GyvxwetoSN4Guox4k8fTpGPU8qqsfyRWGjo3DivusJP7nFtD1AQC+cYgK3gICbIXOnqH
e5TcVY8k+RiVwEp3JpRuhD8LOW+lUzxiZi+XwtwEd2bnZHSYWBUIDxdnZ1JYXEknoPropipU118Y
Y827StuopaHEGnSmLt3LGP/psS6Gqxo9rSWQZToECmpYkp20EVi08wFmv3OF2rDhKFcG6Y/Dg8Op
WtJQVZyjbZGQ6CF+LZgzLx9DlH5zVuJb7hiIfR01s2jGIzawRrmjdaZv3rZ9LMkZXASW4cKGy+ZP
fYRDun2rI12KEg6B9KGGSUMDPLc2wkisfqERwdDdSDZtrxMi2ArOTMb6IkRgO1VOk5aYsYchFiGf
y24GSf4DtLdV9rTE520szcc2B96UYtt300Yc9No9rVUBXC25xWJJAQJpuR/njDN8D7l4rjR/zhm5
hrn9ZoJEtkxIdb09+QkAvPxspjWquYtKq6wVXKdZ7s+fzFhYSHE0V/0+woKjCVLygeiF0tWQv77V
4IA5hqDEEj4IMHXibzH4Q7LLlh7fH7gLXxBH43i7dPAMU1v2+hipR4/+iG6B15kIJoGre1CnjKpd
uVGKuoUM7l0TCa/T1I1tfo+68hEGyaRjF0qGZ1smvw9FGQBcCHnxnl9dk9YfDKuzr/dOpCCcZduo
zXWQCHJFjf7UfvUvNmXTW7+chuOMe8+wisV6TjL0/yWQgHoKw9/31W+D8zcpNVifStjpaL2slJXj
URCtNLp3ke2tF7ztFoHthaQ7c5RJpAyWCEjeq+FLVLYL1beMAsB/6kJmzZ95B56jO16ZHHx4TpDp
6omMT6GIRyr+dfIf1KiWl5sBbTtpIj93Skz7+QzRknhQFH6TtousedGotYeROFGf1vBC4Za2lzP5
kjAAjrs245pT9oBis1HlUQUYs2mwDHZFzroi6pwPeJpBlrOrKZeU1nTtmkx/QXI3MdtMoe0hIAdV
wYRCrVs6Pb1TwMJZt3YdVpAgPnQ08kCKEQ07ygBloS3AzXW0Ji9/0iuWaf4WM4l4hdw+vngzHApv
Wc8U3flgPwBMazxq/mnCk0y3IVSwBNWahMDFWjtyezn+MZ+C+gPvfnbCqIBVMtROen4JCF99wGhP
CAdgE+0gz02EDvJAhfBuBMPmhX0V+91Ziib6XVZ6hLNpDODUSXCNHP2eM9xO14sHJdqwRqMQ3PKx
yDxcrzOfl0CRkTT77EF5mrE9totlA8bDy65AB4GLSemZ7PrUUhbQSiQPkyG4RdpwlQDWoCPeVYc5
MMMO7kQkvDdpuvVh3GKZ/tWHgMf1Wwgsb7HoY1LtC45iKOkeCvUB1LEok7/bJMD1MtwvTjXY8+q4
RLlJjAa0Jt1WUusTvowqyT3n6mE1uIssTXulB/qPn83fuKHV7bOddMOz2IQi/iUpPVLcgJc0tJ/i
kQ0MKEHMMS70zen9T9n0Cz/h1W1cBKd6hy2KAvgspLztENL6p26I5EZFVUNYReOilX1k7fQTP/xX
Nymit32kuDf26KNX2Erba0GGKzLRdKrLJnT9nLV8MMt+FjkyA+un8CDhIhg6saUbVLtuj1ejS6EZ
hsczlUOIdbg4ZUqNle0dZR2gRHDp/nKrwGgCcZcR7mxWvGI+HHCCvBnvwdNAxo0XfKkx/Dj761Fr
xchs81hldh79FfZRamvhV9zi+90lmh21L3DcDJ5fyvamiJm98THq1Ca1ifuJKGO9TraqDcdqoiiZ
wKsRZEX4D5WLPsyhGITB5Hf0V+Eyd91nBNVwkxlNKFxhJnlmhKP1FV0cCS4ynyPTBpVCClYAAauz
hHsWOt293nCo5QJCTVB6A9mGkWylnQUq1w6nmA7poSfcMpl0XzM8hjApfl/2IXvivyqRGsBUcts2
NJ83YUFrkyueJeuaUYpDxyRn/MFK1B1TY1Ire87V7gNgo7P8hvXHlq0p+sM+F72rOJW5Rvv/McLB
AXCvR+9Gd773oW+uGWk+VvTY96WIXdnp2D1oIzfWJAwVAhh2Y4xrdc8NMJBZd9HzdqROIu8VilDC
6h1umPwCRvWxMw6P5YFYq2DoJ2DLkkpC9kw3CSohQ3JJW5BlVFDZYMXw3lubVl9Ju5uxyLMUtd55
MpRU9kD5GlyersUMKnUwBmSsuPEmP2gcerPQdxkgpqBSRgfxQKsMurvRXSLyQjTwroWoDhbI2JOU
fRzB/CSLsa1QjSdlye3tXWqC+MtDmrtuFf2EbJ+bLYHLguGubmVvDfnmrGu0y1RfKCUv3RAAbBND
YLii/5ReO3XIowT7THI89GHoi+Qz10KmtkvKovOCdKuNn+O0Q4rucIdhITmCJeZkyBy31VFRGG9q
IU5pGde2t2DT56qitbO2N40AmXgH0KskJynLdNof16enI3XeanIe/DQeClpWhfQY/BFxf6Ex7I8T
b5u7Q/Jj5LO3AoJmsVATi3xbG9W2nAnhcIgHgBKKlTC9+Yh1duV20c9V2UY4HLHGZrcYt/L+01tn
A5DxqlrgZ83NTa6NQVF59pTzn6rk4GUWaX4YZGsyvUgAxgxirNoAMZfp4KI6CcsdQQmZM0iH6qSO
7MYNRv/Xq11shU9oqVOHk7pPs6t43FeRXnCJaVXKizneJLlUJc8qd72054B4JqikpKLW2O4RN8qD
QbmIMp1+8ArX57Z3aI4Vv4KnqRmgEwLsV+AksTbgGiwJg/N4rNKDthuggxSOHQIlPb2WMmXdwc3a
uI7pYq9BIXTU67QYZTxHLDYibOdtReKIOXmszT4aQjqMjXkCMe1/NO+hxyUV9hHPCyhEY1RM0aVL
1pwAlTO1qNfe7tFxY2UlhXcA28iT0gzMGUHuDsi5BjxgtDH15wsqbsHj/uLWO5U2CE/EJCIprMHA
GrbC7z1QJFtQuKMd+F3bALfQqMge/0+d4NrRGji5iJId9yPBt7f5GVyw75VUHiAAirjQKGqHykxe
qG2vb0NqZTAJxGmnrmp/i33pBAQ3SKS2aDoWSumdW2m7PF2QYJVlm6XJyIVTu34ZhXN30dTvahCV
LAoMibfUyu5vTjfDHJJ0w514DC9EQiHicjyDpvvYFquPp7PcgCPVvdUrvbsB2l6lNXYAWiaB/Le0
iumhTnjdUPf3PnX6eLDkNiIS2l3bhEPoDlV8lMVlDHteG8bG+lk9rH9wY5JWhls1P5FfgzrysGFg
aaBWzwKGahYqFI0SxOCcERxnWGyh2bZ1uGIAfk+mGYQPi8daiRHPu6OSKnZzWombvOyavgJO3NQu
YxU/PYVh+WJz8i+xr07JNLzKn5258Zm8JN8ukys0MM9YxQdcQBiGLofloS3NlzTBv26AuVWEJlSy
DCiikm/Sp0H4GtShK9xi1iHm5I4v4u5C4aqg0CB30YFLkhAxPsmOKJutwFhiBbRiVnJHg9CXmmP4
fpsAZuEW/z4ODd3EQRq9uE/TYFwplNiyJLUB2lFLdawFK5DT2tK0XwO8do2Gn7gPe5myHpOVzCxU
NgG9goLHmhPbcVRxSKq3sNbZ/yOcadkkmGLlGydQYqvNuBX/shoSZC6FhuEiTK4YZyqr6T/HJyrW
yeHlj/vAZu1iE51rJJUOpw32B5s/gOnUEPllNbluv1zrD9QgC+JuCSl5b3P2ccdS3r+1rGemQig1
EJP1OQndfOLamNg2wnC+E4ZoWwP9RcVixEpsShYsfjRcM/lJJv03Hy3gcx3lCrmHhMTCdIBGof3v
TtyWd1AS6fTP0SAasokZv1n/yI0DYzaRRYA6pv/hA2nRPirGz0XTBJybsozdW37bgpwGE/rryywu
JN5yrmC02F1ExPMMRzPCIjVr7LNIxba0dFC1FXqzKraRhysVDnEMlN8MzsdrXzri+ynAqDzNTJH+
x4u74T/r/svzLxSPq5qUfhGGwIX6Sw37njSXx19KPGjJHfAZfEMOyrpQf1Ex+t7PAaQ3Sr3QonSY
VlTfaSDKUSq4Htfg5/r+lTFD+yPUMgahPszkQ0YbUC1rAwGhArWE4e5SV2LEPbcAlxSEd+WnQFN+
Tvif2Pnw92lJrWtXduQGiOnA3MFA2ksM5gsW/Y1HDSeVpx7MSA4gRNPmjs0z5IP/4HKxIhQ0Je0d
5dztgwGU0xrYYnlVJfxmc/nWA8bSgM73fxN4PbEULw0ywYqRYvmCnXzkZFCy+o61OxnhS2vDT92l
4Wag58gmWAq0Mu1GyDPi6hCszVRV13Ad9xuZ68kI1koWjEFbzZVBKsCNI20lzy/NZnaU3V7tMFrb
7PDGBMiNODGEXf+aIidx/pKUY1BKpb8GePQAC/ZiU0XggHpheLEsBau7do/mWBoZI87MSei2Rxtb
PupIFI/JjMG5zHGQB8+QS0wNExEif/Wj+9jfc7rpQdYlwibzh404cNNVd1+6nZCZbZqgbHS5BsOn
WVR6SaUQVZrDf5DnjABk8Y8/DROuyBPe131BqbMemf0fT2AmuC1HN0ITuw3XIP9Zb8FJ0f8+Y44D
tuBNYpgGok1b/daj3ZLJ37R045q/lAr5KER+zXlphaZnqi940rGO60duaUgR66ztd5iPYLePf2LC
uTQ9kr/dPV4/tr8MXkqa/uPOKOx8N5rk4xvAfsrX41o+BZNgjldBLS9sTGsg5Sb0kxxmK77q0g8f
e2encAIJnHlrc/6F8QMmbUn7ffklYZHqxTvyKxX2DWg95mlLY+WTX0iotv5j9Wx+ebXtCM9X6qyg
QNI3iiKBH8Or1T/l4/t0w/0/5BMg8/jVjNI5ct00L78irOdiNkPH44wCs4Dw82bxraWD1p0aJkcO
+P5fbwThzaSopIh2RA56pK53O0XCEJvN7w5wm68QbYZ1RG5v1ysgf09T5hBbv8C/tY0KholCOXCl
geucSJ+2c6aTzP8RoLctKa2lkA1SU6Tv0rzHzMEQPTsf8rLBcivdf2cMe1N8rropGgyJSVq2E1Gk
X/UbHTV9KLop32S30mU3L5YcoEYO+yalJiGxCq4Y6IdK0K/XCTBz6IL3TU4TijE/GvFgY00IgwrG
88d+tGD2MsUHrWFJphW6fQXpgQkENgC5PLOkma+f/Ab9Mr6OE8xjf+jQhT5vNST1ncErLy8y2gIU
NqPb6CtYbHIeGuPRvHh+Xq1I2DBmmILBw3j8VeEfCc7VbVWfv0qOUk+GXzhVFn+seraOti32lXvg
4M0AO3SkvScW5qL8YUnqOc/Wu6/8LJn9i+aEHiHkKgNNxIttxMBv5EMLPHf3xZxSxP+WMteHeS9O
ycUVGtxVNZUuh99hV52Gz+l121njvNz7iS8Duweg2tpD4yiwGKuBKzNrnO6+xGxqJCSzDoDc5yU6
9zYeigYXGdWn2rZmUyiEoWzsUQqwLjt1QEljfRclKp3DBhBJzE8HKfDUxl2eQ7GpS9MHUmKdU9I6
oPcbPcQDbBL1D2ZOwWVmh9+YCQKTonb5LARjTnHnbkx1VVo0uvwG5v6EOrEfMChYSM5a1nZs3e8u
3VpZZMF0zrHPnF5lQWLGI3q/19ERhLUqMeao1xywRbpc7EuctbOFcRWRQv9M+2UIdnYJmn+AVlj9
dcuUMZcVVFRFgqbrUy96RzygoWQWUepQJebQvFfZbw7yft9Yh9xabuJs7g3+XP3aPdIk+mKYLmiu
jfLXfKY9+PPsrqaCo/IZmpwtI1foL2FZwfARd6q3G69PyWu7CpsPZM7/Tf1clGX0w4VZH72Yq8T2
EoJyxbelCv76PJCPC9B7gWrJT9OPwPnBRaGGO+EiBQv4zc6+5WRrxQNBnVBktfJjTIf/HEbsNVvr
TCv47LVQDrN+56kXwvDmGDsrD3/3W1t7LK4k2UJ77t5MLWN2WA9HQmaH7iMd3A1Kdeh4QSUoBOoP
3szWID/5CAl+0Dz1ZBumk4u2pSxg1h99Dko96/wm65Fur/rfIrE0TJALRN7XiSptJgwwlinULjEC
oMXHJJ7nwXh+cWx0ARpouHuwxB+OTbeE5jkwgvl8TskyEecIV/YowJE3fRdTL8Aoe/OcR7bIBDfI
mIXOsexdzG0KJjEtCJHGB3p1c/s2HOUKne67r0HQZTz5NWONL8U7lWQugcPwtOj9fuItuV3ZyjAE
O3HRRnlb41wV7uy6XOK88CSWKmFwcHh5+AbrScG/e0dwH0JgPqnxAR3U+ZsP0fCdBHZd/0N0556L
Ey1LD5N4iZIjqX+AT1MUKWignHBCHcDhIp/7KgbsizVH393QaH4K4QW9eMdfyJ5VRjo/hgkPx45y
N4U9ORtxBRgBXo1zxPw1zX1Qod4OHE/awfnSEiUP/X3L9m1Pfgx3Qu0PUf0cJBgWHYTrE1U/bOxP
gtlb7VDgs3O2PiEL4GNfQ5kOJgnJtBNnfcTSdQlkqgpQ/u2PF0nubCDyBojUPxisfXqLyZlqNftd
h4ttbb5aNXEtOA+pgCOQk7PgPx/urcKYCiQaum+nMqziclYFIEjO1juRE1gUX/W9OFM4rDnngPQ4
POw/xy6jILkUB/7JmehQmhbzIJGnYNDtWUg3FAdB3juyDxfPSsc4LBcz240eBeZvwPnD6BJmldbo
jx0i3lkRWofA3+IHfqhRE6laIVh6HP6itMM0wm91rO2gR/08PmoEBpIiopollirx1yWR4DCRxY4U
ULJ2dzsz/sho/8qt9gCCkqwOSP9OxBdXLiDukSvedni5Zkwg8Ttgl7NpqncvDVjTysiU7DYnUQ+3
4Yf3kKJeHn8eHN2nJSspCarbx7HZnkJ0I8PYvBbc52tZ9r3TReWwZbDky/BSH/tLHBXyqUqZt0/Z
H/SFRd9uJz2IeIBej3RxtWI5RVxd9oinratb/aBgBcjU42stot5k8fjz+R7GyMwantBayGb2hxTv
HdeOSo+NaZNPSlkvct2vgFj0XlhGblmEg9tqpHK2wsC2VPNqAAG58rcfIsYTHXbiUSkLZLsQlHa4
czeCCkJnqO06LG8cDZyDfBeTnqSwbd/QCu9g3IPTe6U2+8lUUj2FZ8hwHBH7C0w+LIMbE1RXjO5f
4RSyAoUp1R+qE5U2lP57+EqMasCrFOkUlK5KwoMgWsE+hvpQ+J+kRgwtkJhm9hrtyF7L9Sdba4aF
uqMI9Eq6Q5yShdgmib9TXbNcQqCeMit+qSLwRU1m+LN7mUtxEYzyPWxTbwmdPspL9rn1+MMwULNf
QCpz7gR+09W7HOLH5R3+BR3GQuWahR6HiJYToKnOCA/XjSp6i5pSLP01ttbi5JzmMLIHBdoA6fzT
pz20rB761PjYtWuzRQ5zfon9+PZkxi8Wbn4CrP+Zjga3V2jp+3TIMTTI2eMI/JJ0BK7znfSX57V7
iRW9uGbb5vNMleMvqX2292akDlZD1eREdpetPeZSDWDWquaDkPZNXiTYG3uF+ELfTQgGAXKK7O98
Yr/AesOdJkR7oci7LwOJex+7D4py70JmN5e0S8xVar2krb5ecH8tmCw/xT1cu2KZ5uLh/B3kb7C7
oI3NpUksWNZ8inC2CVbtg9MqSWSFLB30UouOi7+ShrKIHg7zZ9HKRRg0DdvY/AJgp1jBmKzzITy3
0f8BcxI00i+cmQqKN8PbaOJzQpXifpNGMkslHKk2FnCa+WQwCW+21PrfNQBV7e6+wA397cSblqyV
wC8OFjPxFi6GawtewZf/3o8nwlTl4qlBOCr+32PtMqRyB0GvlzPz7VhVwTvSZaBL8DVbN2nnuR0t
PaAtl5WA9XFbZfC+zCEmCRl2mwG4KyeHfcn7iZX5JwjegagHLF38rsbhZ1kk/4MI0HCgdC5094u5
+C7bb+ipcq+uuY+RXl8HndlrVcJgg4qkO0K3hucNnzzsvTdRu+eE+v49EKt9OIXIteWpC47kQWH7
xTABSHhD0dtuFdz7VLRDPN6IZpQfeCYkhdosVDEZei4tzyxVGzsLm9vhheN1nnWuHhLi7gok5RiF
c4UmuY15BzmYRYraOwJTyPEmuHPgUPo7Mgpus2NCGxbTo25XGfaXLC6KCZNc3+4LdUk82Fx+Gxkt
4lkU/MP9sF5ac7AIv3IzFHp89yMVUoPCwBnV4n6G8NB5qjqlo5zqdvs8miVQHHzRRSgiTg2Kwn4P
22M5FrdPfboG48/fVYK2koR8By9ttVLwSgARpWw1Ba4MYqTY2kZYRXaJdSb6pyO9gYjBSDGDEXK4
q6YLyRqWQ6zqomEHIsHRRX/HCAQ5d0U9g1JsQb5tqYVVOCVna33y1bNN7LLZQTLBv40dPTuFKWCU
cnhkk6hnCOWrxAJZFtMAxlwPgViuDmmUGiZnXwCuRQFjwkqz76RPXRFtQw0d9ET+YNw66OjSrEvK
27EFcUZqsG8QO2fYi4Cld5FskYXdHXl0/bqRo/BjvCmmAanF2vg6g/dYA7u89628ZpXXUH/rQmHt
EtIcW6v9Y9/woiTgSspwWEmv5Cn3aXQEqf6v73hUtG8CIYLrR1FNLYLkNRwQhlvczywEoVsiPxk7
EcOaZqXZoX1Jaw+4mk2yLlH0jxLYn7VkJBE5EOJGmtCUK9usIVri3QiCFv06QtmjCTAUXsPuf7j1
HFSSjmJ/kfO9w8h2J3rhUqjqiLS8Bn5FD+c5GPzI3qlCljqWWtdw4IuoUXv9B8LW71BLMM5eHP+m
6pr2M36XEDg5JJaDNK4DezI+GQrhS06I8KwhIESthyoj1jAxiaalmtXlQQhVL1g+tD7S0RfALPrt
Y9iiU42mUrW3Ay+weX+fM+IOSStg7CP4BcRsfg5/brWMqtEUmr5MOfaNHa6KBA8kb52f5vL7RD0x
v4ObReazlVseM31tYFmYypbPeBRpJjKqZbfYH76g9N0+I3y5C6NIlBg7WlmI+rsSV1fIxlAg1jiB
LR06C4Ni0iDNNf8dx3HQAg+vc2wwMucWJfMBzrq3TvaxLdKUHSkoGrk69Mgfa7DqEKuNvq+7JLhO
cDdu3RybMRSNwl5i7oLB7MkjTlqfkcOYs1bBD1mQ/pLV2PpNFBFufCN+aqwC7IyTuShfmd3MFO9T
AnUyLaNqupTPApCatRdhbW9j+0ZMmuRPUndY5v3uOXS/6aSPVT1YafR5rbG1yELxtyOAfrr/uluj
Pn62qUbHfoRul2Zvw8IP0k3Lk0acvGSAXwUJUBDwLYvd89kg+l4+yzH3GfXlLIDRVvhQ0UYAl2+j
5m6UWnbcl6iYBl409OzVBUDzHMQnJojiSmh51nKR7wt5Y0FdakrGgCZv7lKWR9ELQSElr7djLXYK
RPi8KT3QtKeQbwvuvCkrJ/upkmjOSkzUnP5Y8E+sfqxMWVEuVXxg/g0dlwd/sdCzc6AUBsczkTjj
+txZMYXYvPOswl6pcCjdWMyFmSQflErFOjY41JOXM/4smEGuONSsWDJKT58POVpv3Mjb3JpMU00/
HpQGzev8lCtt4BL+hF+jwJFry5r4Jy3loolrrgiJJkSH5j7j8N7FQHomm+KnM2b5lv2hz0gP2Liw
kz/5RW51UaUEX6m5LCOhoEr4p2MWiYAvzQFTJcktAP6RCNjmJ8SE68WAJT/kUgcGFA0PXWzLOxeD
uJnLfXFWTpOANtbkz/WqXQ4SRPE667eldMDHE+h+elMgsf/5k+0TFkfKwuxbwN0fI1cqWVVEdZm3
MdSPw8B4EcI9w0L37Npu7O6rL9DAGmCvBYn6vt67YzFJ8sbJrrz2wFsnKIGok6snMHWKLBlCY0Se
gBREqTve5VS+NZVA+Pc9rWAtFUomv0ATZosDGMnH5KWqqyrQhhXsOvVgenardpHPoHOW1bt6KrK2
cpkVKoNoyPt8zx97h1pcgbHMQtp7D03uKh7zbJFzs7BEpyClMsvM4lietRJaX0ycls3ZzXgtc1vy
MzW+phk47MMwFa3zCoWGMW3TAZYpfO7MvldC/2cNRphIhyJdZIV/OoegoPnl+KGaJQKIBs4T5pnc
tFvXUlrzQF+DMystOW739xoD/Y/fVa2B5Ug20/nKxkOGBeMdrwtr5wZZhBIIsqUymdKmHANnYtJL
9uZGaep/bUPh0qY+cMnsJkjYgtktSF/ciavirAg79cfLkd+n1qQs1KLLyBYTgeoasBk1ovfy97w0
TdSjebNF6Y5Z6xwHyb7SxCeNWStUix5SbxvrL0ag8CbgeFMuTjZABSeI1+99eHvr2Yz64Ad0436E
yP3MhAQ/z3KzYQHhThnafP69WwVpQRB7Z6bExWp6rmVz2+Tw76RUbQSXcHWamz6w8QtxNiBLiG26
ogGLhMpWTtDk2hRpoB5JUbKwa4dpnp9hPq32KO7sZ2k7lTFrxUQWjMx3CCBizi6+xW730zy3mvbx
ZodZfzTsmw1fPfplPtpjolh5ZkQtxC7Bw4CYmXgj4Z3zLiSSbg6mGJ8Zxt/fdAwhjwsvCcMI62tL
bS+fpr+eg0rr7qGoyAQiJkMrzkt1JZn0JOX+vBk+QaW4ho3QVo7cubVKcDjDwMB+BqAcWI/cS4BE
oLxSvf3rBCjP+QPH9ujRDUbXn80A6SR8Np1LFA1IZBL9p6mGH4RfUP0ub3BpTQDovQIzgpPDjcLX
vK9o/eWxnYUiegtAfVG0FlP01G7VTBYiusCbZnOxeulZ8Lw4i+TeR56XQyvsEQ4tnUYhbuTbcn3E
uGifTFDzMUterPM1QrX9PB0II3AbJ1jeTWn+cGp4tFdZi2a/HkswGZawGha/AD2DuL5COBMVOUFl
mVPECO71GpEw+mYmietA527+FyuIUgC/X3IzzUAFYoAKTdNf3ndnM5JjIWv3bRA6yz8mPJ5T00lk
fsBiF1Mdjo8bb06vkMkH1IGRYYdUb0/c5bSGE6b1zVB6EqgoSbiwusYK/qyKRWHnApsJ86hiFnzI
toz9FyBgzkt7EO6b71UHpo+ZvlzEZjO9/QXcvjE4cEiC/Gnk2rPnZKFZyBLdhVKQtPdx79qNxDBX
dx9zBnD+AxYwTUnVh5L0yxctijuc7N5XYH2Yj9T6LHt8l3wcbZ9d79+gftygtsxivBjHznFpvrYA
ZaLzLnCYNxwHENpAiWK5XSq/tfgK+lYZ1MlfIIxA7JsjWqetjSqKTXf9oCav0TwHZ5jMF1OcHfib
UKM4+2bn1789i8cPIeC4vZ0F6PwBMhcnQ3z89SHPpuD/mEIf5r7dAUmd3K2bQg9/s/tjejw53DUz
DCIRclRgoBrakkM6EmWrmgY+9Go4EMMIMa0rJtV6h44YroRAS8N2p23tnHzzoDCWK2qW7/p2qX+H
aWaMC9w/rpqIAppmzFY1By5+3bzXBr+5Uhp5zfMz9CO7E3hv6XN1v9XHX6U+IcZJE02ULASOn2nz
cp7Xrg7NczXFGeYsMYpS7tFs8E8GUHjivBKunNhDk+EEzF49Jk2a3yTibeq+FCeoXOqNVQ2U48pi
3hiYPNcfDq8aTmSBJqL2oTfaGjDwQN+8TR5YAQpKobGFyJ8SmbKnBFUHjasls08b6Hb8yCXweEol
yu9jYvCz66UX9Lt6mYHoJAiJwF1C5SA351EVrsdevW0dH4FLtcsMJ2JYbIp6RgfdaoofoB0CwnMV
tpnaHYZ8OAqCK+cDvp6GY5bvL0QXJtgyDQVM6OG2lLBAn8qdf8v5s9MUovYn38Ccs6v5MgG69LAK
k6+37X3wKnfeDx76gK9Dww3aLOa4glB+C9mtn7/INwSHLAvPdrJ7m7ZDDrGdutZKAzJHtHo3Lf/T
GEXdU5t0aejeFH1O3ldr+HRVef3DfSaDh5pRLpNGDX3DIHkH/gfB8GFVHCpYIXA0oL/eaSElu+us
d5Pq5Vx1MDGbxVMHsq782pdRjIKTNRaYSwmduQdpvQDYbjIVN+owHKbTxtVha35I0C/zdxcMtir6
zle4jwv+xADhsfC29hREuQDF7SAi8qKex5cP2RdvkRLFXmER8OLFXvpdfcxAhfC3xAK7tjJX3SDm
LvkSJkPY3HFo0WVE4Q6AA3hmAUFss0hDo9xGeXATALttOy+wKfm3EBAjzjyFXNIaSjuFptF+lekb
YctCbvrHEmVhdpZnJdYQK92+qpqt/TfpMZnisA0EbbDeCHszO/Ssg7elHhrtgfQGeUNb1alXVGpY
4TtuASJcsSR+Xmc1Nv1dxIdG6KVbjZCJdPawU79nSvvxBw9j7aBmtwDzIEga9uoyJPCOMY90d8WO
eex8KgGLE70oQAM/u0+1aaya+aF+xf32WJ5Rgq0vxwHfQO1Mtv71MJTWPx/JiKa/uiTW9O50rGqh
Mh/vydstdKaAKaic/sp/+PAdmRjjEwaBYVCauZDAjsfw8O9wEGunPbtvxxhhoMIsYHjqenYNWiqT
mAwOe/uCU1kywVmsg3+bdu7VOfcwNrWdXxWFFl/w13Sc39o4yOyYqfIuerVbGtOHhumt4pqeYH7x
6mzyc5cAN8N7xhhH8XPozmFoaPEoVgTqRNkuloSQbI6Aj2GMC66RTezYFIOfDoOktk+lLZFMYtF5
uX9PjaKfaDyAjX8/2+BZQKEdWAi1+ijGZznQ0Bu1/TKbPBxs9n8Qli1wo8zvfR2CJJMeSX/e4Zdf
WNQvehJfnRs+h0C8unc103yKZMEJFiA/rmCsJikAg7DCymsZSpph+WOwEjJkTu7gs9iBAP7mhanB
w03fsQVN7Wik6L8avIuchQzgM43eJ7umymaccjm9g5T6gGGU/LKiCWJRrMyw6jLaLXnQFgG2q7Y7
5YPwYv7C+MxBZW22zEJEXmFSdFYteDyW0bdrEovfW0Ig7k+CMzX3xU280o2ZypM9mKT5/JDvK0lf
vY18vq/kIE/obVS7Ka+eg9RPDcs3R7hg8CtdFA6GJSbwrAyICoEiyeOGlfi2H/5mwyQUibdOx3hm
nd1hdgNxIJPj3qkjGJBFhqMAoPzyvG7FchOZHX5ZzlPXqxBZzAokiTZHRUr+jHFqoxDVmeXUKBtP
Amnc2PsRU0U2qgn4WcOl4fqkjSorNoiJ/Ny2WSqRSGzGphcIzWC3qZonIRM/31nh6xHzWoTnAcD7
NGvrZkJCk2f5LWgvmzqEmj2gHVXdMHKQZhNNSNQemPIY/JyzGGXbPivVcJaFAXFw8liXaoTbzhfC
cPU/Vdz9H3IZ5JgAlhJa4tpg/R+2JK7RwqP4w7DoVf7YanvXMhvi8Y7JBu0CtaZaAolfEWu9fhqY
8Z4g6QnAaQRbsJD/ASWe7Snl4laTfbLRS2Lnf3SBMKgtdt/l55K0+XCSW3PBhQ4zHtBeQCE5qaLp
PuJe3mpayWQDiADN2RFmlGbaJdBFpV4jhIiQZgQkwHd+Mi93SrPsxVTavvazaflG/zTEpAgB6VR9
HkYLbGkzS0wGtpQW5l6W2uQyvnwmk4qNRhUUqgqvNqHjb+Pk8XxSyKoOkzEnMrOjGwncphXDpgvK
Z9aToIal82q60BsqptAataubkw60ORRQg7v7j+7nygxywkuzPnamseWXOv7AQCBHatGqVodeaunv
M+kX/fMtG1HIb80w+3wSyAmT3dXDqMqoZaHSJtX1vbZnDI4mDxed9VszvsW0G0Ha4wbO1hpZAr93
MsP4L3ZcbfgNnyKm7VD/wmz3d//I0lvzchXSLJ5A/QShfb9VYwXFKqEClfh9EMPiy9C0bOracCq2
M5CVPKXc7sT8l2DWhIBnnEHKu1t8tGVLmiWRivTZ1uXcvTrX1chuRU/mMNXXnF3cMfoO38Plg7id
yzTd7VSwd1oxSmhd2TfHYZL1AbTMFCeJlbdl07eyuJkvHLmvNaXH04D7C+N+FeDTPHUXrwlb5jpv
a77Aksizrn+uDNI1LobfBROtqUXfN4w+sIFjE/xFfe0X4YB5d5rtAsRbc2tRLR4q0b13tlIf2ojC
J2QxnSZVKuR3iPzWxOTy1+5/anbDqjgv8hjJxLqt1Zxf0ps2KHFSpKlLXHsCCcjzGKm5IdOHAHb4
UUF8L7bxwAeF87898HbArF81Vud1awKboCSUnLkpRtdDTLqqHCEBCIjiIF1Yo+HWbm6kfJJnOG/H
hqMEZH0YX0FUyRB8kPnNlCA7LuqiiU9kXiIdF+HG6UdMZ5Eo/RBFz1vxqH2g/9uQVYZoaUd6WU61
wnkUkqWTn+yg37BE9w2gAp0fhIWbddo/1xsY8F3JiQu+av7d8hgv2yl0gIW4rLLrVGZdeC+cht3+
DmXCj5FLAAEoCtPLfl2VBujgYMcu34tNHgQrRZWrmr7TQguwPqvxb8wb/AgGEuyysc/4/kHR62DY
h0lXJJc13Cskl49KxO/fbI5HSgxxiBlp4WRCuKRR6EpWAKoBc4X7i0S/V3QYwtlsqFTJ87YQqXlt
fD3yoLQgrMDPywEbeKUO15+n2hzHXeCJGHYQHa9HpZasfhr9tjpMeNBsUczkOKwZK9y1ktsMEBhE
c7eWyapvIBsAWxPVu7L6N8YAZVtkICYL3d8H473oz7hf5YXVR7Vpa39W404dFaHfWNI4EZU6rRL1
+ifKTMOBnNr0kvqrXxBJG7gUzXnIwWLJiu/NkZTt3c7mBsCpsTbbtq1EdU418EGPgQdb5kFsLiCD
NhcH4uT5G9edaNTxn6TjNoJO4IEW9vKT8frgnrw7FzKuIe2LX3p0miCKMv6kvbzFd+x2PlJ6xCaq
9cuF1iqwO5YfOa6AKAb5jMNGuuPwzgnuVjln83pL5sV0Gfo/GuzH15uC0C5VV5hrRYYvt/qGgyOw
Ymml7MBAcNU5OAIbowjR/27wKaGqO1tpyR9+kS8XOD9lew9IjbDu7VtZhpuNrJfIBde/misV1plX
AmgxvfT6wMYKtPzx3DdaV0e3vGdHhZPybPT3CE/6tmmF7/C3H4zPjWUSmvAsl9celONgQychpibF
Rte36kf1FKi27M12yK6u1fXWrLQRQcKPAJaP7W7+jlLHs7G2ptXBRx1W2yf6Sr4x+HJVsMgJAhSw
iU7cbstuOo/v3l9cZSjfkSX8BIaetm3YMztQeaxUH99QjbqGlERduJ67Ii9Q8B/j49V/xm4YNfJ1
raO9kJtNHQlrxyEdiKtAWhYILPOCR1zv+MRIJjH5vLUZ4amOByiWrs7E1J04QQFOl4hyfqBGshnr
HWRQ9lwLRLdleMV3HsB0TSrxGfO3JEn4eFKSoAHj9MltrpY/NRDjE2iyNIjUfOrOPK/H8atRyWen
mY6tNbZ5nXp9+3oTg66o8sA1isSPYRF3nWpO3KJX6qaBWBp1FQDZlEolbmCOIWNxMeDubJUEh47c
3YHiERdTuB9aMnGhglxXTkqZt8kH9HzhRmwkiduZGm8z1gdjSJjtjMY3f6nEG55zSCJnHEv5lhpH
+72QZZsCfke4N8UD7N9QEFWBgZsw/2bhdtIgenx5WBuUpbr24g9uOpG7cCUqYF3z7ZlZmjIXJ3lq
zeU+/p+LzmmvTmWCAR/LewRo8o2A7s77kfNOIaYcvYGIxs/OyD/dOcpkDsgGlYjjpGjfWZ+0pPLe
2+HiNRi0KxI0GzBERyv0Pl+gvFOKJWaUvjVbNSeo5d5lAHK6e+q7H3OcG/Mv+NsMePb4w+vvAvSX
cjlDjwf0troQv3SrmdSWot78C3BsAn9Z/p5ePwduykcQKmdjkMEUk2/nJMrY9ZnYt0ymTRkgYr2U
4CsEZfqia6yEIytKuH4S/ofx2bRt8E47wkQcIWJS2p3epeVipNAOS5E0R/SAXr4SBijwebFCLhGH
hI3IJPfrUCExs3pgAJAphinHiOLA1qyJUGFCXVkIvVxWAQbbdyFIxzUAcANz7ssKSy9K/BC3NWwP
U3Go5z4rltcvKAaXrb8a/UAAmhkrCdFWprIYJKe331tQWAa5vlXOz/CIaYHondapoBWSz8zRCRQL
AF6Yp0cGXka6PBV+PtH09eyXUL3Kq95lnwhMoREaQ9udN1YPbrUNjc2Awo//daQDhGTbMWC3o5QW
9B4/tWs0Z++NRQDcdNMoD4xV5t1uk/5H+0i2y9eQbVimLZds7vRE5RxDSr3cZufyEXRhNiy6peIA
YwaHjyGRpExhIFFyJZ86oPQebGgHiSkPYbXa7UOT9QVatOXXGFk++LQbiZwNNKOIEZyKlKfBzQ1f
mBFcfJ73DTzrJNf6b9Qe02qPgQwW02J7hiWBENESOzatKUa9WKpKy1i4x1A95DiY/fImlk93v6m/
BcQdkC/YC18w+9TEebWprr3E6mr9xEKiz7CCYSfEaRtlVizWcOEleRHrnlbPiwAHNaG63p/FCjOD
AajXZXSwY2gG6+mTWm6BBlweJUnuEkU3NuqB3tCDigmQufkPOOr+liAoUPtMbhipH1hVCSGRGTQv
UNCa71JdbXWwIrx0Xe/Xru8f3bnYpjg/E7GYPGRXf05CfHUN3ivRbtFEdsv+Tv8WsBIF9qE+iaxG
1x3skBoUVaOJ9NyFEp9UvlojOjFJm3d4cPt1/SthOtPvlQqLVFGvcQvSmNH/Nj/npUo8bu9FonmK
7BUMycEbCLXpLHOa+sJN4Vix+qwDo4pN3iBajMSXmRW2Mbj/2s7u9X1+nfF1BmjIgp68SvGjh83z
v9YcOut2OJMMGVf1hR/gHc5sv/MHCGjlT17/ClqJpOxJz3+m/vEhscTD1TFkyBuPVU6F8KdYlU27
S28Un7NMRJUeSgOdLGAzTLC0pZkVPTB8sd/r8eVS2vhLGT6bHdMOhvrZjerbAzJAJ2SBv1zbfmH4
Wx/gtsvfkwskJGDR12mFHB3paZ+1tc5gZFg2zKGuPYCxUpNXaGGKuuXXJFxJcIIyLSdIQ8CVJXAM
0pWPrnjyVCVC/ajhk8cPbcu56dIS5oatTOzssL/z/tBKg6JjOFzcLW+FHE5jUK5SQMVOZVODRIka
fK0P/P69MeP6ITpd8KiratnPPUGwCxobftx7fl6DylfZlW5cTSSvR1aNAN+ZPbhzT6IqPSpKub82
IX9J0NgPK7C2T1s16UiKnTy7fGlHoC+eZxzOjtsRmkisAKMMc82kYpTboDOPLLeybCWFIAhaKCSt
F1XS616e9a7nF5zj5wo0RDG+2t7zrheLBYgRMFqzoZXuj6Wx8AKlG0araO6YLPZYMgBejc86yJig
VkMS5z7mSB2vqeCc2EDfkbSFbe/biXKK9SU1b9w3ZjCbj0UfWDdF5tEEBjGO3kSAhF/aDCYitEUz
nqNQ6nAq2z6DHbQmV8e1sM+mgmBct24BXVAfJMvTIMeynGlwiRDkj09kL+1OWCUByfiTxv/gL63G
kMC7kfjLG8eH8Fqy/NagsHDhuKUgrUN9hgggmAIfankx+NPhN7NdWo0HpPRu4bidFya17uWa3R4Y
I5ig4Snp8sMzB7U7zYKzwJCOuoIm0JeEygT2V5gYLUtfsUKwhzpzak6N5ELa352XW+8VuU/ficXP
Qx6xAFZQ41VL7+8OTl4M3Ut9kJvtR2EB0pw5IyEvlpdnRDLaswMU6gHslDVPUKrupYXb9MiyvgVg
iIbDfZKYbB8y3E2X2c6bS3XpiWe0Z3iI5KR8+cq4Flr0CaK1nQIQ0Gm2V3YEllDB75XPQb3Pqkkr
baO6p0bXD4eY0BghSo80H4xHVNQS2B51k7ZN/b8FDBynQ4sqHjqpY8Du5YTkNqMsPZ8xbeelh8vz
scSXPn0hGR6ps3RRAFwADz+qAuTePLuMkBoXx5k6vmm32gZtrfZhPXUIJEHuq5iu8a0E0GjvYqjy
Xss2PSeAxtUZ9TlLHRfatYayawB2Nj4LRjzn5NG3oU50rW72KgiEhHHl3HjtUfKfaqtEXbMYG4Jz
QpS5rm+YnIfHLkgvUJ+HcfzeEidka4i+NzpzP73jaZYHmVx1yo5AFpaLpBZhUUYS5+SuvFjfDGju
uKCMlJrDF+o4fEAfo030zvAu3LGGB/ewehfzzMFJC9ehA9nVm38QKH81u3fk/PmwiBhGiX4qczkE
93YrcKt7etr2M2pcNM8Rnl38U9eKMSo8+uai1fJ8diEZvfMy59xxX/3C6LNJeJXLjBEb+hWZCe0W
uZLpbjZjCgnNgcQ+13pcknfKB33r9tfjD/y+lov3uf7AUZfnI+fdROox1/uHGWJAvEqC+ivPsSaP
VqoMjUR9evZxHXODu9qASaD+8z7TagEGGzlBe5oQd+UyfPc88/h/Tz715HtPVCRMNXNG/jrdznTn
UHZU2Uf61lFAEgaqHPS5/1QIW+0LmG61SInVY0hWfPT5r8z+HwyyyVuWjG7y3miBzlCpqX4Auc5v
PH1ynnY4fYlYb+WUNo0ygjxV/oFJVKTnYdeIZMzLM2EQRWlgJ7Ewoy+qhfAACjIG3hxJkBuV5Qxl
ImeZrFSkqslyUhkRgE7LYysz43ztqEpZGW+eoxcKeSCcQuWWwhfpBtVpFQAQjEHuzehVlhONzjt8
WNPZEoTiw6dGh6grgvQg//FQnJ87SmH+tbMWfnCOT5ymAf7e3wFG1kMBkhfJ48phDADNENhS4HMq
b4u+8rhZ0ZHaRN0W1/wFOrbq4W1Yw29YAQ7J1mMtXTdJcVrrJeuzVhZGFqsYgYGtUpMGL+UOzEE0
unDL/6QKGT+9vIYBicF8ux3bv8oMTgpXCEyiBXRFYTEuP95Rdiqem5v5e8VnQ8Z4njlRdZ6Rr8s5
2Fs4VA8Ra2QZFBwAwmVTfq5MGm/CPYSgwlnRRnKU8i/b9gGRxq5JQv61Bz9tJXhgzLure+cn36WR
it+3WeG9SKDc1tB+yT7g6RKVhWsXYKrJH5K+bDiKNcr7hN1Dgedik1m9aNhVXsbo+Mk6/Evhz/2A
1TgOFxOA3xFYspqc/D85bR7PpE9kUiCH+tSj3JDvuujptfe1c4IwavwuMUlJACogm8+ZfcWUVrUl
wcuHyChiadn3Yx1gwidQj8s7TkJw41H42tl555zCmVHMbVJ8vXTloT7v5IexnnQ85pigaweXqZn6
oGPbJPHFPqi45aUuZCSzVvsEa1K78hOWhIB4elPrqqX0UZGwYUhMnl5dppqjwnIOKNkI//8d+epC
ZeRSNT+dFMX7kZxhScgLJk0exBcQU2YhWDwDetbD046EznHgS5/A6wCKgSPkzCvGMjIjskmP/zAW
vCUHsK0mLF7OVEgAJ91SifgqGda3eGwP39uMvbZsoMMHZP/vTsP1yvDtyyzsXhkb55rmU6wj/grV
WVJjDJxHEyiOOoJupoH8onpbQHasd+R0ODT9xOIqsO+EIyjhdEaOWKmNXciG9W1LNcv3XW2est9v
bVex2cb5O5AXSkSUCsnitoEp5ang2H8SKohyl7R1QJV/Q32my22F3XvH9+nHMWMbS1YKK+oq6QDf
LP89/gbJ/zz1VZ8mX3ecfwu92HeHWSQoiCNUsDV/mInDUBErXgT/7mHDfbyLvzNOJ4IZs8l3kmRS
6/Up9FWN1b60jb2ut3K/lrHEYdWQZfX/sSClA8ch+wig2fXWDZm/V7/QIB4UUNx6Sw6XbT2Vs6gG
YfbAOD7euvsPItgEQa5XJmUAZ0kfco94uOakEhTFNP7TRDxRCMJJSY7hDAGA22e5sh9kdOFjM9CT
QqcdADpwavUFaYkNffdFIY/AM5WAg736V/BujZ/CwXXokyC8HnHchwOBmKQg5p3vDGBVBB28JRH+
EJEzBrRR+Rh9IngAdAHS7heMIL5Jl+jzqZs+POSuW2vvgJf9qTYdG0WnKDtASwZ1GvwqAZK8t3Fu
AZxA4RLt/NiD7rbzr9hq4fu1FBAkXQuc1HAswViFy2TgQ2mTHpgDDh/KCuR6VcTq/PN1r3UrPlDR
WRft1LHUQKsT8xyaRbsJh1DPvStCGHH3veZqNjCyd5iIfLes8MSMoNIIKOhFz61zQhGb9ldKvDTh
U2ZAIZHEIYFY15IdkhB3p6KIPQWIEzKH+oNOnS+COX8QnB6Z71m9WovbmCVEED5Ta/mwMXxH4YT+
hxwQyrnkXfL8ETRWrq4UrsdN3W2QNsXgbto2HwehD1BIrZDaQTbsCQ5+rQ8D5JTk4rY7rblUH+bc
PTtPEMtSF/3l17N/KR7gsuZIbjx2OUMskAZwUcnKRw4NYFXPQJDploEia+xgbIBszaBlhUvzOg6p
G+TPN0hivi4+vLgP5en7XiFM/kYpgergx/LZ5DXv9JEoxuGnmZf0aJIHj8qv7b13x6na3RBYtpoc
3q3D2fuqXHeiPH+cOfKJWQTFqhPK5OxFOLj+v4QRhkdGifOU6+W6kl3oN/rtn8Isni4UeatY+IKu
iUBFqgLDlOYlO1tdrFJ7PsYIpNBz5rlVbR4baUZWPqaDmpKtTQ+P5j887fjJDQh7MtPpOafo+jhX
fb3pY4L9v0QGVXDO4tmEvmqCHZrqIJ732H5qJ3KcAFU6zm0LcUOljoNTN3supO/3HiQ6GprAviaY
m7bKZ2MHZRv/LLR3f3NhBjzYccVvu7ahnXpj3cOMOXqKn5wQqAQzQGJTwDXA+shFASOCDAVlUm0e
FG28q6oTlM2kRymbsxLAJm8mWZKLQ34stvCSxBNSwlh6VEUgD5zfpITa38XFiq480LPBbTJ3ghSC
KsGu6cFFl8mvvFLvARlcoo1KjXPifUWILWzaLMaVQmAB3AG5ywHYJD41neCljeS5iXpIFIG1KlRX
qG3a1KSnITq25nBkm4UwNbu69SMssFL2dW/wlP8T0dpU9/Canukl9jtpj2MDGuLH7omEEFebmsq3
eOzp0soCRgcJ8rSlE433DA+agXsU+o9iThCB4tkyrDhNhrq3VhTuCdanfpihWTodaK9aIH0YyLvu
nA5plkEm+3zGYwAHQsi8u15S21+sxQvNIPz0lvwURQ5kE0429f+9TdhgQgAZReZN7ES19qF0VuCx
Wu/FvPOe0pv7ykTKxvpQveR/l8a5kCx/ieC59I7wA38W72/WR0sUkC4XTHhdvks+vB0wjJwOuHb1
zebXe7FaWgu0AgC40b74QVudjNtvy6gD2WFWcQNL0QFy0TzUmrjT3UBt1LgVuSnprcJZolEX5jcY
qnWz58+O5RyJw5gF1O/Sn3vYkCH99uwNLAoUi+Un+gKmRxil+KXIgQUb+wN6bCKE9ZcJIp50wGSw
f+BnvDRGosRkuaz+yf7is3UxQsNoE/Fl9hHfSTixOj9twjFLR2mE2e1GELhNSKY9zKoVf6Ay96+n
w/XULQp2y2bC69KPlY/Ab249Vs9ZqDHD65r6LMEbbARJIPppj80UFgYPxrfKWlLTEgRAkChPGvTK
2KEuBeXTpu4yHE21EYvXxeYS+45YRNpbjJcC5NgYFGSb+jmgVokYyiM9O3jf7NXvVm1R8FGTzG4o
tinzgatng2iMxe20fRressCml5lUv5RwgIiXs7AEit6fZ2abqBPBRZsynQPlCsOKPtLhXrimEWW4
7vIEoWSeGWQzBjlr4IZ9QFZBmFiiYX6iCKPIM75bNzkMTa6O0Bh9t+iu2kDcd/7u9zPRwB4aA2bP
l1b1CSAN5N2iLJvcz9QCOPGQ4iz9GtLY5Fv/NbYTOP08t53Tj48EV2u2nRaKHWpZ/v3/JFHny1fM
lbpB8JD8RAXKDoZP57z0ZjMHB7NAoY0nlmVJPsXdHS9BMAhgbQ/u3iHR4a0pEvIH5/TcL6d4ItJ9
aVlIxbG1rLKdW95GwiOGu61b/ipn1u42QkVS+GZzU5QAHqgk/rE4hGEb4tmVQAIPkABm1IoQIoON
ggQW2CCTDn5XRS8yXGkLNp321CVCBhESrTnQDEt4UHC8wH0Fs0Ioqs1cXzvl8jqArncHmoCsJxWD
yoHj2OHAVs/A+IgP8Rs1LBh9kLsP7Pypmi13n8GN+K1aVonLPNfOSXxbhyaTqKyOfI9HYyTnL+YN
R9FNNkzJCB05LOy/yLGZUEZECJGUn+8mnltz5JNxdHQkw0HjwjC/hhX563wUZoO2iroYyC56S/72
P6hg6TxAfoNIkevshnyE0PJ/t4fy4PaNKJzWrHgPOAZnrEUI+EdIGZZo2zCIeoIqyZ7Dkp4jtyqO
BhMzvO56bU3JA8KgRcoYWqZW/vSiROmod1Xnr217B5DHv7/EUHYMr+IaD1ISEbmguYxYR/P4YkP7
MZFCBG/xqhOGUYpcB1+pe9AOg0+cnteDyEVUKMdPY9Z7LgrQtPqjxrP5QHUDXDGZ5xBv2lCb3G91
s4XcOCm0PFLUlwUfJcbssyI5GTyV5gyzGquGPWX2pmX2eZe54xafpABw/Om5e8Rf3UhLwuNmA+rf
4wV9n7l3G5rkbGMYTANt0xF6eDtYPLlNXp2kY88oj51kFeGYkY9nEzownX56e02HZ6CvDkWmPwsQ
O2twkOqa7HvarfB/Xg0UDwy91wayYMchJttdYSAgT/og0CCBFnzc1fyluJlCEgI13Oy0q8+LfIkQ
CBFMMHjKJQNcAXsm6JhB2yUAs3NFj40ibZ/ptwdgWyEbjucgPSHVurvzKfpM+giY25Jev1pfgk1t
o1+1gXAkYHaqexA1GLDB5Lrhk6MOTaVd+jxm7BFvi+YdKIowBAAq7arc7Isz2CuEAV+U1ZWSOuR6
NzDiFzC2Fv35G+6rtwljfkrL8oSA0x97DYzzv/yuPEIVCdot3CAVnD5cx9GoNaIEIlrJlMjzje/h
8956cYzvu2mTSbxaaD7ZxwxahDXGonJWPqgvIvQPj+a7Z3pqNeuv/76nhMMLULHL7bOIebQblzx2
NunTUddMgpJA7JO5pR2K5DSFEG227Uua4k8no2FUB2dS1ESXdfMbzngrpnCiyYKCMeMDIn4T/rVm
7yk5puU2arJk/+eJB+QZ+19SqWK3p2rGPQrBRVRRkqoxTSh59kRdN/fm9o8GO5g4gkABj4fUrKed
GNws1uc0FHiyGUL5HbdHMRxalwq7d3oyF7T2g+zRSg0Sy03p+AdgZPAWUm+9IklHpzh82dVTdQXf
LriTHKWR5CstgOr13Jj1t4OolZhVLPbjlnWMDIsfNLVDKiIUbMSI9Ro1NqbH+MaeASSCk4+ngKsA
ufTFvyyXAi3w36ybPq2r3dLp5Kk7Cr4Au6LYTZ09ec0eTedpQBWpT23f5zhrRkT9wApCwvwW43xm
Lzj4KvXQabMQe+XixYbY9tB53wuzDKycliIeQMJH2t0RFeqBFzIxmZDuHjRbzNgo16JJ8QQzrYSx
L0Ple9QvhtBqJV3lWgmzepi9V4T2CaL4/nh7Je3jvg+WC2jQLJ404kBVzAswhy9+vPeKqUnR8udc
M0gEye0fQW/8OA7W0Z612VaL35NA1Pd47DpcnNN2Ol21Tj+5Lhxopg15jp8kydELRi6xFqJv0wov
5MI903mmCC4+ODfpCY0GYcvv04WdKl7J5htJo+e5rPT9kWO6p1vRdyhkMGUSlp+0ljhOz572FsCn
JzGZ0+vg4pFcfgSOjkQ5szWV3fEZokUWu+8ve23xUd6ZQzcAliGwqEn+rNrr28J8o07XKbKgsAHY
D8j7bm4SD0iGfid46p++8suAtbsh+bls5i6bUEwAoNfKgLgZ9YkQIdA9rql3weTxIBYWwxeNbD2i
8V/THQN+xF52YHcbs5/f4OnBYsfPUUkjbVjhk3YN0d3q0KSp5zE6oBbxiOMSAf8uuq+g8AUAWzMh
/ltrgf4wLEz8nGA/1KyDoCo4xLX138eeebf5mgtYSM0kGMfUCDX1k+34UWs1Rbqv27NYvS9KYsZC
bohrl6cVTzMtKTnwT+r8fHm+nw3MvtnbFMnLfmKH4rzpK9wIFP9bvutqjawNkfHhvIIYWF8mppLn
6XTA/rHkpafM7NMmcj1NKxV91LQgod4beIRW4HxjqdUtXN4w4sOwsToIyWAR5GeG6bVGPH86He2a
76BIvloc8r2kJVqViWy2pu1R0TzfhttoqMTd9k1bC/B4lEpNimQeGmja/ZRofcozUFl4gXRU5jYc
jxifVOPNX15WG2DcYmi4XoqjacI7g0Ibl+x523vUSAuxjBF6YT0uLwQ9CKlRVNLqcqS5F5bVCmeV
k6lM71hHaLghs0hDT/P3tUfZN4b3ypnMm9+YFDJ1iF4cPSwEAik3rKjhj60J9QPnIFq/mzoCC15w
pGdlV1P15s8aR2sYIyCfmT8aNeCkPr4NuGNMeJiyAUDTC8V01KGDstjnizpmJSXCCz5SeSjX0agP
kMKGjrbBXD9QzXMJ4J5KzC3HSRF9v1mG58kB9y5t9caVSmqXEjkQXT5WnjZCzz0fzrGiXlL8xgZM
YrIbiR9QrTqgGoTn8EYJ4pFqJn1GHyJiLRq9OUAI7QT1J2hcu9UC0V5FH3/NJ23+rGVkBvWRv9Zl
PXB5hOltKzjnAG2H+X3+9/Wd14nx0YYefTCRuxuXq2GoWBsvOfIHpu729uR2gcPzdrV1usYEHW9v
6BUhakEBygOj9xAs9AkMtcZrOAekzRcrTgvrHhdkBIUZewUm6lBYK+jMBUK8fNhkDu4g+KhmG8Xe
j7HFKUKC36h1yBuOKQ7AvQ1ctCvbzDLggMQ9/+cefT+jRSu1ABx70c/pfvoGvKuIS98eKCzNAdl9
4NuIfdqTUAKPgsh34ILpGvxnlmBtkzIj+nGqDVpn6Ilpy7NaWr25nc/RD0dPPsfBDuU/pQQfxLJ2
we42iKE5NmL8/ru084Z6VZ/CMAowuOW01ho42C/+ElJ3DF+WdNTfZTH5F+5RCD1w2h4qpftEvJDX
wrN32FMlsIkAAB4Lm4kQFHtb4/47hW2ZRfzqTqikRTmoK8Z34IqaHerRfsRn3vYm+s1PF2QlGKNk
OpD33Rq74PQ1mRUv12m5NGDiz9mmW4fWvS1wCu4SLmWxbt1Km76MQnzODKLr2QCkU0Z34if9CGS3
UM2a91KozanzHAzPkEIE+ra3PZmqiLIh74leGpbFhE2IcTwtBgQI+96Q+d5wjAAnD5/J9YvAr5o+
z2q0e2jxO3toO+QJx386VkvKf5P7N3PwPq4bGjjO2Tpl90fEYc0xFZ5Ww86UnQC8rTPd7gc/KUhz
5yAR+C3DGhj3QivDGvECybnRB4O+4nPwGHSHDS4CVwycSWWtzqxRcTWYGqsz8D8VGV4ClLbyOypg
3vy7DFwdHK/g25FyiX0pVglSTO9mJZWq2fTpusp+Jp12X+L/tMgs+QzOynr75/J5e1WXjoFhkdaL
bnQdHauoN3EctREgLkw0ZJhrGem5SGLh5QPA3prhwvViUv8b5WBkMtZ59rYVCbMOgLNlJcW5PT4C
aeIyg/e9bod7pzg2jbMHBBYkz1ptJS2AmysYmO6dzEJMP9+/QysB5aldVRDHUpekBzNsiCy0GdLA
dNRJA4CSJs9ojHa0GNxXzIVAw+Q+4qUm9EQ5TyMQf2wNKmRrBe7tEaQbB/jQKQqrKJAn6N9sVpC+
HMmjh6WHRIqbD6c3gvdWN57OY5Cj/yj47Y80pYpHyjdbzHbmoSt+dI0f16z/o3NzlT0u2Na7nGjQ
3iBaC4Cq6ku+DjpzsFgxHeLw3n5yQt/obfE2iDvHpgt8Hm3qN/J+9Pp/ZO+2SUXlKGimCQfmnnVz
L6FsBzujvXDD2gGAHAjVR9tOXYAMrdOQz/m9HYf7yb4kLKhox2cKwoQT4P1egf58qUe8vBaXxCHa
Wg/ZcqYOohI4vPt3nhnCggi6I9R4NDx0/31FbU/cF0fF8R4X7mgcb7R/swP8L59oFGXUDTOadozK
GqxKpMlkiSt8gJzb7gG6BjpBJW7b8ZU+co1W/uabmMh/YtJqbOJWLWjxt+01reBmaPWva0355U5g
I7mvxJ1a0gxdWXVGQAq272vTMw+jlU16jWcNcsEcQFBECUy/tNyJm6T0hAiSzUJ+CxBnbTzfT0T0
tWy/5BWU64uglkIuYP7HovEs8IVpnnFui2lCIwKZX74fYM0onsAzMQVnoQyfDYbIKmzd2nnyyMwJ
eb1s8DJbqyf5vlXxRPYqjp+vHiLZTCP6d12wNcce8OBQgydSZGueJfY1iYSDrjhiPzAzg94alg2p
4xdayGaalhzz8z8so+sTDPgFUqrg5U72GndSoe8uN5GoPFsxioHDwv0m1SZDZH7Nriiuj1C3z1zt
Cfc/ufTpS4Nxw25rPc2XuZKPaJsrGmIpusi0IE4QQ4c210Cgitdp/+Dv8/kXx/eRZt/YbBVoSOGH
ofzxqkVQ5AVT+pYx+HqOzr8bRnNeZRjJsrxBxIXGiKZ3Lt0uis4mYH3fHxcNAXNezZM2Jn+U+HRx
LEaBC7o45AjZpoXk8b1RqE3kR2F0NFQK+0yHHrF67G+cwj2dGUqcUSU0qbP3k8aNpCYKTCmv2wvI
438U2XLi7zvIUt3/6ya581rfI6fy+wLzTWp5f77QNlHSTmmawMY+WPhpJdYWu+YevnlAWh+4LKHB
4SK3Ss1JrjEAtDcQYOWO7uoPlnl5J/eIAXNvwfI155rqBaX30ASzv5A+0ML22zwvC3mZ53YkvwSf
5Xxp/bdGLyWUm4VE/I6nomRJb9Zys1nQwlAG8Kc6F6OvZK364CXsifyzqMpliCdQGAkF8BqSjUZD
IVrV8xcm0MCeyLJE/TIsiZLdTfTbw4brmfE3IysHJEn7/B1MeG3Ybc15x21O0M5GTvAz/gwiY97U
ltljUuOmfAzsRLzKTayPO2fcuIBEpjhKmFE+Xkfki5uez1OyWP3QP1icv15YDBXWWu5BEZ81/hLY
HYj3nd/EAnsntpQyhqozAou+VaOoDn8ywp4mBgCT6SSP4wtNZOl5V63ZQRZViYuKHE/yA3xuzHrY
slXXX30L4LqQBAIbM9rCVfyjTwm9NZz+VwPJec5XZrN//n2B4UA+EFfzG0xVu93LgGkjzLPKeJS+
0Dr+qqKlz1zpcW2burj5zCh2H0MZuXNV6rllfOWJob2Dhl7lq7IZxSuMYkazIIH6wdcRxqKv93nf
CVi1y3HCDb5GIJBVcCkyVKnfkbZCafYgm59HRvDq0OCz/rjAnvN19R14qgCOqXrKbeY/Path/0sN
JtZFGMHrrAl7xoAzGSdfpIK8KsnRWfYRKU6zaijDSVGsnQ62etlnHUlyHA852BWvUkpewpzTubFu
EeutgQJ15d2xaZLY54cJKA3pjlknpm7HYsLh/VwpMIgMJNpXEVvraB1Pp0TFwgF4wbXu0V+wrnGd
pPNVXPLpqRd3V7RvPuOzEbTsC0FJE7PFuMtljdrM2rmDBNUH5ujsCqicdTxy2BrcDOvN04saPI1Q
uAZlvy7NWqp795MxFBBUEczqlOAvrkDV67N6FL+n51LoCQmTUmLDqrhaLKW87AbnZoEz/3krOebY
BC+riyuXecY4hJ7patAir+OjIRnQYqSINyBMkxLR1Tzl7IGrg0vYdD6a28zwW0Km1C/NB1Qk9JRM
hyYhMdGLQTa1NXNFAzeCPerNFq/KWFIWtK5ghE/N5r1NkFRrJQSLjULdXWN1NY1AEi1AjFfnH9Al
2B3YKCVahZRQRYIib37ltebIIt/Tcdxe3ajHpyfHmga0OCougiU4IDLDh7heQmUcM46ayM9OLyP9
YUD/PMYXylwIIy1n9UWzbja/x5x+KRfydCTWHpEWzVeCHLKbpjZsR/uagjW861dQRWAr24fl6a31
dLZmLgu5LryVtDXd9GcphYhlVVM9gJaluUnu3MbRr+cIZnKcKDR/6v/QZyXLf5N4HQY7BEY3gkg4
36I4beA0TckpgWJeD+vHo3q37dqAu1dUs8jj+9kS6zBKOuEPjbPluPrtPQN0OLix0AUBJb40cAkY
7P4J2M0jvXMONAgLTLJTTGy0pGxtgYLjRmKEBpmcuPaC51YUWNTNxMyyvfUzSrNGmzGtpHThFGQY
WlcOPqkjW+cObOe9GOpnWurvbY8Qttr9vCmhxVq1iUeslLbhXGUPCtoNuxVd6VYj+dUUERwZc4Ml
TEMgixYYmodQIvW3Flp9/ODw3jcNNkzdayKf9wzljeLWN/dhPIFZ/Nm4AVjsIKsz90Bqdin+wQgh
iT5EIXIyS3Ojli1Ar76eUvUaXJB3BBLoxvLLrZcBH4wXcjyNzUVjqb6B3FVZ1H4dwbbHV+2Krurb
taFf5PPIx7cv4OkZZVxgIkxOTq17IO1A+EZ3pmNmA5IlnsNPnmyWvbZNGnGlAoDrRSJdiCTOphmu
2WITL6uD9Cc97pwglhpBu7jMYc8HQ9ZHiBIP8U8vUQs4HgH+FQr9Vd2yHiaq236v3bQbrkPRn2QP
B86tCi3URTsy3ugHi0GHDJclgaXkTRQgT4fe/ikL1ckpZv1Qm3gmo0LITUYViYMExTMwr4ztdqg0
mCmGfkiWK8iBVIp1kSl0cWX3UilQ9cs+sd/0B2+wUgZ/1Wa9jVb0OCrfrQOvVVNqO/szR146UaYh
skWVrHfTjhGje3hNbKAcb71tM+A3CEkIvGhAzgMczEaqja/G0pRgcR7PhfBtQ6+xxNErFIp6Mcwi
vRUPFh1FO9M635adUYUpL5p1YJ0zHmxolcxrOdaZtUbcPLza+Cs2bhGcaeZU0zRgJ2h4doT+kXzf
rZWxHN3WQZMlquws261joqNopgmOpiSuVBWWNCRjoJLHqPES+2T6V4u0jGiHyocG0rQOyzEk/WIo
sWNaBo8mIpgxJtXpQZxjfS4Lc6sKFv7rRokgNwHce9qprSxXwEOKPgRb33JwgPCFqjcHF0UC/xxl
+pIW+AMQ01mbNFsfk77VDy2uSuGmIV1habIpnrthJ98VaWXaZPu/1VVeeELfZ23YM9wgcwqnLYj5
GsmN/4omyXyjFN7zYNnUeyOE5DMyRYkqRAlYudAyrNjk4va242+eZQ0BPH9m2cDY1MCsl2lQ/k/A
2rSy1tI//N3GxArMZnr679YB24xDxl6cp0S8EHCkUupQNfvaHoANVxgRCjZjO/A9xifDaMbm9NMC
3HVlH01YFmzhjYqsVEr+U4y914simjq8toznSAXJD9ndWuKv6bHo6P1vEuP+tmQEBVilm57Msjct
NfNwoWu18d3eXgRWsDRkSpzpaibVfjByQBkVPqbNsMTIe9rp+kU+cVLVrxQIE1Cf3xyL0ljIy6kN
5dRnazDHWSRzWRNlvE0K1QIZ2vMF8+Cvx+jord0Mfvqp2HoxhyXFE5s7THAny1ML7Yx11xcZHUlC
VSQHf8b1CdY7SugQZ3YZJJ8no5gZysOo9Y4C1JeJKwufUPJmslnwhTaorInP5gdKP6HyC/rckgK6
TzeuDeTNoaHWdmy2RMEGsaCuw3YuDNVQ+3e+TYX51T0kbvkJX7Esr6jMHWRbfxmYpP5hCVVWwGlN
ariN7nXUJULekJWoE1c0WMcvg6fvYWGV5dMWEN7CdQjLufzwf4sXguTLpFjBaqvmQ/wEYBIC3CFf
wsjDuLiuJX66IHyqueZzrMN1g0+qk5Xc9MQ8T2JTVMVEoo1uxvhFRN61Qs69pILofpI+R5oyPB69
i83IU1JMxik4lSXNjvnHXGKVFSiu/dHaQU0RcITp1MM5QtrgwZ7CgDFwNbNHI+FSId+GFB4dNkVn
Zv62UxVUbk+VIBWWJcrIzHBFftY1OQ+CELrxSnU+KLOXqZBIyEkvEu1kfPZDaGfcM9fM1hZxDQ/J
kPrKx+UBUnPhnm3bpOwgRIYudexehirPGkYU87o+Iu4y4D2pNkWKWzH5avIXR/QjFC0tvVMU2rLP
i3DIN0Au3cYsO5BY5tzflxewaTYMTSul10g55TVvVb7aZZeebgpt/Dj+G+ZOILKFuEZsuhMkh47x
+K2uMMEJBQfvueNTOTqVdSLwJyxr9LayPkoQDMIziOt3MXu6EgLSVB79RTqHn++8O1zh6UUnP1Je
9TZPCCUMQt6B2M3JUYPYxT9WUaWWth6+o30OxwfnbgoYl1IF6FM+JXu20QN9vwWFja/048ZPikbg
M5iC33OLwtSi/nSoVPm1Du7hwZDCU+oEnVetFPe1Za+2XAz9RoH+CahDEPsCYponS4ZpqhfH3KYg
ObjydOiJBJquvl3tqQm2e1nvVwy1d+dsGPiwYAVWX3MSyVdwHy12qbNwwe8htEi28DSxPlcfMLX1
b3qpTFt7j7ZM+/7SfAiauPLxpCP837bUGsJQEOy42qMwD/1uLmMRcOgMasZBdy+6O+zCCW7HFZW6
GyeekyQEO9y7cQmm63AiZC3Rg0HlC+4I0g9vPb+DrjRVqh/pRr8b8UQ9nRb41ESsSxSA1FTlQJBw
myYXBk1AQM09+svFABkRe9UWXsPcosgpuRI6FJoYDg2ITgmZf99ShoNh7rxPnj8XVMwEchu+YOF7
gtmbBwercn1WCnCMrdrDxEN+2ZE8ceXJQOSnPtjq46B9XvFluNn/K6EfNlW9nkrGqsUieS7sMGpL
YX9CHi33H+vTkVP/6XS0Cdqz/4a1XtBanMn8O8NcaN8O/hLN3emQDeTcTi0wPp4Fj3oJ+j1Bigvj
tygd3fkqeFPyE3DXFUswfkHh6I4Be5Y2/2H0In2KbQb6bZ9A+CHDfcmj/E56y+mkhk8P6D0kqzXK
A3ZYtmpoHIgDIVTkIl6id7XAdc6lpSymnwtiV9m1UniT7bkte2w97XQoy/4QhX0XavPluIU2Zxs8
HxVpqPUKutqoZH7waEDVyQG8mT+HP8H6BZ6sFTIg1eWkSlsEJIHN/ChNvuLlCKaBmR4cVa6Huy3B
uahsc6/8audUrABqpzHBOZYIjp8B6MZIj4FmsQCbtvKGkmjlHCBHPBkAsrnb8O1Jl5mF0Gd8PDBq
mep4QkEI7+kS5++wbiUPX6KQXMkxkgmukNTKMwB4jbtum5qbIL51tPQjc0MWNAaTkWdjXQWc+9Mr
BneliPphzqw4ja2njxR1JFKIYmENxjWB2A6OR646qzFhUk/+1k9aXu0CpFV1tR8Qzg4O6x2Xu+VJ
wesss5IyKpKHTZgEGCjQ68hQxzltl37BjL3WubxhJcjGArT2LWDxi+yklWgSr7T6DKVGfvxmcZFa
bCA4R3hLHcxCWk6FcJFS/4NXG8ENf/iXMno8PeGnwmf9KXov1c4FRLQvRvvocYWUtlE4aiQhzFO5
QWunsD8lozBIeOxG4e22eDNDmGFSAms+qgVGLraJrsZYW6vnNvGxcvtynU445B3b3gXyofRE+wj/
rYo61N7KF8YUNvc0FA8aSM2NFmJ9kqrq5xEt18uy4ZKU838+rzFPdgy3T44NGkCQyajE/IHBp+ZK
V7ux6+UZGMtrQqbngvHLr2OzTqzno0f2lRruJw4oJMmpIHIBQBYodNC2IKYuC8XMOfvWihHFpNxf
RSIa4flezmhFf4qbcoIIn2lWXj8NyjYGT6gDvjzP+8/jnRUJPtJFjnaCvR245TlXuv+8j3GtAchS
HEaP2nlHxNawFTol0rt87s89X/fiyjjrRFS6o5wPO+hQlncvhQOqBOD8q8+B5ozqldQx0BO5jsll
lYuMBUCVWO4GZCbLMpdEaNJiayEsyS22VzxMhIfkoGRb4oeAdFApuMfVA7yJTsynwywB1MfCmLNg
ZqfeFymj4vwekXCL1GPsFPG8pPtxsy8i20yQp9gOuvfxHEVDliYvAbXs3TcdGudbyPOO+zJchRaj
TMfm/3Z04c+jfKE5BXGfHz4i/zK+Es60He3h+IoUTsrsEbQ7WpEFUmGnkV6Rz/20Ts9Zv7ifMqtS
AjboFBuSWVE/jJfe3QOGcWiCUXTxDC+9cj6qa/pkz8T1R/D/X7yfLG7zg9+Xz8jPa670DjtF/7o1
lEW0j0naxxPtJ4aHorzPVWst/WP6oplHU1NdbjB5SLurRStHVbN93GPv81qCMNnRpU4seb/ZScsE
0V4V9WEPk0wjOJWw9e1HauHecPUXZ8g9WN5XtU40Xu1wcbB6CdrMjaM0kVi4nM3v+qvkAd6702qs
MNmNr1sd2bjlYY6EwDyYvhW2K/24Is47Q+H9Me8fu3WwLEYc6utaqLA/eGmHmuynUiRWzzRTBqNR
+XvhELZAzfRWsnFmse1cxnpQtmIavakIaii6gIBjX286dgfYGV3/O2Xo4eVXxB+oyXEKX2oqTlfY
WIkOmzAoqqa5X56hwuUkHP7nNZeZM6xx2ml1CcLPGtSkENGp3hccj22PGtOOAvlX7SFQpnrNJ36F
JskdAjXnN+Vj0Hrmvj69ePcm5t3+xNP9GQbp8mbKsYbbK0mPqZgnSCslP+bsCl7QdiHV5zfd0wpn
zbThGTeyaucs15lzGL6rTwCEaaOmrwmeDKbhJS9VyftPPhrJcyHPfcVW77irnvuqdP/zjGZSkFG1
IjDGGQAWc65peXdYuRA1Jxt6FI2eKuZlo60dSunpu3weJ7WcckVh8kM7Spx+D4LLBsQg4VP9/hKf
YieEPWWL5ErBHBhRF2+K7KGPaLYFsYGvQsr+8kB4Dfn7SnxXvPhgg3MF8vLih5ELvt97qYTrB7tq
g9CJfwOswV27qD9idzR61+B6vRLNPR22Ei5X64xXgKwGR+XKwIx4FqZt/s/82EzOSagRzu3RJpaq
FbOwcUX7HQJeou9vRp1+n4QvTP7wFWiK5EIxTN11zcu8Sc2cz3wioSrZARfnLuuk4GoUEDMVd/Kj
QbN1YfqClc3Q0VfIE/KLhl8tmeGZEBL59zvXrdZ+KNI56TrDQGoCTEqFSBbqT4DFh1Sy5hOkfKQM
+dFozDPcy3+ylbLYVsxceoxZWmafrwq0sS1RbMTWJ0urB6wmrRMa+gMI1vmyDSlKl1YHNx046Wu2
/1K5EzeQUe09AQ7T5aVj9tI99ZyG5Gasj0RS973J+hu8atzPzZC0QacLVXaTWql596Exf22WARxu
pkJ0q3KfgBY52hxqpX12SzeMkWKLvFtFYqS/dtlK69ClrDQ6ilq5CauHaZsN1Z7cGL6yE9bqym0h
r2FDqyBd7RBemUUiAILwG/16otIMiwfsOEuiOGKLEP40oHb1Ymt/y+SeTvKy1usV2B1om9eYt+rh
o5EkyB49wMwkbdI6nYYa/ttNILtGS/xVPqjtRrvBBMzIwr4tKTnYwUY0/N2GlgNlsQWc0A8pdfcQ
6iVDXkpOtO2H1mqE29xHtU0T1eB3CPITiALGSDgNilwgAxWsEfurwQAexovJjq6iRxaFrx7KmiVs
zXUho+7rsPci23jRIRDtWp9UUxUGijvOgj50oudqiSsG3MlcnzWMmYDpF6UpEn4vlsBgyUvxkymA
f5GU7GCg3N6nomDX35ZUsE3CbwFxH6PtW/pxaq9FvSYUogdI+1UiKYKiFmR1Y7h+JlazYSBawJle
idO74htsUlU7pPnYO7Zxe9W+0ewp98wepuXR6XWcs3HaUcNdFGuKpxHm6Lgm3oBbthQ0ADUzxrbV
b7gg6COOkoLmTe46BtCLJK2V86XrHUB7WkLUln8cxwYI1/6zVf6bIlTMj+Cgkr3Tx+mbgcuDUdn5
wwbFpqMUb9yGDdRDvxxHJf9I/sTG3zsdIfDNq8Y3KTk5jFmpFrWd+L/0/j0SMPxwSg5ynSmLCQsu
b7+9ye7JVFQSVoIxy4N82NHxbCAjyAcQwCqGDSJ9p66qvrXM5XNLkIasDE0dA3t1d3ujXCRVJfRh
NCtgeKhhlWoUSLsL+sNQ8hP/qVSRJ5NiWtE501G003SVPTo/E8gG4/sx0TSVRcy9r8Lv2Hc6Y2Mt
W+ISEaWJ5bsEGp+KapQn0WZIp1+J2PShXUEZI0QQfq9FA5OGMtGTou/CAlQekboUdfwydb0ZG15A
HN+XcX0JJNuMCc2IB0osY9yO4cv/e8wIQNMdyMy616GHCUjt/QjNwY8ImN+OoGuUCdvc6lWV858i
kYaZs0x3jBgRUc9Zy9/3GwQ4eIEsyZRh/uwLtNZtksPdGcN8re01d8DiK9+kX87i6STEJnul0pG2
4q3zCvRH5U5830Hluj0/rz9FYZTIjGnEJRp3dCz2B3Oe7kodhlt6L3ujpDcEZ5cfA10+Mha8HR6Z
AJVjabh0FKWtHyawZY5/sWOi98zYmwcxIvduC/M55xFGeSLP7W3BeywaLq2Tx8HyYPHjsz1+ylUy
sDMauEObymCeML8PJXWdhcxUleNbd0tre6s/N9GoQwWygxRieMxbKQrCpM7298TgYLM7aFG6raKj
nK/+evqm1LkH8hncJyf8nCoQc/IEhuIJoSgDp5ttbQBvy98wsLOorVxA6GVe+6PlGImMbamiloTm
IBjrFMXsN3s9SZm+oGFZmLi/E963oHKIH1dvGf8YNzAoxDn/ImPl1ia7zHvnonreWl2MbZc2g+0/
q8aJM5cSkg+p5aciC8x938JtdWjbyYpsAstr+aDiOZnu2M4s30dEWE0ZfhjFms/65d1sWxJupBLL
AkWo/Sanye566V+h13S40N68QmwVhEEow9xuUsmjhaVslXaszRXlYc6EARG2iqeKE2e1jPSLz4ui
LV2CKhEKRCl32QzxZyJbjzbz68grje4BvbFihpgDSRoBJnt9E7Ud49ZpjrVY5sGOjJAUqgmdvVs4
ohvbfbmyEqWtcBu/1YdhY/h23joyRNIdQnrjRt2nhxOBO1stkTXKHnAUem5opQO00RUr5YMMueVR
ab1Q9kkbkfbYSptvmXubT2hd7N9LCSP2CL/8X7/lpWTJpPa5h6EkqAo9KafNGAeuJG8GAb41J/Wf
roDeviHg0BGGJfquXQH28p1ItpL67mkxD/zFaG1WLZCW6U+y3pWujGkSzRpuvxVpWT0NSk16CMD8
ENfX2wJF9Kq03znep8OiEFbJNhb8hvDXJowaYY9vqY3ue2XLp/af7rpGo/1gm9UV2+3ctKW8Z41G
hS2m4bWfjLV3+MYmLMWfQ6qgQQNe/Q6iU0ZG4nmFrOuF5P4lLeuF9AxAPVV8ANIzbIDWyYPNABGk
u/NFDXHa582xc7mLmUcMxFwfNuVB4fkYQJ9/58VX7Vl7xc3OQ0dmqRr4r9GXX8zuAQH52zfTexEw
ro12MRZXIcGGSesGktyRZk3cmj0k+Dwm7Hn88DRZwYUsDcy8Zdth+SBvs+RWUMD58BuR/VFr4V9n
fX2hYHtU5f6KKfvl5iMuNT1a5w2An98WqpLBgMLh+bWCE8+PcHnAYiY4poJWU6gsHUIOTGoAWf7e
qezn9+BeTVWj3sbqFL7JrSFAur64UC1yjNdZiWmZSVYdXKSWO5yvmgjodwP6sjK1zZG4oqyyZtX8
NndL4ZY+LDjVQAd+z8ayl4dvbNnT6ywBPgR4mO7aZhkLDnnNH5qIu/wyylddGxu5NqBoRmyqXva3
iqznYxXyauZk2GIhXRmXqu3nw7jY1K9jtOta2Ij+ynS/KHiRokxQwTrq3wQgnieZOaFVZAh0I+0f
pPqJTL++SyHQcfZCi3Qa+voDc8VhB6NxApw511wKQCauWsKnU5bXbxO8THK9Yp9g8b5k1NbPJFkJ
kjhCx81mZKoi4P8b9u5IArMUKu1k8Px3Q1o8cNDxn17rp5tsU2JgPAfy44j8WVP14r6araagiJhp
Gp1PFOWa2pXJD91ro7tWzkwq7tOIrR/3NesyPdHbJmLkk469nFZoKLkR+js0paEGpwKmr66y2I8c
P1uJP47ctRkC7KLAnzG8/hmqvNXd6jPTJJ6nF38xiWNSNMiF8awx9bhjdUkbiI3C4bO5jYCxSF8R
hQGMZMjVUPdM2h17ys3vU62O8TabkSPlS3gDtVf+A1Y0w5GVZojMYCgKsbpOTpbIuUYkjpnQm5zF
4SDStXz0Hq16+1d7KGJr00HOV7saIk9TX73C2WciBsaxXEJ2wyUhC4kM+LFxbrBvdRJ9qUL3G29/
nRURJeEbtr8loxms96THIbmQzSYd1GAc/NnvksNBFMt+MAGVuWWnPoZryltp418dxSjiLk2bVsBe
Pig5zv0t8XaIM648IXkI/xuDt+DT+OoBp/lmjUs2GK4ZTtnZ9cZaZzcOHwTlgtLB3o/31O7uGcPE
9Ra+yyOL0YIPHumuUtYPAYtqKPaBdHGGpUCjHFMviy1FFHynWxgn2vGeUKsR8uWr6tO+06o/2X3E
E53Be3ThVKPjI47JM7bHWhjiFLG017Udfr9XFWwGx6lo65uwhiqAjVXPNukFp/sh+TlpqH77GTLX
REuEjlpwV+MndB4ZNYy5pPFTjNpzxw1/YrkM4PItYRBycjUEbu6vM1ve14Hm0OjW5MgUsTkmhVuT
PLGuKb91df0I1VpmggwiKfhC5gJomc43NosVFphDOrM6KsCLS4DaNNb7qNl4hipbAP8M5EpwWmNp
Lvkbuc3kqdaNRe8OcEzuTEtSYvl7peHIt3VBz7HO157F4t+0JtwAevuXvnYB0iJ7BP7wjgIeZuBb
wrLfZihEmXdGvD4+p8XvYDxvRP2xZ7RRqByCYuMqYT3uGBa5bYqFejRR/zfS9YUvd/7UaqCLiuWY
LquYamsduhZi+mrIOpR4tlJYjMb+gW4oWV18AxKpqiiJYIunmXd4dVAwgAYyxyA3MKcRxS5t4+iS
jRObhC4QnyrqyajzxEgcwucU0ZGZLhNanYSS6RCUbRaESO/OunNkT9ZWxcAARSuVYeJZLEHE1In5
yrIPZjD5U0UMdZ64KtMsjVGLNrhzRtQuc2c+i+sL6Z6SERYBgp1ugRwdazv7YOui9O7MnyjWDJFh
3wbtI7a/rjja1qq3llFti0okMA3sv8BF3zjtX9eotuuT8wa3U4ica+M1KmQNX5jtzZmhg3TRtVnm
ca4vLcf7S4Xt9Z8/7kOqbLNBuiXgTEjFxljr8XNzV1iT4tjKEcmkWLVKWj4foqRYhM9FO8bAuC25
tG8nOk4I9m06bGM7LvcbXgjK6njW6ZBx94ZwkIiGiPL9kEjrMqVBAq1vXlLEJyYdUI7PHyWgCYNG
w/dN1XnaMt2miaC0RS+Jp9JFRVzlxBqbmm/UshgqKmWuXQd9GJMuNzZ78fz9lw1Ht5UhPUZu/M2b
9IkzFTwyjf5Rlb/yI1L2n+SCp2bNDvNb2MPs5M5FSwSsggCwy4nzq+78Mqle1jCnPlLifzFwej9e
+EwSFOz9JZpiQp9iN8uprRDCAHMLXJ5wFqd52XEsSm1pPr7suBr8vAOLtd8YqBz2eFQylq9wu4xU
UjsIG44S+JfNcICa0pawT/BSvM5sQxdoDowQrLfPJ02kPbWHkslh8W4bImitGZFX5/DNCWeAzhjj
PTI5Q35XbLdwYwDEM7iUhzl7cwdTP9MEV0d2y2W4jYr179bbNIoAzRWzpwsjkoMkf+EL/86jx02Z
j3v/E1ng/fXBB19WY88NHC6o6ACsGv6VnOLUZsyKSL+qHesk5o2AAy1rF9l5STj67i9mOy1idTvO
DyOtEEkjHVnvjR/mk0Cx8OcQWnFb72uVnGhN/as5hwEW8zBHxtccGRt5k6iNAGM95yn26Bn0lBgT
nXRCKuTd0O6v4zZoXkiAaRLGS3kQqXt+b8oesB4ZJ7q/iW+DrOrnpb5zPh+kx6IzRa3j3alGf/Qe
NPPlpNa/Mkadp0Atz/sy/r+wN1WLuS4PPJEwXL4OlRopMQriL+nqTgAleo7sKlxBR2msMPrmK5eQ
UTUvuV1m238qeYJymi0uQL7mvCZjVKvaToHBkALz9mVxt6a4YV8Fd2N4T1xhbtG5wAhEmaf3fE+g
YE+grVgt6+e7Nb1d8OfbuamDXGT2Vw2q++yTu5HM/2z/Zs9kfAzx2LTB284yhGAMO1MN1qsMpUrx
/MmykL4WImsrx8EHbDfL2ItUYty89VR31aln6jBR7XIrRoaj0BRzm6+wRJVsn1OJzXINDmkel0z/
yDUuoODT2qBbzmTme9YqhD1eEW0bY/1DhZ8aalqtapU7vZLe5QKqJWUPyqqhOcD8sPITHTsagK+s
ZHStER7w5KcYOqtlaS5ewCuOWMR6LyDP7IQUeq8RXVfmLamkFPOULrcKwl3QqP3EMo3g6VI4ByU8
9NDvuaDFIKrTRCD6S2d0kmtb0rhNSnYmZHvmRYUhszuebba3nBscqqjvxCkBOXfKTQRj9PLQecFR
lZNdRf0IPawhDdXj/HJ2Bu19rro+G6rtF+rEgQkStW63VIHJfRcyR95FEvokpLpdoTFqnW/eGTbY
WBPvn8Gni8poi/p8HSNb0EW5Q14xbhGldIIcvDIbj0XeIPey8De5wHCr+dAtC+ZNMryk3ETUwbG6
tuYrP9SfwXeaavonj+yikkVbBHZoY8S4Dro0TeZeDlIXU/fPwOC5w/TS89Xa1F1ErTaZ26bK7O7X
Gbglw24mMnh0Qov8G6NiNGIYDbD8KG8YrmvniopeBZQ2V3IcxJbDwCw8p1+Nj/Qezjd+Nk8b3xIw
JWeeXhgJ+go3lfw55CSgdJp857xY/cVAC1xORPaLvgZ0y0mpc9cudl+9zy63Gg8qkKmDhHBc22rK
m8V+hJrfUrD++REjHG5bwG8Z8ZWbQbX4yNbWA63oYMzn9fA7o8FlilNgQ4m0Lbx+IihygnDPax9X
oK8MiyPuTqRo6IFnCHu8gmHAkr04/tqugVWNaQWpdTBrlhOP1U99NBmSLnlAF4o4nhixx2YQxNhu
OjzrBOVkAGMS2Dw7qgCmA+0nxI6lSvu5mHxE/I1Enb6SYa970AIq675/h3bmnFDuqmvr95Q42mBh
6TPgssefvGeJ9ZBJ1XrhmG2L/Ad5bcKWuNnN66n66H5sZHBXgme19i2Y4oivWx9dQhXOLQldBokt
ZhPGtUg3eWE5slljtN3VMF/PsfaLKauJFE6OKKcAsF4gmeQchS0PB8znrkmSKcl82VchVigK9D08
/zxyCS3dLk0qZvpW7/EUoROwjO5PN4QcMGOm+WNK8wYhhs+UtX6Rve1fZ5Qe8nPyAN9tytc6CHvZ
TsZT51O8eMBaLFHpNKqNL6puuEaK3rELJXHd1dfEn5vSJSCfOWioGYhAw1TNsgPebnSvCsUi3/Od
k2X08VlrJAVLJVJbLWUxqVuPzzzlqhu/6lkEj0xkyWv1I41MyPC2gKeLgnXTugDXe7PS+lpsgOpF
Faq/QpboSOix26WR3dE8ugSP+IMa7DidQy3kXbPnlMX+xEJabem2T9j2s4GJxg4jNLvsmp6j4GOI
cKjxln3MBgakYhvV78vKXJkliZVuOcxmTPPjicKKmmkYENhYw5EaytsYPqI+6U4/wM16bqihnVDA
If0RJ00Oy0ltbpMqT++OPUcQmHkIgYkuZvoDp1ZYqF+7kFuyfyJSA1h3r28VaU7Lg1nlIDyLCKBp
fjcCoO8655pSpAvK6/y330J5Yat1th+RxtQZj2+hHvviIPtCDj/2awKke91YFMe93fxdl9fqsQdo
o5d/jX3v4FvClxGLAiFxBdvhT1B2WJtvgNmwTICeR3uKw/UxYRjHk8eetAmiLyUENZWj3LWhkABi
+krHt3V/po6ynZZme0zz83YInO0pLF+aDm+Kl6XqE8hPP0hYgfgslrGT63IR/nfBC3aG4g63lxAd
9OP3xqWZibnGKw57mRiG/YC9nVaXs0OBCWOT3ExZUbPHR3J/b0kGJz3r66H1TzJ/yTWuNJE14SWa
BZUYJJsV5nV1bAWoPtBbXnhaNgJPVLUqp8JaMLe/fNmwF1PxDQXPqErsd8GTkgrbktuJdeHn8ojn
A4iz+mmSVhB61Wwbnre/X71YERQToMIcnJAcL5rXOJMFKaoT9pn2hK1wgKiLxT4vScYXZxQJV2aR
A3YTtrKDPNZ3P77OBRsl1lQX9E+DbBYtsathCOWKm8dwwGbUUo+PIn2Dp2UF4/lVsZHRhXyyuZVL
VUYhXc6pQtAka804CxQ9ZjP7OOF68r3nZSezTHDeK7BGaqA8M8rrFW4K6fe729DebYHotMxvPOgQ
NO7E6u96xufVdY7qfofSLG167b0jBV9jbXKNNdUa87B4vBlydWhplxojTVpjHy6GeIgscPHiuozU
WZFpnZXOVb3fIOtbgqRG4eh1IFSpTgkZRhRnhDubqaKFTjm49zpCuuFpnACPg1bg5RlVi4ISpaN4
c6VwWZBJVOgJgxc6so6zGZXtRvYAnMhAIdGQ1ra3pble+GGr6NimCiyueb1h+bSBDLioRIt9p0uv
ZuIh92kgGH3ahtIFDaqibwP60Ir5O6Daw4u7kk0whXIq8mLlLabNjgbS3Yrv4mASxYd3OHIk2C5j
yptIy/rGcNBaFThEMiO1eMfPkIQmFwOmb70z9xfwtU8cyG9BRiNuFykbLnaYY54Bft+5OXCFt+43
p/D4O7mqLy7Yyf+N4mlamO98oFT0N7cwddd32CQwzpqeOLX8pXqmVqLqPIQ7athkarsxiibIyWm8
nUUJJJFoHowu0RwjFKJxwpAtWpeAkxt2J1pjByq0Sv4s3amo9u6QbIqemUkKIW3SXqMYXcCnbgus
wG1Lk3VyxFZnU0oa3SjcODfTBap1qsVOuAQgeJipCjCp6W5rrxyWKx6axo/k1rrv9yAvt1tOocxV
Z7KIWac0pOBiG2ZfYlwPXr56xgTa2CGj72DlYWgKYDyyHvDyXg8lu2FkpapMheTTgQhMTS0XVZp8
GRQvROWudUfEXKXd+w2vONn21RL5w/JiVbTGP+1lMEIKcmeA4SHh/2pCCuei+1oh8zev48SZAi45
NjKRiMfbXp090tfrfr/SXXf0HLhBAVkjMyXDOZEUYeTd1zothNPeWHgMQSm2R6knIU+BfhqwVshe
cuCqSNjOeZbEb1Ztcnf59pZw6vC48ORpeMNxcxDAiapMHlPNAtfV3O83uoA54wCH45VbP+2Q706Q
/oC7dFDOEkiiRzhmkiwj16n9cgkBtwWrwpGTP7RxShcF3B309XQHwqJBjQbB3ZJwQfeu4fRwa17x
NmkBtmU7TQ1pqt6DX/UUIgofrqCZbchv54U6dM6tsIGMU3POj30ClUCWoDe+0gjm18g97kP66wQ8
vbga2yuV/Ysl+BGaLmvABRsQL/jdMSHzJYWAVTUlOqWBeG49lRcnCxRIxlKSJeop+SoZASasMeg5
EE247lYhJlrmB/uYAr6ZTGma4tnZSnzx9w40f62itJviJ4Z7XMGfbJlSRYrqldovdYwKXvNr+E1J
aqQatfnbaisdc5re0CeOpfyM5/E5dWkl7sDOxMp1+Uo3ByJDyWm5k22y2Hb8YCOw3O0R5O7Nn3xq
G2iZIkLZDpaAPT6cqXLWjf/HAKZaMnNXDlb0VdKgRCd+vvUNA/hPs0o7DqhyQzDnvxIMLfLJtJgY
nUFq2t5oww+XyI8TEr668FixwnwlQk/h+bvaQ+VizLtFXCtX7QiAahu3lQl400DTqUEzot0dNAYD
Cu4G5Qt1hwpquqfrqsORdapW4FCiHzULQVBKSwcBkF2F7CXnaQi+qikG05Yfk1bnNw1NzdJb+vUK
SuFDPzU14avHfBW3ZsSsiz0wXr0E2NP0WqTfkuPp3EJxEyt5irTyQyy/3/93kbEtuQAWdIHpk6Cv
8jxAWNSp4lbanRqyH9xuuNkqUubD6aA0cuiKHQgz9uq6jEyhw+XTbuduMgB0u8DyEKv65orKwHxH
izQiksViPaVAHSbotlB4+8bu1KTNW1oNW3rE6MWN3T/TiwTrcKgU9T/YXBhz8zQdDchXc252AfPn
3uksY4x1DBQWhcf8G7/7Us1am98fdQuheEIBEpbEo45IMguJr2VbXO1OHTCmym/hU7uCwJXR6klv
j5JhNeCxXNWWgS+vAThQ9w6QhcFIObDLRkhZwkeCdQDeJlmKAUAu6gQUURcqcjdMy+7oQr61dUwM
28mTGISlNdYu9gKospfpiuAhDaw210zTaHupgAj/DSY9U4EtKktnyMkZSXE5TXMCPL1neyfANe8+
1gC5CJv9jgNbWxfdzI+M4FpzspXNU1n8BzkLkX+6AbRVRKBCwqXa4GqiET/RX07LpRkt+n90kmhW
w/w+ldP0zfnniEc+TpH7e5NGM6swgR3Zp/asNNGguHnWQL4PuyHU1RlweoqipZbO+B9jXGvFE14z
Hjhz6l3zk+4StndH+ZwsAyi2GcmYAmXVHe3uHmKDSJwIPMW7BXmBLwLY28JvV9cum69bzI52V6JM
/D47+R/pa33DY6cQnccQKA0TsLYnCyfxsdxj1zQZqij64EdS8rjVOFDl6lnTEo63H+a2my3YjG8b
yoYt43YtVKtxeOS+QO4TUtaeDt59SsKgJ0M0b/NAcoTSZ6nKt/skLD6xRT8dBYmg7jwzvWftAgz4
GN6MnzMcs093Gpyf6JFNXrQ9bOp1qpagMJAoff8Ny7aN4a+wdkFVmxOBQwgnKnB2Eh/3XOfWBUER
KfhcHiICeeJ7JyV5FaHimx28vH+RWbqdvKnWJOe/9bG5o3mfX+qgnin2dIvcJ5Zwtg3DQjf+uvaa
qmSA7b12amqZsshWnlsgW8ZVqKSqfVAAuuIxr6QuQwTBYaPlAbsNRJns0zeBB97axjskJhasZecV
6lZyaA8GsqJyVKIvtpDUOmfLL/Wi7EnKcfd7b/fGXEllimxq+gHqJOSaJz2h1H2X1UwogDVXkV4N
p2NBRzhrA/XSOYbXips4z2nUpXP6s6umem1hC46vb2EDXG5KvbHjtxTure4Q3mkIjeOzPWea7nOv
YT9Dt2x84/9jL6MyeNEDfyfJNV+KdC03S3rU6ZQ54zRPhgLft45XFxJF2KnXsWxzZ3Ixcfjyy+G2
P2kSRwvKsZwTaEHPXiZktXRFzPRGfk3+nzr+Nt1Xu/WkLPvyWma1bZo99cmWjyMkYc2rCTnCVnr7
BgC7zxV0vpkEfCGDolK9hDxcXb8hLTBeZuxNdxkkdvOQCgtmtovF9NjZeYPzrMQumwV5Vaaou7PF
sEZBoi/WSJlV6HvkycRWGPmXkMSzeZhghPvvCiY5scBCdZYIzS9smfZqQ7KFXBObq2qbhdkYmHa2
A+o/r3hbDb5ILyRs+w3de7Kt+sEoDP5+dNM5G/DYa3Va6wsKXNslzAArLG4nYsxGtPdaSVRQTz/o
RCpHEeO9Il5FMMvx07ZWfNzN+QF3DEjdYmbrvSX8NrWwdmSGy3W23Lt11d0gx0H7TUE0w890iiU4
ljF7SWil6wyheYRaGxCMOswLgkh2eApf05jA+v2jXWKaBYg3ejuJtFGPnKvsZeRTKtOmfw+bdvL4
FVzKkCWcZWrQdfY4Mu14wkI2oKu9JxN2ZqV3ZOLQIc/EIrgdPWgxp9bodFfltJRjSlRWxMIskccD
M18DSUpsB7DRG1rM2V4Uror42Qbx1vyvzrVgzymJ+13KPtPT1jIMhsaoTDOnGja2FAq5v06gEugD
h1y62ahMO0KLB/CWbmd3oI+HC07WYQaVVUPD4sMyvfPLvDayHfGKKKG/EwSYCxMryKkT3CPA+hLY
MDa4JsleLambQo1HPdskPlldLqE3adxO5E2WHwMc6CqLUIT/caXN79ClnKjagoSsNxYEXNHpitNk
QJCLOATg5c0WKeo4B+QRkoDkp/Abmny5RSO+nPnhW9y+KDfQfua91cTSbrGt2he7HC+UVq8nmIog
FWwzQ9sUXpD45wwm+xHpI6jc4yXDHR+TIz6jAIctghgqlCTHJ+RSg/x1dEhEPOl4svFVftPWQU//
MsbP6bupJwTXWMXiHj/KItQmdvZxODDceI1lwjVTB2XZoKKoU1DaGs2VKgOFqCpUXE8ZU9f5hgx+
J0o9bBB84pndcykziQplxptkQ49TXPOlqccObzfbA+Zu0Yc9j2XCyKLbtkdY5UY58Iqg48LL9D9V
aTfxjkcG/GiGi6/u6tht0PUaNrjfbC5Vtc1DDu0COQPuYaHuTwwQgnPmfpD8YLR6YWC0UX5e8q/n
eNPN2zyqjw5fyN5eRsFLWJwEM4Sv0NmO3V61KeSAoabh6Rr9PZlAeUlMEDZlhiFPhDSMWKsrxJsm
INRK+1Dlubv2j4wzWG5kLKNkoyWt/eHVCuZHFWwHY97NVnNrA6MumAMtZ/h9tT6Xj2PpXb69LBA5
59g/QbOX3lHbVqs9Gw+OMWyFD6NWaw5/Eu3hzdL75j1LXUPocOAQKCfhJv+2RwHNgJZICX5kibQb
3Qw4p1xAyWKxvc48yNpKo1VpUKze5ABIeYWT54NSd7QdPILITTw7x3S+qojYIpWCrs2T3OGMwPYa
rva6mwTlTJL7pdu8v42zVazDFXOfNK5Ni27kHbmdgLjxTJBCBWXOZHTu20U46kpIoJKCupCYGZBQ
kJbzrezk1g07xtC6YrLk8WiJlXecIwSCQQEZmKaWK49A6OxzQFyk4NoFCYV/71IBDTm3eIR08rJO
Mz78kG8nVRypZV4GISdAMk5U0ZjrhjS3vzWZbgn7ViYtocLqGAL/IcPjkIam+NyCDfuLpCUBpDTi
k/FZOZAoZ1hn6nDBLHgKxWHKwGrcgl82XDB87//UOnT+8U/xmIdnvsw4cPp/eg5i+GyyrTz9u8no
WC4NcWTzUr+qH7DHgq6nHceoTQPkdfcUg0RxG90xVIi31KYEHzXDJnqIKTONGhY07qJRRoX7Hh8v
36PkXdfDDXDpQkoObqVzhmxh8+dAU5YfH+ruE/2wXE9Tzeah8/rlAfc+QAaG6LaihUB9n2RDkyWr
311oSEjqwUmxRu6m07M2Glome0q0ky3qsLx9zf+BK/7erXxO8nlB9HUBNeS8XjkGU5WGfbfO70Tv
UE1cgyy4d1BeD5NVeH8DXPYZMdo6tjSWaHn92/UbyuMnE2DzFXx+Y0h0LBH+OQ/uNDyL8PIX3sNs
BnpdgAbXX/aSswkLLLQUeJ+1QxdDEbFAt8jmhwtACSl6UOUIUlOIsrVlhlAfkt6gjeZB9jbI+d2R
4SBTvutAvjgE6DwQ2vhvhP2hKuP0Ji1efkVSFT2pZ5inPQaLaQOIi2GaBndsGPkAcTCkouo6e22s
BGH3YjcjjNcPqI1tV+BaDuk/acTKRchGLMSaOCEqfdgThJHYCxEC7PY2OwIQWfApyZgK0+QeUB0o
D6FFolFiAfWosatcVVK0Qe212rLFB4QpfbmJM4+MvSp7NAk20XvgBNbc/d4gdHjmUUEyGAxTUToJ
0kmGvpKlVIv+emm8BekJxl6/x9ApBawG3GYHqO3XPh90t5RkEAO7u22u9OxnCyOVC6zL4TfMWnSu
hocves6cI7vMTGjj4osE/X3+PqN6z1KC9tfcnW3xCZ4l44eidPYoW/IRkQCkYFlnqhp6eCIf/4Or
I0IPfwDAthrMpP9qhlpFKRJwa5TaJ6fjHhuXONEJ1VK31kp7MYSSmFuWcT2XQd0DnNYJDmuKyOw7
eNAuwVY9vuk7PdZth0ifHBeTXxNT8KHKKPu1n4ZLtJ1v0WqUiXrHyh41roKabszIgQT0P4QOyEMy
z+IlO7Z+e8YOkG3CRtAib4SuNtcBrz4e+u6ykNbNgY7OZE3LfwkXq4Et3qzGhfoXzotCpvHmoTxo
IbU4fpxL5hs/a1FUZ2BiPBpkrRIVFf8NMHrUFu6w2h9idElvcEgj+RroS2GLzKMexW1MLg+GE/Dr
DVdXXRWFjbLib7jnsuCXw9nnqywZIxbsgNLqV8KGUZ5PLOfS+NhjXTJOw8h26VVQvLfDHpqT+mqU
jyLAt0qpW77sjCh/L/JQ8UkGnGgmShoj5StqG6Xz9LmOLIe7UQ6L7cVrQgNhm4XdEqAtIMKUZFyw
V66t0OpBP5JHwM5+6td18To7hIvzFpmGT2pVKkXQ+OK1nrN4eMxXYTTFoGCWZi+pk9dTZPogrvE1
/pXH9AGqh/byQ5HYhMREufXxEsyU4OLRFHhlx+XjwtCUkzTcRpt1SMR1OsgkUmgyTB849XK/VF/t
xafoJhpjZs1TMKrpNG/Cr8J++1P6jeZzbnKh3eU4DMr04adnLuCWUdhVtvrQ14IUfKV1Y40UQsaA
Bu5U8ReUZMchIZ+lPoZrCgxVtc2iDwwWzH6L97xed1UL8YeiX0ZVox0mZ+mSH/VdNTeGov2sW0RY
1I2dqBcrsnH9Hi8Qyy/J5RRC2qgYYA6jpYviK0Fhqtt5+okkh/inpurmdKJUssHjAIeUK26Qp6On
oYpzzGJyl0x4EgwFZRVnX8jblZY3tvBaqHcdMtlnMyBCGOzwQYZrcayu9JlUozmxqT24LE4Mu5wM
dbpCFAUsqCI63YlyUBUX4Asm8UYjuIwq/rlHiNm+H0Fx2bhjmBVrClciu0/E4yaqH3+yMv0Zbszf
uTvNCdTUaanZOTJ7iNiyWNblqbQmxggUPUgXujqtoHq/ODWjwpoeAi3yLYO4bXoVXVJLKJMqRskC
6n8b1XKncYSgD9m1zqoy00veUZrKWo7CQZY6McU7C+v3cXWIQV0o03BkFuqUJZRVd9AwFJaute0S
eOsnel6vblbvUqqCS3LCjFgNgzfPmtGR6RPSIUm6/OFpLLTKRDAmdXQPCyELuvC9W73t74KoXfjF
cALZbZIa9qlC/k9fcQ9r8HWr37qKE3iqJh2/nMG4zNEvjkV169H/NyZ6nKsPVrurWPgUPlFoU07x
N5FCKpICWr0trlNiRbtrt1JpXXEg4PJlWMw922HtPnJzAoYdionskY1bQGyDMbOPVNSRJaRX3Upi
pWpGPbIs0hzqnF7JtWX9OP9x6LR5Y9EmuVe9gGSghBhTBepmZ64DYZBe8dOXazALRcMwUK4KbQuZ
uxi5fA81lDiFJ0DvrH85Wqc1XJ/jxcmjF7RfPKSAA3pg3azZ4nJV7NUrDRr5yU4En9bzHhvUk/21
r81x8km4xBJ3MFWwmk93ucevukxCVOyYE9zSC/h9KdHyFu9oH3A5WwYaVLmavxObjOh6ZLTBDItZ
V/oCD99pkAErJO4qJBGhYayOy1i6iozky1XBndVKoc83OFXSvVT23edqsoKO/KbbAHXzccktgKj8
OHxVphUaKTJPm3YADFh+uSwzbRq1UvsXbgqVVjtNpa6WcZkUEK73R6iDftZlAaJSDzNYHmj0uHSV
DZfD6VIHVqq5PGvImRysm+v4+cf+ABAQXkzg89lv4bIKYKLZmAp8xNclts1PcnTFNj/8wsXZLda2
lVgh3evtV1vAJf3Uunkn51ULc4w8bVVmTolfEUvIpaPLOl3fkor4XqwCr7x5N5metTcWJW6GAsnj
MB6uNRN6X9pq1QZXh0YieKVKhMriW+Ds/kadohyNBHf0jUgTEH7XPkByuzxgr50Q9c+eDdQS3YVg
r1/PIHd+DHYZZnIeR9HUaaPU0mU4XK29dBnqJLrpQEx2FBULLoo2BurBGczxE2ncp4fakTfPvfHu
9gW1CWI1Cytmcjts4Ko0kMvgP9KRciom9ei7TE+YiRlCA6zBdOQNdt2fJKIlxPBRVl5fOagWenCS
A4lZsHjqrb4j9tQlQ0J3vaUoSqUXrtOugVD1Q+Y1WNCzJCdG300uuVAOE/koJpPpFOKCk4OQcT9A
HRtX5zOXq5vmFd+Kgm7dZdQqSoar17uBrTA2PBo/DpZriLJr32vnWAqT2LJ2ghjyOwx+4b9EKfTJ
X2J1MIXPpxfm8P+ReXnuzlFEsUO0rW7YMMAkU4A6s5pv4SJUf6xHNfYz1p4RA0hDdMmngbdRkTnm
XmPJHe+gkb1Vb+28fO4V8AWmorHcauQKRbPJoJrXhPJKKUbR7mrwr5PVBq8AzaoZqv5MJYWdz75x
umxBDiQ4bnqOdirIdNmqIkjfL9ZE0BOOUWIVh69hFpaaWEcC0yM+lJ/IoqtFG9qUyUxUfHn4PZvM
aGCU8mcN88yGOKG3+Wt0Kvnf7Ox4jVDjQHDgkkqBBeBD99X5Wq9MwaiQWjdPvpuyTwWvuQHSli9a
rd76tpi9RI57MbUWpVa1ioZ+KJbtpO2oOWnBYn5n7zQYbfq+D005ScsUXuYdURTj4GOoTpZoTkL3
SMgM/hoPK6etZwx+DLQMNSqBo9LjOC+HtkC6GsUXZHIrq7yEmjnQ92VDYt/MdkEt1/QDbcsDGSW3
smGELNmwAP98q5JT1KNmUPFHGuUpl41uEwUVB2Na62Se/bM8KRdEPLrIyMBw3Lh20XkOzCZ3Y338
7w2S3aqucSN5CbVW57MVBSjAW33qAhY1Nnuj7GOsPXh0eej9fr2skxVlDH1+So7Iwqo/9pO9Gopo
wV18j4qCq6flr0o0lrnIW64GpLldVqT/4p7Ak8U6KEtc+7W1V5zM05Ror/MJ9xbnDti8Vq80JFe4
fKLIF+LuZarUfbr7oUWuTW2/vdJg4st28hX4yoUKBdk1+sA5BQf+i2jTFHaIAbyHmBDudc+odYkx
HNnPrtow3Ktu3NEjvb/TBMMmLX5Vic68m+F+B5I8JQwUelpT6potrd+GarHxKuuGm6DMRHICIsXF
ofGpSRaEXftK6MaBHu/0tq3pDVpsW7joiqx+y616aeUcOwij9fbKYK7gV+AunkeI6lHNZntqJS++
14b5LfVlJFfj/P/9cKVu9dgBmROLrTSs3cXM2psLLcQPb/7rRFeLwrp+JOvSkkSvK2F00RDpsxYf
uy4fgQ9SnUBvk+XtxgomGVLK268Td++C67Kh1yqjcQIC7rH4KYbL7PmOrHWDtRvnHC5aOyMWR0hm
d2AGIYtV0SE4U6E1TMIxjSIBKNuicQOHgDWoabZO9tGdV/hmjjAzDinuOMAyd1edf4i34OOvIazX
I6dh0/CHkKgpe49S6TeNOW4aJtUbDkpdzobCIDGDx0GjHOM48FPmmTTBSFyznuteYkjA/Lkqm/Fq
dxQvYZTknQLeeLUvPltsBmyre5jVvJ/mths6d/T4HglydeTTuL0k4eXOLqasWeUdNy6MCIaJwqey
c54qeCeP1tSFSSmqw6UtGo3Ht0PJgV3pl8rrKoM9NbcFEeXFVH2coJZN7jB7Bh89InDdZRWIz4vD
wz1Ra+ppAxEEZ6qR31lKjvT4QLGenogSeN0aRaPGM7Ao/DwUCqyV4MEtFYmut5ZURBehDEkJ+lDw
BC1gIswTatKpaJMKj+gOh9n4GrkBOnWY1TPpnFNKn6Po+lDxl7NcT6DtMmSuZNQNa0I7Sdalzd4t
klG3KQvhB8Zd3RNuH9zHbc1s8+DJD0m5wKfYzTliNBFAJLILm+0LvJI5XRfZ8++tR4OxcqlXBtpv
8ZBVgVW2h/pSOZJMNL/+yeDsl/74JxpjvRn5riR0cDCOWQgJSwxpKDXMGw9ZDkh2pk7VS8hAeT4M
mdeWfDdMDyghl399pWbwf7HbzTtybnfjY2q45GmibUB0J4kJv4htMSXpLKHZp/j79MD6RR27n13M
mdrOCX54mGsXMn9LjRsXNcK/3yrXQS6AikZPVDMavWmUC5KrimKm381DFojqPC1lerqXHxjDiEej
4/+Zfum6kdkUU7mn8djXybScBEaanwnRSaHAYmjcpv9Ns2VvzA18DOYpjGDQLbtoSJpjxtHGrrMg
/OYWAfTHtrccALhmkXxh9F3KYipFAvebpsblKIQByUE+95tvhuRXyiFtcgyyQiQAm8Q5EEeGUyXP
9KIFRHfni04EBQdhJhhL5PUm0zd2VdqQyMHGdHYrUHqKW5yexjxIbRLxd1xHeVlgmkgtfOHu4mrQ
agF5k4lRaB29Lgs+/xFDPIHxGx4wxz6qUM2chKuzco/Za8bYf7X6uTUBqdeEnmTRFsJXDt8c+Ek5
WcUQZtvbX0EX702Fl4tpgn3fHmdI21SXhKnrLDuUFJqirJ/QoggI4v7NwhaXVYswDfhsq44ao9Cz
QAltm0kybH6E/lapoOHcnVMCUlGGl4a+Y8TQ5CzBYPeWkfrSBL1cMD+LJS+3kWCz54QufndpIVeL
WoSFcrvDKNQonQLGG4RGwl5I+tuB3uvTFu2EBLJThVp5NVqhidUsWZkPclWoFXgfk46syPjstQfl
qOCBq+P/nvuWOZlG4E5COmiGKRxEmjOxRcr4wREu6mnnoK5zPtcJcARCg/H6LXCDhzEh8P7f4889
JW1CHboB0gvgLxUmF9akbjUboLEm1fbUUd61eCun5g+2DDwCLN0LvrXTaMuj55shOMRbpaZesQxY
VFkAdZRHRsVwdtiNxJbUTjh7nSLgRu7I/QRmGzmsgUoADhApiCjLVp1zfvkdw6rb7RISO8g83Ajj
b+rG/N1drAIa0pbP409xqZ0wkdWTaalHo1XfVysX7wFeBHKRgmkbURRJ/2AqT+iDUEcHN+6X3z33
eilIdgDghnF1vaQgRGsd4P8oGT99BW2IWZMbfVq5r/G8m+btPJNvo7I75rZ0vCjoCFhD3T8gNDlz
zAvfqsL4T6rSobKF/r1/4FXO+3MIPYFFwrwBHrJyG/+imooVJHjJ2f5SrjZqc/d0fpO55Ps2nqzs
mW3xjzfqNr+YI2QG+/Z/bhYBRn96EOZ0LAZpykKFa2rw/No2J0gLJXDz1F/YSFMfAGCUh8Q6fr42
ybRHkRjkBiHJP1bZuSdWKQGl9EfXWaC1LsBJekN9uiUSUT5dLg6Q+ho4hUb/5P62OmEBfL5mwHi2
TLPA8eFzb1waxr0m/O9YPjwUes9VuY9uWydAS5JPirUlywLvkFOIS2ZSsfxap/xJC9Seizc4iN4X
ErqhKzdCKGUskzJJ4j0qfvr8d8J+MZoBRi4wGQAUCm06hoYOFu5dCFC1tX1LcNbJQTrp5qt1juD4
rjqi6kBam8dlbySMcZnTLZnuyyNLseNimlLtQoFRqlATJUmXwUXzOmYLp1UzYTl/KCfCHELlH5z4
R9mitwgV2es5PaziaKa7jPceKza5vhtZ6htYvnSClUd/YBoHOGnMtUviauqU6FXrvlOe6Bg4h07y
CEpF0t9JDL3pteHWfoGQwNJ0NRDfSe9XvThExA4ob21lX1IdgaEoX0LWQsFUjEzECPJs7tl/i4vw
xOIFZ9CiAnzh7E/71z3mud//wBXJmZQ6ouOC/jmfCGjTtmD12sCMytTG6G/EnqswVofQPyUDoeor
TJjVyg2y/BYf7x0PRZiwrcK3+S06wH+qVOHdgGYvHA43+K6AF64ZBb0fU3iZSt3xMnxrpVaTiWtz
oGcGku51EksAz4vyS4PL6MsG0oR8k2aKl+5EiqGMIP3K3zYiJs44YCP9U3YmmT8REw2P4tWoRZzc
MIUWADlNCrc8JuVg7efGqjS7IwlTDMwwIpaLtgPdsfK8HWYQwwcv6viA66xfJR4HwZB6lsJuBDzd
TaaN/ZRQfs7Io01CTzAqruMlhRO9CZv9HpkLsS4y3tmIZErLgg6mIhlRe+H5xUebxedyv5eaiouX
eo/4SbsQQ50VEPfM0h1tu7h8j3ay2udbBu/hfaDPjX6B8kjDW76lwuH5hhPy4MpZVMU+qofGRORq
FCeo/VJiUrTeD59MBxQuCPZrW2v0FJicGU8tDr8zbCCu+jQm14/YMy0+koU2EvHlB5aE/iQhhggb
28LEvCWA4MiTtswhz0e5puP29SVkNEChuVUtvFXV2FnE68YYtR8zecarYpoebMyxDTakAcwPn//D
ZvGFW26IUah4SAcDLhYGdK325djb3DASJZKwv8dOTioIK39OzgLRLBsTlsWXi0/YoimmWqaxNtAB
kLz8JI1x7QHNPij1hLw9xqHq1pS+RDMgo9hTVDM5Ousla+/ENYmKRMOejTKdYU1msy27iSp+Uhc4
DGU5mYR/QZii+lAfR0ONYMGNJe0yHgpLuTA2A5JPgHbL0P2AEhuTJyRIzro1Iqf+sZhmmmm4O/l2
QnrnYp2CcqGBosOyHo4RE+qgOvx0DJWJfiGP4VMZv6C72VxPGZWLBSTnm6yrB6vTU1fHUy6tDmq8
9AtCNZzni6IECunDiT3Yb026hkYkBhSbksf6B8aY1EVeGjPKB4xUIU6sdxaaIy4YtJfg3I1z5zxR
eBClyZ82OdKSF2Zz5PDV3lGkNnbykfV1/lAJGrkpynPrYhPofK+4I9jDrzNUAN5ATXi13jTos19E
qJYDp+gza2iMV+9MtSs3h0XcRHo5nK/lkdj+E4G8rKe8ibypQYog34khNH/zFgqeiR394vKXEzGp
D2jk7Dw/R4YREcjsD4v6EzoM7b270XHx5PRYFt6n+e6vlaXvNiWkOxckYfDrm3QdL1FPG24PYZe5
YbbguMXtoxvcdPF3l7SZRvQmZ5aQG3utQOvXXaC/OTfnfqtl81fwcxJdBDyf0qnE+B+WyNfhpTnF
zBSTxfgtcAXzw4J7jyvTZwfKNBhaTbc9+aiVReyKW/ja+qdoIiZSQlnLDcU6peDo3M+yK8egEoXd
7hprLELFuhq0Jdp2a6l/0MmQVK5eBSdpovf9wMDqonTgyaPrgIZOaz5kSysk3bWTn/XVvy902ck2
roihfhC9/w8epdJVRuWUUyYGa1AChazhYXvk60jYLzvVEBpAT1Y6gzu65O9P8Sq/Jwn6n7MJDIQc
EZfcx13KzU0Wnfnmq6sSPCaeJnibHNUDrUL2oMZ+VqQvin6aRBEIRWXV+acSoFMt6IEtE5nxqxvX
kM3cK/UywUNwVmtWB+JskYwue+ztohbfWp+PUs2PNWzd49uu95Qsw8H6asuKMnylK0Ef2GOzPLKm
b0kUXqDfqukB2m0dp4P5wJIMDAmws96gGAtynmlcOCvAaP4RN4kkVHUczNyGfmhAoaWHnhTDzznn
dmMJLjlv+GopLZwIJwfvBxlMI3eqWH2xz9X3fjFEqayLQE5SXC9cNWPhO4hmmJbvKP1JPprPJI15
nFY9P9UHZThCCIw489ZbfICUnvPhE4PQlAEWrwKfL+KO+bmBmkK7CwgU44y4cJB1RuMBgdSmQ1R1
2wKyUIxoh87GVdyebTRBbQKvSbvqiUE4+IsIUtq+K2+M/kpEx4ap8I9jJByKzXM9MWIYNrjF7vb/
+PwxbV+aH0joA0DGmkJHk/1nD5CDlqy7d3FX2sS8erTfIDaNdRsI/TDWOL/UKAGoOEUNDZTdhYPq
D3XuvbmlRjfQGthtUEDDTcXSMW4LajR4BCsVpkpD0nUezrLvHXNdns3gB4SAIYiQf8ukMiQb4tpG
h09hIF488NWANOLIr83xwfw3ljn2NqLrXlPcEp74U8t6SoGdIL5XSelgzNvolaUzBxv50SiLuqFj
eKtEgMnuY7L1bN5J+REGQBmysH+2DA1jY42/Pf2d2EH7x6yoQkKlMNdmPtlulKicVDUoA2bIUO2y
QRh+PzfFeYXK0VSpSG/q494CATu4yHTQY7V91XR6gJiwUR74vUAuIAX3hK7MjYj06BETpGs2pCj5
9fLIF6YeSwBWjM0d0eO84CbITTLlspPk7g+86HGI71iAEOb7awjck4WNVMWWfav1AY65fACZmO3F
a5Qo/OsfHEiD2ESVC1bz5a2wT5ympnJaN8iFGOTE1sRXg3wIS39EW9A6KlIjCh65oeOl/jnQzQsj
Z3jJ335XSVJmF+x/K1FpCLjE3SrCAoPJSSUlqug0OgP0wuCjWAV8w3CPV9z7Dh5NN4NJWKOQNK0v
jkqT4wzNF2EM3hr+9Ordwfgz7+dEPw9Ormw494/ak2DjCOK4+kAFFGF3IYIXNqZXtGkQnVLmDmLl
vkqeLYCaEnczB56ZH7bmWfTbnz7dwFwNj8vIL3HHjq/XGftmkW+PyGhUHDTMfE5qP3wvfCiI18ND
n9+COqtvzLGZIxuUaYMROS9dwiJ02B1ibvzagYmSGCZYqSkwJ4YIUQxqwSgSYgh0c5UzjCeADhBF
ZT8we2tZE8rZ2o+UEZRa+1TKm9PRKoN3asBhkbEGJv73xfkx7S8MwBIt65ZsTXen4/KIhxzD259y
YhVPCeSZSB6uVYmTWBzL42NFUyGEC59XDVMdKdXbIo1fgfZrpViRdlKwl/2Noox7FReX11TvMwFy
qkG3kZ7yiVBcFZjJK6N+yb4/2QpJsOHLh742tNv7aZlsY5mKfoLhNzENBIULkwgfWDz1DGGocbPg
ihAEOn2gWpooAKfnlb86HdddiRHWlMUIw3ba8mUWrOO+6AB2ILs/pUlgllRyPIiJxc7vWa/z344M
zj+JYPNCwecCEBKgeNPXjt9B7MVNo1GosA6krm6T2ON0ratuZPVKqyQ+c63ivrZQ4eqd80JxY8AL
LfF1yqgxMzsDg0EDb7uT2XOj1pGEuYdt7JeFe5gnq9zePhNtXerO0J6/n9H7pLJjWHnQ62y0ES8z
YJVf3XoZZWHPLLJyyL5c1StODzDOXWE2aNHKt1z2qO8wRdN46eReihbKn4XFbLiZhBDdSqHoRNIa
0S9QI7ADKRUI9vkAt7mivTTrNmirXfpvk3eE2GdxlHxhJM05ozK6Amr+u7r3Dz5gO+Jw+QyXMpPh
PPDsM5pWxZ0baC9MCgxdgfBacMwMZa/lxov/nVDwVXlgVmPvCU7LdeBono7x2m+nWd55avuW3DUA
HKNwZmukAHP3yCOMOMoaxzxySwXG4YZJBgQENEDvEndrh32OvtHPdfEkiPjjUDzCjPGlgYUhOT52
XmBDi2+ev/p0V01dPmHns0awsWRJFypPj1fRHPaJ/t+nppvIhD74uWlsJ/BIYAQx87Oa2YC+UyqF
Fe0Pt/Tp8SAoRG1kXxVBPodQgti8d6eo+JJOlkn3R9TkH4igOnHdWEO21evltJbMAuT9mEMTga7C
bz0XiHLQO7+CUCypExwH+umzEpa6pfEaZA02wCZ5lIvgK80KOqVyG2/uN0UWcsi9b5QGKqLqBepU
wzCQ+ZEE5Vq/pAgE6MeC0ctgkZwPZgdzcIRdMNwzjRCFFCZTD81ehCp9F01T/DaFJRg9v9uBPwvK
IKtThLmOYMZPX8XREaBF4fwaTGdUQlG7YsoDR91epg1IrBWg/e16g4Gggy2nITCdnhswOQrUIJQp
BSLjWHJWzDxXQnx0ifFk+b3vyI9ZOu8W0p0AWCTORgwtEdf9qH1bsYH7cVT1GrH7XJycjSiZqIZS
FREns+zfug9kkKYQhXmEFWqhgJFKvg7lTCSPHuibcAkM5Z9DKT6yT9VKPGdMlxEeWF5cOzc++UTS
zjfITtsBrRxsHw9aT7KFW1/2n4I9l1h0p/YwzAey+rrV+r5YpfC8Dz51hBpWi+rl7T8aAh1TEJWj
KgMMZDewnrlQfPq978qKGMDycH9VgZTaHveIABMuy6jh1Wg0T1NOHRVmaHWa7HZEne17Pw8my+UD
hpZ5Ezx3AbhzxSlL1FqNjNiSM9KG4qqIW0/Sz/3Tjdkm3CIICoitPZO7i28Vj8IsDmt58SOIjpLC
MRlKAYNJwQ0FUzHhLcHcOobxkSsLxjjjejT+RRlT5LgNlyaZTTTbx0k6/q+0Gi9vRbEP4O5ItTKQ
FY23yX5FhT4Nh5FVLu9qb5NoHYAZeZ6xYWEgV+q/qk2gLd0peM0OsG3py8ioy7NIilxZ/J2UWYB9
jIgZhdmMzFPmtDbQ6OcpsKjBf61PQtAoiOIv0OWibbrRr5YFX/KBdI+V3gDQ//NEr1dNB1O93EBv
1eDXuO15vso55l++4KbBgQzWvwJtANxhr7ysrYyMcp9dgpTh5L/Hdi8vZlHRpNtoreXP3DEgEk21
8qmtpMFj2zs8X0qWlh5vqM3hTCByKC4NU6KTV3oHyLIykaOMEAMpRn0g6vaVFFp2kOjiz39lcSvx
T4NbDZJIbd01GEAPNjEvnR2Zzhk/GJyHF6C4SJLICzx9ipIFYe3GuTRRN1Mpiy+V3qodTclSThp5
Oge+AT89Ox855CSzo2abQDfcgVo3nuMrpz7nl434FcKMg/4p8zllmulJnlhX+Dlv5/gHtWng9GxB
9KdLJgwF+q1h5PjoOycknEWjA5ieUuWsTKp10sm66lI0IsTnIaPVmgaZURMtDiz/+gHIeebhBhjG
2hTgjBC0KPLHsXeuWm8sQmlGgwTVjgLkDwbm4dt8FeW0W7DP7KiNodoFP4ETbl0pEpukdlEVsBR4
IE/uVgPj5HPZBWQcaniOarv0rhL9hRLgjLcJXkNaTm3oal3ZQ9Z2RM0fUQseDsdnj9xrGlFimZ5z
5J1Kf9vjpzx9P8+nCLhCoodpqI8AcuIuNvFQwuW1PWlbo9XVVs1hd/V9ktdj6Ip8y7IRzWuQIqE1
1iJYoJbriM5u2tHX4nj+EaNrEqmbAF3cVRrF0FJMRjUKgO899FFNNoyMytTqk2LgnUZya9Gv2N6m
icP0kbl13pmtw4EYvdPFRKflT2atY8JujOEhipFHO36W36c3YI+z2jTJTF/xQx1wfBa5L2lQ5d/F
FntJgE88qG26QgO+i/AFsaOjItlQhC4UyupFJuAvrQuuc2nzBYrfjVfp1/YQZ43GFBRMTtXX9UHp
4IGBFbWuhcxXIdYW36UCFSZ+S59wbK+F/D2+46nUKfbpikga59NDpbfkuPAq1FL/psO04Edly6n8
f3lcmiBTMZmEs0YFlkZMe+bAkH45TNONgQ5qJok72s7rFYBMvXnLq/E/BeT42+SdeYpG3KO1H/zi
z6UxOtoTA1bysmT57y1hL86XkUmMq+8FWzh6nACFCAjkT/CHgfQ+yy0BlFsIh8j0vtdXJCYeiJeb
QQc2T+4+IXkPjDnhqbDWjEgPKYSGj4vWMLiIEhgEzUwgGUvr3U3xZdkz76mO66mA5VEyJrYvSkjJ
K5/JXutAwXc42UQFtBjG3gH5zOpDukI9CpB7RH0050fetnu/72FgEPy5lQHMn+YW7/2JxBQWqP8Z
ExZrGkITQZEsFKLycoWm08bd6ekrnAKQdI3GmXOkU86paIdI+JW1JrviI9IYLjLk6iLBmxMKy20s
6rdIFPq5QAK1evLb2D4vRnOX6ENKOOsKdsE8z5WfV1Y9G8AD8pVBhHYLNdSaxDJWoU/IQiMlCrle
j+LcZnHfXs90oaVTWXU5egqBi0dng4KN2aZ+MWAowan0ErW+vyrXhYeW3+a6uSASLXqhYOaC2fVJ
mArvtwpuY+szsbvl9aP02iGdb7fzo+pyEkWeZgVxkjAj5m2P+WKMakwt5FfZuoc3AFJWjWTn49rx
6QKdMeunH/GEnWVhscpKsm/TXxR0VqbX8SCGvhVkCEvHFHfCW3N/XsXR//QYTx1kHjJkOx0gK+hr
IrB7zAVnKTT1DKaEVFA8jiLLCEe2mfLePC6A32z0cb32SGPwfnWqNo1K8jx1LPOkvRKy2cJ5mmnG
G4CiBYUZWAoLO3x0dufefIQMzALe8BCQivWMQ0mbl85fYrWFSmc/cIwgG06JcTasBdYpvNFI4kVH
m0v+6t3bAY2FsMHkjOndVLDJzhH1GqiCWRC6qqW1v2u0/TCF3BQ6v813xh74wqB7USy1yjCVjYrP
x2V9fFQsImlOSSpaxyR43jypyFLLpZIqJWILtbCqYz0/EhqID4Wp486LCooeAX46NlPoPz6iOrcY
4YWi7iRq/A918TK+5iQ/GZJ+rvRP3mdbtX2IbMd1ZH9qQ3H1a4MocjNjsmxZVgFAAQ7dRREd+vYv
Gx+kz3E6q14j9scQUe5kIQyg0T756Rzqekyeo8zGeWxPog54DuG34TPcqfjVJp3+YOIGeYaqVSwH
Wka+nxb0PWWFdGe0bbBu7wm3ASmYoB8KMKABJSTgf8YqoB9iOVdUGMcZthCKKI9JjctlXvxKC57p
HQaTKnCL6MqWejtQoL8skojx2EktYTFTwb78ycidxelyAcEfPfyxOEIDdGorSHqcrv9puAh088CY
DQmCzZukX3K9YdYeWDTLtd8WI9BbRnbsstO47LWMwlm8u/7Du2FXJSs+mW4HnyZrAjwSlFIKSyKX
hnPZqTTGWOpBr3/hAii+C7O38n9pRkoKYJXBDwX7nw81/+JABAgCgPObHHr2BEPse310GHjcz606
XfivSxleb3A+/AvJKDbhAlet0eW1tfBufcXTNDhAZUATHdQaYAcQEQXBEBRPEivSbPF/hcsiWHM3
kqskNHeQlw3TYavROEGqka1To8vFm9MR2CYmfbAmCZxyi4CQhXyLXh/S2W80/dH3NTzTEpd1hva9
Dfo+rcRR4kGfgszQ3Cyag0X2GMVJrV63JTPGaH4y+W6NsRI8KYsU0prEiOzoeectk3aNsVBgZ2W/
/TwT3E7Q5F7tk4rutGtrjoLIbvCmhsZFSbKoL29Ucwn+Ab8BTkQBVi1rx1MVnd+AY6QWIB1d6tjT
WDILqcWZkCjvhzpide9avPuPD+uNqj8GqKWSDk+rr9d2PeLt2giCZ2KCg2EwwXj0s9jt9C04xYui
vtNHr2Q6zvcZm4c/HUR9wazSvlpOBDW5Qa0Pux3ZFnhO/K6M+1jQbRbGereJLHHohPX2FdO+sAym
MEnEkPkuTkbjH3B+g6Ye7jdL+oTHfEJW8//VNw9l2x5sC88ZVM73bWz3aw573f77E6WJP56ogY0N
y5BHyG7da9XJ+ZgH60QHdo0/afEL8bk6yeCfIqwUGxFUsnWrGL1vqNiSlvOAGTGESyc0ESo7nHKC
iOlcWw5XN7nq49Mq9nELYXa4ly+QkDy5eBWLn2zDH1QweGEBBhviNuha37R15vxJ2VjoWPLbPqbB
OJd4EDsJZn/mQNBj+pdzdEdb09iylFu6ZLO5N8zo7IucywV+lwOC9KDnl9HfW5KZZqx13YKUQ96d
osp328LLO0Jnwyxspnoxale7ygVL8w0aOFFZBIUD9AdgLNtFMPMswFzWfGhmyFMp3wpnhQYRh594
PylyiOOGEOehokku8pBitN4cvuswIbdGvgvuum/sHIR4hNttik+1lHLsa+EB2egULCha76vMofdV
7prCTWsiQHjvnSsZI2q0tATfppLVRXzD4k0IJoKNhUo4iQSdAIy70DfW7x5gv0FBm3qVPxurM9lj
4CUIRj/JEYR2J+O8NnWilbzS7u5XfV9MIhga2KIsHJ72PBJjW+44tAeJt7ku0cEO9Aw23dtt1gSr
Lb+O/NHOjKXZuUL9Hiz8hs0qkZHbqahmrXSESHl4NvadlfI4Jejklv2gJdh8fXbDgXnMVTYI7NXk
/wMOkkvwmUCw+1fiuQt2kh5r7HTL1qSz6IWDcwQ6UiQH11h0XE/ESyh2QIvrmOMVFGZ+mPo2tcQl
+SZNqCoiZiso0wwXB2HlgBkphFLU2HNidDtNgjWw8UoIK7NjoDnku2qxebD5OhawLgnhE2H40ECB
aKaEw99QkM5Ayadgc8M/up1gtRMid/6N41amMUzsBdu25364vAX/tBMUKOCLapfyahIBlOrgl7nB
MTQ7GFrJ3Bb+MMThmfFIkWu5U3omIq6rwXqLblCz5E7vB+5lRZpaoxaiMX8/OaIpQr7zKrMXbYgd
PMW070oRIRKCb2lP4TLAG0cDucGkySrx0InlhC6uPLFhNHJQrpypyM3pgunJ4KokuOpLksdSyKu5
aSKIfhoYLtcfXiqELcjrLkE66K0taTyvTate48AXL8LEgqGyd+X0UECCRTLjo0hXmXMdULFaIhud
AK3/VwkORXpC/5p3iQNm/g3UHs06ZN0wQGP+7PCfrFRtBTr+X3ty2OqC3AqqAWNsMykF1gn2b0lI
Iq6ZG/cSVq7inqNYTFhxarPo2Tr5nnpnc89ZMDUcFdZZoSL+v64k+9amlRFiS/+CTaUyhDqfReIH
HYK1J8kc07AhrxfQRLMVXyxolzMKE6EJOfDuG59tkqZ9G4KEslB72jGpHff4fDehxtvL6NY9ZPHT
xg0Ct6CONaeCx2yYcT3iAW+9q/L0LCXdRvCihUsVXz73x/ZnWn5vowHu5yYLwT0BuSFbJBZzQ+tW
FgIhMtspLmQi4rTPCk8cAtZ3j8WMxrP2OOny2Nl58GOCFHjCKz7LwJyIjBmUx6Rr9/OIWzPr84rn
mk5IalnCvtw8q4YmsCT4CUUksdpmCsJ7bLkHXmc/ldSkpyXq+viqLlWdJi5MHGsa46xpWn5X6Dd4
q8oTX+tVpCDVhuBMpJkuE8/2ozS2kGVwRUdvcZUoKmfWXdUvxr86Lr5QBDDPBRofkdQN9fgzxUvQ
93s9FHIdWojug+6baJ8UtWSe79YEMkfJr3T2FWJDT8QBTDk8p28NamtaTLyrlRVHSJEJ71m8jln7
oUcBi3lPYlayMMHWPfM05NLFzzMauYt/NzEp5Fb5uovdW7lL/ofcia6uE8K0fr4YDycJ6M5moSxC
lEY8OvuqDhNkfzHYvIxP/8yTZDsPMMxycFE2OmVGOz3QCWSLEnO8UyULSxc+/jfMxowTvLh8BMr+
eSnjh60GTQaEIP2mzzabrA1SNxxQI3ZkrCE4L2XMF7v0RSVEg/q2IJpH2nAuKslVebaFrgH8FDBb
iUCCgNnLpgTAJLuiWaWa/fwP0DINNhSfskBliSrL4GCyQ1Z4o7loeqitbMSSFHUy5pM0G8J4n8Ws
41mRtAwFtJ8A9rNIbS0KYFc7acltln32SD7kMV6k6vU4nWA1UTADDSzSkGVHRTlLkGM4Ru0CBVT7
qjblnjGNXki1yuXj6Xutp/gE3JAYQ7SiTl84DFtYS3eoLeTgJQBgJRaBc/EkfJ5rCk2YudlIAsOp
+o6Cm7TCJg2/ezfwiNKhXzPQkj+0+t4VUNTPh4s3OWjA0P7phU4kPXowj9fyHelNJ82QUcQPzTtP
xMp+zh7wFWyM9mA7Jlm/e1VlBh7AaJkh+C5YI1+Dvx1vijDDEbRryN0+Z5x4l0Lpg1Ie/iT3OqYL
ZsHmssV5gNdAzdCEKylmtz8trMWEzB+EOHKAIw7awzg5dtTIsEBRudQwjhGoRi56BBOebCmZMhJ/
ta9mKjU6iGswq/9Ruu94dcXAfzCyxGy5lW7aa5ToVX8iWHBg0GHmmXfXiaeTDQGffsALj1MfU2ay
iXGqmkZSvE2b76P31QYLCE13+gbUsiYpg89IJHjpms3xm0v2fHw0qFUTUyhF+Le3clJpj0d8f4X6
eTsd0/IQHPqUWJ0kCRvli6XhnQDmrOeir+tKOzH/zFaWoWT3QLXvV5e3cRpjfWKSjEncCu5DUf32
ZkQkZClggMX3gHKcDXclNM40twsojfiNBpHTX2SmVIArdHHZmP+6KAJwmEZIh+7EYVX+gTYJYJUE
tHRC2CmRjHOG0X999x3tQern4rZp4v2MxidM3Zao77PgvFmrcv1Q2mXPW9DdkWrVNgbJVM4ocFbg
YlcXMpa2CeCsx8F0C+gZMRxDKFQVG+koy/4GhML7J4n+6cDip9LZ9No0q6k2l4rjaxlXOyy4mouT
OcPrXw3+MnV1wU81nvDttIzZKXe4fdOIuhozpyQ+YK+OEiMAx+SehQlLBRf2rH75xFiCehzo5llr
aqfhZf30i8omjUalCoDorvIe0eK7A/ibFDbJKRZSuEdeXCoCKvSXtfMzDZldprBMc3oa2m8NxviH
uxI/CCRVseoh4IzfeRnnvJrGnnHuCmeiXZx8mJ3MNW0AuJyyZ398z5d5EbKf1xgl+D7dMvvVAJ61
erwsbaqGPaXLPAykHppO/GRu6ir4wHCJTsfL53y7UW2wfCxz3ZrtZ2i8HkWEb7dqvEGqeOucemx3
NQ+FBYnYHA6dnSP3/UqHlIL2PquzMt4seclT/fO/fe2ICcJAYz73ranXUmcUiZzHd2toJVXyce4J
zW9WcySEuZ4KTwGugzUPviqINwB1w/HK+gE/onu96udhRd+9NlrdF0RQXxcxDR5jjDwMkMk8cyVP
c/lBulCLwXHlJ+CYJhY78zSntHqeT9Z2cEBAZlw9Ly+wCk1DWhz18sVX8VuxZp6DsldBRP9kwZwP
U8xtR55Cep9OhStQ5UvCEJPkAoY2dyrR/SkJ/+AhZq/gFJoMEZoDrV4rcdT1Rbkgu46rIWB5ZykY
ot1cl6GOuvNbQc+16jTPLuGqWOYGUv7pzjP1BGiKQDqOWYERJI6PULcwqXaBrHnIra/xHpRTVZoM
PdJxS6HH2WA2dX7lipWAOZqQp66D0fLoCbFZmSujDmeoZgiQi0j2iyeGs4qNCofOHZeGjtwZITek
5vN/RRbDvVyb083JOUR3SviQZPMZTenMaNjbIHXqA8xeohU0LyzhOA9NodA+cRM5ikd9H/Riw22v
RhJ1QFJtAOvEuokjaLhwwPOgN9jLZY6IMJVTD/UnrTnb4CTFdefpTdXHX+jGyMiOykoS2tRCz7IR
aDr0jxfHOylBr/bVnCMdhWRzS/0a2VVdTTke5LjKx5z2KGmi8CRLdnzGR2Ym2ebi8DewKSoF2LT4
b9iBCyS5UHZCUqIpFICvc1pgbOpGknnkS/5g/58pS3lGpFGqgrjb9Vd82zjA46hkXtqg5KpO7pje
aiUi+kBTqaYnv/RxgB8WZPnDdJ1lPgLjpbXID0UeSzXqHt43N4ticdi/vl1vDmdF1UYZZLXe3v4r
djmDSwZR4b8TljPWT4NuDvRvU8fJHvrCyZvHDe7zKAveddXUKaBhgHNK1fpcYhpx41NisF6LaKkV
ZuPz/wDs1qs/EXnyvpyJ6hx3J0c7UKoOA7HMn7D4nefhvArBk4tc0rhu21Kccdplf+LzIHa4TQv7
3rsrXiZCOt7L1nX/Sr425b9MIdE3NdpiwMhcIpwlHZrlLbI0Tk2DZOZn4rxuYcUtV/jrt7Gzshjj
xNrnvvIybbWxlv86HxTMfpRc7ZXpKwnWK5Ebb5gqkvnOZJnKmHHbBChcC8C/R+T4fLxbGd2SndJg
EwNdu5IL7lyrd/qLeY0e5pJGidQhBA0ciimgNhZ+SnmAPfEsms1Rx2bYmbIsJASVzTnkNwzygaJH
hPGt33zKMVH5OB7pNf/4qct9xVutw0mU3huWyTDDo0eDs04ip+Kfs0CFAskO+ERSeajNc73asP6W
g0uLkVFAWeTfTMObbv4sUZEGIqpLwbHu4vi5SOkT/cf4N4mvcQ19kRMR3+cWM+c3QCo/7hR+rQyh
taCeUfVRKdVTXiiKdgIFXr/aAfoHlPu9zFtjFf6kezo1ps84wsUar5CKLr+oF0hSA8FbxSnRYY17
8lIj6wRD7I8SDYwAH2rsd+PMMk7kTjZyPeIVlTDJEfJ190XQI9hw4GN/hMNxS+reGYr2CaHhsOZ4
nFPIOfxzjldHx9T3QoRZwy3LlhXqUoldI11OCXWrvjmuXEWGEcyvZW80g3vUfX8iLJmjeqElSRMk
yDxUjhlX8uVI+5LZo9tUYVIc9yQTblJmNWVyEBFxoxNle1RMluVq7fSr3so9GlLVIPdnYWJp/5QR
R3mK0HX2xgsVa4qn4+utUihCiaMVM2GZdgwG248UttINODstRD67I9gwthJob3hs1XQ6qStAYZmZ
TTA7pXGBjvkHxOi0h3VbAmNamluRBF8wXutNCPsduwzmye0vv62FhhOlvQ+HGnPy/ItBLYDvR3LG
eTu1KXnsXHBd3IUT5wTKoRdtCRkEOwiHiKCZurgZCTjQscg5FJyqRh6f76UAfkZIqwXN8Iz+ZZ6E
e9xIy2kJtCCwvS5Jp2Na6EoHAm9kVaFqhp0QMREtboq8Lg6jBpW+wEH/5eo0tW4hHbpKQtghlgKX
QipjUzeTw6eigJB45ww/tZ+7tyii+AEGh9gRaYwH/Ffo/Q+G/bye/eQ8GBz+CO7rGGDyI6CZti8W
z6TEwko5n8XcTGMWXyYGev9NNLh/lrUN7ZfF8oHduPeGeavP6Rm96XnqpHTS+7KdjVLPA0936doF
sC2OwAu6EW/jQixLc6tcenWH0qwPYa2Y+zgjnkZXMMVI0uoM8UizZkGPHNvTA2A48JcxHJi+V5BQ
u2Xswua1tXMaY6XYyYcjGnoEoZ1I2aBqzfwE+enr8GfZxQPwTeYRpq2ZHs/oPzOxgOpTjc1EX0vC
OucAQsIp9sgiqTAMRW4lSTe5q4QWYzjzPzWavGZvH1GCD11IcN+NgDBPzwAkH9+VxE6bq/QHMn6F
SMaGrThBnAwywsycTQHdGgEgr1W6XzUylAs3WBMn8nh04s01W8BVcfH/JTSGCsoF5j6CDS7AJe1c
J2lm6lnH7Cw7HMqM8LoTiIgXS0A72B/GaJQlR9jr28Jg+9vgaLzajbIK4HBIqFy2RocTpxjfyr6c
S3E4ArBoK22fa0FeHK0vlEpg0njhX317Yr1Qq3GpS3cJlay6gu0ZSrGYWGgFlej98e6Mq5ShyN5o
KbsOSoiySbzYOKBfASHXy/gPnMyLFXZ5d+om7vt/Xbk5N2aSNb213aFr/xl+1MrZ4SIwj77yLSc/
4V38Xd4N+nmaJLMjRc+8iEMAoWFiowk8KxyWGhxVmXGUNyMvY4iIWsum0ioVase6+Dk+BBKCtzDq
zpBCURxbrOROzP4CMH4wzCkfuHtgDoPHrb6Tjqb/xbWi1k3SEGRb+onO5h5hBCQvLmD3LYbxHYBf
GxXfzU/9IJ98Lvv/0HtUc79osND5e6WAoZCO5bJ/Gb8e95lmZxiOVgD7EHz7VCu0MXyFq7E3LYi3
fjJXqXeoLgMt52luJvdZQKN7qd8Ci1N/trJTU/mgm+IhjU1sUTnJJ8UeACC9UZZrF3J7DNbIXUa2
Woi6PcLaNwI7hsPQPRypjtpiNb9UPgMhjs9BDZJwYi3dD/GxCO2WyDDg6vy1zRg0VNL0Qhy15X6d
0gzsbRztn6/DsIE0tkwcT65eE0r0SBvkClsZePw0gXPzLVia0uFLhtLgV9pyotojAFY4PXiioWYC
XcejI1xG81C0eEHKqOh0dHJGEiqXFEI6IHgTTQTfQW+TZkSrgRiJOzbT+d3WMzGoYhaOAEf0WJBN
Q5El4P+XOqsfq3uMq9UxJ/w5ocE7CFRyVSq4vWYKUMgw5IUUhTWtaYfO5LgHgFyDYBp+zyyooRLL
jH5eUzjezAe+XaZwvorZEbCi/NbjR2XaY0sLTkemtLRLIQcIGqu0NW9jiLyUFrT2oJO0B4PidG7g
Xt3oWfA0hnTGRXSp5qSU0mCct0argRxAk6MNgWE0hYxpvgyHzjSELgegBkFgn0bdQy/DFxXUSI7J
/3rdZF38FqNg+L5XTQXp963lR8wsV8Ep5zd9fzH1hDal6Hml6UpNRbqhDWjkSLEqroivMLlSp4yZ
9uKTCzJurAEKqYFyxQRITCUbVvm5K83XgMffqJcjjaiBegoui+hfConcOr282dZ8sppCUrOGnGEv
BjF4UnxxyuiGAx6YxcvLa4alcSdOjWzhjNFPZ1jSjZIYT5T32Kj8YWkNr3pnxmI+1Xe8Xy+zkk5z
mTyg08LjVFxVezA01oBnnUTzzsOxl49i0Qp7W3OkrGMLsBBPXKhOAWMwGZyGV8BzCAA4myVdBCLz
gDtkeChoecKCy6z9raZd+uuxpfWcQ3CEd1VvPW8qQK4tJdCz6ms0gaVlhPH5UHqR6KBJmAlf36RJ
BbVo5lgx6Au4OTj9XGL3vLMsm5kUZBnLpksN8oE56UlJ3Fw+ud/5L+VRBYV9SD4vND4YUlWSkQuZ
axsKzCFKiptvqd+deNEkJ37+Mrl0zGZJ2MXjrfYZDGQW54a9rNYtPau91433NQ+i31fdM3LhhWNI
cuW7qJAG9mbfKsB+3DCxzvx9xcFZz/QqC+rCandcweKuQrciytU1ciFEwmqTSFGntF+bC4bQP6A4
0D2xw++VHx/oKtpNHuxjQ/SZlOaHAOgNSPNHP7m7Z3I+Sn7h5rkF8Am2Nfal6K62RJRvqMjFdkJB
wM77n+54peC5K9o/hyl/xevwXXthl7pwPIWRlmmBRDe8tNO4lz/hTGGLL1HS+u+509GIQ3T7rNh5
9KG1HUebfuBc97oXKeN4s/3MLj3+nKEKZeF1AYSSozav3za44ZTOvxIhJL3m0YlBIDeejpZEnIF0
VDVYL7Qp7QIoJZP+TmRFGGF34sEKE9O0uh305wSjSEi0rc68bpCZ6HvXazIKs+XXSqmiR6ZsgHVh
lnrvLqHtOgZbpDPKcTRu1CU8bpceMW+wPDnEuk0nvuYyvLnPcBKwF2fS4rT033d/hspKstWM2NPz
x6A2JZjo+60iwCLoCTl4P1BxlvP5MJTrcEDHhC2nB67wbRFGW/Lz5voVm3dfmvgrZwwQgcN7/uVE
ot7d4t7/FpI1prQXhbkSzQY7bbd3EH0MV3voygNHzSPesxevT+S26g0DoTwth2eeIwNFaycvFEW2
b3M/xxEdkYdpaIP4cHLlpr8Gh7jbknwqG0zToH7oYDzEyYKHrVYIlLObrwtiKx2Y3dYLTsdDrn9z
/Txhc6/CdjTGkxbGBMNL+oPAZXkmRrbzQrR03lVGubAmd5ph2IP/KgM1IYCJ0EYtaYFsWg/VBqcC
gy0GgaoX8TjVAuStc65meQd4+/hAv0XPSGuJsPBHjjvzEKWuoer5GaXNQu78Kcx1Uo55niOLqZgf
oNulMG7O5kAt4+89xWUbgttJcn6iWG2/hoQwV7o7uE8XZOWcCgrdZK7YiFq5XfjfHwZCDngEo+RZ
pV1jznrmVW/1YCLq2aXOnMg0K6+N7rKI1H3z0cHl/Hl5hH6F+f6NckAYDpuHPNnxTt/TBDMSekL9
NjJaXI4LAw4K8z4FbwcXCvYti087z95ZocQOonoh4BTRislHGALDC09w+rTTkGFi9ZBWHh53Z13X
s5txwjhorS3QBl8lRYAN/C/f9Dq4KA5zu5+ifUJzj3itVJKMZQTQIzcVuDcYw3TNqLVAwLO6a6YY
/8K3gV0iRieA77pB9DfdtUdv5Y7C6Xcyva1z4mS2CaJsiRR63AN3SaOKPUGwtqbMvzR/778rs0T/
ofuJvdRMfkQEFN44oUin2zCbHQM8w8/RMkDMduF+wZQF+e4wDtoDqBaYHQ4ykD4+WjUXUadl2w/W
2ZXpSTrVJhsUAJMdxBSo0uFuj9T7jufy14XSYj9YkH1PUIf7BFGaOLbQlSnLDZIxARpfAf/TtGcD
J/PVewyI/ZYa/xjMUa3fI0+Wr/HsOF6wTowYa5qFgF0kukUt0DucN6rPwVPzBJkJpNfrRbPuJpSn
xvQ8di6FWhH0p+GJzuCsY9UYf5FjriQNFYv8ESaN+nHciVagk+4xB9y7GGt9wMFMmfTl2+IRFfXr
SVV7vZlmibFDOSJ2ONqaMsXXtOP2dSpADKK4b1qS0Oxh/ZRPytYYr3r6xU6lUh6U9oNT6l9mcT08
GYsUITtx9K9s8WPyiDystR+cNbTttuhOb5bRNiSnMgJGgxgtrW2nS/cM1XFoDMCqgizXUNgY//31
7Npm12Gd8x5BnAQ6x+Xc+t3FrjpTYu/YCXVgigXc+z4fPxsHikpQbn1RnabKN1e4qXfRC4toKTXL
jPcGsTLii2jK6PnnovEBTcROA2ecJW0aSPZdc88uZRKPCJiFV3LReDgOB6/tULz+p9djiQj8sIhv
5GvHiEQatrnc0/M1uCPWIX7FCvPmwE8RpxsUuYy4LE8I+FeoZ33bC/OUVGYbT6/MEuZlwrG06mTq
r9PEQPuznkvEPpk1gVkAh3/LK64+GFM6RgUH9AW28rFgxzseYfwUIWN7s3OAfb8l8ie3a+gqP9uE
YaHgNzxy08utpAM/igUU6i5mNI+pE+N8MBy4YPAj8EDdVYWuctEJrDvUy6ZnsWy7EOCqv9KiYkzW
bOQOVwIwXcORAq/JgIa5NPxDdhrYOCfQU0Am4AUI2L8a/KVKIX5BWHjnEePSXMVBvTIocVlaZoaw
6UKi5EbrEwg1ma5fRvVl4ubBWyU3tzT3wHM+VroqvvEClNV003jcTXTciqrJ6pkTK1K19lPe5b5+
Yli0zGQA5eqRdKNx5h63X2XWxCPFK+quX57RA7JxI0xl97hjkVGwfod+Ryk5xDgphvsXPaxC8lHl
GRehGqxAG3sbrhVSRnU2qssJcibnP1Iq9Pp523gpi3RpiELjdmpRdL8ZFENBgHv//TSkJwP0y8Wg
SUDPZobtNSRJ5xIvpHGK2vD61FDYgzGaXlYxsy2DCoqa4PYZX0yDoDyNzVylbsxmdMlfiAg3DlvK
KJnVSWNC3Ome2cLdq9wZwsbuq3rWCN54IHXpjg4khs+hZQLU5b7+anst31hdkkQmBS+vcH7gCGtf
JcQGu6zmDsJHnjrU7y61O+SaxE+8MYbhEESyyARLu89WURiAN+HZd1jANniBqcFg0bFWJXAc2Bya
OpAg2hII138rvTCmOLtoCiBjIt7YbWPuhKVlnVT/4FJmtrnv6r62A6Rwm7bROc4HxZFUT+5KKWCY
m2sd2rcrNsgJYwSMnXV32dAs/Imr20HVHC0tmMIxxquK1Riaeku+I48vdcHfphcoWEumhV5IGDwm
ZBRVyuY6pwSZaA9BjgOT51T1N0xn/3CzHiGFuF7M7SloDSgc8uetULEmL7wf8RP56doULFbRxhCd
Tal4vVgOxaYEPoxjfWhRWVEPvRKFN8ApcWD4ZCw4Tsj6+9YPnL657fXRl3E6CngYV42t9GLMVGwl
rmbZfbjQq4hkl4dTDeogml81irXs/PC5LOpoh7zt2t9IpE+Bx/LsHwuzUMA+Y+yYZE+nhKMwm5SE
h8sY1+jS2x6+S6SmSzqdLEBtnLbGLzwPsHltU27+PBa2Wj+vxFMGEpDc4GZVE3QXvW2ETweKPnvr
2K2Y539rzEUxtO6OPVLT/TdXLk8qxCQSSJm1hnCc+yvUOfryb/rcgCAh6c4aXgT76xJwU5WW6hK/
OIbwNPhx6ySSZ6gRD4Qj2YuvSXZCtMNfr+5IK5nyatiHWaJdWKtqNe9Jgua8rdSv7c7WlJZIocbi
d4ubxVs2ivb/JPPgYjnx9sA1W/m9f5alxT667hA407VibCwZ1orsMWyv5qmNN48ArC6x/gNZY19G
t8XXuzX1rYFZSZcg3KYYncDNzKz+WJp31wN+YLIuwaro7qwTMbPrbk0bu4SchfvlgnV5CG4Q9HGR
fU28xJeCvxfWry6gjyDjG+XesRnWtSHJtxFMxz2AzJQUbWru4eGYIG1BprUQ3azIkpZfDJTiSgsL
VG1qL4zemvzJiakl6Mie1W0SmlF8UiEbyK/bPF8kZK7z+miogsqVfBI6ozlDna1ACfn7z/lDjuTb
kRvr/agTD13ZK7JkIG7m27BzX+RChbYDynQRgiLgUcj9HGc4p92rK7a/pUziPxpF9EN1vG+SDVH5
G+V1XOIG9bbp6MO93ONNa2i8XwgHMbDBJzqlgnbrYi68iv8on+xlkMp4CFWm8sJkgG5m9FhlRwe5
3hAKCzVse7SXsdiuL5G73aLRoEYkBjzNqHYaYCZkiXQPChWwr6NT1pZfdNsfcV4ZmMel26hoWqOc
B6QgoNHUHLMj2tOzYOZDi+pe5JZoTYn3VCrXoUC4AZugWSMAdUB1J4eUBTZXPs2Pk4b/jkkzW7mK
aW8FIe3BLQSQb/cXq38El0tim9zaey7wo5zLJjwaFpnrqP3OO1AB24onjpD29bT54GBPXZJDwhZU
EaGpPRBwcrqO/FkX72WwgQt93pI6RI5N6ggSwD9iR4BpgVFGaG6W0DgnfQDXpcyFgP9AScYmEmHM
geajMfSovoXDb+amTjbgU5gufUq3mRah9fLsQosj4rHrrVx7L5xHrJfudehDZswUGYfFl5KVnKbi
1pIp/GZE40kpv6qu3AiS8UyvumUTW8WB2WtDVMxvlo+rL0D184Lecdd8hAQ5I2EIT/ACTy9WO5nk
H+an2wSu2lscJlgfdoXRe9q+CPWUqw7nGMafUPEukOiyZ76i89tyJ4be0WySix8vIvvYzDTO9R0r
TSELMZkNyTGvTJtkvSMsq4m9i6Ixxr1gdmsodPSVy2+sZxdZV4gKi3Cn56Abm6Py65JK2884WM2e
QP6P+N4Kn4sy+jIzrv1KZtc/TJM7zvvtUokbsc67hydAon303y5eQfNt/x/vdHtCU5ule2pHYvq9
eZ0YoDTw8MgQF0dx677q4OPoGgP6qOn6i0yUsVIUyx4QOcOprdm6/zeM2nwfnAmQOxUb/jYHc9un
UFqg6fZDp4Sjq6jPtnHJl6nZe8b5BPIOHlTv+dDx1HIIB0HuwRCeLhGjCxa9qHS0UZK5pEh7hO3h
WgmasWwuxqKcjxCIicZq7ECn6m7V77wosQ/N5APQOOxlVtBPJwzHXHzuiqxb4clSu87nCcXvOU6S
2dzNEGRnURMz3XCG5nuDPwn39Javt3jB39NzmhHieL7IAwlVyFmBoBYzLgnPTRQNMAUtFAPj3UZj
Sibb3xUkArnItyZXPBOhnvEKe9mLymzuWzHtqdRbhSaEUvEZ/BMUQbtr3WjrfYUO0fo1H464b7rw
rYGO1CgGygUK0EQsdHAfcZ1ycLvI5+EVcQcgidXO5jvptoEH+qbhg7QQoeK33PFl2rHVRVZnvizS
MKhIWzu4YhPC0fYwbcg8GpJmZjfKcBHGZBrEv/svbWbF4RpsmNnz83l9tWMHZVwkBhy+PtSSNSbK
lfGKEh0Sz2vWo7Oz3shl8PI7v8uPua1+JZRTQ8DHDWqngJT933NIS5GH09SraCJOsZe8gaeYSFKG
jFFRCx0kyT44MEpxS/s2Tws4EzWRDt1drqJTlUnlFuAeivikX3pIlaVHbcDgmcLDU0j0zCNHq+1o
q60cLHlCvvfRXuFv5gSdRHq9mGYTN6ERMXcL2gCKGQlyVT+eadz+/BKfoosTAXrUhO82m6KUoK6Z
/noUo2SkBHKImm0lfbtH1hw88ANNvmBTC+9xVSefAYFVA9HMo0zhJw9tUqj9GOPnxgpwJbNIavI5
o0RqgEKrQIIsf4rGnsOvE9tod1qg15vKwrAtHVCzYOiGffmYz8I4vOSUXToX6XKG8FtLQd/S9KxP
ML/Er5WMRGZa60eUJZIIjx1K3VHchzxI3tK65WFwKm6/vlq6uknw9+KKBysrvCi9+1DiSph0QGIS
ApLjvk8ZEfiaGJEQtINLqKWRW/OGNqRZJm1XWdtVcKTyA8tbnwirq8uwP+Cb/fwUTT9XyyT6zzjd
b5ZO/OvbzK5EZXc0fdgdldMqYAASqPuHrtAkmbAGtPmGq8iKoChKIiI8zA7WmlQVBV3fbusLl4iu
gxlY0IycOhNTrjrDmV8JDLhPr7WyNU0PZE3yp8x08INu9quCfSyhwaD3hLBVeljvOpmk8ghFWqRc
bV5X5yR9ZvKRPVZ7ENaDLsj997Hjl2Zgr0Wis/TtH22NA9gA/7I2LxftRmYXWMotVNMlcB/AOVpX
cW2Lv8mhucqIr5hmTtt8eu1lTIa8m+j72Rjm2pPskkByRcfRtnSqHZsA+v8vJWlogG3wXyi7zoV8
fX+B08RKVcOLGnqF8zC8wm9ywhRm/0I5CqM/0rEpdJ+eOd5ylMjrZ4077zyo21h9atbTz5jxr8no
qG+HiSDo5Z5Jcx3EHOfcpd8MeR4AX9neu7h5nMEIDouiM0LZ9XMkHPAr/nHPX5Y0rRojteezbPd7
C+ETCeBLaaFage6zlxemszad1ykRHRtH3+yQ7BMw9qF09ZAUwwLtRH8pi9thI/8VOR9Xpq1kJymO
B81sVsnS55IK2xGcqZSblW9RFzlxClGZ8+Z1EnikTCz6KOV9cYvNqA7jdg+YVjLx0Q01dcnU6lrG
cRvb4aVPxHdXmbaOtDxKCbYKVFA5Oa0eB/SQRc2C9RcXSUUl2CZ9GSXk3bBobAOYLShYAtqyT53o
qT2v691q00G50uCLOq5UBTxp2OkDywhiUPl9C2DFNqJr0p62qoZmirihntdRUWXjRC0HYtKFgGFl
qaYmVlqya/2kK7rwm00rfwg0Gr70+uj0VA5NYy1pNLyex81JHiokrF5Kb/dBO74UdHhlN+lMOJhw
JC0metvwqMF1epqgPxqWfoL65N/JihVaY5x1I0tvM2DkdujCVGkIq66yT2qcIm29EUCU51kuHYdz
5qiYYoUd+mERVpOM8LPalmZ6eVxbH9Nu7iA6qmHx9mOmTUxDwF4MaokmmgAKnXk0cf2r47fSKqAQ
lrhj8e5eyJphLOEmFNwAHxL+OMn0QUrJE1dxiQv3kr8lA83Hxbe/8uCC+DM51kBYBGhMb//4HxPt
T+xEHP4D+d5EwVccxA4T1zQq6xtJSmekRFohKNRrh3VD+NzS41YK9t08lCoGpGZn6LF9yHsz6MNc
GVxMri1zm+CDZTca6un+wyN5COBypvhx8/ZfW9K9qa3p2QmP856adxb8BvA2ZmWH5wDgNxVjaHpZ
bu86pmjazgpDMT1LWhj76zg30aKS4Lcn7YMnfGYQ7OGOggNCD8DblfVZoQxGWJSatyhE+XzJGnh+
GKYtEJutHgaPgAheTV/5tM7lzczs/QwFn+BtceKtDf7JV/GpSAwRgj0gPSCf1XhPCyHWQpJtzIfA
y8JEYn5XkMH5JhOFKZqdGkalGSLwGvvqWoLoPV9CAIQCqUzUqX/GT3tbrtvy/mIa4UOsjCc9Zq7T
LoB0lUGEv95+PagJ6pRB1Twi1no3WkEEh8FGd9vZOXhLSiT47KdTXw0T4GcBersTDgu1QKleLU37
cmH+YhMIgTzVeWco5OvcAbYpQmqrQiSoPGK3kXeI2ScA5FCgQRIxk6ChosRRTdnsaHZB51swWNpv
gIejD/HZ70gl+ggmulC7SstTfmqFZH9SAinr1vXrd7L3ZQcJVHKN/fHnCE0qzFd8Rn3f2yf4X5R7
uhTAgpodLiHN/uZaFQxVzQuoQW6duYmNafKpfJ3cy1WDAR5HY4avi2EZVkhc04DAr/Yr8BLgqCda
W/SqoldrS1TP1LcE7kc7Y3m2/UuxpkeQqakpOSkksiDQWULkjneYUx8pzgPp/0UQi3qkZVKbSHcU
LlXL3mt39ErtL4ySufhEFQ1XpDGp9pbV3CcbdRYksNNEMvztmPOm9MF2hPtBKjfaHo4v8nkLT6WK
GQS6CBc3GPIozpImaB76B6PUqKDNhTwhWJAwCT9b/UEhwt+aMivx2r5882dnZNL+idbgrTIMmZm8
lef4P1GKHhQP8PaC23pp8chTbhXCD7dWz/fwhA837lj9vNeBXedjVYNklatiCN9Zbwy9N4Uf0HJl
TgbfYfFWz8eULMQZgYewq08QG+2DH9mJWA35stKd6H+aHclx+aWovxGkbxtxEtHFjdOEfVbaCy8J
35LJZq+ALmcTe/iLyi5fViMEfRdKKvyW3/rTaTWHiAFjLGPTxYpVoUnfBYhokHct+1Bn8goR4xDC
3clTRACIWoqQm8ODc7F6u6DgKgq2mw1yvz62WUvVvkDxfPXlVzdnOrE0w1bPiaOW8H11WkULm/1T
bni3ZdT+lry4IztgnTVL90S/pxbA12nKftrblxj2Po7PgP3ncyb4CyoFAAU5clJ0h0Yc/VTjZYfk
VFgWpHG/k5zXDNMCNJ5NSRFK3TeOUS/9pua7UsW1PAtD96xSQpnRWq0fiFxSnECjper0AUM5CzFO
bHbNpBAw73OLZESDEuW31oORUOodq1Yu3aMEHVJFVsTex6SdF5n/JnW6R+SlAcefe36OeSQCtSIz
0cjjqAzRvChOVjLSWYmb8svueaqTti2yu3imvS0ol0klt8LL0c4hWgQEznmyNJT14K0Batt8fAX/
LGo1VeqZo4Stp93KPs2VtuPSjDbL13sjw6CofvdKnGEndLjIIdxIMN1KIhlvwVDswmEpMCi6V3yX
Z5Vhaynaiy/mxiXPb4MNmD+4iS1Re2v71lPRBjM86wenud4qlOWyi8pV2hLTyZCkEWccP1AGNc0e
N1Z8FRPOnlmqYdYV5p077Ns5LBdzTOwk0+fbfnu0rc7SxdJGo6v4WLDo56j0bePmsZFnKRu3F0CX
yjHLgbqjbNQymmi4ss5ebOsFSgLrwKDHrecXW0HqUO5fViaf6uFnuWLsfu8IG1Aqjk6/8b0Y2pju
DWxDCvyWAx3JO74HRMEK+fi1E8pNf+qfbKnUsEGrBIO94KcgTYsu+iOm8rwWBTyk03mvQonOcfB3
L3heNFITriIB90rJ9myFFJXtIUdGv0FnBRGXNr6J4/xURXnAVJ6P1gu80I6EGOs5hzFnGhDloYyZ
wz0CwE6z9lETm/HqrzgS7TVu2o8bI6caL00y5XNWr+nIxr+ltzxI3Zf1rXumRuN9DlkASh42lHjA
dr9/QuOpG8GzvP8gZJt404giI5i0xmQj1S3jztcUja3GhQpv+jum8Q1moEiNXWnmb/7SrPi/qvRV
Ow+xwoh9FCbzB5wCjOpRwwWw07/6Qvd9yJIna8QRiscMNaA82cv4B61n7wz/NOLH5kc9rW2zb/rk
gVbApDFlUok/N3BA9ThnwLKOFHkov4OJFRvDujKZo76epjKE4hdfzvYLfyZbg4oMcG/xAvbQ21Jl
yKzQXs8ERlWN8GfWgcR1hbJX9NsQ/pk7ykTJGPT0LhVnJNEjdNeLZaqr4HX3tcOZopptRH9stPVc
zNXePFqyk5CwYXLoKfyAH9R41tlF5w9wU+5HO9gRnvgeM64IVDSgfU4ivlxbiDeqEX+vgxODfaD8
Qn8qGvSNLoRA0EkYLd8fcsStHgtTLmQz0LmMTfrD7uBITqyNboTl6Jsjn5fmKOUoJgI9S/GKeTy4
KE9SWg2FWp9CIUbdcKjJu7muuJc9k7IWcFInnsysCzwFqjpVy947m9OwxBZT5LA3IAgYu1quRzip
2yCHsI1pWLLV3EkCzP/ifN03P86oougzUHFOpuHaIwyVsGDQF3UooFTMAJLbwGLvHEZ8GhO0zyql
KMbFWL/blRoEIoVunYfWJqCj+pQa3OPIEawm1aoQSXnwWRsjTqGZwNsLucFzlxJMZ/tZYQmwiMPu
Buz1qc9oBDKFbGh+KhqxWOZN9WfjVVGfmASZUkr8bFpKYCDJcUgXh1zitEvzwJUIDIqAC3L1v/vv
+fegZxsn2iB4LZFtoVojUtcLB7qIpVrw0vkGYy7wkJlTCnGLcjQwrDkM/SK5Z1hiRn/oid2Bus/4
z3qS7/mmJiR4yXf160aYRTd5k8pjpCPSySG3piDQDXMRizrSh2NTsrB/bW1tgbnutbc8LhCpPVsx
8XM5XPXbqFaf5smhCxCKeLu65LdW0TFxYkHAm+sRFhZk8KINog3RPV0ZPGLopQVtyaJfjdXILogS
OYYqzAnLL55l6tMtb2C+AuT3a/x2lF5ti8kbv+cs9U99mrDpns4yCFMohy2ri/VNnCjQqLKF2vf+
FYNGGXgGQioUc3jdGfytAp97lyHy4rfQQzhQrgQAmQffLW9r4XuMqlLTPyYVeqVTln2690O4MImw
UCQ4iVNdB4kSHMJo+e0XfYt/NfHUHPPgkvbPSQ/r0FJqnpK0b/INesnDoMRSb/nbZWLNMTBCuPoA
kY1fKhVT56N0IOIaTqRNoJ+gP+H/BTOTNfm+Py5/NpS/xIoR2kZYSBu/+4xGnYCQqB3dbTHeefoZ
N2YntnnsUiQowaTE5xr2ydguEWjVpvQCmnvTOAG3eGysn7FZ5pdkXvhfg4nC4M8QS9H4j0AtGhI6
wyBU3DLP2wP293RZkToRPPsCX7AKaOFcLAOxHtHmm/oFIdbP5vk4s9xAXoAD4/V8/hWgy6DQ1Gzi
sHvuOXYyWMEP2dqtaWBttgnUw9gnO7j6RfkTUqmujXvSOkKzPJvvSFOCBj/jEzcTd8M7Vt6ZuwpY
xLhvkx/gWnD3l9i+3SGjlP7F3AfCjfmdLaBBqZqowiKTL5WLUS1C48Z/9aXlz4yTC7ObVD9LvaXS
gUEjfPpUYbmqHjIHL740JE5lp04jobL51DJdXSyRf6U7n+FyE2Dm1Q9sIFOG7CtFglfnyxbjQK5o
QxXR/otpKCNMDaxuWLHrrlALZHIsV2pp12Q4Cw26w6LbIXFnCNcPiTI8YJ1e/fz1vD6SZm3tuQOS
DkldvYaYhj4TaEOBSoAv0dCUrNM8TN6tGR+IFpXLG0eaBvKLPKrRnplAfo6zZywjB4hcFfI1PbCh
tnX4OZTyRAEWKh/gHCiDlYLmj9jpc6pv6EktPHkTgyOmaHOw3bxWmrp797wUFfJ1Nl0k7fYKuo+K
96rsLZWOUOvjdIokt/LKvZ2hzfnEjq9uPQdHKzXI/Y7JDvhybuVJ6HzL9Fh1G7yFGlnLY56lE+I4
SLvu39pIItGS8zsXZxzxTlV0UyeMGGOzxiCqjZKIOVxPP9/wh5359S2E5chcp17Cqh8j7K/q/00Z
FsrxgGxO85K+7jMc0wspuPUSrThIk6CYtBl5FDu4M8ygYZMuXA6rn1QOL0Q3YiNUstrSmn31O771
Osb4k3Wtb/EnOP1F4lzlsY7qXlMuS8LZPLt1kKxedbhdFM+JqiJvwg+kN2aBS5TgII7KcOhuT7XN
ZuJ3ep5zfP876tLCKJf2TuSGGq9P/E/J6QNbZUys80Od7gVwOS9Uku0U22Yv7oAMC8cYKV1HirMn
iPWvb7MecvtWcbuufpo99C99Y8h1+m24lJuVKabYUsvZ0HAyIr9fnysuIKnzQb/8Tf8uQbY4amKe
R2XbfMh60Jn9nDQ09lV9NbRW/CIuRFCf11ZOtvZnRKqm1MjylYl7GSSrPs2mRmUoVZswSrvDtaJW
cIgi5VAAWPNH5ZD1clkJbi6IbWHVqaDRpPOmrS2iPXOJUeOWJEUWcQuMwjAGP1G1PJ5ewhpDUMyj
CLbek6DzByfa4afQWm6Y0pPolB0DnemdHNyaSxOkZrrWUIGM9dzsKfCZgywR2MBTEuudNpxtLJ0s
1p3/PM5w0VimU7HX7dVJQVIP4S1XFCTkVf77uoTr8D2VY7swgBWdBpkLr0WZDBd4htKSoBJYieEm
O9jJn+kUBzNyFG8Rb/IqkTd9BDkCDxta4VQjlJcwmBXFvSqZ7EPE92Zz2ae2GxP2YKlPx5lbXgG5
Bw1H4G9mkfnXW9z5aOSV5eCiJO0PnxTvQLwK8n72XQXXP1Gt0ihYpGRCCoGN5/cMx8BCrGNzjAfI
qunZxWwBtaidhXxWF9oBUdb8eKUUDCy/rh6rq21iNZ9nep6nucSiYrZDCIWqWFbqhmaLD1MrlBij
Tla7bI4PTVa0Vt6MZNvc5Vi+SmX226JR/0A27ZlW1o2UsAiemOTdUscD+J10tbrCXKmK6dKAjM5s
w0HvzovFEuRuMMQOoGFpsd+zVqTez0k4W+NmpNFjHi4Q0rm7BMgkvibaIZK8z03Z8aSnolHq6G7t
3ry4SXlP2a2Or+/gCZ1bK4+XQVWCu+ncDn/ovO4iq//C9vQxteignOnM/66nPxEIZVjNtVzpnXvi
7jykMpHgO9zRya2ob9ec/vI1A18E4aJhRL35thJkzjy90jZ416eFV+Q+N0/GQuI56nMW4KPjWTey
iY0QixYWJDBlcb4oSIoKcVtI2ByNipz9yR3nt47xcm77HiSLoD7jmUmasn9bvABCR+B4x4BBsgHW
+8RHEWaWrRmwHy98YBAzFB/1Ug19jvT9GJ6Sw1dHgpIFcNpDZDKUGvKetqhwwR/7h3cIjXQUTp9z
tpQ5KTtPHelGZvl8VmghWMPv98KNru8qy/uF6vDlQz6dM598jar+iNpA1c+Wo5o//JXHbHl9wlvS
ylE3eVKtwR85RgbWjbBTZpk+X1oVHKOX6cfLZQUEBzTBNjXQKnMPA1C/OiPRD/YvQqA9HAhcUfw+
k11ld0EIoX91HZwJKGKCBJ94ST6pD8B6M+D78ZDadkW00ec7SogxqkRyA/mmdnHHBzGwYR6kdyq0
XcU8ZBAJq/9CWeVnKpQ5nA+t8EiJeG9qX6774kd4b40s/jaJt4KdEBaWhYTnJ/EwkOhgzQgYYozZ
iw/JrTBVKyjUjRifL3NRUmWlmxkm7fO4jNOiJxKtm3A11+NCLvmIzoEpybqbAN52PNAra6wpc97H
pnydbU1U6F6hPBXlbc6nj8r1wI0idxtWKtixNTWjGzsTZDoRm2JOGGIUr7m/TY1jTzpWHKU2cI2J
XZi4fP06pXgqrmjtd2xMOd2DwBoJ7ENH2FRKUiCxDpNcWb05rbxR/avijD3/eBnRVWBB81tbV/o4
TfNgZ/fSgRgdNticcFsX6dluP/mftX61zunXAgxm9kIQroe/n0Nsb0mgPJcKWeIg6CjirS8j1Xjx
Cy+740U4TI7ulbJHmCl/zcFDGqzA09JdA3iqHGH0dR5wAqFAXUCejeSwm38gQGZjtvzNxTcgNbsH
B/EobJvrJ9f0HCGb4fBG4GN91ePZySJORyq3Kq1rY065ZGJz0NVgSuDYTsN46GprX0htUjhS8AU6
e+qgDcoddCeIepu31jRWTwRqMevlNh1DdVZV8jNb+d9mJcIuE0CC5Z/qNiiwcJzRuyK2G+Xu3fPy
xnd9QRJvLeLp0TEWQq/xVnuaLBPaWTypirSr5D27ZbR92W2y9lNid7wFueHDlAMAVyELSefy6FbQ
XVaDswFYF9r00nB347R7UhChE5Y+w2/xHf1R0vuYP5MwzXrogyKC0YUzx93ok2e9Hnn0t9YEEtFl
U/6XAMmlnGRnEaZL+Z1tVPpRDqaVVFHU012TnV6IDfTmUI71bYEi3nbdBTthKOR7DB5QAChma405
9qcR3yBJPUsUyBe+XTeYyNBi6OUhJPOkEyJN7mgZrxuyTxHcIEmXOiYFKBgk+mZta7uo6b6kkM8t
rb3C7Yk2T74OS5O9SHdDFntnpcmz9znx8sqs7OZ5GcPn2oBWbeRrxkOKgDCdBSzStWeIRf/EgUG5
AukF/G5mf/o6IW7aI4cTtAttRTOMg+hYEp7k0QGO54zyfabbydGUMHNqevdmBK7xJXUGENSAZvH9
IG8MLK3WJH4BKU+R1vXJUGJfLYq9jHfOogIM4/h85Rv8GAzO/AV38q3urJoGc6CRxKAZydOQYrWY
MlukJ5W9BOrbrIGG8pmiZ7J6xRkpyNbSLpbxrBdIqhc/1ZK3UMJs3FajPQw9gQVySzJnYBxii+Zd
cWZoe+/tsWAaxq+7DUqsW717I9yzHog9wFbDRoSBm8jJ/hFxnQ0N8tweRbU3wuO1r9pn+IwhkLHB
eTrlS/LZYJ2ddxrsqfBW7BBw6XKfmPIwSlJdBy+5MlV/2nRhn9XdNrU6j/Szb+OFm0bLaxlrl0Ns
hrZrU6ZVJxvzRpL+2LMFsX0nIpYglEBG4IWxCqvDhFsvNQEeQCeRkUa6BhBJZXF/1bzQzKI6OpQX
rLy8eb4jso7IgXtleGpgdc2XoQmnddF8TpzrizoNos9C8vcNDjHrFnk8kZ6MzY5ljxxr6xfirqLl
W0cHDhx8CbifPHIoApZDJ19EQUpy2oMFNXl0jSmt1574EXw1BksFYNxNtV5rhD/pV6V9+Z7QwZEL
HGTiGEnceq7FsLiTBK6JnyH45M6y5cnwqFPiiUwqWDqwdOEOafzKOd09ugMn9Wz0CmjBlIrceG5q
HgmIni6bN4H7o3dGuy8DyanEYzZdWEB7XcOttQ20T/XhdIzf05/tBLVaAYtm20XtaWhrSBaucy39
+pxoiptDYKyrPiMBVLpQ7KSQdrtrkaqfQfEj1z6zk1cjJ+UaT8l+w3CWyzQEWn/53UiVuDRenVxl
0uHFoeSgPRDBDyKX03J77fhgQZMg/cwaXzP6LqL/RUzYVvze5phxQpiepEYoiuc97JAZZqSo3pYV
59+jeTzrjzUQ59n/h077ssPax9jhyCaFCNh02EMgRs/a6aihe5Pct/YcLgyyqWxa8UJ2kppQAJzW
8F7Vd71Gw2h4NwU3FD69kG5YGLcgvulLpABk59MYgA6JvvAi7aeOelCpebZ1ZYoZASABp2oqJuaK
vEof9/FBcMi2yB0kFJMatsaV57ME56hUFviw9dxrriFZ9Mrn/ejULMdpB/ykOERa6YwOVUwncryk
Rufn5/sMoGN/rzSmHfGhD74ddpZMEvg3DH4Ij8VKvqaeBGbABYSW+e6bcTggpLAFryY0sJgZx8r0
MdVyonRR7xp7lTSvDB1XGZaOEKzriOFzmbe4apVyiAURB0tvS6BCQ0GLj02wUAhoGviQupylFacB
7e3Nhv6JtfJKp5gzN2lObe9GiCLpKv8BenNkzUBkYTF4v6L6vH79K5++itXRJZoTVXtW+t7yRLl2
lJ2TPaQ8SuZs8rDvN7M4zXXN68OLlLQXSb5Dgsa8Cf/ACO8vsPgb+wVwaU6+sxjjHNyadr5gSkGX
ItH7Pn4JR+gH4denMIXRgE7rdJGv3NGa3LA8NjcEjkHvpt4uGAezI/cBzyiXvEUelP0D2zzgYv34
6PR19La7yPNRXaW6lcPz8avqETACgE6PXYj9rGTo6w0LDLDW6QQtg/yogXGgLJOr8XxqD8AeJ1j3
s3eln6MWG8ZqG+t5g48QeVZaUx2ZHiDW5HYJXxxLCinqooFLIcyJp1yebOrfl+QyID0T3WAnd5pw
8rvaNuyVI419A8L3GIXF1UC16H83akeUgD46kqf1DzeDXZene4jIp2yj/owB56noO7/0fw+7tNsr
G+QoHzRTF8nQdH+7tMLAALD0rQsNvkJ/gV7rj4E6aeFCm9rKgirGS/lshFupKC4GyF+QjUY/kzcR
vAvznt+Ptaa+LcHO8QEZ5DPefvc9/fkEIEr9HqtPM/XEGqx8iB7f+zYfQ8fBBZrmCvgZrTEy1QlJ
R9QAECGJkQSHpKUyLcV3AuptwdL0ellovcz2Tf/wymrMuhE5Q6LZ2mBm38UiWOxIn+IIPepie8v9
tc+SZdHA14F+3vV4sTPQgnAJGbUIoyPJ/3CD5uwX6IQfmlvUuEKGdHK5oB4YeDLwAca6lLKOul/n
Ku98yH76WA+7juKJo3dKD42XDycczw6sjp1TnFc+anGV3falsjhoxfct0ZpBPMILYNQC418W1utN
YM7zPVa3g77IB/tqW4+oNWS0Yy04p5/0PoU4wWFiKzNp1uJO5e3v2S85oBPPu0KNvSvpLVq7JFAH
43fSmPYZqrh1LGFIxVkQYiHkwSB6l35kKxHZWW6pj2fnIL0VvIsmbRjtkbimqmhw86xMYa9synJ8
hCVdaA327I076G7s/KSqDo4g5ZaCqov8ySQr1ByxwREuuanonnWmDoMGB+v3WJt6ZLqvo46gKiQC
h+o0hMu86sYqbQA7Ku94ZXxRwp+9CS6sZPUheV+kWdGRyuE5WH54rewePIOWrFWS9fF47c6sQVgk
GdJ9m7Z+eoj4/mWFsbs8+YE6F4AsL0TUiNOuYJnJsSqvT1UznqrpoLBoaYDSwL+Vf7Aml18lMGnU
7/xiZ22/wCfk7qhV5p+P72zLoVShGe3ujctlJE2jFr9cleLixtFp8Oc4RZjxljWggZmjQr3n115E
W4k6LWw2STXwQMfp4+4mQE5aNU7KFtOpXBOjYzE5dfMjDKGFS8gOLzlnRzjIy1tlZoI/jdKrx/Uk
sbKRYPXGbgMBpzI9BEEKrV76u3o1cxsFR+xi9oaKQxJnqe6ODu/JCNZdOuYWuUs7puQQNuKxzpNC
jW6SC8GbaUe4jVgue72aQVU5ujZr9sMG3exRXJDVxwUU33+7+9syyasG8os0+VTwDjiizkCA/nmI
K8ccmTs6Me0Ua016C0TktAfip//PHuKax0whaNkjQIDltNyqdoqK1iFhcFFNCxroGReVf90sawIE
C69slcagQQ49te6HM8HM74TQCEkCS9Qbh2uePrUk+f1pdiN50vVx3Og/yAhHL0q34kVUCGSxNpOh
5mhzO2MJ7KVGswq23ADDH81dUsk06G8gNyBywqKf31iPdsIH5p8CIn1kMqF6FZ6iXnSN5yU2o55b
N304NAtis0VK34Qp9+peGfEXgFiLQd7gLbgRoRwnlSAgRzUGJKS9sKMpKZppmClkeeeHqKCD4v30
CONJNXepyQXxV8/N9yts7uKbaaSrL5sYU2VttqLEOpfDdLJZsX0adNOt0APbErGc1YnD26lQMqE+
hSempdqgInRppE+Lr60pqUyCZ0UERRiVQ0lIFnYbBuxb8j73nSCw4TpiPWx2ZMvCwfB5Zy5FZGZU
+lf2HGUs8o/GpHpl1uKNRYQRyRrVhdhSYIkgxeINe96+7ZF2krNFVC7S3QWQmsC6o8RHrMuVXOE0
7KSbDokhkIrLZIjxZzSO0fZjanjQitX+abSwW6f5zN7xj5I69wTAkMMp+Pelf4k/x6kHSQeE1fh6
Lq+GcqpUyOjrB4D/GAjb+tHKmvTg3U9y0204+Dnp5ZQVTxdRLpx2PXswbfh5WvLi7ltAf1XboZso
7bu/qVEtYcKwSpDr3v3BYt0cIr5R3fXvybxSb073atFwgzYmo9oUg7SsLL6TMfOGvC2dYZe9wUcF
f+Gw7nh1t8z5chPboFgmbSbgfDoEBHop4op+EfuRDApsQ3OnozCuK3AJXkXESCNySCmVV5B55tKj
2vmxoKc5Z1AZh5UCGcNDBo8XVp44MVe4cyKck6O7+FtTE+S0tNnMk9c6WZeoZyMwcnn9K0xFIV1f
ZheQ8BAQOfHf+vBwsu1Lxhr4a2ukdliyqHSETRu65pi96ti9S4nuI1VNYYd5xblfGzuUnHnyiBCb
MNkaryZRYv0wdibO3iBhtYH8/VwqfjA+KKEfORNK9DD9jMJJFhDcXpxgKPRKSKjoy6ZiOIyuKu/+
UDqwRFlbbbifBLR6ezoNsHtU53allamT6dWX1qNILicZuSaKHZ47bs80q7jtkeXk38CGpWYmCO3Y
GA/tVtdwUSfcZEbdhCvz27KBpiF6bVDHgdGFT3+Ka3nqg5tY+iprhq5n/H+OwHx4Xg7zF51mlYRL
LjuHzhLJn1RPg1kYMcamv2gkwc8eDzChpWgejf7kIWOwgVKh/60buf5rMWMcCrpl8oWE2aNjrB0W
ETizM7v+U9XVHyvLRm3Dy5PlQhRhzazKiuKDbdH/7AYu5OiUZF+5MvBQdzuqnHOc6Y/KVO9e46z4
Qdas1VDaBm3srMI1ht80rmmJZWLXobAFHsJN1mM5ndrYsw+AJc82+iYbeVcIbOWuEP7e0mrfL8zN
RYTFQ7WagJSvntpuTkulnkUZWMvZtlPY3DNW4+hkRx3WK9knjX+5aU7RCGu/d/rND4Xf7bRG3vkn
pfrImpd9/ZDQrLcZ2EFFRXqLWhL1vN7tktLnKdwrV4z2BaM92+Cb3B2h4cLv4WmVsUzX5FuAHlBD
J9dEpsMIe77DhYbjRT7LOClg69HYeeJeztDfy+lH2G0XkfxzO/nYEsuUYQaY4rvhDLCO5Qolr85E
OQqCsCfbHwKi7jt2Yjo2Rb+G7Web/gBu3nWFrYVNiJ/nNHubpsCmk2XLMi/AJxCg0RqwPHC5bEMv
Hn/8pmW7zFS8tSkWK/j8jQdfziH2o3RaWvwv6Ni9mdmpPrjr5qM6OCFEsZO2mZU8T9kW89Gp9sC+
7vLv9i0Qv9dzpJBkmL4VDA67JWwNEnpApEvJbAJqdLX6tK0S4n3YNGvsunh89zTx/LQAjbShASYK
7eNOTqampNXePBR9RpQPEn8RvKuGqYVkUfqpDTIJrFtLVB63Sqd/Z0QGaQ9L31Qi5Fg12GV3+Gnx
gezlTbPXPD7rO2T2kIfuPFWiLXYGqbRrchd5jCus/L/HllT9dnjN5dz3lpz2TI53pPeC5oWGqDdt
Mvyfk0HeLfnvIKRoaz0KXV6E0TpYyZ1DTnODeg5HMcxFR+BF7x1zfr9vl2btegc+89SHoV16JmWI
i7jKbPGxvGeSHLmw48tnZnHEGZQTHH0Q1dj2yUds6mRPvESOqC7mOMspy8d760CGGkkT+Liu8wKz
LZoxBY/N0IPNAjK8hDkr56VYksHsp5t7IQFkY4+jPSVXevE1jUv1y6FFg2FjUnxAFP6/kj9o/nil
8CYfveJWCEmVxlRl9tJZulho4H2RtaJU4lqoDfWp60xB1na3z4VMLLdqyeg7RGQhy8FyPy7TTp3n
CJ1rPDtCt2QaRmOArmARszQtUiYJJDQeOfJqUblgCrV6rz/kzBBMpVHXtaGxX+gImA+IGVru+8IA
8QODANTSGXmuEZx3/i8/iPiJoX1GxyS98k4/VekqjzJDThuQePi1BXXEjsFK1I49wN5jCVXQYqhC
r0dA6sr/DDCaG6OmnTuh5f6ShtaVSpym8vmSiFTyRXUgmcEttC1PkqDwhuGh72eWk38/3JfTEWVx
n81LK6HxDB4rA8D/lCXgLkxmeW7CnFhQWxsffZC0WT6IJnSLR0i5VaOh5vvOg1an14KQbxdczdRt
GFs/qzpvLTvIiBQ8MQ55E/013OFi8Nev47y1ZE+ENYKfkPs5lUpr7buasLm3iLwTpxWOAunMehbb
wwLJ+0ktwOwA4C5qYZyzFT2bYZqVjYJtkVEthqdw2NZMbuCTIFlbdc9gnFJrM9l+GMLmvKBZKYsZ
UudVqyjBHk72rZa1XW6CnFM0JAjO6+cDZqB4EYEoIwoeWLZvJ4CYY/spwOIAQPn5zUgc8X9j7EIF
nbRqGpkzjkBAjmHjYh8LIeIJMInAtoM08MtxzfvgayYpHhV8R876xlmKqDCKMSjn1cSf2hWkaFN1
FPxy6TOM4Xpia9gln6gUjolgLelAD88O8v/BI9TCe+OLRn9Zd/Krb+k+cA2m+MFEL5l5CT/kp6dO
1/YZaUNbJ6SFci2PIiQQfS5QqldsloEJc/RaOq5D8bnYTUal8ZIi2h7mRwKFoa5VuF1KdWjUUB98
Yluhny+P/cJUiHVDINuw1iVdMzlvEFkPXiW4sBz8OrqvQRNoP84li4TMWBOLNREP8cJ5dLDZBXLg
DS25W/lYtwf9LIiuMmg/lKdRABDSE9e/wGujn8Tur8fbV66RJNjUVQqq1TcerBRoBujLVxosJTJv
liMTV6z9rAbCnbXmysmo3zqoTwmjqZiL8YAqyRGLYx2vFnOt3ZlV3IzaWwWlTmzPim6sRcTwvXTv
SrL5ChNoSdEek8s2d5x1xNLQidGlF1sIGTASNmSK/rOw/AXitf0xtTphcDQumeDaFjY1fBip4Eij
61kI+i0L9gQ9499hrn56itaBN3GJ/xZFzgL14XsZdHv1yq/UpxmmWccZP5cnP8OFb/cKyU1iNoVK
CkB3mGiHzgZHPA7B2EZeHB+mtnC+7IwvgW/32K0Ka3UnBk19psWNVeG0JDPL9NfpgWfVIczKiYXZ
ZDipMmiV1FlmJZxpxhILUcfGw2sBKEntYlE7FkHjzwtnb2trlsVq9zGAzVB69gAtRWpwRKWZiRMA
c0nYv+XsF7K3QoU2q+jZBtzJczU/C1dGGcpT55JBh2tKYDJMnBh1toF4vIjgb4OZLUThGFMh0BmD
y6hlkzuojsBBnVQTwGxbAmYFdi1NWSAXQ9hNRl4QQXglPpDjJ0mA6P/IDaLLy+Uo2cZNlMZRJgaV
l99bjm8ggOXU7G+qAzoUafV/tYW2eVjaku7msUb399A+BOf9mCQWhrqRQHwum+kZUb+XWbDy/qgQ
tcPtDJiotRt/4PBQSYqXafj6NzQmwowDY7rEhO63lZgPDceDeagjbEdCi46qsltcfe14PCF2euJI
wd1caE7VvoaC0dfwr4UWLXfMOIjMOqvQWWFMPsYN3GL4V7ijsFz9NmyEmYyjgdCTiava2y1zojN7
7ydx3LWkaUjLds/1zqCRDDTbVOwS+VGi0eFg9OCx0+BDi17FpvPrg5hopVAhpYnfl4M1wzKotlnW
S0bfq7TTL323m3puEY2B7uoV0kUVzLknCNXmvAFWIUKHudzF7nw7LuyqnCXerG1zVcp/6ssyMKWz
LTdz6cpnSR9UFMSQNzav9NcZ1mjRdvOPf0azU1n9ss7OYvFLPGD8mHwpvFfT1Ok0N8UHN004QQ4Y
9MvzbHuzPJbcEeNROwBXbU3roZYJUJCHLypUDTsb/4SncZepjT3PVtIn9IGES3oDAcN0pfH+PV6h
svYDg1AgHr4TZjen1475aBYjlR4FLUcEU06lLqmQDzqu9S2B8eDquhnAArlnXPZCYNMOAUnJI6IH
2oqnvpIxmMrl6lsCJ6leTcPSDgtj29OzObN6uH1ltR8MX4oKlDHqWRmsayA17J7NFV/vgzrL1cTv
2FDmi1aH5+OpEoslRKTiMCQE65/Y8y2jHSsQHgqnOP34RU79VdLZkqcu2zTGNItdCkdjgPpKgQ3I
PKNNWNdPUTAkWelNTsuqv8TeRE3GjPwHAEx8kP9ulIY0GrhNtJx7RZbKQhjE/EE/G3KVdUah6+2G
Diuu7UxxNkN5G83OBls9UNHYFp3QM31xzYXZpE0/VkBqnfyZJejp3px0pJ2bvPKi7nyKLr3CU45o
d9Y15usnDMalNZSvlwXuvuv2MBeSCS/y1VYVNr2HpIV3neqAZa5iuKieNgXRZ+i/kfXGBCF1DbZI
uPzl9RZljgnIZfSjCRRw5MuJ4ikp5ZWH4KmGAsYPYHS3xr+w7yWqKfEAUGa/tyZJp1m+4E8FalTV
Tnyf5m6aG7bkphkP2te5Cw8yb1cmAa0aa1yh/KszAvJHwuxFjZj1fBMHboqLZSWI4PrqiJ3c82AN
WpQrZ2nHXzFlruhHg/UF7+qNj1EuTOPxNxgiwXsG2DEi3xZuClVGe7qv3T4C7zE9KT70Zvyz0oOr
NVKsULwRFAoF6skvjtIOL3UCdFZmDim17l3qMCQ5WefNp2mY72m9z/DtZMXu1/7OyYVKi8+ZLchX
U/O7cGME2CP+zpzDccXXbfOhN37uOufuzv5gsPhhATHhubqRKkuzm5PxFlBeETS4kzgFtF+YNaJX
YwimRGyvZw5LUi9HA3eWX8kKZa6MAfDzIgGg461q68VjdsXzhwsWM2/pziWUSj6eELOzVyEYwC54
4tFT1aOTTNE0LyeQ+e9SunbJL9c8qxGxDKMe+mUQ556nxvbCaGFBM6yidg4ID/5yL5PLOwbulmbK
59OeabHGkTSZQ68dCpBeBlnLvGRp8SOTcckjRdjsc5vdQd0MRLfMBZirYejGReVzKaaBpPQEHaCB
K9dx1s3WrrM/zh6cWLWrsFkKHhGEp/0dTL6SIfuXhKw3TAWvpfhev9H/ODEH4diXnO3qFO6eRX2D
eFx8XXOTq0wYT7s0p1DbUU0HH+CqjrI7gzrcv8ONnQIFAu0rTUGqvwjCGXVsV7MlCbcviYAVBBCC
CoCzrWB9fgmEuW4Q0XRE7g4m4TBHaGx5uK4ZHZOdh3c3q0qpJfoFqz/c3TKMZu3qq2EaiCud4f+A
oyi7C1WVhFViiC/JwXyWg00AZWnrH6igL9MN52azGHhF9Ee2LB24PT9QN6SJVUfnjmcBdpG6n6Wq
9jltk7Zq6++2VjWT11USDKtz+VvVu4mKzyIGRhus+ju/ropEeP+C5yy3faCdh11u62M5eMU1nYh+
TOTujXezY4C3jIlARmOKKHUn1nywLnxT7CanTAMO5UxMjcslQVjIDDWg7A55RQ8lrzFhID8+OIkx
0JtroeDtz6OYlN4/4c7/GC1UrzeJ6CGTCOt4MeEu8ZPhWN/O+XI9o6YKwkJY4OXctrp87uyD5JNR
Lm15KnrUclhoIUxF6A1JIuPGyLRJY3ZlKEhAXVF2RDjoxTgeWCbmp6wIbGZEFGrzzCRsgh3JeR6v
Q0gtbS1bdVHF5BN+iJuA9mqrilNV1A0JETFWNqiUhzyeZmZV/HqyRHnweDACyy0jkwzTS6ZtvEKv
ypz1GkZ+VsIvSEX/UU/3s4MGSIxTIWccqiM7oOYY07wSdJRLkLFbLyalJPxrPg3EmoEw2BXKZDjz
UG1hQupniPRBPXsxjNBU4DpgaWXnKZofTeZhK5Wun7x8lP2y88rbzzGW9x3hf4lJcUjpnNJv9Ja/
hBz9eC/5Yq9jbBqb5dx1LVFr/DUup3FL4e0O64Val+r78awYy0Ip1Qmx1GTC4OUHoiKk88HHMdyi
DtphHoQa54G6L96wV32eYIpkFjQacUdSdQ/P/NKXwlFJ9L4UItwVrONCr0VZGIZCT/IoHaJHBHLf
aPBjsMhjBrtrdRJiY7pybG21yab/xK4eg/VQNECddaoX9dDF9kLG0LFdJNKU4copsl1g2Lt35YQ/
USIbeVx9tAZoOonk+IniwVX/Hwa1zsgZuoErqREFUa+0glilPULf6HJi+JXPKtPIuL7jV9KShb3B
o3sy5T+9WuvAyd5U8ZNPYEnFl+b0iKSfP9BC208ZEo4QfsBUs+ARStBJGq3Pjgkn7q8H5qwRKZeu
N9m9Yy7iDqVyM4CUDeJPRNWqfIffdtNwzQZaN/aS65B/Ca8i/tZzgvyuarXVfsAI7u/j3vVdkjEQ
4S0JKHiOFBZsFHFHzhrQ/9+qeyoGaqjimjsCQfvuHrpkz0sT2Wf1AHnv1c5vSo8bKrc6wWQMwRjm
w1LaLcZ8aSY9vyf1dWs2WgrdNngw+VcJG5GuXc4VzCCcR3S2/o8R/B/gnFpjvv5kOYLLOXAUtK+M
fhm5FDaEO6N+wkKIjH/9SfuPvCB2Y15BqTQHOrcPRnXXCS1MV/Kw3wFrp17UVaOy2mVytuqUVRz5
F9wJud3BWCgyDrrLMYYCbtTvwM78o5c8gTgYhqcOuvJUe1rrLtZ+7eASKaFb/0RTmO4z3ge9BQ0V
HO2ZsSZbWb/PZ5LXY/+yiIyJbyCpffuqu04snATzpkOBuxuwJEDnAZYg4iEAU03+NS2Y80X6F5jF
5OMbj5JVxQViTg9cIvDh6V5bl2PZ
`protect end_protected


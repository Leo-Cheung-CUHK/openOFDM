

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JyzzRYOPvALd1+n0h6OhFLeJWpZqai+m9G1gTt1+XdvmSl8CM8+DESDkmdo/iSod4UV7qKGdzREk
xhurZL7CdA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Uh3HQ9MYQCOnfgfbo0Xs+fYfRhBW7I6lM6nFARWXzDWJdbXLdQDXYmHQftz1C1OLUQQE7C4dUBXq
dT00dZogf4QehqG4RWPk6d7F3tn7Y75QCE0Hwxa6uqjs7+oXdQh65YYvgBS5EKqouNQgbBWirj2A
/O6p3Dk3LXi1PDC7sQ4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
b03Avj+lw247JKbbtrBPcXCg9zTXOiu8jwj1jF3NjD1nO9GHqik84DfX0V58lqrsrH0D+SmqG4qs
ZDsMe6f9LVCTEnKWmYthPlt9PzVWNYgDu6L6HesLNnRMV9TjJ/scQsgpJN8+vWZSpWvbmzJa4V5/
YDFQAUnzZN4qlNwPAYykHK+zBkPF2e9FhnRcpGZL4OYtDTLMY0EDdOYsRLxL+5sELUgEdaIZNLVt
5nK+WNStkO1LGCDby8DvvdpJtFQVJIrmH5/ZqUcp+qSSoiyx85R/9j2BwYYfh5iQMUgbKoJOVJpl
AwOZ6sQzKTlp5Jo9k7AJXzWasteEYtt1y2LrcQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dZgv5mGQWdpc0b+WNxvFkdblBIFCaMTgSCbDL6OPVir/NIFh2mbMpEDlagVKrhDqtUspl2WJUIvK
WVCPokONeoUQUX2YXU/2M6cJDMwC9P0Cta9LirDQcX+m9xLP4zUi6s6d2phb20vdT7exxgjE27i/
OiMCLmraNlYn3IoSn6WxMekR9xOwc6NwqOntFAL8EPrhs2mFUXBlDxxGUDMmRoSX3KAf1Yljpkq1
ElzH13NNaQAj8EwskvhUKS06GtHycaKS0PJI6BoqZfR8wmI6OLlnwaBnwBU1OexxsuJZqD4RpnV/
AtyK2U9g8WHHDknhaF7VrWI03dPT+QRjMi2HTg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rGXoZHxEO9Sud7P1xF0JTgZMXtKljokTOQnslaFqfRTOADB2sm5nTbILbXiltCqL1pe3cX4d94Sk
hrk5vUjtSQvqWbw7xf+zcJNMMCTjilITlhm8G03/LWTrsTqgRt8HrZdU+IC6OfIUepPii7PxiHNh
LSn3VdihGfW2lp+slugMVUgGhwaAcblMBx9ti6RsCd3s5Cb4HQk5v6vch3DiAY5nxOR9DJupzHSf
5GPg7NkhFZ4zURPoH59I7BKfTTajBiQtJpQ3hL5INjQgkXuEonEgqG1GCqWtIhgc+RMEM17xgyxT
z8LRfywYV7oG66kJ7LM7+8ZeYA7iE7OC5ZR7cQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pFWUSIOr/mjqQ/PncvQ9tWAvzGUR0DluRbBMvWIA7v2v0EJSSwnYhoaiAfEa68QQ64JJWT1n47jd
yiDijsjOmFtJUeMTIbdZh/G2f1y71CaxbIPYCemOdxRf0RG53R1jYD+fpC9nHJTFNthGKbZV5FX+
Y2OeUQ85RLl/kbY+d04=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UcEibmP3nx2gTMiM13z/i1fcD0mpE0oSpX4V73bMBV4RliRtcJpTK9bJsaH8pNKFxCIffkbWSF83
bl4CMGv63U0uDX+XJnOXqBkNH38mqh3WF9bOqwyETCVmEfkjWqeWxwnq7Of5JY7xuUwX6hqf78Sy
YjyiaBwhQcFiwyxfeheXGDNCAxLDxKUe9RJLUilmwCUXjHTTFKzPIU6/TYxmMvhlhSgZU4iWRNSu
6T3hrxHvHM3h3FEsvqNIwCzPVIVfAS7ZURK8qWlUz3TipTnEiACdWQ6rhMUN+JygWCHp36uogquR
oUhba41/v/CLPaJ9RrBJUItxOGKAjzptwAB3Zg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23056)
`protect data_block
RYb4x3ZVPTiDwF0hyFNOGYb30K7gIljLdseRYjoeIC7iTDZn8LZmYwzWYr7d/rOVU7JZlSZ9JMOr
b+vbzd8EVNx5f8v2MjPcBkNS6fZrlGHnEnCHqH7az1h9gY4sXohQ4hSqAAeDq6IBEDVcxWAQBFX9
PRUfvAuiwCeSMykkRHnLqm+hWJa9JcMENTE3eVIXQ9BO2XPSOU6P0GoZ7lQcqNao+MpW0dxTLQpp
KCWvmMY3PsDPN6ph0oeNCj9+MG4TOcVfgj1A6I5YLtbannbPfAxtrPnl7X2FJX5g/UBwSrFP2v6m
CvAj3XTJysHQWVC6aekSTBx8u7A5+j2yHsCvkyIDLXsNHdl0oI/YBvLeMy4d3c6yrWiLnKBXnEsA
1K/Uwk2E9BkyP0pr72nwkNvOQGz76jvhc/Xjo0oGYve46eJ88Kn/jgSYCwF4RvvtaaN+dsoKzzwN
ovw2dhzyVXLY7DVunrM2m6JRK6/nL2Mw2CCDitB2XpImVzdt4RjVlupEyyrZZYjtZFHXBYp2tTP9
0e6Cc4xsP6t06h1wA/JCLHi9LRMK64qLxV6JvOkvpfzh7CJn7AjGXgK+rx8aKBiHEVH/Kc/0fjZC
+6A3VvisdNV+zaw2MQdLngMcRoLZhksYRYkYZf5NGLTPFHvnv9VLvDlEtBGPD8eQKvfjRTKWpyI0
9Aqhmaynje0x43N9uNFhaDEcuKSWaSKShUEeXYv933EvQOXdSQlAy/JC6Pk4UgPj9nE9hoUzKgkr
7eLQ1PK9/6WyG1ieXaKyew5Ig3jqTz3zCqqmWUfhZF0t5uH5fffhApfcm6/jBRHVZ+CuOWF/UuaX
AEmyX1HsHem/gJPUC6i7YaJ+FylO+EZqnTeiMhtUq1YAKWkZed8yyySHt4CK8UtRBWsBKBjiU7SZ
lTOrtnWjiPIEROCoU1MXPivJ5PDEzoteHgNGyVIJqYqqzfUBWQYafUXDioPJ+BL7wiFyzMQd0l0R
qKVxMm20S8VClE+BChKF7ZS+uskMhvLQkDouhe66YOlUdRp4UBmC+J2nc79iuDCpJk2N8n1W6L5U
Y2FkJPucMaIlAcgiW0s91Z1sGZHLZQddO6L3TGkvJMW47OCrFuEP9c35/5D7z1xZrTlkX9wIUkg0
7+9X63vGvW9O9jRamx7EMHVdjub8pIrcegUqhpU0aqDBf43kxO19i/rJ1des1BOMxS9C4zpDozGJ
uQI6bbhJ4kp+Sa2WMRbkzFPHmSTNNPhOm3Yhac225x9YMQtUjtcBdhIgOy3XGNaoN3yLT9wpBONc
99WTxSInsJ59CYUX1YNj5V1r8yR5Xsus7B2Y73anqGTYLTR8UtlYd0pMWKy9rXhnnnaeL17Hk/ic
dc3N5n+TlPEQEBFUw7QfgPl7I8/hKQD/lw6XRiISVfRT9fxarUR/PLXzsc1FWXTNu9D1H9+kljHl
LD+eDP2gcW0zwy6/2C+JhyVthaSjOd2jY767upTL30yWMCDowB6iB74xZ4CILx2JLUjIVYSxXsaH
m1n9GcVGutCqma/L8AW4yhOJ2jkoyHkyqPVPXfxZZRyXe635pA9kTNEOvD8KKmAb8b4oIMoyN83U
Q3H3lQhKZRwunlLevwWAHYF0MPXIyTmZzB0CU1/i+xsrZ5sLir0xWX/VswjIBc2grmhLZm0FhFw/
6iMfZuTJDcVmKkR47sQ40IgNOemZq0FpZtd/n3AD3E7BIwQvJABi7oGB3FbnZD1MWWY27o89Z0kh
bN/nNTtxs1BaHYx57kwBwdgvPaY/ZOGeuiVW2yEWOZRrGFJ6qC/896CzgAp/gdf2dfwc3BDLQ0V5
yOR03c2I877eTy2zrLyklR2H8DN0RG1apDbuvr1L5ibV1uqEesRBO9oUAdQRrsWSw3GO4nP2B29b
52MfW7g7e05pNmFDO4if88WmwvRH18xMQEcZr98kBfixwN9Y1s1P8jVY5/G2jHL+z+qLMBiUBQSD
8NrzbEXnByOiebrnfPeyCwug0D6pLBXBqEjHCjYV3mAPqB205POZghMa0Rc1GLjzba3SPws3gRhP
AgPC3tMtuRwP1MDj4rO1bFzYqrQEbpVk7kN3x9g6Rl/iqhYFmEGkvsR28JfuzqQpq/BvsVPV4OvF
JTD4TTJPe0mieq+bTsY4eR7m8Zd/+i6IrhHZT4Y3SfAhEUoS/rFJDTD0tCq6sr2IWzWt2W2//dtL
r+nNc/ux7mOQSOHWXZFv5CEfuGO9baN0zb0fwElZQ1xyToVWOlOTUbM2lnOKTJEy9ch6j8qVLpNh
rllVJ5Xn/1Aw8a/hwN/qp8i4UgohLLA9PrK2GSQQW7AwbpST9hHyrC4s0eQlS+GLT8pqWWS+XHLV
FytJlUQpA3l9l9Owb4sOB5EZSufVYbPC3I+s2pawtp/Cq3Q2CsEQ9UgxxLHFPCAy3AEcMCIF0Ioz
lrvoKyyS6WgsZ2EIvDse/Wsh2wU+JqNAftjvAUtDJhdKRN4p64Hp9BJmdoDjSImsZHvp1i08/0W/
kMSufhYOwSMZ6UYvCWbnDQNW+3breXZAdHy2dhP40Y3DxUsItGPdaN65AUMH+3W7Yln8wAywKOG4
W/6q/lv7t8E91Ubg9gqfBvpMAAGTaXBjkDzGvHacWZdW9X8uVAHyw58PaJ8VnFGardbkf/S5i6gb
xYGCvTwiyC0amHG9tZnDQ6Rsduhd9AQR1P6h+2VMkIdSBBrMMhnCoR+w9yNr8+aoTbVJDiAT3IGs
23LcyudUaalwxsQdr9qsUmZZbCnepN9BvLI5j6bDNiwo3r3sza4cooJycu0f9BcppiCkfgbIgOp1
p79D/hW9YMvH3NJrfjAOEn9P0gr9PNqo9/Qw8a4i0g/xp3r9Hdtw+hHez/ILEbyFFRgyaD+KxNRi
lzBZvuZY4rRpSOdy31Dl5RMNLNwSRjsDBHv2TygkHsVFJ93ArrwXfQcS7KOr7xH0+Aoxnh3c0oJK
MY1o8wj9432HUeMCUjouRnL9IqDMFF1kwSgD7OzVQQNqg52lAjIHxmBk/iOokXP62U8VbczwnuVb
Ov70oMdaEH/eDkfYkUemlqeu+mxiEFKLTTUpyR2F4/MHKZr54SQDh7LrAhKi+avizeGWK5WdMbmX
73H4XVyGa51Kl5d5Av7HWghKBTFhMi4nc3Fd6D0jL837aK2gwG9vM1Ms0wISMZDNP7GLed1CDBlf
ri3mzVdkFSOXnYfcbNMiaLbiNc2jjLsrIjhi+B4eFQvAnbwfR9eBKOk0LEvzXgHtoD7WLBnhhbx5
E032zlQrjHoUJRP8mUH9cVDS78EreTElLVYIzTuaTmHHBH0Ng05iX9WjOtuT/f3MKEnLZVgXpoKG
19lBogx6qn0U/QVAKTQ502XCVUXrFjjX9bEATrZ3eZYzM8F1o/1KHXoRUTppy1OmERw+uqkD2iaX
0EpDejWouAgk8CNOBsouFZzkHnzdHIIbJ/cqssHn5FIfYm1hC5EY1FLi2JnSKrOLhuQoxn2GAeOV
kNH/TKd/6MA7ea3hQn848rqTjZwSCLzELOYEHRlINYgiYzskqhKwLWeLbtKSmgL8gq5WsNQiINXi
uP+G5CNmP3dCC8M8A11HS3DuL8EZday6UjU8okgfSW+Ai6EAJcNlpzoJtZxeyyd29Dquut2c1JFY
0t9ViMzIuE5GgUMQt2zlLW8UsgSg7RnVW0K6lJJw0RgMfz2u6+ZiAomJWHc751V17hglGpJFa0el
YCHnBpnMf4Xt8fU6q6TjGCVMgetinbJvDcNSW4thE4K8EugDDpFKhtapT9VQ1Y/DDAPk21RC1DuA
wmM5Be9iTbNgJmpZp+zsEJMr8ebK0p7Ijw14LFbMQUezaPUymHSIaJOQBk8j1DrsolDV0lnmZToe
abuvdhtcDeiy374cvjnTytoGrsL3yaRwIr9s0f8xW8G+CpBRqPFT4YFmgmX/jukP/NnZ8BccqaPj
Gwbl9ov1hTryOv9qWZfJqxf3t0/q4ZSEYdrN2TZDatBikBlBrWhTAUKTXApXbylQFTtqzG2IaGRI
vNgx7u7s8LBbWsumFxNH3b9/7RI0tEDPVZD2cuK3eDzfgOWd4iYUmhqcN27WLpslzrrfkOJmTR0u
rQGbCIzvJ/oSFVl91NVKSAVlNC5yDPPjj918E1yUJdAe3Fzg88zGECPcdHlJbDlaQFYGxCCnFBar
VnctQGqboUdwV7saG521gvYmjH/oTJm3iv1w6umdT3Y8F6vP0fD2NlqedcPKZWU34joGeFc49QjL
qQXa01wJ1u8qqkK9nAgQULnPL5uqEGf3v1iyYHh+F5ENFHG26MrOr0Hd4V8b57346Z6UjavV47VE
mepTUbquQfm1IedDDu+tP4U+7Loa4n2hiTZeCqaPgRwlH/odPkehHZPBRdLz9f6YrtfZImZv9kmW
ePbQ+Z1H4SruePuo/guoYzPK4dGSBGMQawFkWjDdOrm533Tl3pSV+EV95ffwt6aLB+xPUCo6psK6
Gp6kESiy46UxSl+nhSfUPZ01lwak+tTPHxFpV608uzuoo0Z6aqR2onAa7SUGlTh6SqlIDq19ahMd
+YpgfDP9mMi/D4bFDW++ktZ9AiogWndsw2kgeyur9b+8ecJQLhEv+1rYjiZq0QjaUTJ7OFQT/FrR
1Axul7/OaCd7U1ydss+RS61v9bepQTzhINPBG8AeOAinoNlb8ZZ7jAe8idbYxYEqylwWRAJI7k5G
4lQlMsUpkOq6EzlnfLYkukEJvYZlHaX+lUUAe4ijm6mSF2SIAmZ4yD2xsPDC6xxHEXWTMJj7VJWt
eTZ7PZCM7FGqqJjYLxMf+5lCQR/RrshO0/veAC4dNNBQ5ZVPbtocuAqUX+uPSko1mvJrCgbi1GVA
hx6SSYBmY7jBhkqbdklUbOnAs4Crgu0Jh0M0wCQ4nEJihPq0dC5hUVkw5q7Pr43CZzV88Q3gcMIe
Fx7NG2HS6LuaOvAfcgTMaUR/hFQQOXSRj+EYzHd1GZkN2ZJtsCUZT6EWXhTubMxO9Ds/CIzxSnYs
pBIA77v2sAOfmF/MzAE574L53ZiugqtYlq3eQVpHtLt+tAx6NLq7/SP1I92VH2dfMyKXhuoZ50Va
y1gA7mCh5vRoS9Mpy2VRk+U3g3VNNTzTFevkqF9P5l86wzr1qTHtKD0+MMtaiizB6inqPkUzgcjm
UwI+zEEHC3cr83SzA6y5ZFjEUkfY9H4aRcD31EzuIvLKbvho16f0pLnq9Mmu+m2inMJlymeTE6jn
MCd5fawfpCGyigtfhtn2HD1IawWd8eNW6gT6WsgYhPymm0w+3wEJYzUc8lesvt8oRUmUIVhT7kJ0
URlaYN9ramJ5MwmGX4cDyZDO5ch+MTPHdD8m1iwhFrRxgvypVoPpAgiqKt0zcFamQoRPDRGkJBJW
chkJxhBKmrdoRmYvz/vRO7qfo/ZwOoyauMa1a3gzNFyiGp94MgUoQpdq6/KQG2DVqXmsUMQ54rTJ
b1GklGLYLhXBLUvIyRyDvvd7dQ5ZbPqH6AhBmzfqjXHqpx29/Pu4yFCOPCpxalLAzeqGOAx0xekz
lZ8w/XYp1E+65WJ3LvCy1gXcNqB0wGTnb5Qi1ew3u/Kvq/fO7bDDOAi9LZlVdFlljUPMosCtBaUw
eLW9Zhb0JF1HsvreoXZ2RilgO4dVXO1O8EAdBQAp1FVjNZ17V0KXUbLRFCC4L85ffOaTjY7LMldL
NUvJCOmyF0h6bAgdkZoIyDYBbrlJBvvOeZMRa4x9GPr5oYUOcHBVuGqPf1AI2AkAlyJrTg9zyglZ
dKoxdypmx7HJ0Od6n6BVj0dZKqcMJfVozMbrcMc/uWexoI4HUNnGMJCEBcMt6dJIJbOBOK5+ctoZ
SwPdDs2gZhoM/TSQ89lcarmf4Q067L/y3ud2aTJx2IM0rzmjnZShzyf5ifY9uUnu8JcKluYXyWYs
WUX9WoSh9O/5NyPLPw3DgVsmziuX9xBFtYRXfhOhDyR165qMTn6h4kYdsaDtlrdcAnde6V0H21n+
i1RwnGpajFcua2xBrrj+F17tl2TOoWTklHSSObIaNH30gCVppj88XNJWe+X4NyMkNN+qDX+JMOVb
7fRiMEzdtBzpPYOvtyaM7JTOpaqJpVKldOik2AkvZ7HGNbrhV1VKFe6xCd9FirUE7pZPZjIY9zV4
CA1tia8gxyPbklqdazM0m3d2qLUjAxKPf8NZ45xhQDIxYOAPD2rEjDs/GXcOrlvQQMB/wKo9FX68
StONqYiEcgyUEkdq2sXxfJYkDY0CY7t2SpkRsJp9MAB578LBfLU4a/5GIOlLOvRqXREGf0CFgLhX
Kndjj7r/R8QLJvkekOUIr7nzMew1QodemXePxksP1XAVBC266u2F9KvneihkfCi2ElYg+LnzKgoG
74mNaFZah7d+mmNimyx1uuc08X4a98aQqYNLa86ahICS2T0OX6lLZMlhteTDMlw948EmFi7RmlEq
XtWvK/Z8ZaBu5rgeF3tP+yTPaiMXSoYEQbAbmNy0FI/s2L3XzAOLvpuisAQ9+djqhukfPh87IByi
R+TeeXD9SOANoJIYt/CQDwikHGTTlcj5kVB68DVJYYBA8mO+F6Xbj+lVJ0fROMdStzfdAZgOrEdj
iv1SaHeor9wfoDQ1rRZNEYeMVrV9TdWcyoyi176KuB5H3lZ0nI2D6aSBhceVoRw3fSFmBE/KkST0
4q/cEB236L3QEWW2mdCJpFHS26IIa2l0TPi4z9hehH0m8bZDGDHwzJU45eSIHuYPlxSXyderAsSr
mGkBFQcOJMZGsiFupNRMdxzJANbAOHoAaPrUy3OWQ01uW7/+wOqSF7IFRHidgcZltMYgCNOeJcsS
S2q79qzXDKlQHAy5I7/6u4jRrguDTiTAF+KU2Jblc/NNXZkZb9LuoENdey7dYvHflnEa4/ojnnEw
SfHfULhcUKDsPTS46HyC8qUZxxYRCvrrImUFOKwgx5vVaP6njoxscT5cVyFSWnECJRVnV/lthfnW
KC7hQX3ihhDLlhBeA9zGqwX78VEoZU3BCQdke4z9aEi2l6yGvqLODqToNjOpYtRaZp4PisOzAxKk
qqWxVR2rX3sVfoht5cxYz5pNacoWrOopUiTqE2cgsxzevFQxplrBgyuhWFfyOqoNZngGJbp6dKwQ
YeCE45NtuiFbZ0yG17yIUPE+q8hBlMRquI2eEID4ELWCSGmM6mNWz5yNSb/06p2ElKDXjJpnA+9/
TfwpZX4G6u3Fj38nTd7QOzJ1N8ldIvrYtzqrKhWPlC/YlmsEgAh5ZgchOpZw+Q2GIVsopLi46W+Q
aM9p4z9FI78dfvL/oyjKzfpspFzBUjcYKG3sK/788F/cZJKFTVlkMLjPythkgirVwE0eFOr2eGZT
ERCkfZ6AzoT2DpWrL569vRKUKRB7q28xeVHp8CGSZyjyQJegtyrXcwyet7o32mSVNeBMq8rz/zS4
qTc8l0u/ytTV0eZDWIPOGZ3WHId21K/lbuTKwrycdgppfabk4p0W7VBOlkyo8MSE1jZcehWUj+CW
6DMXkxXqKEH8d3eKyiCpICJd4Yfa7aaGQucpY2Q3o6cAyGfzpl7wUTslwNYXKHjpPpyt0kOj6f1q
/eRWN8+GNlg7wt51Z35LN4q2l5iMP5QLW+yiA2NY6cVrAlRlpQTIXmVvIIQrkNThzCzY5s4hfoKI
DlbGyziqLSgFSx/3hkh9Sw7Hq6ZzydOYIs3APMw1rZq34rNRC7nHAay/IkK0wKKR0E0jNgN+vsLa
jgWRz+dD/i8mMZYUOviXY2YKeHw8n593fMdoONcq+8ODl0S6NDxHjkUAThgNa7ofqyWETOwJtETb
YJRwToV3fECZhj6OKnGKtweMJm6ARH0ZSz/ZC8XqL/pI/idqiUvgHNGO6aIhvHDrXXvH58PmwGoU
psIAEJYgQTbvq4KAF5MGG5er9yzBzvD9TETTZuO30TcGLjhxXorTPi0tkLx4mcys4n1SLr3z3wPG
Pmi1wvj8RGDXhYv51rbFMRmRMUYqE9xZAssx78VXc2o+oIO7ZNBDZqm2LULx2ciUu6GMkswocSlg
HirZGhPxiVSdSdbVRMCHjaN6o+Pkfzm+Wj+yN2c1hR2C8hRKegzT5tblb0dus7ESXbuNsq6+Q8qK
Zo4b/Y4M/AjpF8AKFF0SvKQaNQrRaEr4I92Z3HncgoI0UxQQxp11E44TVWMbAVd34UBIMLgy+5m+
JRniNtU2VGKvCK8sBdO/vUngXczsHO1ARjsYAaZ/GU9UXmu8kwaz7LTIJ9OJ+dj/mnGTWgrxfbQ0
8NtIpCS2CHcmeQ6pt+G3BfWq0F+Z4RUfSUaQMb8f5K0hYWupappW7ZkVW7Ppm8lZwiThdo8GKCmd
e+lbkzBAnZP0B1p/ofwN4g+lnKGAHZKKjsUjdzfenqLgFbhlCdzPsMpY4y/XQxJU9iZqpaB+y2tX
F7D/+s90S5+Ti+oqDg8I8EHCQu92Qhb08W7MESgdXz7e8iPbMrHlGlZyJwveWY7+fpOvJMomss4r
AYCmhs5azv3zR2Go0EHnC8+LqZqjQqGGT4KBMvAqorI1NJgCNyflaWoFxGQGVs4muResCeL90iHR
Y8mPKw7G+8JoqYpDmDPfMLPcSdj5J26uY3zuSQj028S7brsEdrjCT/4OGfv8l0gLdC5WYwSTPj/I
P07odEgbaLavI7bba53ElBzBt1XSI4FIUMT6WakLwriZLIDhfWT5sHKl6OdJtsTVRqr228qN9yUI
E53toRJqQ3w3E4BCa+mmnDMXQSsqtaMfjJmF187zRhcgUeIOM01XcVKMyhVvAsNSAcWI36H43khf
nEhw/HKmk+D+RME3pSHcBhU7DH5K6/yviOIqkxyv2nONZ0VaL89NeDI8et0+mbymkyRVNTneHIS+
fErBiUwgEqTgy9gNcclM6h4Cm0PUQn2LFPczpL5ySh9nkXEv6NRgDqKuddnqX/hPiBbyKrwyijYy
ynQmGdHdfg6fjLKXN7q0Buo9Xl3oKlr8G0Pio2fvhRK6HvRkNgejv+lMYbWDtJEXwEXr3A/UR5gQ
i6gMacKNfH1ueZzdddAZRPYRTIaYquU78hFYX66/FjwNCZrnE4Nx0DBokJM/IF92oc8fs7DIrCjl
tEODDMMLtwVoIb1S/nAiQLdTbNiqsfWjUQlk0fxxxabfHILrgivRrYmiQ+NLLR+JUVRvyHhNr6si
f9zFernrfm8/9S+ZpJj2YMMs0lqg9SaScotvj7+8g4TGGzX3DELTUhy1bR4fB/tPGj0k13ihrCBL
JuXpsi/ehtGmNnCgzRqsksiW/Jr98bLo3jqz2vCi+f7ylOYR8oLTpLAwE5VkoRyVH+qNA3mEX84G
KmsPca4zboPxsx2/85J5cGgO0weO8PpC0hYdPv1I5tA3O030nyG3Hlk+z1vgBwFIjYs24K7V+pGa
J2y4RoG19QbvCQYG0HjEhnZCBaIOQYv+CscNsvd1gn/amP2dvfnMy0R2miUGYwaEMe+yM6SqYNXI
G75jVNr5RG4OUXzXewbcWvWZw5VxFCmL8m3eGVe6S7OciAUfeOigIzOqJlbpi92iAfLLxXmkJ17J
cDTggHOcT5EjbeO7gb5U+tGCWKUvKet3DH+F0eChdghav6U8gPvm0tWB6+jWkRdVXF76CadEHBcz
AjVs4jMUGRzyq0J691GH++hUIDmWkZ73Bt/HwmpjDqcoN2AZpgnHd+jp5Z0Fk0yx9+N7zQtMdrQh
i3H0zHBQ6M/YsTkT6H5/EjLAfdkdZmsRbWw/9L6Tnalcl9AiW6r8K5MTSkNcZahhqpeSmyZ2NXk9
51f7fnbVRnx7qnNjgtEt6g80PFE92JMeXxLkm/gfqE4vYKOExEdWqDwTY9unqBVwQR6qU541OFzg
K9H7Et6HzHghN7ZsBeg2Us1MYYyIId1xeBN/YxvE2Umt9mq8jc8OM/4XQU+PiscrZd3rA6ADvHVh
zr6npmAAZtKHA3BAaLV6Z6NPRpjYmOVKqwqf4QMAewjkrbusc4YXSI7+DU6RY3fnKv4lvICbZmY3
YB6Y4P82w7L38VtrZP/QjG+oatyjbCaX4TKjR+sJm8epRV6xwRivlpMCtmL/DtYQoEhghXD3hK/m
pHeTopWA8DByeDweQs61FFqbniJQ11rtV+U17s3lCuOb4DvuwWLy+jJy0e6cNQCYBE0xY4w9IM3U
QZN/M1hA4miDqdnff0cKAZuHErB3puB3SmdIHfl3JVSy0F0pKqK4bHJ3I2K3baJVCIpvDqM+SDPF
G9AY1ohuhLGlDgU5Sf6FlZ+8xk+arDfJvU7lm0aMQELf8KL1m59mejbSuW+x5P/S+jbDRR9HD6i/
5mVxZUiK6FpAejWPQ5kvQ+liGiVHy47NxoMcPG45ic25qawYeHvjx+nhdT8IvoqaiI15b5IeNuiU
GZaMnlzw5wHxb8d0OXG69MnYxVVKTiPV8sT2mJ9VkNhHQQ9f8xHV4luy3D9/JoYzvqwMoSpVXfLE
J4fm5p2ixFsjoZ2B0prcpfIePt53VRQc8poTLjOJNT7IGHvrIk549ENfiOshW/8jFJTViKGN2Nu9
e6uLWbiomuDNEsU27wPwDDQe3RZ2PR2Gj0U6usId6ht9lXBo5HpQFIBVWWvz/ySzv0mb8mYqD6X/
PPUW8AR1hYgD+VPE65vKgnakLScLbAj94Rmr62GkK9OEWmn/gBETIeSzruVZhMR1+VEju8/73uY3
dLkyNJ5VvsVlg5goKL1+RHPmTDD2qXhgbx1r25NkOdXQwLkPmNE71ktdjRFm/vpIBN1YRXopRG+N
+jK0yuQG68kPMzXNNCDvnIL4m9o5uXBHPth84ohPlgHJiUzVB8tN/VlEp1AN/ADjK16EG7t9pbsq
hdjVvAabKesE27UHP9btmU27cDdZ01490KdAAbnjl9olTo2DLEu4/Lg7MAKwEe+7/or6hMEEfz9v
LpW4cKmL7JjybKJEIhVUakroRwPzZjCUE9JiaqV6NoCcqV4Ih/E4Zh/i6MwjMztjOT3uw2Yp8l2V
UlYZ5xiZnZIu9DtAX7xYZUmACkVKUB40+xLEeP+XR94L0pfayE0z0uec/sxdPdq9DV979ouJSqdt
mEvp38sQH4vhvomFJWKQMCHEQk23gVZagE8v44Mf26vRjAVazMLjP24zLnd11FZrUSo+gt03VEFB
me2OHT2M8VCA3KHvuhPJrOLSeFEw5ZUqrEVZAJVupcWbRxowBeyfPIwJxpzeWWePY2Xp9qOWL/oa
b21C64huYgoivYipk9vIt2x1bzETE2cHe5hvDWkUssLdIaP+u6C3hH6YPLhyrrSrvp4squNsJqqx
ug3Lvk5/1RJtGtI8y1/XUJhvLYj+agena/QOKVU3lgxRUmJB1Ok/nIX8Tm5lFpD+rEOfucxxFd3d
le7EDyIlNSRIV2TXkQ97IVkSaaXB17zTz4GeGJSaZxxwHPJ/rL7c7FkJ85BDjiWe/jyZ7BNVsY/7
8K9b2sm/HKnN1YANcrOvqr/jAPgh8f8tAiuCb8ui0a5VzA0SYrelVM1Utf8reFCENgNRYVf0MzCy
na+QvCqoH5XZAcixzVQCyELdMNq8iFe6QEzTu9ujLdXkuu9VLu1APjP9OIlcZAru/9SoGIGGWOOu
Adv//L0rDscdRAqNvZXxfq0p90S4TRC83JpblusXf1tJfu04AqN3Ck9g69qOBcvmpo59Jo2hLlTh
g9hmApiZ318ssjDA2a5nbqja+q+HLtvMx2RhtMztMT2+2RPzZplj7duntVxlNDj7kSkhEPxBO/1y
hXdff9DQygz3PI9jTLcCEwzG2DAndFfxHR021h0+SOfmGvuqoUp9O26jjq1C6ciB6E/Ksg9e46tH
DZBg3qTcGC5VmOMHQqVZ02cTWGOmstTArNzOsFa4DkgBfo2cSAVTF6IHoyXEKcYOqc7kRJ+wl2Z9
7QMAqM3LIGiOoQ+RJLT0nxuGzv8dTttYyDyt/IcEtGqJmGOLAwgzvbxZTOc3fY2lT/ZL/7yV0bOG
gdk4hXz0rBjaXiujn/xuR9ZYk9nHBcpNKP+1SAhtwMYeGBmBZ79zFRfTtJWOKUnF8ojsd/TLTJbS
3xPmqKLolpYvz1qHmhy2W9N6gvWf3Y22sc2qCEAUfWNRZZlUst9HEzg3RGUaEZaD4Zqm97BVWLQM
QzX2FI0OdZsyHePPUFPwPEquKyUFlplo+WHQZl/F7/g6zfjI094MJ01b9/bmp2XPVf++Z/t3YKNr
1VjwOg268S76OT+h5utY1ZycZDteNgE6h91TH1GQ+0B+ysDBbOu/SYu/wom3Put3uHtNfJjkGLRB
xx6fFpPzR29czoDOw8EOUeyAfu9NTN6gNFI1c1reOXR3mfQyBbK9A9XKAqFXhp8L6iWZ5ycKWqrb
mD+HgmWAA4gr2RpIcQfsPLI9ieDbcSnSXAcTvh/dOYq/Uf02XhZ0znvZ9DfMrDW0+T/UWbnUWk2a
u3Zw445rxNIytlZvwfMdgliRK6qiOgALeTe7ylVhra7ZQIdap1qcaFZQVMvAxh5xP3vXKZPPe9hN
Zz2HK1H3KjTjagZJSJfJnZOuVxHjp1TAom0De4rAQHmnxsU77KLjCu6PSPZad2BpPuzBbQk0XVC2
V2BoipuIbVhbtMLQJhOgIXvPwQbetwWJvN4dEQzFHIPF26WCEXZ0gaRylOhaN5dZyjfhrWx12GrK
CONcR7i6F8C13k+kwUJpmQhl+2+fVYWbc0iK2Mi68S+VAz+vG1cI20hIeAz68nskTmarbXgEzopQ
x7MNJR2KXYlWZljBoxhcggYSpCFh705EpCKC0gI1TKmpqvJhXcKOTUbOcVG7Y/F4sLMu+aJmStpC
z6TSM9RD8GrYQkX5RPV/BuPzkdziDlqDbmdFBE6LJ/wkWXPXrp8831Gzv//C+ffZkskbOXoPF4+5
hV0YQyBCk/TaCXQi9BmbTXk28m+1ZNJcgxbccWhvYLL13VXk5wN1rjV12T90vtaHLGZ+65PWV4Mg
TZjqTBkXeHj6kbCp3hZahDCZEH3+lrUP1p/7qApFGqPauM8CuDQa6o+tzyoltZ5Nuv722JZ5yhiD
g5ZkrZTRotf4z0Qoy9ECqVZ2PmcXz3lhpSXiiw1rU9P0MlMRCRchj5ChRwlzvSrfu4mryy7gmrkR
HYEgdAB9CcaFe2fD5uS/InN5vS8aAbUEMpu6v19oKQttZw/abGQpPGt1+lUEXw0D2/QZ/djj/NBu
Z7nekNXyALY/fmAFB5md1p63OtolcsnW0HEn3mz336+G0jp4L2f+ZH+NkDM9pMfaVYKa64EO4UeZ
1UbmOOiSllEW082+/aXJqxi59OqqzqetQLIaEM30xgUnAyHP4ys53yeYUWjMrtKvxmBV2rnEbe4X
Z0X7QxBYNa868tK63VIh9cZr6QXyyFR6ddQj1c4JUPwFteJfUJkxjS6GztQ6vxfSZb1T2Xw3LfDe
X0VhtU0JAB3tBuwDHpVD9sFdsaoCm+yUTnxn8FdymJ1xh9sKi2uJdJPjgQeNw6+o4hqBkDmIQYKB
eClY2Ov0zqsQSboxonr9sj8kJCUvz+4um+kU52reiZcKuq+W197bDd2uVCs+MaOCl1RArTJjGteF
YXJO6075XPV9YwnnaqSPpECL0Sl0JkpxKlLHZC8JUnWHDa0azVKvo7HU92QeNUwWjKDDjjbOAvre
auzMAH2mnFzucprMgjDtlCWHGZjvCKRNGM0bGlQjXZlqZrjXZdexriO9Nbk9YUXsWJQbpkTsyA86
R2GjHCpHpC/TQEFQg8JwkbHMy4SjsfGis860P9frgyp2pXnR3lFZPTa+JUWHQYZTsvErzWQwBJMP
J7nH2ulmHX04sDjfvSFIr1wkqDbTrMkWqCk3s1DS5tJ/5YpyEaDFGAuoTzLGFai9e6E16RZRbOo8
vce5KA8iOOEXa+52ITEN/t0TeWw3lFNmA6QH+k9A9+g0nu3tM+p/4JW7nhbzM9LgmSJtFAqx+Ufk
mg00y7uZh2doZG4kUsnUigZmecqIoZnRSIwbThvg5EDH/MfjIc0F8scXA2CUP7cM0M3mt4Uexu6T
GsasXVHSOv5X6teR9vMdNGWX3WTI17Axi64eFFBPyzDsDv4cK26GEM82kT7wYeCln8Oc0lVVzxjj
o8Bv7/mz8iHJd7wQD/fMAszG92ZtBOsrQ1PRePlOrBP8EOgXD7k3vW8ZkwYpB007s0CtCdfygpPa
yOzsAHqNFQqoENPy9pgiUu8ka8atd1FelnO1n8fkxKpbT4+20yrk60ErXZDWy67SPQWs9wPCeicT
A1Fa4+ejrOoxXG5RTD5uSIqCnI0MPlT88ISzN2V9z+k4j/4+lCEwHbikh2NDiUx8RtH6SRVowuJN
IDArRgf+t8x4351OtfR2DZEmBIYJqciVlzUWfDleKUXO1ukIJYGZqhuQQHtP/UaqjW1I+Fd8UORf
6pbxF9Nwdo3Pz3Yqzl8xHj5ZYbOKXNkezwiblStXC2KMvJPWBmQkClNBVzPfKllkh5ILcoT4wj6e
/WA1Mrk53sLdKl0yPMsjxSLTXxFZPuloIB9xOoIzVxF4cwDXgFgs0pX9ViclN4/VxFKTEQUY0L7o
0JvCUkIUV3lMTWXHZoHdHe1xYQe+AHnKyZP3OqXr6bADFR61Z9o0ThjogK8/tYGE84xHHMeh0qLk
PGsZAPn9zJaR0X48EeV6TUY25cKgkh5XUKCJeXoNZMKp6avt00n443vF4VzOf5mSPM6ZOVlREqfi
u4aSZileUd0TZpxRgHBWtWkjI+9GUKHoaTSTfoNZTYAXtYsn0QpsnbIcZtRUF+YGnt9IMrXcKt5A
MNM74eecO2y/UPCcTpeQIAxeEDSxDPL+du5Y+hDoJwvzY9Nsv6nPHcH0m9ElfajsPa2pUUh286xu
Vdtf+ShOMmO8/6+/YwrW+4uCsZJdNc8HnETqtOj9KvMCWe9c7MvBqzNovay9ENA+AO2d+lBETKjP
NEBSHNDVtbQI+hx5wdPnMOtExi+fHQ6j2IUKjwNRPaYK4/+qHMU3pPd/aWnrszkTWy7JJsSFPu62
+NrwdSItdAPKjIbi9hxMSN42Z7KmWygz67rYAUH5IMeR0S35rpzZ+oqHaKKL7XJDl0t5Ffo6SsZO
r4wmBprb/IdOgyomLj7mqdkrhwWpcw63YB+lUcRmGmn3ynzmAJofx+gnw9XEhRkCRuhwa2Rd9P3n
BBpANns39BSghrDuG49llFJtLl6zTBItPTBRpVfO4NlEA9GYDOZdXFOw0953/xaej6Lk2DRiHwTn
2vgTZyl6TZ/OvuSHv4dqJWawmNxtflAqBHZNGYPPKHboyw9lU8suoyHmIg3Zypci2meb7q0uadCg
l3yRQvLkeGXNu+Qqknw2ZLlMG/fPEtu8hdhmYxqqBQXX5JUbSFeAfkrhFglc5W995sLnXTRp9CxI
Uxk/VlO1glMZEXtlIlzSes1tK13ClXp9dLcgg2lxMed/0AjCF4ZT4QEmxqNDuRHOm8qiZmv32L8v
NrZ2zgVXpz+7Wh+yLHik9d6n/NnKm8+NVQfih6bdF9yDzrBus1JEq91sAvciQ3DQ5LKQCZja2WqP
g/+sW0lEKCPYD+YZjGAczedoqGtKgMY2SgqJ/Hf5sZmiRWopE/3YnZslf7z2TCKJ3MkpUC77Wyiu
yIIl/SnMr0OyLKvlzaINoKfjqX0zHdLe5VIk29UabSlwU18jlDatWShwHKwtR/R14fomNpID8leP
V4kauSA5z2FuXb4rbqZt9rWJ35C1O+6N883r1xCerQKzYA2sIxe45FJ0eX+YLcFMZqCI6M4AjjwL
2mtJUbmCBkQ8cfCRcaRh645z678CEYDHpulbdCzEDDI0eUGKSlLiBOCx7I23iXYx4kg24QBSnAI5
6vitWZpzAgftx4gkNKrb2+IAZGzT/Ffc2Npx6ptOiSBLiZic9vJTxxMD0NPS1yDUpsGVADfpMUgs
JqjrDBDcuIcodmEz/2BavX+Z3jvzic/fsbnp26ORtmi674mJswMxFGPLQbFtHF408aal04FazGhc
IY6Y8UsE6bpm6+tX8oy0+UISj7SlTmPmR2Pw0cQkOD7GguUbUEITbYlWX90X3MGQtY9oQ5I5vtJO
mkAIyUvBX6DW0/6avXnfg8AoJUtwQBuKDbhYTgmWP4M1mZ+ROAZNb8BYxJX2CSaEb9BUqbPtEb9w
8QEA3s2FrLM71HgXCxWdQLgQmMB8czlEMKAlkzKHBbW5BF91slb2FO93fLLPdk2VbllMwpPploJr
jSDFTiA7Pdel1dRoEdyXxWAabD1GxJTwh1+Af3HnpVJmBdrOodAahfrqif23S+tl/+Utje2Tf4fj
7uf73xi0Hwx+zqniBMMJhbIxXRFl6fN3FXaDucYfVsqnbci8RSbs2qAkcUPBZgz6CzxGVWRSDPKT
OSklVqTVpMqmcLKshcqL6Zfun6goQNSD/zHUIqB6/2DssQYazSxfCL4hkQbZWNPCMY2Pjz1J3Yq8
nKECgVE88VR2aZNAUHvWWrtxDRL7MsQzxsiG4LFh5EoLeSN0IAbQ2jiBrBg8GhWZwwdKvx7Fjdud
s4S60lzXhxVEPPrNJS9cP/3zo6Wz+xPaE6fMZJjNXhuaNEU2ihlItD9I56KgQUVG71ZIF5nGfZoP
q2SMy7JmHUeoUFHYvP8AkL0IfyD1zPrArAMPmjclrReLAXxbxVqEuGdC/SCD2aHyqXEFxVxmR7Zi
qhrqRfJfAIu+JVEHtFQrS5XrrjkIMfILfiQwV2tdzgAFq54NqyplIbIHpb9w5JCJg2yqma62WOaK
R+7TDKmLjkAsl7fRyKQ2fFVFKA7IYc9Ic4AVG5z5IzSUUvq9c0weyVNTHT8jSAzu9ntFsQpNcA7P
UDO1S1qHIWCBUn4jS8IQ618NCE7UU3yqxO6AUvVx+PIJk0lPo20PYGa+XSA4rlk6od/olD9KjRmR
L4wNTJnrvlfzDBBG5gCxm7+8FKwH5wbDlEyjC9BfxEBGWdWI+mY8JlMPR5vodyF7Jf+X3F/QvSNZ
I9hccxdMIQljzKALnzUV9gAoVhxFLQH6FPC2UJQdh4vvEH0HZ7eX4wz5PVUQdtpZw0BmkJpvciN5
vV9gYqIMX+yL7RBSpD+RLyIpPjixDR3XsJIO0Z/NqDmAmePVSOnGU9SHVMxJ0Tqj0lN+cwGiP6Hk
cEgVQiM/0sHewi56KDg1h1lXTsg1EwcQNwahOlf7/cLOHq3XwAalhDTyS20PWMNvHhqR06/GvDU0
DHwxhSFoXmPaBJ3kYJrfaaE07J3/u234YrH/ncgqNz10ytLVat38TiBaCrgLocx3pV27CBY6bIyS
t4GPVgB3g4q9YglrLy1jeo+VhpeqVcJ40DvI4OgjNc/sjmofl5vIDpLn31JKHE4cD72ZslivgrFe
CCXKCasNxAFINU1Dyh+tHXkwJX79diGADMA/OER/ky8JlDGJUrcbG66viRAXklGVqt0lp4le1ePp
XcesRouSqvMoz1F+AELxIOLfR+JrbKYP7uWeY9wgVYkLSDUvHGGjXzosv2JeNHizNGQBdnqTU1Se
GwRZNIEoduWmkdm75jz0fAm5YgLZ0OaYBYYcaBBl6ee/5F04P4qgK1ed/x882ziPkiPeDhCP58Uo
6UN2T8owjyJZeLBVQ0NFNCAorP3Qlm5xWxbD0W21DOLiI+kZCfnelD/S12fhe8WNy9DhIRfEV+jk
O/OzaPYZ1qIMnCQQ6GdzBep4fugtq0DkMErEQ2397lpwUWxbxGYhXOF++q9t7ddAAsaGOPDZ7IbJ
9VAgc0m2cLWlZhAwQek2fjYNtWLKwTFbL6CNEljf7d7uPcHECMeQMfDQtDBjgstktHgZDVmXtJiq
yYZ1sbVMXNPWD5kqRIiNXn0/CCLQqKobk5eto0SB46tQS6xlk6nGUQ/ZtsFts84aoSUgD9QWg3vD
XKx8lGU8dvjl99Lw37cDaN2dDyptPwtCXMXIUfpK3eiBISV1dtW6lstE09XMPGHRXMT0P+5ZumV3
ddV2JKJqF5X3QFcvv52nTeaoO7+ZeeXCL0XTrnOMgbu5ECb/nw5sDO3t3xzdl+GJ1g+L6ttcZMPT
MzxQgoVmBBj8tjgv1fol+38+dNIROUojwQH6I9Plo4wvlpI+2ZDuZAPP+kpeimUDB6mBNx+vWKTI
7tg6oFHh6Xz5vKLkz4gJdW2lon64r8O/t+9TjKbolUTRQJUtxjursr6u1q/PZOIJXeTZ2EV+Jx8y
j3eBP1FBO1wq2lYdw6AmP1RtsozcbbbB7L7vapkqtpiOuSdd6aOcAVEDkmdW2JaLsJHTaaeyA2eW
ytTxSQ3kGEwPCnDGKX10G2CEFUlAwEWDNOZDwN2qPLBAF0Z/A1zMDXDN8OxO9kQTQju0uh2sEhy8
JUU1zWK29NcgbaU5SuaocItM0XJDpC3mg6GwTEUCp0AHNzZcizoCMwXH+7vm80QgC5aAp11TZnr4
r59l3ukpo9F9eFKu1rWyseRSInebx7RgfZ2i7QDYs+099VQQbNMUm9aj3UPykxh9KG2ln3sb+Rd6
E1E+8+fgwS45NPUA3xznYwxgiqYgKwvbID/mjt8qZ2/OGA0nSXZsWhYPtUcih6UQjwYPX1ro6+ON
4LrLIhzWNhIkfHuFdOO5NycEq2gHE+W6BcDxKQRwKsVQSCmLpp2lYugkum2IdLRGqEtdUGPrFJjm
sr+fAnPgW9iQeOer5L2xRemDPZPhw9aPe3eCz40GlezjuIt0u9eOP6mlgS0ZbQ6oKrys99ONBvDW
9bHeYWsgNZwYIsdj0Tw1kwegoOxJWH4MtrfLwA8LygllO3vQpTfRpkXZYPpz3C05EOLxviAyQO89
IkY+rdxHMPYfwXTMxf6m1aMJ5bTsqxMqPDhzR7a4K4pJzrqJ3AVBLtS4ISSzr6Fs6B7xybiyUkkk
oC9gmfqb/LiYTnU6QX2PpxIGKjjx9VqJkZZ3B7fa2nNqEYsC8C1J1zAPf+og7qnGh+NRmvl9WAXe
fDGPSWbRDHcpTswpC1tlsYfovkk8mW5Uitnpeuk4Uxij0YxnJPfOoKOgDx6d6VkATnnOGnRl/MsI
iT+JT0ahcc6lruMP8yCmR/cMzc0ubpZYX0gti4FEshppQj5VLcLOuMQWIcIHKb5tKS3dos9LZfZj
lErzkEHNlpSJ5ewllCSVaTiYYXUbqS6vffPPer9juhutWhyhCfn33IjAYkZtSZJfnJP8t9EfPFTE
Wh5IDvMGlNdDEGqyYvi+Q9mPt9wlH5xWkkRA+EMioxmvjrMUYMIG2IyFLuyQp7S8kOP+z2NZVeTs
XZ6e4U9oZJxvzyonrEh/syleVAxApKgP0lMXcuaRvoBD7Jpb80pMOiwxsEy/SFjJBdC+ju2wQGyC
Y0CN7aHRkgSx4k3p90MaiZdFS6uDi3fmDJvLyYLJu8664MLhuj1f40WAshu9gHdzPRRRkdwISHBd
kwcNsHm0KZkk+Xj9hTcGsmThC6LouSUGe3oAcs3wqAP3L6sQ4y4ktw69NLF7BUJHHoopVP5VXhS9
BauIfMaStkHVoxTvs5mskohF/obKhOYvLCmCUE5U8LOma5rHtnd4ZMlqSc6tmBZom9w8UXUSB5m4
RW0Gb7Lx+ujbha0VjjCOaujvuq6t5fxNLXidXdCVCNlBbTlKMSu9S8bPKPKtITzU4vBvx3k6OY7k
liO5KwCMPm4THvPxwOJjdY2+Jp4DsD7Jec1LN+kpSCH/xj4pZsJO7GRFL3ocuigj3ENZw4pqq3iV
91GwRQ9J24unX7njvQ6zO/mxoKTgxlvcsLO3R3zANnAnyxhrLFYdD8TlB3jVQlYJyqd++UZRMHFF
ONHV2FQUJory32DwLoSQ8kol92vccs/bBnYg4ct1AxKVd66kb0zWT2R9Cd9OnF5hjO0Fk1+Hx7f4
RKAtj972nnmBBkZZUf+LFiyv6CGqTIqB/HyvoeNyNlaFhGLbEXNEgMvUYn/2O6gkM758Ow/821VB
XRn3Iwpo+/thLBnzincc4UfYc02GXVj3e7W9nOoeE+CZtonMrNFKl80tUL0Koq3msq+CU+558kJJ
zEEHY44f7hJY0x0EMtbypbAOGvwKnTz1CHNYU5sQptYYbRMYGaP2K2U76TqX+eeyNIOdBC1vafdm
HR2/kcM4FiZzcyfeR7wk3ATvF4KHsul4XPqjv7Rfl/EMQAwBrZ9HYqUsKMtUN8bd9kzT12orR3xs
CC2qv2/DP5eHqvvUv+rOgc3moowWKdPmwpmK+mRUS0mt1WJ41dBZPyWcwNA0DVGPI/VEBs6JGXNW
WgOV0fJ6y2aRTYw11v6PWq4sgLyySm4lO+n9bwwm67Z5gPQhIUKJRCjE3bCXFeFbHdP3hqn97DC5
t2WImrRDPQR98S3sKzJ8s9dnYGV8AHrXilXHOrU5j39ukY+XGGPxU5bxGhm6aMtH20nPO0ev/6Ki
h95rgCkBveDkqM8UWRXCtnIIHyXlU+Jo1hcxpLE3vVtvjYUHcnSpWHTwD7dwOBtf6A260jfjFCjg
ZTbrsstE/gtoPyVDSPTjlBS9hh75YV3PYrhUmtADTevrhElW3rY7N6lYTHcXaDSZEF/0c2A1Zqtt
b3pg4SIflvqjnbEDdY5Q9/BVL4F0sH8mzi92kl3usqzoS6byQgwvmTgsmJOPsu/dBJ8j8iXAJ91i
S5bUJImXnXGKiaWPxKHlTx+HgFSRPo2EREDe0uo0WFQLm93co9LwjaRfS9PUqxyU4M7Co2GvCuoj
T9TfvHfsD8ErxpW0G6JtJxOrLUSNceFyA8U8MlDgAsW4mw1jEjy8500Ni4CUQwITKsw/vR2iMRRS
V5t1mdeB57AzbKm070aLjqloZN9SF7wOqI3fKC54TafvVCqoEagCMNLFYyGnKZX6OyVIsGW5qvPi
3N+CwgnXPAQPyZqDtd6ht4zL3FR1HAkEji98jLp8Jr2Ldfch4ZcITZvJLnI04EWm27IgPU18c2KV
mRUeZkKwj/Z4rEMFdpbmlG+0a3KB5gtgGfptyqLEdjhz9unvX1Qa5Uc0DRifn5ZP6P9zWD5dcABs
JVPkjIqiYXM8vE6GYEUDhIXSbRm05sVu1Cae1BePChEwtvUMYD9Zq0rbppBcfbTXT/+XdVtqkwKL
dnP46M9bTtsXYINjqo5tJJuj0rFbpLoMaxle9Z3fsi5HAtxRBi49vG+BvvO/XxQk1KI8st9ZQOrF
YqLg+qoqx+zVvVmJCKpo93cd1Uvd0QSGSd8CsW9iILnB5AaG10c1I7YEsv1EIsNdLmCGFMgWntGw
hgDhzEstWkcaN9el0PtiXn4NMuTINZc2HeTa9zPkjeS7NZVX5/My2nPsxgz8vgGnllVIOtoXZCzz
YX7RTWdRcCgVL3B5QFF++a4cGPBnD/JAGU4pjHtIfbbEZqs3TH5yNgN1gF6CM79vlz+FpCDqh0ts
3nSazWJdmBfRX8SVtKoicpiDsnuVtQ7mqVZa02wEGYlavmL5ey4ayL6JlS6/eCW4jHOYBCBPWXQ3
V4LNfxGHD+bsQ6sV50WFnfsOZRdl/u3KBVXSrTdhAo9XgaoHW6nVmwFBCRGvvsK4Dr6Q9seXzpZj
LOnfsDsV51d0WgTyi4Iwmce/OYFCFyt1kncNvwwtTDwThxPB8cLA66BxjOm7qIqHZ+XsBtelGrBe
YuFM3KSzhu6dklWQMnPFZIoCDYp/cuB6NksuavV5w6NdqIH7LDewBjJaXBstpeFr1qCkvw6Ohqf+
KSzh3Gaigq2hmE3uIf/qlVQvce6US/8pDXeLSopPGLRewjXpfJfpSFwVp+ZKdqZr6y9VQvhcGXH7
Dt832c+iqRiXJlLL/o8PQyrlafIM+pPCd9fw+lhv/kBV/47HGVAdnrhtSSO1CbBsj61YMqVk1jmu
TIjHfCs+GumEQjNejp+Tz6+YKzy+1B/ylgDdXYKxygtZzxpJbCqvY3GJ9uCDVNZs5CLw5EX+5JBu
zPyemBd03JOsC4ldRNdED45xJd5zXFFACTvS09PrGtnrvZC0priX7q0IMaTQNhqUM8LgobJAAVBK
XlHIkqgbFQanWeS4/rIJ3UrgtoTtttpHLPSOTyfC/8grMInuBtQMgKO7Vbv4tFHB7BbSP4kMARQc
KdxKJksXqQRchKcYRcVL5dI8aNlI4uGyMmG4AzZ80z6s0tHeb83VLhkMA9rq9LMGhdYS6e9El23H
q65tp0k23y/Xf8bYpbazq3KzVKHjTzuTjwBt5ciBL5z2xMwO+C5b6Rs6NcfmlMpZ2JFTAov3b43v
0szGI6iNw/nXmHY+GOg+95di0n0XXxdMDYwFayKrY2FYqLOQsjuxV+4U3UBKKb0yEx5ilJ2gO7Z7
tGirqwiECmJCJGGCJUqvdxoLq015n3gjisVnxMNJHmMxp2BBGcJPMkjNlEpbaaeoRFMYCw3bnKDo
ARKdJdWxbOgTy6AhCk5ePLDlyrkR8Tr6WnfHsXiJc1n1BRVkI4Bk1CEc6rK013SHfWzhgJjQm/HS
GP1s6MjW9+H9JKjBwmOCfi8hr9496y+q6FoNWlaa7ehMLChxucsXvpb7E4p11i1aoGIC791GWtaH
HFBMJprZ4nyuNzkySYFUMQ0nNsTInEwIAjt4MTA6t2e+XnVoWrQHOVMmRUXIzYEUIA1N59eqGrte
XoGadTyysor9p9IR1FjuSsExvNlFE3gSi46EVpxcL1aBQ1PJvG1eX6XVsJSjVgZ8k4lxcElwtxaP
B/a9peApbDSED2Gbogm84ctdBXhZ+vt4GfQuvYtpyD0Y3eIpm5l2T/KRWmaJOwXDrZ+ZBYM6vhKH
K8Z8gtknBoj3zgsrh+I6y3/ANj+5pfw+41X3LyzI2Zw7xjBzJBjas+P4vt6wy4+94IJG6KK8hPYp
/JCHOeu0jZE8uFMSxdSJf+O7DIh2ipKm2qatoB6Wc6E637Ql7FDFJqUr6Q3dIQhyFQ2AEkU2LsIl
cFGfHn1Q4AFwrHwooz8Y1lexRwoutcxNLr+gckxjiVdrX92a1BMiTNXD9g0mxizgkTgcJX7GXFpX
SfcCd3ADliAsCt60pW106lWWWtg5eos911swkVzPgzcM2TJcNUK7pFmo+IgQ2LYuN7ejhEVuDT+l
HIpcubsOssx13ByyZpVWKRBSRIXAaKIQL8wfrsEz56X/9VuhQUZvyRrV6OAVVkYnq99TnEIfd6zx
k66zYLKEZJeHkxGwfJMv/3Y8iZVS5ynHX+jkPCYi7llYA52HB7gistZga9dIrcOu6suA23Eppk0z
/RuFfAwoRPnV/dQOafMmDySke1XtWfJQ5AY4cJYt1aegVkKOZvaFZK3dskiwiHoKlMB4t35eVi0X
b0lSZObvPEtApnm2J3XsXHU7S+I/0nlR/3SNrhN3VMGLA4w/DNN2MPu2NX7QTZRztK5uUDorQX7c
DYnH9bkU0LDvZny4S+bN2OnmKHsBgmZq8SYNKVJQcsBsBmJ70rB6+dSulxQgtBnio39lcAr63c4P
tiUcCPgim+fybLWNxrDWbeGtH+WwVHuheCTyiRoeyO7HCGbw9KeinJIp9LDkILMQ918chfwmDEgJ
1ss17Drwh4ncrSBXamcheVupj/oLcu+sEnYR4EkmrpmznFY06S/qk3w7m/2OQPPTbcpPpCG4tQzC
wicwjkiPdoYMcYmqjcKh/Aq6pkmgcJ/GLh7lSSEvcBC812WgxTirrgNBIdtgWeVHH7azMWhSDaye
K3wkLk48eQYdts5yxSMI4v+AX4w7SnJNtrgm0NSeOUTWxwIrqEuLetP186Hefp9p91Pf1wPF7w79
mxejMbhNaFOYMaUALSv8fpZNoOHx15ClVxoGhF2A8sVlmSOGo+3ji1hDOMVlQP3Skawerp7moSoK
NgpOO+6ovudu47MsfgvqqzGsWtY4uy9pySUam4+iqG81mpvjV7skT4J1XUD1bFPdkfWan+eU50pO
gHdK+5kanoP8DNUTfRs+BiWdPylWj1NBehBD3j8LQ5BL9wTCLYxl9B37PNHrO7FNgb6+aQMzuJC3
diTYgN9zU1LDw3YHkZ/gH1sPuwEtbQ0TXtPcWk3M6UTs09c/iBomQABFqP+JOGpnrs69C+1+avb/
d4YoGtyAAmoIUbn7YVXFPxZpV34TpiA5j2GS0N+ySw0kWjQnJ5ZXY58xamW0okfnJtIoyaMII9p/
vuT8nrftRr4jfM/I4xPf1qWZ1PHD59Bc+rD2UYzxhCCgM0FsZGmYr3MyehDqrN4jZ35HE2e9zNgQ
ZoWfefbl3pCo/SQ3ryJFrcTE5rjNN4DPpz+qH83JG37LnGn+Ug6gzT5BQ9xpy5hjqY7bQ8EI0wco
EsUlXyjXw6KLzRDDCKgMOM+kyNk2ffiUMoU0z+ACGFgC5UHDR4DzylMsdCtLJ3UYz1a4tIjNlubF
RxWRkgJIatRPzNp4Oq8rRMoCb25y/2CmSu7HZOGXBXbeKB9rGuPwBGhupxC6feYnVjlbbYtOIfa7
LyuQDTCEfu+rjoM1v7sKHk+TWp+Ap8J12pG25+WWP9oEIakakVRHi/Oyz5JtvKfIDRVzIRLGcZvP
jYDPiZgBTqTCvvBX4Sqp80xD6JQzJV4veeyitE1dG0Gyi6ZdmaoB27tHWvkQ9dAQaxoD40NbgRZI
E8ZtpdrkhmC5TAV+7aJs6xWFQe1l9cUScjLkO77TzaJDh9GQdlPX1zYYSGgUQzw8RttIJzZb3gPu
81/93XlQBbw++0spPk+kySU4QNgtxFX6Wr/zwUcqFxxfsKVnNY/nJFh/m4LxGjveKoWhVurHDw+d
s+lRnhnpG7fnwF2OqOmFezPm4sphnHUMl3rYJajLdR+7oNktvx92OJIhJ5tY3krC9gApTsIcgOrp
lOUCezLjiyEh8ui2KcY1pqFcFOMbtdRwd+2HtKRWzfji6b3KeFF5M1nB33SzOulojTJNUhsqlI7B
FVr1mEFXdqmmLpFqorlAu4Zj+XDoQ8lZ+z1G6qYRlDDwrtHjvreA3W8XBe/po9a0ObcD8n7LkOOX
7MQoct9g/GtsME767xWt/YKcQF1O4asJmFdVOnv1fcqWj0vPTQkdARvhWh/KrOWhDtJJqLnQ8lhs
1QPJI/R6eWkJG1QjBQuc5vCYzhQDi+leX3AcfdN1td9vv4ICvNiddfozJ4xHDBpCbgB2aHzqinyP
5DDVxBkvP6ZHzj6srYCqhULL5juNuKGm8Dh6P1zxWN6HZELQ7CY3+8WsXZFS03s7QJ1mRzBj3ksD
PGqjDB+pVaDbbphj1pBv3hNb9lzEWyc/kaAJRTUqIz6OPQe7fu8JIJ0WExRlA8ZzdT1RpO6AT/l0
PzZolKJIr00DYZm94m3C5K1ZbRGwf0b5cNFhtLlC4rwSvaTavTLtN5yupDJjpOjes4V3Ga3v9pUm
oKxGpqJtH+CchHEP7oxBcT/OLcXSF71zEcUooeoiHfEMuIebNUtD69ERgRdncYW1vgbTIFD+xvVJ
f1h5hLMyOM0+ApxYJy/B1n22dbaRS7blGYGLrDvr80IBUFyF6C03wKx0ylfndIFmAw0HiiL/sXyH
l530pRPKkGd7zQWLv8U0DZkJyHOUJCxlt5wJrg5o3E9de5lgxSqBnmEF6JBnrE6l+y4lUofe5Fse
d8nQvkIjlL9+wz1A777QqMAbbLekhkm7FTiix08lLjqzcmun7poHLTzHdrUzy0by2khw5v1snwFZ
B4A670JpYp7txpNSiEixg6SJH8CTUi7Ho8bR0I6grYHOdQTTjbkLjnI14Bq8/eR6jn0/xyGKbmr1
GdbND6XVAMtSEwkWvUx/JQp4ldb5K8O/RoHOefo1GXeD4mL07+1oS7AzExeeoIc81jDdp67JKlkX
FQK6bF7jH0B18Yv+rYPzB1XdKDnfYm+Dl021Q64EEIsMlLovZjqYeqA3Q/nOZJyarV6fvCaMxXba
EMrIJ5oFspA5xb3dLn0MBSOizJAFnic8EXi7rvTs4MV1eie85k1CYuVtMM0N86STPDVCBiwIrRXW
27/aHov5v0TSyLgyZ2QzQY4BiwS5jviaLJ3TR7Tz2rKV/dxiDx5i5PwidjqvSmB8Oq9zAcd1/Nmd
JKQOmnA/PpMvPw6HcOW0kBVti7YmVXRplVmd33MH/EwsOQtVKxUgQSSRhaWCFEdHy0bfLjPWk3T2
S0rwCfdAhT1TjGI/Zw6qUxcz3ZcLbPYP2x95er/GbBDG+N3E7Bo7l4dFQ7+wNQwXWdTNaVijZ7JV
pp8pOg+YAJcc5CZE/4W19M4fivy6VkvsGwSiEiXbN4IzX29L51WB1O7bJrgXfvtVqQ22kv0+VBp4
Hk72ZgjnU31y/zX9QqpDZ0Aq2ccXK1bvtEMQ/7XC9iq6heAMJgjXLSShZ1nlCrz4R7JnCNcwrzNi
lBIB6LprNvdm9nPZzDRYOfs8F5+i9wJ3v/dJdEMyEgXaPj+rFV0wq+lC9FoRWgJHMUXnSY4zlZnr
88LxUSELTwwfeSkdh7pCMRnMYAc2MvvpjfjMQx6YqLdOSTHXnyOyf04A9cgEOkpn6U8MvWK+i0T5
UN1lh3zYk/6CC4X136DRcA7BX+eKQOOsMMyXSjANnnA/K6Yvh5UNPFxZbig4lO65lef3ZelEItxb
3r6XXNbjkg48lNliQo3ipGx73v6AtSmORtIwjq4eOBxh3CGMncgqKg0CiAISJ8wB7F8xakv83u+b
0y1BAZPX75SvzaJICubhy+GpiAn0PQDAwo5rqKLTh/VosezorbsJu/t3ANjXENcK+KXOy7dfnZdC
vkmqw6vjZHmZjJXio8zZWNlX08v4xsTgO2SnpRmW8Y/hHGJFH6XhmwCjDM1fSW2Qh3GHlK26RylM
SKQCcQfiyj6U8nwZDEkT8kex8opX9mg9DI2TS+nfotpsa8XfxdzuL5uoM24R4EporPlxqbV9hOGr
dMTlvUAUjEB6puiAP6rckSGr6aYlUw9vyslql1oI49OAc+7V2Xh8kxCI/CQgHp0aL+SeonZrES7M
hX+ZSVZXqBFAnM7Nj3TzxsUatb5VSENhEiZHk8yMuRN8wnI3+7XG/vMPq6PgoserLMmKD3psMdw7
G9xeSoN/+2tlWtWZ1i5sNYkYbMn96kBzakGeJ4Cv6PJtKVCiQ74XvFGVzNASQeK5Jho5jZ7Ubot+
E5j+q0S8W6A+Eeo0fRhyKl+wvsUpfiYPgZe0/OEpdHOtoklIRBBHtVazp2r+M9ecQjOpMxXyG3l8
7P/IdJkBm4JmszLYMZO60QHVMQc/pqTlEI+nzjsLGhEES2RIs2AvJIZqnMR1M3pALJVvsfwpJEc4
F3ZFST25bMsjjfYzK2GPyXFrLv/WSA6bdAzElaSpPOcVuw3e5WmSGIzJQvJqCxfHRHUUJnl08fo8
RVkXIZeuhuTjfsgFZjf6dj8lk/W/uwxWhR3NhQV8hwXPqDtpGoh/IxdUHyqwmXfXnQjJAnYMLeRK
Pt37ohPazHRf6vyRfXaK4qez/MWqATLxQi6qB7MvRNoqkYgXm0e3d/JZ1WKOLUnOVn+cUaz/cIC7
HZcE9ayTWGH2k5D+XErowDVCB4R6/mDYN65cc5y8+BNJtqS5O+1EPBY/IojMfvKQQfQywPafa6DA
OKJSAZiCUu2JErEFfkF2Kcb3iW+pDpkKx/pHEDNUeLBtD8n8ITyCSpSPJGyxPRuDvrIs5ySoQ14f
1Ol4tgCYEv+DG8inOYtBuEBhsBMyr7r/w1yJuSK52MPJ/+ZK14Gc6DtSr5TBlbkLIcOAi68Xgl0L
rE5zcCxdTfWlk+66ytDLfRS4w0JOJ5aOasRWORQ6mXcTV5iFcQ4sCl1jRB9jh0yTXt8D9/4XL+Pb
t/123thh02YQCZn0nUk4jmTrnt2VeCwrJiKyy05c2MKt5UumHYg6EsZ3GEf8lZTSQkCbzkgpHWys
KPAcyLqqgcILR+r/p+kg+f/A7g5qMHdVnSLqjZy0iDH0XPaA4d6QZy7kTm7/o3T3JzE0WZMqGpKn
L2uAdY7FpJ7o6K4Ht/JsoUVy5S8zbhb0TcKR1DRIt5SB/mrQ4K6Vl0TRSj0G4i+SdbueUxYDd8El
/LaksF2/NbENHzoBsxdO5FbUBlU/N4Jz23jw5WNNJ8I/5qDF42pUGe0demOfK6+sV9P1lVY7rjMe
UdGG0sMS2vfyokl3ih9UMLm3zhd5NGsTRlSlmHhPtsuJQ/LMOgdQkFjNvFrDLF+6wieqOUyo37sK
DAf4EUVaAVJiyJHbzr+NMjlwMJgNJPYf9Nd2nVD63GIrx2REOQIMKPSPOtIc9y5vWPby06wCxdd6
bn28s7yrI5KlLIfQpE3fFG0naJGgwiDb6P67FwNUdZftGrdj90ned7c+9Nu3XRQnRoEmupr/Zm3I
abYdiJBtcpnaEWVl0M1ch8p6IupIQQ5lckBvUpvFUBVkOsKAp6lwkNvsGGOBx82mUos7W4bO06Y/
6hGgXFqpnk4BzUIpVTzRwif1TrUX6+G4MVlxAJ7WjKsOIZOlpt6oHDPhu0Lkh8OazzNpp3N/NtGP
bsCXoBaw4pS0xi6cLUpWbr7hTSoNrsApyW2lvdnIll1ohyGG7yFbslinelMMfz7W88HD9RCfrOAS
ddFHy/nJL6wN3GmelxmROnRGC8GfrCqoiPO/J+Gw44QkaFeo/WwiMJbtkvEcMBZLuq5iDuucoj/B
azkSvCcv8k/K5sjgjotOlcMviHuM3oTPPi4XmmZmKR23jF5K8lhemvzTeCucRrORvuYIl4yuVwAR
XWN5DsfH+ZYxCxJurFF1Ttv8Fm0uqhtr/1nX5AVo+gyOvDG0hwJxcH8Da/ssdiqDWvfIPfKCIBci
6uYXcr+/yFsBbTLvlKNn6Jn8LpB5enM1eHsKVOJGbnBzpN878P/ucNEvggGzGFX60QrVX8GgXSa+
Lq2S4dwphJ9ZaF3TIx8Ev8RXjYCd6fDNj44EhDW2Dhi+9IS/4N7n5vbB817acGPZ6fax+aPQo8xA
PpL0PafVItnmqyzZMQdGaAvVGOIyeGluYz/LmJLwnSSCjekTsd4H2Wj4PRdF96ySqShTZqb9ZI2v
oDPKHGOUHsvnPqi/cycPnYOHxkmecMtL4rBCcwlccV4hQFHQqapadDP1RQ20jf42hnUoHoqqxjfJ
ioz7hIZF8n6koJOmDVA9pZSDlBP67GrAqGB3OQ8nsy9/OA6P6imMwl3X7L1up4W9GSgqph8kFbbt
VirLNVcoZKzhqJplP3YwdExEVYyNq9XDwd9JI0G/KtqxFlMxegKHagdiQasFsUnd0ZErY7uAH7lM
fvAc0ov7hXAhEYyl+TErIikOgvokU/HX9+Xip2wxo+27TCvuhd8f6ljly2T8C1yTLogTkY0jOApj
ySKV0nn8qT3ok+/03DdlvaBSrBd+RZoxNBxMQ/p01pnOGFpvBWuCe3mn3vYvTqNaUgILLoAU/2UL
McTBes7bDe0etiL59OAGp13g4OTj0AUOaK3Gok7/+NRnGxp9XGZ0yhKFkIohq7FGE/8p1oaBzfG5
wt9baeD8GPubmb9hxQ4c2zUf82SauvcyoIzDHOKj/HSO4aV3DnJWcTpkr/Qc1pbKUG1elqAwuq2s
AtNjQW9K/SUPnRWz5csJPZVaHtABeYBO4czLGpQkt50dGhMJHC4LFvmQHkcZKJjkscaWd6a+tAf5
8M6WNP6y6G5Rr7buzZaetyMPNsAIHHvy8+YtXc3QEp6XCyNFg6KK4wnRgiczjVJsoe9l8F3pNdRR
N7Njegt+V4SRuH5p6eRhXcKhViyftnD6FMoXi0JVJ2jqR5EoUUapCe/z4amuj9E7tUXgozCQPh00
mBj271CAIkPnS+qYR7+M796DYpw/mZLnweLi4qS7G1i6oKpfndu486Sp9NrqVue+zfVF+lP7jqj+
YE6mBpsjR9K5Fn0mp2vkwj5fe1hyheyL/jPiCa/h3WfGYKNEr20UFXufNvoI+NDHy6l+/vOYatbB
1bh6uWPlS+Fxymn5PMycOL7d1tjA8Pp3JffqbODO4vqb2mAX6I3YZJEhkmbr1hlovwwQiC7cPCVI
YvnXiUo0L1PoPnC8r1JmXigXy20w1dY7/b9C4kayMW0cfloA+tDrraHNLxTbhgutXg3raO6bfl/8
yeYg946OdEnbsef3hpsRLIevSnIx3KN2H7bqdQiztAGB7uBwCuOygPSnLQNw4LdJc8bA7mpy4ZvP
6SZuWmfDz8KyrKKBrxelYnvDKkFaSET87bYXHiTTOpodQC9R1hkNADKjsJ9BZNxVUFNmAt+ELHhB
K+Tl8X3W0h1FFVbW8VpKDHusynyWKNG6J4bwHyGxrIvPx7WIdYPgGww1uhbaHRQbE0N4sF2/jQKP
7KqfGkEVSTT+qvHmKswWkohz1Rs95VtrYktBLqV1SZpsdCJIfCgkMeSpjV3G/xf+HZXmWOMHH/qa
b8DFJm5R+sKC+kTv5HK0AYWvKRibrnSpa5zF/bk+mqqH4OSDEgDbfsoWNDNZT/GFEuDg26q8CtFi
VfkBrIZq2AR+vH4bKbMxSwNhoYAjGqwXjC81eG1MMNw1NsHmjt84StfkSVbMqVxPR/Se9T6FJ5Y8
Xk/f0ph6FhxNTinMoKjBDQrQZiKz2izwXzBBrFSy1AEra879AY/a+Z+J4qmn7UlvRHbv9lCqScmD
d55EVKLCfN2rs4/pu3IXB5R7A3R2I1JHcENaHk3vDepBiadNkI6WjCMO8c+lc4YsFEgetrJgqOFL
K5G/lWnW281joeN8kb1QQxLlPUcB3draZghXmw==
`protect end_protected




`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BnodqyFl3Jbpp2KgMyJuM2OCn2YGP5F2npuvYqlGXHDr8HrGajiFtP2B0FmojgyGA1opckWm0pFk
Sgov35jO4Q==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fF53X+IZ4lYG1k2atmCt7+4+pDiHZhx05zMzyvHAO6WJRF25pevNJc9Eo4ozuy0PRr8NHY8MDqyo
C8gPnutWqb6Auzp7Kvy9EZnVnmu36ceptW6463FM9Jgq0LCEtVNtI2xbqd72UdYtsvWmXhFHxcuJ
CykLvw5LTz7pfVjPdfc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pqfkmBE1VLyI90TMQ632dYOafqVwGNxO7obezGgCAa2MsN4JgXptLMwxR28EjgPxWLTH+11rDnmR
rMN5ApLbO7z5vgxw8yIW5jvVzvzShCtHi24+FontT+2IJMtuZN6dq9vrZ8qjCo9uX3S038oDuUpc
HhLCq6XWrAnT9BgtPAYh3TkQEODM3d22sg8MFnhYNetbpz3sdlVgDOHCgEOOW/rK8Gzba+ZqhQMc
tHvpoyQPgaeWJjrEiTQO+hOvWJqEjEkkqcMthMjxqnu2tR2rCL2O/3DObpL8RSUVQyekDGvA3p92
HVmxH7Yxqt2qY0+JAwj5+pZCxOYUscEgmVJBsg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hdLJlDvMWBMFhcm34e17WvdE6Fvr5iVwqmSV472vyX8fBVhUCF11F/WqYeHMMhImgzihtZRu3dY6
30ZMnV/A/hBBfLfWF/EAWhvsk6DdddqxhrfMP0ytvK8Lbw/iWf0EmEQS9FWT0BA0beTqvjzan9XS
8rVo8B9ft9Bdk/Y98FlNML0rD3Qd1rR79w9gNTMof3nSVSKfDWcGH6pYmnVO+IFLU5pizxJCPPKt
StOeWjb6UQ7Cljp56cXgdX0FTNrLeEkEsIcXA9jvKeUoY0/9xEz/7j/VXLpLnc0VpEqn7XJwZvLX
7Pw3W5MTW7w/oR4QVHlxKu0+I6DGgn+vI+YFvA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vwR11XBXNoXXRZrk1qoqgWGQJjd4RMSAKh2Wu7NLlUErPEvrlv557zVUd/blhhL/6TK8vFt+wR8r
UIFb7sydRYOxq+I2Ru07npwIZsnpbhOaEZBmgLWAkmANDZQS8MGQSWXFf3UsKQhsnpOMGU3wUF6e
Z2SA6OMe2fTtHOJYXoGax4teu/Q8Qi5NS7cAoQVLuWZkP6ZNu5pQjTQDqhBz7LiXu2HghBGRsdNo
Y+cSw6ZgNyL8qswmpS/0/qI3zhtsC0vXytJw3Uz1Cz7AMj/xrk1wcHq8n6gp7sfJ5AhM8KJa2+BR
L3IYh/Jy0d854jYSF3LC9LvvgFfqBV07rKm5yw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kY59hDfRjDFMT+S9blS7LjNpEVZoTf2MVOpjm9NxSxBL6su1G47llonz+N1BxkHdpinNbuGaFw5n
IkTRqmxSB/TM+VHDcS3XKhqjkI4/R7VBX8TcvzJ71Rc4slnsVcbr3OwKRNx41f73IUgGcofU79fa
yhbMPQfsgZ044+/fOyc=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fczWmPU2/9l5BVashWvpYijZACkjqZoirngpfBUA8cmVm08bwu+NScJTnAPlLYsUIwBFEgHfnQre
3no0D4oNW3WGDieB8z3zZdytFJPsqaq7/5Xy/FqnE/YD77wAUiiJQfleM/4ZpOtgZwnPcWoGL2W0
M2ZrVnmAUbCegoTbL9GY+js4WtfKL+hIufIYVWnxWSfvGhXNNJgX+2LrwD89m590y7Qwu0b6hTs7
C3hMSPPrU8yQIHHPeAdvXkLHVIsLq+Q96TXfWhUArKCgYuZTvovLWfxt2x4jshD23FlLEpheeqcq
RAoNdz23cUvKUCLIKnBFWXNSfVrXanXc9IrIGA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 121856)
`protect data_block
WOj6oVwJ1rJn3WtAYbla9qgBtklXC2DuwUWrGTCOBWqNYKaa9Qmc1hW9oTPMKdaVnFTPixuImGj7
yZHnl/JOQw8OGpXssE5tACUAd0hGbhebmOXSLt9drOR0Hy+RYZTg3kOoEJM/6OFhFMW9oKrLhkCe
Aa/yv/b9/9veEQFgmdtn+qOsrrK5jAsBuzqNXz+c0v3/EnkfX3UPLdUL+ME+jQB6IhR3S8H70r9D
57qka2cVa3d0doBehz0KpKDifRGW7FEaBzngVoWNkvc++QY77vWnZWtViGYWYB10ywU9kXZ9Dqal
rXvirM+GSq8nT1FZF4R3RRDrZtElvQzleAcsvtn/AYnJRMeRizwV7ZuAudMrYUa8Le8/z1ba+enn
DK3uJcgnN7PMMD/OqeWO99wb7/x/Ny+Kg0Pxri98NqM0EqCCQNqjCoo1wrBGLsAqgYxfc2kGJmlk
hy4CYo9InV2OVLsGMHCVdWVr6HWyfYX8LnezBpThN9hO38u4vy490+hTl8daVMyHa10pqh7kXSMX
RlIjUsh5VIUR8nNR8qjvnTw2klrfSTtImYiEcoGSij4GmCwTxvL7l7DrXYfI2naT+2elobYRSOkC
ehAWoeEJ9tjy8vizeHNJUXb/d+yCe8K5ONtGFRZcb1MZZar77KqJZY0OeWOXpE5ijn1rKz+tx1ix
DA5hUXLdK1qWNgCC/F07u3WThqa3iNMQ/Bcneq5lYxiTj9n37P+4Jxyc7WIap7xhwUlXUQHduFOh
kTA06C1KP0An3A/xyIU2/iI0/wYEKsELJnXT9HJHwVdJFIyW+ug+eZs5MR179QaqeDfL0n4BQ5fV
dVsxEYIhWTzUSau8SWAdqCY3ji+qofwBUqd8x8Eb9NR80qSRg+/OVQshVJdYR3Bg2d8GgDcZG6Os
DgfdQhJnf8P/gnnBlfe8JeGgdeF3DvTK7CEpxNPSQjyKIq3okLOxMZAWNvIZK7JNbKgrceGq5PRZ
MMdlhyJxf/A3TckB9BGTWstxYjiG5bz1+ud+3Z9SrSB+DVmwHpCkpE6Fdy6BW8L4UZFYzjMo/qpu
eE7W7yhZ24yA0EeBvG0JIlu6cTPrhiaXeHHKFJY90l7O0Nnmvxllj3fvlS6nDCz6Ks2upr/innn4
tPHR0Bdq42nmlXpDau+Sq8ANvYtEiXDPZWp4R3C9vXEtIhVYdt3xnMpx2s8KYZSmK7fwSIwkFM3y
d79HtoHciIJKkHwqAyXnAtV9ym2E+NvZRXBI+8LHUVLdLKdN7HqdC6POk4xR+3IL1d4WKteGkFQM
h8UfSWcOdvDd8EHcPXsS2k8o328dI9wR5FbV6HTejPHqvWvQhwiDaxFMD6ruXTWVrwx5imDVXsoL
LMUKEOrgXEb9r4bXby3JsiarOvVpyZycx5QpYuWE3MjQiGPdz07jQSlCSiK9GJ1D8bmSDTxK4oi3
BVildVek5zns3BCaYLoNHbj8yCtLRYtHJk2WhcA6zYiu6wHPZ6FGDMRNXkyUr/gYPkC5sehI092J
eEiA2YKkYram8GiRyX0M8K7UCTLs564tiDiOzxvbS3j/UAAht37H8WQ2uiU88Lfgq5gYXv3qtP3t
0rHiFxJZgHzqqiCtLX0xSJTYJnpSEQCoNpPL6PMSbH6KzrfmiLnPcrU7eelKtKv7iXVpf34tHySf
yIhh6byfAW9ZDcN3pTC9ylXR04CDWgXDRbUw4R5M/LiUNtn7qrKck7K06cdwby0NSTUsCOGX8Zb3
oPpRqKg6CunPos9pZPXZo5EMDF6L49KOxhj94coSgm3kKBOXDbUjnYB43ROWrhZb0NRhQ4SDVQHF
Ae3MgU4i8rVfxsE3aQ4OhoW6wdEX9bamnycfM15gBkv8B29wMrQC6fQpub9aoTSIbKU5v+uOwZqz
WoYMNWJ8LQBpkQEvImZprguuMehrLETS60RWDS517avD+/DyoDNIOKUwhQtkvebfjXW1uBr2dBqi
qSWmwAmZSuUWCDz7umcuvyo0dKU86ylIfVGa5Ow2Oo7A8Q0aBeurluTv6pF3tNsLAJ8QyJU63IVp
GwcFGhGqKQNu8RbhRoFZcZxgmjU5cSAH3r4gKOgeA/syz6zQ125KnHBASLB/u0tQ3ziCBDhLLM4Y
40ccHGuZEdSFk+1DC+Z5D0ObYRaZJLfh3ThjpdbzT0n2PyujbHAbtCY21NVFpJTeSis90f/43Aon
SvCk+KRWOD8+hut/H5RgnKw1c6ph4w37DVWrpoobdpiuurwoXAIT/yt55wMdr1FV0x1NPDab1niD
TnEbc1Jf1ATF07srdwOIwj7kQVXqpB9Ua9/9wn6Ca6JNcvyCtg59anhIv2IjzZA/mG9B+1fz7/FX
/M2Nd2S8OODiuWr3Q1aifdgPhe3vSUqrS/lDaNwV+auTNdFGyk2OqGgxZoK+9ybxurS05IPsUAmP
0c7BrtuvpTuphlyz2U94oPBiW2XugTvnp0V/RqCQ2L9yZAaQHB6IHdimJz4RvLqcIZtimo+B7TyY
y/brYMsFiY2WqZJMHHLa5ti5M9U8yAw1khXZoUp4SwXvB8jX0u9vaaxorck2qWQkdI+c5wZcPNqo
CeA0HAAQQ8IBVRXsHeZgyLpspnglqQgYwTyRLhfJ5+296svUa+81i2nxFG0oSBueIPZwzpNH24QP
I5oMZHUhLyJP9Tl4VEnMpOBZYYFxzHJJR9gdFKypuP4SazaATVhYM7u1KumcuA74FljpWkmApugo
oCTu/dnhQ7UAE9nutRIQk/AyjmaUSdOutU6Wny5XkHEvLV8mDbO4jqFYV7TVF7uh38b947MTvOTZ
m6ycmnNK9fFAh/Indz0lL9RFJ1IVnzZbyd7+5UbPeSTm4/ISbMRjORaP/5LTHB5Os0sUhBP3elE7
1zGQlZrBVf9m4iDwB03SRmeb2oymrjjF9P+SJGF2AgzRGXjjSkA/zHgRzU4iskMVgfbccPZFqlZz
JiXPKgwj33IkvRqMldIOmMyps7WRev44gRIGbgWsH2n+P0meRibKyuWhwQ1I6vy2lzQaGex8+lrC
h4Y16d9+e6UlmpScr+b1tJbIx2eikMMdAuWcWeV1TlX4FuYvm8+jOmSqGpn1+BA4k3TItCfJmj5J
2wW5ONG5QtnK3msYsXRh7kFp4KrDLppTFNsiYDJ2OFmfH21oJZeO3Y6Oa60UEgWhJXhXjd5fKtbg
NWd/XzKantgIbSKRzJcBuY+5sv4798vMzfPGFONb0d9Fb0Omh5mQ7BeBO+GlVWs+XSDmIjwUsDz4
blHQz3ZtRAL23MnbCIN1SURwhHVUlFzz4PnrJ1d8xoGdO+Q52Kofi+IMerv6k0cCasESQGrjmN9l
mQFV02lsUXltq3yIW/pWAfLx8hCjqm+fv2P/L72HTekt6KEhuz/cz1lDF9NGexXJ1EK2Sypevk2o
sf7I1Vjif3LDky+enf/+VEF49bCwKduXeXQVP9YJNELZixp5Pu8b0GN9g2hq3kb03Si/ZnGpl+7R
SjrvCbKoYP1/jAPVNfTYUvi74F4EXmNeMqTQ6pzTnoMMWD7VAbU4Db45/17FkkTWx/QCINtFohDJ
GLybo5hjFp8IgH6dZiOcLR3GY3H+HZm70/F4yyTgTQzuPMmSKKzaHztnzgCbeGKR23qK7e2/jLGD
MIC5andwi2TQbWYX9w3Cb74df5dyMaPLZnCDmUvBMPagEEogB6vuIm7Vf7Irubh00Hcd/H43zwwn
bkZh+f+Q6hCs0yCqHr0vm3V6yUvYWwm14LKuC0n+LP3rFSpf+iNPSKAFkuQt2f80Q947ZC7AIejv
/yxYaCADA77XrtlqaCk6iEeMjLCC2PW03hON1mj91cVf8G3OgJLxzTSbGZfnr0LqudJzMOjhjjs5
j9h687jf6NJoyRPmtb2XFTzLQ+zwxFqY6edodgHhw3S8FzeqrljJwMyemeIw79uYJJFM+8k6odFC
uy7pNgz1ZeEvIHJ9DGpFZqBF64pBv2HqKiiMregnhB0bUJGL7I06mHCWhCgmhOmCD3AORd3+TGhN
Il2qgORyA4AVgJZ8QA7EOf/xiQqOo62bKD+K5+iLFyUuq0C63/G5PD5DiR8w9lTful4KZiD9T6k9
YRPis1ECjIKa+CGGhL23C6VxqKXsgZmxQohVD4Aaxq3i4DImwyz7MG0CW0Wqo9w3Ouq34+vzYXl5
oRyIQJ4CkniLr2qofnbz4XFwKskCmx/IsU6MhWB8Ib5G+ZrvOiLdICDd63Xe/o0lIMJpxIdcOonw
rE+OtDfL9ZE2dgufkJ4QzfLFHMtzLPQREYkftQv91lPi0nnRmSip2PQr7gaKFiGhfCaiMMrOkfM3
7opMAZYHYh/ovTz9wfRO5vL9L1i3Mtbk8xPvQQYtrUD0EfEuQ1+P1p+w1ZDz8iUZQnbJG6HaOhYn
29GvLeFYUH0kePQozPvjt8uS1v26uDh0zLwYIHCA/0ROJsrq/7n0+h7W6Wr5+4apLSDoALEB8gj5
XcN2tdzv6gbvWZolrK78hRW24KkzWN1cjlsh9KfwL1liDkvJn/g9495YKAn3o+5lUO14OExCIwik
yqEEIp9e+GGIXDj3S8TXO9hIwSpKn44oE675aVJu+sKJDsRFzmLIyycOUPFg0rTXlc9WgoqH2Z1y
rzM6eRdJG23/CcO2uYE/OCwfR7DgDVA06E9qIRcdGhrc843IO+fX3jeHZq9/JC1ZaYteIKxN3G8e
AJnlOicJcFO/qpS2DKf8kC3OwtNSzRue9uNZjoD76tkthepLQqNey6vPrgx1b9mtjrzGFmf8Xd15
qjETlh1msHWBljuUrbBGYST8BVwTcaL4upRgn3x+iM2g6jxVew85yFCaAb5lhIY7l50kbHm9xg+C
9PTvYugRhXTyiIa9jyRn/rU8CmPTCe6OklYgRVhEE+tPhCgs5iYv9/HR+rhB9yGGUSck6RERysnG
cWSI/q5MrtzXxZ5zJ8McRcL5USCpMD31WW9XWAy74YUyQ6eYH3BeslgbbqUtA6zAWzK+L0Ema85R
QtTRE2nnUk/ZzI4pO3Vn6yuVCJuO6vI4baW5ztCMhNKgb++iAXwpv//SOiHk+5rAscrNBtf/6ieG
O55pFd8KffDmBeK/JR15H5xQ1fP6EVv+QYq25QPqW8X8fQwxlY1tXhP25NPY2+mUiHlrlQe5r3PM
ZsyEmDfqXEzeELsrXsfcW3ol7EOkjW0nToQz7+hAL7EqDISqqLDIcPyAMmiX6EmmubXkxiuvalYn
mAcYJYfAw7k3tk+MVlgf30uz1TNCwbIiEMpd8X8Hq9CgEEUR+hLqsya0ALlneyi3QH9HmLJcxc2E
BcyklII5Ad57HqXPkiJzddt/YO5bJ56Bnz+bt4ikGZgJF2d2A56vtSmfMXoQIb9sZLyuWZgpyuqb
PqGZDD7jQ13iIS6QkMEGCrIDkn2rWjY7lNyDJMELgnj6hf3b7ubCmkHFXVNDhqJ0HrrL7URaZIte
9n20FU+CmRLF9CtL9PxghbR76ScgenGLQRGbZWYB4W4XUmnEfXsVhrDKKXRqKTSPOEp6Sa//1lml
YkX6TEc+rWusPMBNzdhvXQv4uYh1OvKycW5rg9IicZYZiigtfQ1msxD/pHTEg1vDs1Js3vpXP4tJ
rEX4g/0yfgWDTlFtY8GOjbCzNqgSz5x1UQEl6B0jaVAYsrZf4qa20I5Q3/sJ1PxtDdzaRKdZEtPk
Y2DC+NdQwXL9IcDnBArI+O7bLRuN4cTZuk38TwuQRNVCZYLn0YOPCV2sDRlg4KKADXTzcU55LHYs
2XuKhDB1HNQ4qr7myuuuw8en6I+aXlRSvPEjJ6SOpj3AZZYSJplMMdq6PNxcSQ0cwGeYQpKgHvm1
SKO6gRa1lms+GgZ/C1RGW/WtwXOCNsV3HnrCkIisGzQeVMmgMOiREl+Xiezao+8/AgoWvAQXbTaN
Kbv9ibToSRHdfxUqEJdG3YzBcvpW2lRRZ8CdTgZdtCBDI1lLbavpnOnnb5oE970cbIRhCBgewJ1N
SimEMANZwHZGj0VGdVsc5K4HHDGuaocu2ChbEJo1uTQ6vrn3dfIAmKyXTgRLg8XnubHiQAiDHVsu
k9/777GzbzVavgQD72oTe5BA+AZLNo2EjVhJBMdI123+a39maJfzcvCg+gzhcp+zeh3yShXwZX0q
XPcEpf7gMO2hhAKk0t54ZozYN4YYJEyoEMUOToSrEgnfDH0N1nUO45A+kdZmC7Artbly1f3m/CYQ
WWXo97S+swNE2Cd5AK9WMUqrh7gHLXHckkHUVAkN4cy9oSUi8vqWY8ttAawzwL81cFXIEG62uQY2
j8VlDATKqcvfBvQYSS4vG2+WIGpg8e5ZKrxjNnQur7a8HBu2lBJDY+wL1f0wgYmIm3HYm62GAYCX
rENcPKoRufJ1CsrUEhWBWNUE2vYHDfsm28ZPdHX0m4zlLGKvx3h8oJ2TtaFdlm1r3ZkNnN7cxlij
WcfOiuVY5dWYXGZ8E7IT28AEkm+w4A5CSnaI0kVx6233UE9TIYcwaG3UKw2ZZhabjMo6TEjL7bYp
5s98bHJRDzw7ygZjpT8Nu7VkcyXzwwKD9Ujjuo6vZueaslIdynHzYu4bGXJlKOSwNhaOr4AjFnA/
6QnM6zq1HOdZbmeho0GiFnIs3U8Y+2ax6Qvjvwl+UI8PR8flSQjzEDGA6Ydkxz7btljfFUHaVd4u
swgvwY80QBCs4DSttOhPeZeBDR+8ZQPkxNt71DRpL918xmYW+//iNkKgovrBfzDRLF6j1cUCDgWD
LMZSFUP21ekQPPmnJrHsHJGqGv3wCFYgBU8Yk5RswhvnDWXdByE7u8i7ZNgq72k7ToG/yAnQzbuw
qIYu4goC6Q26ps4b4wOW0NaFbt43cTHExXAq31xBAJhjLKQlVQFRDP4qhv4NP/srYSrjKrhi2T/9
kgdSOqSpjS8c8EmbbRv8uNiO5etBfoiTSx0oVLQNbyZ16fTDp+GU2CxDdEo1wIAOfwWUIpIo9JIj
3befwFlrPFw25pEWRaR3wFadwtzPivgd/FF2ohSWDsbpqbDJP4zdalT8Jk00IvALl/tzbJdhMBsC
qR/ds8lXJDuzS7aDqtyD7CXuEr7Ihgu8n3K+0R2ove/UerTSsEhkIHAOssKFnnUwHbHglyqt+0qe
v1uxg953XEs8AAjc3rAbvP1c2XI6Hv6YqcrVD7zD+TND48EjjdvGPGy9G5O6FyGLtA4UY1JIFfEC
qTwmlSjv7rpdxWe4c6OdZj+d5WMkredCPO3JW5slzqPH3lblWSb0BgbeifSxK4pVGLpaR2xJ+fdU
INYt2ggHNyHVPvB5lc8QtTxh38gcpOrerFfYdUgiXuDztTD7idL5sme/UCokK7hEDog7ZDHARMeP
OP4UBya63qasPP8TS93UkMwuhfoTjLGKWh+ZoL43G8zVyPoMNqXJ7r3OOdcqJacW3aHE4XjEiK5o
bJp/77rP2px4q8QJ41bGxXBxXViMlbiZJAkU91o3TzrdGsEfU/b6yXVZjK3X5mGdPeCSWOElrEQT
7Kucgn7M0wkHjfMl16gXvpE3+OYfBZHsI5JRj2my7KwPtsRU2upQo7M+Pajof9fMI5pvD4YcIE+h
3BJEDc6MF6q0FjZ30msEWQICO0hFKHM+ZRdFNTiWIeiVH2eIHU49SpGBhVUX/P85JCivY15ETJLR
CJGy7fUpMK1CZMdSXzaaAFkhWzhFbYuH4QvuLNzibqHygflslcDvqHz5p4DI2RXxGb9gVkn505r3
sthQm/1HeBsJ9iXuNSqq1Nr62N382DNqFA8nkjhaRRwKAR/EHNaoy9FNR58cgAiubycgZeGlBlXS
ndzYueKey/lFjgqjdeLVM2D0tljxeSeJ6vx2YxOPuL6UGUP0UC/Ev6gV1hL55A2K3BxZnNZq0XF8
LLDesvDPhijN/wnQzm+ZmmB7npDINg3o50vKcZBIafdPlNOm690+6OSAuS2WhkdBacugQkgEMvnh
A4frUZdIjWM9YMC7KXIVaebR9zOWBGqgi/53mYrHWgZSS4DmyxmiQUYuSmMbyJwOez6yLmXFegdy
BBc4746+obfdJ2auaWk3NH/dmry/oOotWrDAV1QvRd4cu+qrRnvNCBsaUV7luUGfUjNDENhMs25s
tEt3czQJQYwbaV9plE8Px8V/g0rmAqUf0jM8jkudZF9nHx0vcrG3tpGH0e7zdlJpZK25zU8x2Lc6
FYfdX/I3nILSlvBKy4vmMMWpE/alrAt8x/T6l4Mj1jj+9snP3sDKbCEzwzOMrcyAw2p3l35DjMwo
hsaCI3EH8Qwwu8leYrQ+WgbBYsazsywYrjMRgOPIqkzEov5i/ZNOUILsWqsIK/ftSvnY6GUqhmQo
e/4IjKXGfHFeVpgHP4p1Y+yDh3AxOhdO2QGsDKt+rD3KO6jVX7S83Y1w4sBK4WawybHuE2FDHPuj
xbfMPWAD+wlR8Ok7U+AYaJV92hsW1U9JRtPI474f+nC3o30darjdjR8duKD3LumPe6BYGlzLnz+0
oAjYXk/eQzb5veAU9WNKBydWyPU5IZ9jFTVQv2EO2ji2a3F3Ex3k9NkpJfevLhyO5dVy0aWlf7Vy
GyWAyBDH1YD7gVeBSFQAE9kxe9IExDXbmYlvyjQKFkLgbCIb97gCySQWwni4iBzCm9NNsOD+RosO
g8fgruyYLTuqbQLDaAdNLIx+k2nFzcnaBMYJqQ3Pd4iULuAW0q8maTlwAtwojqfzK6ngi/PH/7/d
ye4I3N86GcVlHXjcY1A0FCH13TzJ7i3njjSRH+6bXWDYVxhc+kmT5rNL7X3Yl1v9SQlmZBrk1Wa/
WpYW3RTtVbV0UmEQjwB6GSKuclT9+NtWadNeCTPis0J2Xe6JhdCda/Ssj9/TEwlDdvt5hIM1EG1m
QdmxEYlLKheloPHCX80nDh/TmS/vaqth8tTfla/J7130zh36u27e3K/eOJWanCZZ4XDZ1by/YU7/
xwpleTtuunuamJSfDK1ETBfg2IeAas7AgvuLtmLwqTRrb6esxCiamj4Hc3mVtIITbZlD8Q6rfGxp
Q5Y06w5O96JQqQRHVYy1aOe2zcvQ0UrHwSDR2+lnEbaOEqm2K9rT+VfTxs5p5f2yEKYa7enLSK24
WSj6eGYPmtyou87HeS4yd2+VHw7ObgW1laiQNjqbgmQFjEV4LSjJpPsWuTrkrq2k0QmMSQJwVYCK
29RHww97D82U4YV33i19cDKetQ+ZHvpHcuPgJsx33ZiLcRG4st5F81Q7PU51A7StKBdOOY1UVmsp
0jhKXkGLeXI/1TsDL8WkScFUtFch5txVmWd5biXpXvWnOyBplj9sJVQ5DcL1Z0buw46PsU8+834X
L5A7ZeNeKQecvKyzEsLRXb1IYjOCwPI1AEI19GJCadFpr/gAqTDzNTMo+C31Qlj8jxoy8P4WKnV2
otseGPq2mI2vzAQ4GvWtpVYd5GT18OZGbaMz59VekwdcSWugXUkmQO6r+tJXrTMuiguFGuxmlxoR
iMppUN3A+9007ms7CExyU3nTrxOI+ao1IlYfe8AXgs72WmoRSgYwunqXHp280M7d7vciqV6cO96m
KXLffXqTbCAodo2t7kqbLHKFKuatN5QEqaKC/s9FzWQYxYAP0RG/dGxZS8DaItmzEgjQIqLLoFFl
+xXtpFtbUA+aMtr2Gs/sC2Us5+cxJW1LJDgWdG8PZYloMGUz4QZZNV9Za09TBhbE3pf5iRcYeU1b
lN8ol04Wk3HKQB0UmcvP1Oeu8O1bbcxxFKBoxn9dV+MT/au6enaX17TN9mmrSs5GM0Jcoa/8tG6E
G+yw07Ztaj0qhgpzWE46ZgAQE2A6XBmNM0VBnRKXyOdWXB7Djzpmd8fVBfOhJQxunSzUAhFUI5L8
ghjfrm4lqorN43uIZWR1RQER3qWQomd+BkAb0G8GCcGSRLP2osu5ydvmzNeOBzMHMQw/pFRk8ofS
a2nn+i/LV4QM46bnPUlA1SsOgY/Ol2s8jfwNyeeghUjEVe29mHR5e76n983P2TKv856kFWVHjF1T
qYmvJBWw3L2LshFMXh99tX1l4AUuG4EhDKx63tRqEtHhZKr0+qlhW37lnQUpKHnvA8TVFgnBc0qS
AdxP+bCZrWBn4PTQl++ri8ID/egpqeQjq8l1cKY0uNk/WYvDTKasQg/9noxqtIxtijDic1BVemFB
bQImyeyIX3B+gMDp9Sdbb3fPFvyXAx4I1R6McJn7ttfodEchgWrrPr1axlnbEAW6862Z7QSlFO7m
sSvB3tySeyuJwOxJYA6ke5o2XKd2L2czUplDd8YfIV+YkVkUTNyQA0rTMSyILU61gDmkGjDCM4qI
A1H7P78THwkRolZOc+ivoDvv6smEoNn2VSDbum+8IZS0W0KR0kVe+dJSH1q++Gc0Zqt4dknOUFyo
NbPvWh8zGN1pOL7oKd6gQ1C+NyyOfJL22LdeUEx4fJlUn/+8hd3yvhReE/q5x67FzpZjF54uJIFt
oPbumsrletTfqziNFV4/C6WW+x2NtfD12f9L4M//26hCJgNYLyhZcTzhghnPehKRDxqrIpJonM6Z
Odjs1tz5tomq+KFbWkuNX2y+Ip+a11a21nXK56gWBWflgy13KLATlEECxroHK6FEKqj1hy669ftV
Y8k3zkDxMStamzUlr7unH7DA70IApq7kiX2OVAYgNhaPAi0OUGJEscVDzoFNvDOFlCdDvhfOShcW
Uaui8uXUVhWFmRK9v3NRMQhsMjIYHs9Zd8PBiDpMpXLbBmU8mOheB9vbyA4w/x+ArYf751do5bET
YALaX+Uk8nPOXNz8vzdAc8ROOYgK04l3/PbzTOvWqsyjvV+IQQMSCcxF8JAdyLRhDaSbqQ9qQXzF
eA2NWZqxxGXo9DvbQBc/hz/O2cWWFBxt74HZCOkpXP1XBp6+xl4/dREZQmKWCzLJW/pKN1lJw2cG
/70F6yZJ6z2NkR0DJkd4guhQwf6StofHC3rXvv6ZkxpbEapoiSDNMJxee/leREHKedxynJskWIEH
V90chOYcKN2oHLEXFMbbNt4bksij8+6zXnJCU+Y8pbtzW+Dgeeakl69OsLGxGQEIXg6/bBe4KaA9
JLFMIRD+gz8o/oEtVi0KUHxht30jqIh75ztYS05uZDi8j47icbTBPjrJ5xgdMhJeA5GdOraEAZFt
FtBf4ktjMjVpc3gg4g0TRRCSP3+rvLWM312bwkfOKWWV/V8xbxwvBgHF+EYv3hs4GPzV+DH5rAVC
KUZqeXYQyVd9urN+pAXY0R3BzUgu5NyyvHH7K3e4mr8KKwE85y092NHcmRE8nXBVd0PMod0CdsLC
Ql5vSEB6+EtXkH2+6fr7iFsw9/ecZXmbScUEqYo7VJiREd5Vf7Miwp15wTP0Kgh2eAJmDy6Yxxcn
1yV0NGknskQt31/IrSYL3lmupPsqIYU6Mtyep2eR7BlYCE+IceaSiV35zQ8FFODqJbRg7KVVaPE8
Gp35p5sFCLz49LMWg0XuwhpJo9Ka2gI1f3zdmWUsOtlDm3bY5vTCqLRFjL6Z9cyvnhyekUrpqBdH
6lmJUJrzZFKbtsbVcEBi3YVmFKhVVBElD2tLG/pNG3sNFVzrADEQU7eo3rU3V840BO6iah+0IDpM
tKDUIURhARI7o2F3WgTLsnMcCbYqUvwahW1sDxKqAaRFU6uO8Mf9e5U/TYZ1lL5b85LPiXtMI4zW
qDYl9MVYiGCxioLLHyXrot8n21AjLwBWGf9Hfsq73w7JGHRJ2+fuEcyWvs5sMv9M0ShnoCqGzeG4
g03abQQmiiWBSrJ1GPu+5YLNq2RLH6DRBNg1vOp4AgIWMOYeV3dA6RNn6T+0KSH2J6WkjXopdvXW
MOCNgPwAZ8st1Z3FjHRbDjYPhPU/anJufmX2eRpAy5aLL59eL1b4a91srEu8u3q8xwnqRkW/Bm6L
qITj+ZVFeLBXMzAsTDWE8c+GkuOJy+kCfYN14NRBaTRfi0n8ft+uVAdj0f4PXiDoMtwcu5faOU08
vsZviRObdSlqPfobOU0oZQGYIW4ATxWI0UWDJ0PbihGikI9qKmu7o6SbpsmkbcDWolKtx12w7gTS
t+05eP1cdIZsHi3vIiykfunCOoULc6Tj/MbybzRoAwoD467qcVgfqo2P22EhoiTA/Z0hIpR/1QcF
H/JVDerzNhqHNdMBBReb2/l7EoOxa/r7xljj097czES3ug9U+bX5/32qYJ4pwudEfYVvy2tmLYyD
dVpLXGM3lUK/q74p3d5itmTazokHLV1CQxzerH0Z4kbQ9Bexzz1mwfQsd2Id8UD8lCdUeMeanMEf
uTyGIYuR0RMGyDy2MRlgSssmW53sJoUS/Is+A6YA0tzsCHN1QpVCN4xOlP5nSxY9l9pOtsqTdFk+
qzvO1STrQvRWZXVjQiJ3BjFQwi8h+2w4scl3w2NaOIfk4wEcTxFm4ujD1if8cazaI2j1D/7Sjkqz
uy2unMi2SrwaMZgPNqZADqLsWOgAm/jHbMzwXazXgv8OqP/h7iGNLKPJd9FtYU9itVYtaR2sLgkd
ikJy8ONn38ZkzVVVdqR2B3m04Zg22cCifYDBQa0PDtD/CCFN24iFUWhMWIY6zU03kaza0K5TPQ6H
jMm2846qyqg30fi0MSF2YdJIykk8DAwX00mIDeIxggtfKGvZXp0wbbyUirfhxi9Qb6MdyJabP284
9+5zvxZRQFv0bgyAYZss5jMC57jEPoQFTAvRhBmvgzvvR1Rarct/nH47DA0ddyFW9iccM7JhmNj8
ydEyz0cLeCjTfKFwC9Axld24gdcH/b4hEDK2q4JFUKNwOhdELRu+/lKEBWgVvr7wtR+ZyaW2E+jt
MmSWnBBGY/iVvS48WIgxnR10AWAdbBRkh3OhAuQntRGUxeV9+5ixuXfjmZJT0Sd69QVTK1v073AN
e5fS0Z2jeCE9QF0VLgs/6b7NPc22v5KMKCgg8HHe8MBpaHPWVyLfQVqD5z6cieBccbhAayDbmQYg
dJoNawvWHeBpQkI+znqsZLbY/RIozFlw6O2zOlmzWZ6B+H7gRoMTbOH2xl+eeoWayIC8Sbb1dNrc
sMNoikMZwyMSObmhEKHZ0SnpROQY9kdIXk/fxOZvgMeQXcgWBKJGVNYXn0d3VMABdtjRoJ5LV19Q
IUJyxdBzrSMfrF2Q6DhUdI5BDQJk0gu+DrwRvoAKb7wTo7VaIb/hS4KicGu0ui/oKveilkV6iPyK
BgVnljrmqp7JHdg5XHL3LJtS6n0i/Dl5KOWENPEVxMldvYpQ+QAmIC0vq1Jqforvf9pZSaxnibSy
vtgJMMI+1a42CNNtsi/gvQlJ6A/w4ro7YPFzKXOyKExe7+9PiGarRbvC5VtbwJNqkp6VysviuCny
mKy1wzIsGTrQb2m2IDkO4G5bBG/eKBHbUT2uvznSArW0cWEZoj9VcPw2b3i8C28SYRlrucj8Wvii
xX6rEnV0Eq8LpQ8HBIgWv4iopRElas54cFOqXb9LkdgjWpJeXXNTqMDSpypN/xn7jZ4Tjvbi2vas
pFE0PhV5HyrktZyW6DDd/kG7HgthscZDDtsNua8EDHbm9LApHBXKuAYuEraN6NWggex6oky/8cf+
E4coBav1aFLLLUER/srPu5E2UkQupo851uTFMa1DHI+ZvLTtzJcl7uMKX3M1pgA5yMgJ+ihhCjHx
vnHxmIYasQa/0BfM4Jmjz8yqhUQ7JAdzKe6DYMLmUBrAb8qZ6PYyYAWAHa+u5ZrGk2/cfsmvWFOH
G358XPds0MGpzv318TLyYCWuseDMQOQ7JKCUQ4lstj77/4scZpRDCBS68MzfXVHvnhO7KWy6vowb
uCgltQM/hbsALq2nCoXsm2Fe3LUqj4eH93pHecO8ayeYQjELFtyYIcAba97rOEy4gvOZZMEBsf03
JhyWX26ZR59TGPYb85LSTA8200z3wk8zyN/6TgiQVAUAeUUYguAM2HDR2BHv3UHj1xBSYWWMmg2h
14w8HpIGTggz2VTsDLa5NjKv8SPZH7CVSqVfYZ3aImO8XrVCZhwN00atypwqenBzBFP0uzXTbxfl
l7+HLT5JMlwAwY0rJkvr1bg9TZ4DL+2lVqfziy8J9mWmmovwwX25fDnNHPugUR7olSpPB5TX1aEu
10LTSTE2BYXpPEbjVZ8NbiHzClnygQ/FTUnYmozu6cW/GSX/knzOGU1JeVwo/JtoYuU3QP+qDVGD
CXYgvZFV66gh0hWvFsXCCwrYCoNK/nVgb0yB1qag/Ab5+nOF7h6Lxdr6w8LLosHFECGNu2QlmvVH
Z9sQPQaVoHVMmu1o99xU0zR0mGq0RK6zsGBmfpUL8AuVemePexrB9Kt7PUo1Wu8jhRDqCiFZExns
W95SmjZukagWf7fReoMWl9yRmhbHVlkCoBLiAsMKrU57m8/wJ0Q/FL9pIZB6HqvRyFhQGi6K1YcG
L6Au/VXshxpXeJ/0frLbGogKiiKod6LYlQIImf94BC5a0U8Eyi3e+b2eZHCiKnyGTwjhmyntQ2zE
mTkC+0sHN14c1VtQaJpI1tu8reeq0LinLM+xsgNLZF14bfvuFO47p5cXOo1m5YeR3h/d3z8UnAs/
eEBtWMiHcrUSbOpG4h80HgBtpzPOp7ynhKRWzN7BTpx8ZbBm2o9ZHkWp/JEVXJrMAz9ia/vtpZbo
re4BN3xmC0HFltrXrGk7lJ7CJ3iJlFuV0qUvIkCL2SuK6BiEBtlXUBIo8sluLfD3TnWnpWIxoIhQ
93chz3HJhz0ztTNO4297SkB2ozRbQAzwFH3+G+ykzEmzwp9CYGYjfTrvYtRsK5Y+D7dzlfnJ1kIb
bd+pBUqWEbspxJ6SAS4YmmWYQr9abKAaanlKwdfkIAS8ukNbRwjBMXxfAC1gMvCJ2DXYxT0WDW28
FGqB7FnJMz9FQ/AocH6jcE/r3vUth51P1FLxm2G14eZ0C0Dpb27ir2dXFCP/tKLsUGyFiR0mRi6K
a/l/XXwV4v6XReVbZoCAg4qAC90bnDgumso+GSPGGcrPAjYfBstUQHHGVE+njUbLjTDmVKX08UpK
rV50dQulq1OjAYCpfy7xyxpnNHjEXUyWM+/t8autsZakC1hcrYGzT8pFwVuREF5iQHUFLzjLYqZ3
gcmEYriPubYuY0DFiXN7MX2pH9bGBO71bR12K7nzmK2RqThY3oIe1dhv3T962Zg9IB5fXPf0ziXy
jJ2w1JJTblHMUz8H/om8HtGlL9ZnLjcCoAoptyIJZp41aU4kcgXh3jYL9TRmkOjL4P+rcB84vbmq
Rh1MjWb+yS4KzeyMbn6xDsV5f2BOXouicPenSaBhd9KlvufnL6PI1bWRUxoNhl25YmTK5aVAZJNE
P2Fux0Gug4PlFVOuWqPWKSfNdmVW9lqacnzwfWoWSLRd1z3uxilE33xZ56Y9BwT1PlijqaNcfpj3
7QDsDq922TPeUTVbtRkLAcQ2MOmBbEGbChDI7mGTolrkBYTQcZrRFfSsL33G1TiCRn74IrGJUgOE
gSGWyqcarlutwRZ92cjpZQxr9WRd8mwaPcwxoj8Ys0w+ozhJ1AslPW8R1fGo1tcdE69ncq7QA1sU
EtKpYGa9Pr06PdA4L7lZdRXQLgcsKzxSnhMMZe6m23CZMa2XuAe4xvPK6hmKH1yCPleDT6vF0mDv
O9oJKpjRTTQ4FYGOtebziP9eEB7lfPtjwHUbL7ZNcBMskOgbErIZjQO2HfcEt7BgsqEWS04HHMxD
UA2JsG3+fvjR477g7hya/wMxaPSBTtUkrZaafG7Su+uMQwZ9gde2rZ/2mW7sgT+oZ3QNX611YGXV
b0IRxJdK6XZAMnctceJ3KUuw67KbmtrCHnrd5vX8Mtp46qUpxLX9FdOCtrrKyJeAP38LhWZ30ZVL
YS6sdX/dSgQwW1165M/ZfwsZQJEIfWiTIYVgcUsP/RkHRuA4YBD8vQrTva8SycmmhNIWwf1jdVzx
PtlhcNp0hd7aNgFowoZFEyH2nbz/b/qsInwdatNtj7jFnV9O6mOXpcAAF7F//2Jjk/4Fmsj0EdA7
jlaidYuXZZD13wRdPdq8i3aO0OKhTgAFeCgNQduoCVY4FdTFhr05+yy8omkZpSfKCIiv2ksEhGvA
0Oz2xoGWCV7T/fHVmZjR6kfxRaWSeP0vMKMTfcqCfFtsx9AcVWEhG/01PDe7VnJDbpxYPYB44C73
wptPx7AY7jsQwddHLHZxSM3zEDeEHHDmchUM2Q7sJogH78lbsUeZBIC8fjpbxUPO9iXY0OgQ20oB
I2uAflFrwT4FIdzRc7awWNAqCRVFlFxxizvmpKIJrdpfUHML5EP8+iEw/PtwLwlOd9G8lyxgrOsa
nC5ZsSvBPUA4cq12lspx9U4pYEdPkmUMCuifmi8IEpi4KKcg+LazkEWTU/qkWvcFIgxLexhT6wmW
pV2sq26PNmcEAp2RQhmEDULzhlVceTpAqK5/mwni5JC4hV8IYwEi6Pze0T4RHN6+qO1RSD41YOx/
87842l/haQzmjZrj2HB50ok22PhHlFvOxV6fRoNZIO+2dh+GS0czomoAPuXDiMLsMXUsciEsL2R9
bzHlidDDAtUkCLj08GzDrObC6LYtDqV2eNzplsaCK8YJA2bTEKevPVDjrmRBuHWw7pCLNXagpc4t
w2+oPbLHqDghtagCmBaiW7UIOI+ug2V6azbsOUbo0GNA26kOOs1Ra8mMZryEsCX2YNCKRhue8w+R
1JhjPwApX+ONe4Dvk2AeRQ48uWaCUmN4eBUcXt8Ty+/Fi9r8xt29gIpyaE3WTh1Ey/pmxphb/kT7
zn/uqnUkhtZ810teH38JYPBy+073Uk4Z6RUMpZQkxmtbC1t7xicjgeB+0PKwQ8SI9t5a7s841oe2
n35ps2giho+QOAX7KYzJspg10nvEiYmc40cTksEaCJD96zhfZ8HINk3TErj7VgOKTBolXHfbyM+n
PyaC0AwJ1RY3AU7rXzt49Pv5tRSH52KZNG6g/ecW9o81NCPMpjKIZ8Lpfu6BZgCMqk+hwT9CWAv9
SmWXe5DlefLQq+5tBMmzhe5CaMto2Aysj2+Rk0fTGJ9mBpAKTm7UE2mUlbvwhQfzcT4LykM7jRZG
51V2TG5XAmtZQMFpzNROXvOEh6XvOXeb9Om4YnsQvDHeq0Fk3SCLyI7sVeVaNiOej3KWPZYnq6C/
zXl7j+U2+Q9vaOM229o2WjDBf1xcPlqYf9tCuP0QuZLm3Zc8oZXNPk+hNmfd2mhmGfqecrraCGx6
oU9a8Yg+WjyevkHzjzsuGlj9MXDkBH5ransG2zSUdMvdOaeZdSuxDlDAKONQ+03SMNgUDlBWD06T
KxQK6iM60lN4SbqyhbSTL57rfNFsEpSYQTBsUzWcnz+WRbFyW7OeR6O8YVcwRV/M08PI/oS6ot52
jjrf4eCWAf42RIvvKmmYrTxInyzy9FqE7WXjBuPFRBYpR/zkHIwWoZOvgnVenwQtp7UF33vn4Pk6
4xhKxDwe5N4iwrOI0lyfe8/vKvdfWDTn5SXYswEbIr5D00K0TXfigzNQIAHOxsDxvEezEaUgca8X
R0tcM0B9U2zlPUniSCKvnl9ASuZI+z4PtU/Moi0aOlbM+MzGVNMdSl+3tj4w6vbHSxEa9ehDoeJO
vLetRD2ot1/ohcECP7b9DccdPMWHVfCoTZFeYJhI35U8F5coJFjk2bX+mQucws4AcFMCGg2W2sL8
e6USkmwhSKjPZ0PoQDuamyirgWTq53vBOExvzEdluWOygvII3dWm886hQjWrLlH89QNVrIUwqbQT
U+QcxQ1vCnBMojtG+3NpXcmFx2HXss+msDgHCkqBQejyfvCm5gzgn7v2dl1Y6xbFO25XUscbX3KF
YHPHNU2WBxzZEhr76laN5OsUfmnVgHJke9FABKcdPS+XSk/kKvwouLV7u4XNsy1D6xZr8l2OrfkJ
SAumUnv+OCoZGa+czZolNeWMHGOso3Dtvin/d2VkWH2ixwVRsyze6oe7ql3vSRKWPR901BcF2G0M
3913f/ZK5MUKR59IbmcMJD5SFgvXebyoBm0wtY7Myy88sYyb/nZBxVNBwixAMy1nANDODc1XOcBL
ovD8li/GmjtS3azzTz6P2ovLe5VzeNA/WcvIHJTWfKW4GUmE6g8wNv/aBV1n3l+FYG9MfpDBdCg+
oc9CezmzGMl9lXBvj24qA6qV+Y3oFqoKfmoIyibgjWP6PYKqJqYerdOvHZQSozhtFDS8XyC2IAxu
ZOCfEYDAYj6xHasfcPJ19M4B3xdxmMsEq/2P/djtJsz6AG4fwDnL62ZDj77ZQuBnqLek3+TrGDVJ
oglq6QW75ZizdARGBz87q6UVKu2Gk2TUJ1m327+CWTbBRSTLYRS9A4ebyg8kKVH8iry9Q/Kdd8Fb
DsLTLRvmp8CDCYGIa7BElbIEiPozyBBbQNcrNpJ03szDbcTMjJDr6Q7GazGwnE3AXOyg6RmHO4nV
3hibNadpbtisgJD1VdtIh4KnLmnpqgBK2VmeBlO2Kg/bqE89g3lHEP9AF9NZiVw76D5LgF1dgRg5
lpZhLoivlWLW51v8NqQGXyEds8cmhX0UdkpifFXmD9UL9KLsMwPU023EBov6Z5Dky8VYRrRtRSwV
ITMR1FAmOXS0k/PRTC8+3HoVfLkH2ohvmxPfzBsQs7dxIPTt/N+yUerUdBEIrmc1pviaVJpguBNG
vkDAfttiq3rdCQWO90Bv2n0G4VCAYOzvl80NGMvMmG6WyjQWNBLMVXAuieasWNmqdlNLWGbJuLme
GKJsReyQWGyijKFTQZ04KKrvwXxCDNMtO9BB7+CQ4cYP/HBV7NoxW81yW6MOMqGZlik5uLV7AEUi
qaSppnLf8IzccekiAPUKxwJa48NXrCajzKeZSwxzG0pyxwbl2Iicj9z8Pip+2WFAKkvc8DAWHV8A
XfgDPxDYaFG/UZv5rMnPYf4/KlkqOG45FU24oYl/H+Rc2e/dkm9G+KT7Q7Wd9VD/4FV4qKICUZgp
pT4eDFTa2spH0n2L8jQaCnihQ9l6EOVUAsouYCKbDKmLHJ/X5jiPQOrSa1qeK+qFhgy11h3I4G6F
pSVoAR7HPuTzESRYjrS/BzqwZpS6gvcVtxRAmDycP2ocBJXZaIJvtRk9+xg24T/Nqs9h960ITbT4
CvWM0nWn1E/OHcRm9EOdpF5damhv5o9cYNe5bYTwWebdCJHUkGHNsgTZjZPy0kyiWnItLP+FrbxO
0yKttWNTyjTULIrPICmGoAPcyenHKMHYMEDkajCdklNU+UQ7sKQNoF6zfpXnF9I+d1yLds6eX2Tw
sNjhPqdT/jvLuPYvPYubMhQCiJXb3RlOhpAxbuRgMPeO+DWnkpDNi/4bkbMUVEMompLkCW34UYVt
52/Qpkn69mtKaJRwfXI/iOvfVXJ1w4nmhjfBP6UuUD+xIt9CdrRIZi4I6wiAw5G3D9NpfWlO9U0E
nDks76oWPT3j9XVV9vzprYodPrHSG4rD1/3R374AH8ow8LNQIYeITfPs7s00yQ37FOsqLbofBiap
ajWsgYhjWPxUB9/iqZ2f4BdVzL+u5qs4NZ0AdFpS61Ys4hvDa8J6bCo5DR+s5u3zWEOysZgCJmIY
7wKEy7TL3DigoAxEAmdEkBAwZL8jXv1liDrB1Qmm6M5CWwGb8JD0mMeVulp7KLw5flzZUqPPC9N9
60e+KaAah6BDI6ebooKsTsXkd1IDKeJr4hDNFnPIqqB6xu4vLfAkAGvIoiSGrcQQkGrR/TOC6csW
KF/LglUhGLiSHz6Qo4KtLOnxeIlaqYI5uTpG7pqSJ1HM7Vc0ePhFn/a4z7VFVTrf/S1KePsc6t6k
FuO8Njg6+pFeSYX2G4TEO01CxZRchDh+QBV4oGeS7TWF3nxgsaHpm+l34BESy9RTs03Z1a1IRv+p
P2SBGEiojjbeocr7CJ3vNnvdINO2gOWEBUkppO8G4m3NCEK9oQQpXFja8NcIpf7LlFDwaIXpVz/6
NdvEFmgPybev/javz0/95n4U6kckVywcnvWBouFxXuzDsNdDpFoGILTqqkFhgQG0YdeuSofdLWvP
h1/4cmtHB2YJQCuJUh4VBngBWwk09BMdDFPkMjZ5tdZ9VNSC6nr0C9ie7yMq58FKQlesyV0EEJTB
sK36gWGVGan1HxZBH04q7QtGTDlI8Cyq31jQoHysHQ1tF9nQL6vdMvfo95GlotUrAz0jaRq6kDUH
dM3uhXC2sLeO9Ns2c0gPJr3/aG/JqijRy2ofIpF8SGfJZoxBhH3oWoV7xV3BqMh8rXoO9FWp3l1M
PQqZnzIsCO5Jy9V1XUJmG7dErUVWZH2KveSS0qOgpAds9xwk+1NTUq2w0cgEBCKbhPKiJawlDkHk
3CBHsFW4cFsmq9DADLMKhpSBdFLdpXZsM+AhLItNSOvZRMfCkP2260IpPk/bXYfJMHi6eOXTvhLN
HT3hteoGcLx1URRhIIkLRIYEWlvmloOlNFNwZ0bCfYY7sWdX4nM4QcZo8esA8jYRQZKcRJqvucqQ
q3ZxyYIRSn5LIQMbq0T3aC8WkI5ZHgF+qPeGZYtQYZHnDCy2wIkxbQT7TAXnzeTgFRfvXSIxOxJ4
y6fXH/5s5czrYBSGpnmgn/fUu9NEYgLb+hlGGGEIrWp4Z5KGP9yrYhh2+SKJESbpiVJrbrVQjFLS
4aN1Jicrm5dZwxhPHf1+JybncIYAvsFsdooL6e8QCAmfGKXAwTW5qkudAlgjj+3gFSqiLqW8sL5+
ve9I93RPl2agxpB5RC8wr+XKZi2VDhRm/xcERtTKqAOurrZtk2uFXES3FhR4hsXEmTOfqbQ244tC
aBSmDy6JSzc2igBsJ3POACo4nOrRzTV5WCOxGUoQrJ1EF6DXIkRWPitikoDgUJLoTEIIJzt0JbiT
jQtI+wjDTERX393jgXpFUnLRypbWsX7v3AfEIrEbo4mOmug4TPhiIar328iefzWZP/PSj0bSjHrk
yHmZvj2jfLXpGHU35Txh9bs7ZD1Y1l3dq/zT936qzulL1dfKVbfUK0fTvnvga9Kl1XeFTyZhBgwA
qbmhXpgEF+qzzgiyak0gmZyCxHYrUeb9hbUDVu4J23Z5dwyKOqGQCXKGmSzF9zaV8mRPBhwOGRJr
Vs5l7dZoKNsxJvlI71Svzud07YH9i3bFX+9uoM3HwmwfQPL1A3KV5Texmkpj7yGzOcKRoy/hl4rV
9MIx7+YMYR0ZHtuNIbvKwWZ8PBBdZwb+HbGkF7W9FGPbAwtPg+o1sVTnD/xbWclIGK4f/sBTg/Jg
ToSCUd0V1yQxuIqXrr7q5kOPphP77dvDVKFeKCRKjEhFVhUGenrt3J7OnCVdR5UFS5ShPQezq8w+
pqC2dlCodlklt11kej0GG0OCT1B+m2UzQTU3bMv9eKhU0RCo+x7/NRRqqchDCFJu6nyEYiJyHInK
g1whK25XpScgOqQn9/NveLg4H2/KKvFzf3C7VBK52OD1kLlXcQGy0VW7wZCxsePPizMlr4ylVFrP
6N2zwoKewfmHvk13Fyxt4MIjabJmVtPAbhpfORJLv/zXUFKruZpersFLh1hlODwcsl8eZTYjZtLc
rvhWGGCYhj1LBsVC8Eb6eKgpXHGw3ZJXJil/dctjg/D2zUytcrWstMTpIEkyk/Gt8PRlOd9B41YW
K3pH4nY10WttwnU9pASGE6X/wCae4pM8K6lEFRZRgQYrm4KffqZ3fxJ+4xvbhx3pgQCpQ+f6wj6z
rY2XSp5oaJGD0E93y9brKvG5W1EurPWtRDijEI470UtLw1B+7NxZjzv6u2WOLUAlfTFHbsLGyMlf
5OOYt6yfZ+WHmMBn+cL5X9/ayA7J6Bsus2iRUCGhxBP4eMk6cesBQ5lovX4CVY40uBYMowggGGwB
BzUa4KBEJVq2quETSePJdWKALSKR+aVwUsvQZWQWZ24BxUubreVk7sfpsSJYaAWjPE8gRG2vS2S5
CN0JkC4+gENNW0KSoWOaPFDCRPPlVyp5yRvNbT/uDKsSq26EiDH+CjXpggXThx8J1ZKFRfY+Q/kx
OgoWS37z7AG2J/tOM+2qaeeCGalvV/tsD7xnm1RJKwUetjvrRUCU32QekOBV4inCFcqrqyOD3pVa
dwfpJNzSz6L43KocqYBOM/+sKZLkOudNoT29nLWKZdVesGpmMSTn58/E4iiEf3++YaS+GjQounXl
eR9HGcpBgg7huGWFrdFww/7q3RBC6+Qb6PgprX/iRLdqAG4zY4nOwaBOaJ4MPrXLj5FACVnD2Oom
z5Lrqox7+tRYI8ttBAYrDoYruhJ59+1XzFZ2l8mgTWUI+l2u/AoXdkAnR5Bt38VKVIk4kVoTYUfv
hfGmI/JObvndOFZRY/HOS/Gck17ON6MDyHiUWAHP/auuLkThGo6nA+/+KeoCFR+hTPOggoz/vYVd
ULwYgblD0+GbxXv65r2Wa3nAreDAuvtyjk5NzYcdP1InImSTRBqU2S+qvqEP7uoJqAHIaeN/jWuz
i48BHqOam9KOXG+Ca02BFZ3vWa3IHiaPq/t06kyl3CAHUYkNMr6DqGKq/xcDtn2BtfjCqKQFTRKd
IexVHz4pEinhcawsjysQ3gOBRed6G+gK1hB+ZJhtS+2BoZIcedlljbNmlON3Nu9/EjmKu5ndPCx3
38ZZJCfaGf0nfL/Y1dOL2GrnJmzCTVl14QJiCbSjE+l5gliuqeltvQ0sPZEqjF2beclGvINuGo4a
oPkVi8lSWDpeVb6jNjcK+qpEoMtVfqRT30mWPXO+5Aa820RAF6Ud/R6ttOLkoBzU6/hTejd6FAO3
w3NMxAoHr8Gsx8KH5rQNnYXoAYc0qDUZLsRKPH7/40uJQstKkiO3sJvsdM3qC7bglxuI9VMFscHf
3A5okVu6FD9jhFJ3nxcCu0XazMR9xv+h2faqzdCyzjqBRXWAO3yi1gf4AKdrJQipF4yRhf7RKyVU
aF7yyKjQ5VZVGcCR0WM18bx7+xtdcI/NWIbj/vELJ2/FrPmdPjgo9JKB6J5+mdcUlcFChDRoeBZh
ImKLo8rfYMTlKaY8PFQ35uHoyd0XxxsnHDujXFpcEn5cHypoFWiTCtJfJw7NypP8yPl5xIPYLYN8
z3pCsJxkHZzavtmAxCBSLMBibS0a9oRSt0Z9BcY8uvA45djMKG0mZ4B6x+pSped5btTeHqE6oL3/
C8LfNoa0wUNC8UrNkyjLBQA67hxM1KHYO4anofbTpJ69bCkG8pbmg99+3l5zg8fziEljQIxrDkvK
GkOMaEc8K356rX7NId+kir4ZyHKIgymlZaP4hqrhxexRy+BXAwmCtoSaSJyR8QhOyi66+9EMU0av
y6143q+DI4Iva7EeGIOA9gs7mw4V8UTxu5vsA7ce7QmY7Akh+lExdLNa0G8SsdmGNCgvxywmw3BS
wyHi2TrnQaKq6vxMPqnzd/jUuzRLjEYbmQdko4nMetxTJjgeBNwuNUFGSmrboUtx6brtYNkg4ib4
iaxnBBRfo8kHOED4uoDE6lejdKf4lgOKD5otTXOiMbuUugChfgH1a/OhASsFlGKqwChXBlDEoI9q
L8fgsvmXXYntSsE5oYbKKmMoePoegQouVzzFFNC2eYQaiW1sy2+nYESo774oHMbMAa3nT+QxIgjY
SZCTvMOXnvcF9Ocd4GxYnCCsm+OUrzamML4guKTkv1HRib29ll0xTRXqWSqt+Qmis1EmFGeS3JfL
N5i3m22W7u9kE+d1NrrEHUQbZ9mC8oqr5T/OKavbF5P+34sUcsNUfZhzqDgU75/86UuxEdnYLPVq
pSbT12OYE2yyCQHvc2MetzuDnjYEZCqJEzPJngguJ2Or9JOF0gDqsZ80RrjP8CoJ91udI3+wdn7v
C30NQ2Ewt6Gj0yHxVZ5m98n819o+y9XtUUORmbOdnX3hWFy2UOpCIYN9cZs6k0oOMe38/LsgDLPn
/4/xihZB9e0bLTk8ZpWcsNO8VtDI4fs4N9khrc+Eu3oSUd8GoMC9A7BYYOXfgVk7ua7gyn59kR24
/7ZpPe2ozud4LaCxW236u6Kj/1ctgWNiNdjQ+cSXuHLSnClSYJQEUS+SFZgK24oAC0y2cjyr10Nn
XafG+5czPey7DXHoCmu06HuNe3mfPjEzqdiwCPTdo7Ptr75m5n6qVYtDtZN8JMXRTkjYmwNcbORR
NvFXwhEzaqMz1/vo4fNK+gh0XdbOBnEJvK+mrA61iyfsKdNKyyhZbLjXVk44kWWIATiuP3GpBxSm
oFoHVQKLfl3NNtbHcIM4xO2rqg3X/IWnQFqBdyK2SOwBUoEqz1aDnj7BowDOXdss6bsPprv9bbVu
oPo/YQCcd7OpUr20UacHnHfllkize87Uss/4AMDzoaDi0598k0g6xbqsSEkuqstvsRv7coOYNjDR
qs9ai+LH6TdyORbRVyW+dTsSv1GerJ6+AfhpOVmyTkbhGDhJ7m8RSYzYZuvYb37jLDBaZYjexHZP
UZTAbeFLFymgvbPGfaWfO3qcCBTSeG/CF8gnmbtku6t+eRrdNEeYifGZpBSYcEFNbobiNUPUjCVt
h2zpk7GgQ+qe+mVIr0tYmxob3f8eHfLOfcmop82PrOmTF38zKKLmhKxkuCbLQIXLOKXInLvBGW9o
FEdVS/hZSZHOApEW9M7sYHYYhGyL068LSmU/iCoUbSpa565VjVnPmkO9jHGUbur1v/WzuhEdj+Mm
1BsH2lED0viA7lTORhhvdlR9xBKph4WWtMYQW+W67twwBbWKoaN/sDqA+YEF1hnQpnKT1/hM6cj+
iJzS+aN2/w2VP6rnEY6yJ92CC8giLnyRursfY6UXgOwr2xLpeSgBzfpL2yxFxWybVRlRrOKFj4F+
fW0+wY3YDW8g+oVgf0exs6FmTuCLTrzs1pHM4KNt4fPmg7u0LW6DanPrfMhwbSYqlFbosRHWMCp3
76AWYYXU+cwKZwEkmb68W7MSr5ZRGQnd6hkVbYt2NYYwMncm9Gk03rg/AJCY73vZPiIln4n5ovuj
Mo5XrVQmUhHI5y1vobc9MDQoTO3w+m6UamgXOvdz0PmANIwJf2qqreT7z2G4XxjNgZyuvZAfu8kF
hGDa/LpiUaAi2H7oviFQEAaS5IwIxLH9UvBYLa5G9OfAxR3v1dlOT/nrFBCVeZoS0OY8HS3kvODi
N5qQvTU1dcs2z7J0CxnC6LFzHI9x/LWlaOvAmqwuYssyrwHjBn0FsqXUGDKtcXWRh+qQ3etvyzjj
LlBMYppvB9ND0K6nQ1aspmK0YOOW49uHHLK2I0WpAE+R5G4MtCyH35W6YW5aRmkQBi0dOrnAvrht
zkkP5k2CbuFfVF0gTIAF+8xO6WPtYPRQqx17feLE51oLPYivne59ZhOPhEdhgvyd4i22GsfuLnAU
XTKoxW9IOTJLc7PwnnSQMTECbULFhLJGuHUsf90j2nWjI7sbKMqD96pGq5kN4DaIEvAM2kZmiYWr
oikd4/i5iZh/JsczEwOriC575I8v99wLwfiWLjjv7nLzhjLfI3UX8xgxqyznr4E1B51/kruoEEf7
IGhgUkq+3FRZXe+Jn+dU7xjOfvKD/MAN/Ghb7/JCnvD3NXyqyLSRXRf2+M8jQy8AMyEcCD98euwV
xIgRZChnFLubdirTT7cu0F7r7oV14HQRTQnPg/LobfHx1epy5dTEUtAM0dXI163/64ITV1uZfY67
bBr7Gz19cAzlpyQ6XVhRl6fUl+JUYhgxmu/R3aOfzst1i+wSqY0r9Dkbfn5wWAFM8JckG5xV8CXx
mY/Y6Cx7fLixD6QumNZuTB9SDor8mgak/YPLd38m4SorKAnzAFkTjhqTTBvpybXvlxZH40PSfmuz
W7D6afeqbvvrIgd3n8IlhlFaau6WUecZycZ0mXhNogppSmavBZGPgrroLui0FpityQ47xxVQpXAG
FxBGVFC0KpHXvVWU0duFQe+rfK7pOTXi0i6xsx+3UQk3h9BoXCarBHzblmuo3NdkKKjE4oLIKdMB
AU+zljgoASzalnNVeUkUnYticwcfZmu/Lh6E2TIH2rTDLXjmEd/BC905uUASQZrvfao4hg83eZG8
qRWgsUSyKuZ9yKPFxPTd7XT7FhjxpLpczlpj5aHW+7fSj1MDqzXvJrkKDlJYRxsIr6ExK9FKbuXO
6W1BYyj30I8lyHs9dLtSNRU2XS5fWyv6lUJaS2GJRkI8sxWXxBYnBj1CYkBWhJ6qXK+BYFINeAom
MZvC58AfrB5s0pK5NEeeOo5r3IPUk5T4Vo8GYDDXN3I3T3yB4ysT5GPekTShd0+dN1lAn8Ek2S/E
Ni92gBHkZI9+pYV4grjKWQW8Sgpkk7UnyJ8iuM2VRrxI3BEIcx33MdJu5aiCTBtyQ0c0ut9dXdfe
lcNvwwlY4C2kssovonAKM2qdTXStLCMW3TtD/kQWcCGrgeuflWCgkaGbnD++hEpP5td/Qp5T5zC5
aYoiT97wnaNLr7JI7DhpU6sms6bJvGm745ZTrBIzmf0S4Z0v/VHMKSifW+TXXWA4kOp78tkpxIGv
nH5Ib4hJeYdHLpOQ65UBw2Ic3RKLAb9m/SPRt8J8mMyZPBfwWbp0vzTtkWRDo8gKbwu/I0rtae6U
8fatYn0/ss40Fb8lPGi+p+tYsrhgSou1CUWMbfSkeiQU5271BFDWDQGX30ZQiyuuf3xz0x1SGnnG
VJBkS6RdHALPfLVHDjxNX/LR/a3z23TODp7Fcyn84D1hGSh8RpPodcUtZg7i0cTfptGO4C0zSkXN
44900WB0hFDsdI44mGNdv4BosdJqxf94gerGFIHl7GOw0HdeUm9WeqjqykUaygChgrf/V7xyHyux
ROWPsZ7c7iP2vtjdpqwt9CKADQqt0TqvH46xIOxKZjoy2Xn6wXu3TI3Qr9o+nhJsyNNZs3GHe82J
z9L+UbYe3zPSOgyj4sEE7SbFFMnW9CmwhSiSid9TUal6FeMA0/AQBEO0jDJM578zvrwxRVZuAw8K
7uVQ/Hxjowk03H2I0ZEEKO/debArXCn+RVEJF4octE2ceNFBeHsHlpIzeMac747l19fvhuP65Flx
06k2X4/VgkVdcI4jfZz0vz1pQi+YzPaN/LfWjOI7YksayJ2ZzTCEd7vhtjX0C/tfJHcwbtS03SF+
ds/Kn5ynhZO/n7G4wzbnGj1KkBi88tyOhHEog0L5bABvkD+gJ152+ZuZf5RZ1P6XtpUe99cza2j9
b1QbjfUNTtmfpCjICaMlEQIdPof1ANKEcM+DCbBOGE6ZA8bQ8ra46C6IW/yTjvM6uFmcoinp+FlN
/QamA6zaUPR07NacBA3+VWHmKTPC9KYt+PQZiuONNx/qBc7r5XrILVY4zpbFFWqu97XNox1Hgt5z
9p+1HX/W5S3DOER1iIUuevu7giVqLpr3Cvl1i7KKaD8Rjlk3Hf3tLHvPii0/CaFpdB6r3FqMeahG
vbzHbEw4UCSPp2EspSU4PigKQLpa2Suprxg+t4ViUZJ5VXUo4o7IbDMn2ss8lNlYGrxEJfJ6R430
RYJtNfRFAmhY9DPCuMfaetUJL7FrvJqoqP/4KKl1JEKJmFh3TLQYNVNUV8PjbdqG9nU4z8uj2VBL
6vcCm2TDhnS/+S+akHLjktX/mRTBOxJySTUWUQ62UAWTKKcrBwHsGDEJbrp4+rHc+OIq3cdsQ2Ui
Gp02K4fkJf+tRX41jqxRHP5MDfTiqav7LDJJbt4on2PENVbIoHSD5CF+cHD9Mz9qLyEVFjoaNSR2
CDabGCnGoRf9TTBxi5q4PhKNwoeeHNnvxe2pZdAC0101DNs+sh7J/wLY1UYuG/ni+skYTITL6G+w
hJj+W7rGm7RbyLjkhD/5r2PWYESZJJhGFK/oT2PDPvRBPN3eqLZHygjNTjDElXKrPV1meJYJEYV4
4jXPlm5oI2pX1wsVz09r5CDkNU0i9fhc4dItrK8/m7S5/23ZseNr78IevNQfUxOOtMe72p2z2ooK
4N+0CyL9ytEM+J6+BZyffj5MXlp+DkNfl/gliyEqV5oB/EDRWN+4KEMLwjNd/Dn7ojZSu3WUU/9B
D3X5g35uX0/k98Ov8sZ4C7kB6ATgXuqHf37Xp+zSYa9kUvMWocVWwdNAx+Ex/his+CLmTlEX7K0I
8QXGE6AA7n6WSen8XxsLjwb8jMBQUDtXvQrzyjJXF+IT8/l66bPli4zO6Imcvs5X3+hJ6NnXtXO9
QJ359Ve2n9BV4BHJ3uoevUX7Vr3Z62zdEVTGcOTU2Xki9PcZJmLJMQk6gzhIWRoUiYPLP9BCG6J/
cmtCcuyDuyn9Eage7icgO4MagL5SScCCfsXVT6VKbAr74lP3o2aMHNLRBjmZiWtKlA5IhOov9wSv
IrFDohZfkeJUOtwBODSURir5b4KL8d94nWg8SplYEt+Dx9xk7KhfFIGd0OWYmQ0oFfU02hcQQnd5
qyaQRLu9o4LtIOUZNMX5WDe969jaJkPD5mPsC17JUIRb+3d2utYaww5/Kj9z7yCtxg+uUMdkrQqM
8RZp9RD9AYHTW2SasEDY1bDpyD9RjnMkOKpaizJ8a+JCVtVxRDxErrbL4kkqM9UeLLQyU+hy0byU
hi2oTFLLNnAbwyL00AKgPerS6lrpucAcktHWrvOkqzRcPxZkHCfu4lmTiO+vu5TnbrkK708oRiC4
xHvg4ecnIv4btiHDbje31JWlJ752/mkrSDjunQZcOsDyeMKWxkH97wxH90PAomhrvKvrRfQdrsSW
1ookdp5hDOEgNrckNuCfFrzuEVq2DzVD4gRKng+K9Uz4qSeIwl5+FvpAfsAtRQctPbd7U5/YmMXN
GtgC1gA1XSUMFQVumB+lAF4OUq2ZhWkqUV90fY2HKf4zRfKucqJZjQnLH1i8E2m6HiLTlmQtsWNK
rAAgp45+AbA1sq9n76mXp4W8ReUOSa72DNJbLpVegp7oNT0eBtKuQEjr+ju1vwq6pZnsD5N4vf6O
QZ7zvGkjwGMugGidCw7FGMnQijkk3iGsTFxcEuEKZdW9d2JbKBIcTwZshCNQHld2kSZiDwinA9io
AwO1TG8yR+npLczvrG7DmyaR/n8WP505AxxEq6eHTQrXLCyns93/Q5yQwM7z8k37+4DppDipDYDy
4dk5KTwSt9NQYVMH45gSkHZlxSfuAII40dHQkIwS36hJnMuT0ZVZq1LFuyCcFDW+ntEwbYpQsM0e
feMKp0qtyT61xhlSJRqwoqRd3sm9akUr4j9skrdMMY+Jp2eXE9T6R+V2hAPCeZdGPkR8zelfxzE0
R316FOqG1YNaYouJz1/0CDTZXwxerYThYnfkcQhhUaJiWiSlivb6HKvZNzILd6QQIH7TW5CyA0bv
AX4z1Kx7qYF7zruRrVqtSAolsgf/39eKvudmXqEdHnnSwiUPZIiGi4kJ+lgI9JkPXeMCjK3mcIRH
j8+T29+x2qsZYGo293rCApe7QA8OZO/Rj/mByF9eG9qYl667zJepL1DS7S9bz02PZV6UT5jIhwbz
NiPqvCtIBrJFBjUP+tg3EOm24liwp+oU3/61dbCa9BM/3v5qqwTIMfWgo8v8O+MENGigkXxJ7IHb
J/lcb/GPw15bQ/UIUVKIVJ8KcLBezFOxXgoXkojs+3b1HlnARkFZCN2Kw0w+iaLxCLTN/AOsULxN
5CVd1KWND5w1E2f4H7XdiYJnUYyNmCS0pFRjc8W4SV8IY4jRgstkn5vAaMXAcs3Ax8or61e4B+bA
QLG++ma+I6eDeYg3MnUY32b3u8WwDQR+HcKZESurkpNyCaz3/cyixp19MzM47/xZGuDTS1hq3K+N
MtGW2qHnHo4HM5tRdUkufFqiNlKvXn68DRlpAcFjT8wmBQJt/vtm75ngChOFOMT57RTrU1Y18Ywu
l6JITI2Enc9V69uJvhaa/epwNSgIP933al5qetBAPKQBNyyrWFSKM7jCNharHSMFvDG+f/nDuZ19
CUvoNa5j00ztIoxhrFCZH6nq44hpdflwgsZclAI9qg5OD8ZDHTSpGvRPHBvEE2Wz7Ar1PCzgEmHG
39JwybtQRGVvFPeDAmAy8LhsibKvpHNhCnq7ZoS60BKRmeTCZ1C4mb68V73aPKLW0X3wbk2Qp3Rt
qVxvR8IFyjJCEq9CzyCmpCt98csHCbt52v3wswQgg5hO7RMvti54XPY7f1OuAAmD8IDQWmoNSSLT
bL2cOPNyL9lPgU0DzXTsNhGF4UnOgWioOKGI4Dibg734KgeCNP7rsD2wDH1/pb240CjfGGDkayEi
IEFetaoIsYdWNOzikll8Be/Oc3sBn4VWpm1rY4gbQTcxhCm/mUXWHNqhgahYGm33nl6ju2Og1VzI
I+5CxVQx6EN2mIma00TilWNJBXDFaJVjGNf0ly6wcvz80rRLtYuGxFqyRPD3QGyPhg2LDu0IMuQY
Na91F7LwLMaO3gdVAe/0/lWc3icWOxX7WpW3SDJd6KwfYQM4yuah7mAZoNjA++RFPvTTBDt1MVRP
gOX1J6h6NwK6aPT4v+nuJGKXcKIYdouiGc/DHDbv0JSZKMz75z3E0JTemxA8JHGtKCmljCZZj+mj
LjlQ9WQxBDOUB6FQKxTmWA7syMeJ0POn3SWGDJ/Ri5LCvSOGo1T1v42N1uRh5dYB17Iw9sNyCOX2
9qM//EV+PjONB0AMyGNT2QNHq9dAHxgMbObUEMPLkKjmafgoFjBd3Qovg5/H7mAc6uwPbyOYHcVz
9bLG/XM2YMPHawNXRElObpjwKCKMa6wAXQulx3XTxeroCYylWqJw6Sv3wEChvbE/dNqE7w8iJ4Ll
lVLeIqpgoCop/LtVs72/XZHq2Elpl1GEGV0OFdZBGnoM6fQS40GWXlsQCILwlkNUZj1wkDQ579+W
JdFAi7/quq6+ZTwEMa8hXMPDX5vHTT9dAYyApSccK4rlqt92WWeElmN7F29JtqTbaAk6ESJ1uWW2
Qj4T89JLoj1h7dy0ruam05P1Aoau70oc3L0+QcT+biDT+5eI8ORa8DnFL6MfwIBe44HFFJlaDEtF
eMBglAcwuBpqIRDFQRfmUNqmJWLizkRG+5wMOvhXR1IbFTLr2ORBgvtR17YvxKOR0tFyPRPe/M4/
n871dlsVWF19nQv+rvCNISJzXoDWEHPkibit37BS/aiCjg109fq4Uks5HxNBDOAfFBFqV7f3M96q
DaZg3s5Mdjunu/scCfVaqXNHGu86Dc14yZOSe1/jNnjh2rrwPrmfVqKMDjTfAZmrBsX8auzYpay9
Z9DiJiegKPbA1LZjOdQXFzvU5VX/NQzGVzzQOL9QTuq2fAuEHjqfiy5abNB9b64IOqiMGbpQoBdA
K66Dg+rM2JmD035z57DN69JM3285+hM4b84R08Su+oENMccp0ZXB1gtCQMHPniVZa+6cInmSahOq
bASHcQfch9ki5bufMgrjkW2cLvppLLZxc1Q+wT9+qePpZTSSR/AopTNleQrfXZowFHGNN9iumMAs
7dz24m31IjQoNGkzsBweaaZBtz6DCyZt0uXyMDHunYJQbXV7Kca0U6Ta+9cC7Hs26psZyvlLVryR
dcRG0ts/h8qH0O0tWQgCcbUtlRty9L/zgsO5/UPUjbRt0sd35fgU6N0EpTmaivVrb9AJvm0TnPmI
pO+0d/a2FuR+JM2Bo3tLfBiq5hdKrHpGmrZ+2IsRCXLuUh19hTvSJ7wxAK6td2FPIc8BuL5wiMZJ
TMMRsPqbqpVVFlUv9vLqcccUDiOA+5h5U3ll0STblkPZkK4LEdErXD5CoLZyXnYQDCbjDVv9ryqd
PW590p9lrbEk5+ZZHRL77W0g8c7XmmFFQBCEtfkN7P58XjybWjXIAJ+1LA42TtoTEwqvkBqf0PMG
2/a7WHPW91slMnrS30VYyeEOLd2x9tdlRJXPBX+rRzV+1oTnHFfB43r3hkMzcSC7pYJ6zOR9ahGo
RNnSRhnhFDm6BGabSVYTJPduee/p//2yBBN8GudWKFBGaL05saMF8giYGXThsUskrJ6tMj6NZFmj
GyQp+mzo/bfNOESuk/imMNalnAYuechGnvbsfkZE2z1lZeNJVC119BNAtrneO8TYiYrB67aZfhNs
eynKRLycxnxUpw0pJGvl4aFFPcSOM8au3hDOXgdVAiAnKVRXInYACI/yUwY4UCI4o1HAywLvk6GW
m/VbdWvDX/oZ4dQPNvq9beYtlAGX9uwfzXfHnJaHc1JuMqu6RbMiSMMJv3J62g36J1FZ16AA64Uw
VfxZs5q835RHjfJ19k54x7QdOsTtVw8oE7iguojK+PuELoAjoBbCutPvTpSE//1p6F1uNKZTUTjj
IeCfv8X3JhVyDAgOpTZCw0W5qKS/Tu8FLaNagerH2WU78MgfVSzpvqiMUock1SQ1zfp5VBVNzm4G
DSNrEZb8VQjrlsXIhJr15ZTeu2kQEz4D+xVFKl7i9kXCxDCjZBLKMBA7PGM/kiiXdyvh0sCZswSP
IDJqoGf19okEWUJcslUshqKRwnLXGR9MM40eggM1XdT7g+Ygn3beReHrTzdWUgKkqny1RMBPMWmD
XQrDItQqLhwLXGmCXBSAdOBFTf1bpx7CDcSk4M7Ei8dreRe30w2diQ1VaJyd0koJKjdMOTzL43CY
Lu7WWkPJUVSXlDlojXV7s80xvBL4b0cVv9WLONF/dianKmZ06bC2RKvnaTziVz6MaFAo+9Ekda6v
OqvW8BkCbs0wO/jimavHWN8wgo97NxL6dmy+IOuq+4WU0VeNWmaj8/ykQ2o54y2muUlxJrp/DK32
TMTCAAU96B/wmVdRwZZPJRdKYqfgDo9do5WPn8Zvblef1pdGXbe/O82JLH9TbNIq+t8eg0EXj4sz
K91kz4ihQZDw5o3Cs+g1alcb4LZNVVYr30+zvp7oH+41YpfHrriq/oY5aPlJ1PneZ6FafSfeMl3B
6py82Akk6nRBzC3AqpGTfX3X6vjDIij00/nLrWJok46RljL8oKh78dOxpcLyyPypEqfv3pE8BWi3
accAylm3kCe7Ofs0qRBRBmL9wvVpclz203vfe3VcxZlYGhbdXnC6mKH69Soh3JWWO5/mrSy+ndC5
06oRtQXCE35nYuNI8eZ0nTT9LvQdhYg4xxX5F3vwvCaLqvv4eeakJQHycg57LpgJsRTnOcr8773n
8t+r+e+KZs5BjWWBuXA+sYlwClXS+2vFO9NPucMmanvLfLZn4BieUFL1w6eov5k7wuIKEeVbpMtY
Prn+iqYWzXOxoBWPdPWqva3jQ19aSASFoMwgPPE46yUFjTnWi3XXDhrwz0RnqQUo68kHYCdc99Jb
uwTZFJOdky+q9HHz+H+uT1i/gPX7rrg0jDzVFA5/ZeTv+CTEO3l/qf578Y7681knzt15rutSjD2+
2n2n/eUg+MfZ0l4nIYCXuqDLrWDyX/8Yc5LB6pA+hyeHsXkZoqvwKVCfUVwuL1bNQrSakvpv4B6E
N2gRMCbwkUdbPr5W372nK5WqwTT1qyj+TSl5QeOcdXiOqziAVtDx/OHsQ+AjbGN9yr+l2zQGPHIi
E9ta/Iv/oHM7i41/Z98Xlt2O+EA1y4GaNHRgnpSOunZAD+Uq6LRcmwf7vh866lrLjBWz3l21Oxe1
8ZJmbE6V69pYya8sAnLxizU0eskbVFWxTP2xCswinI3ZhfXHJCF24KgGcgraCIMJEL6T9QmSK+5u
TJu07S4mOKiquZzC3HfthbTPqAVYkrtOkJkvnTkXW0FQnnBNrdgUPJOdv3qIS3u9BNKaVSR7M0gg
JyWigCa34EDBE5dNZ04t5Pym9ZcdZIyK9R7kD92YH9fECfzaDpaeTorKFo7n1JiTRdt7FRBaOKVn
PGJMMQHl9D4NCKjsLVq3TcdSRfRQ8AniWlqUA3AQjhRwBmfupxoyzMoYPGCzECn0jOkOty46bSrk
pEG9u//9uPvE168vCUFnE/Qz9d4K/Q657uM2Rwx/hhlqgo9fP9/AHMB9Mm1Ud/ut5yzntay6MBna
aE8zHakrhqO4uV8WJMG424AP7y1FDgQXYLkPgFfjhV8QNnmsFn3mvpiMLpHPF9/olFWeSYxOCWdi
EgSzRew2bA5ec9D2RHeU8WmC1WcKhhvikbDwhMN1N4UaWbcLNEyQriMMB5l4Lic2h3GLnf6oDCpl
M0Rmu+xXlVdmPh3keSW8sYIde9N8b4EuFoEfjSj6xi9oZdZ0rSl4FD5XxDis9vssjO41rY7wNBT9
8E9xQsyxFJ3NA/8fL8ToZ8iTKEdC80cwxSDh/OguLmOZ0SJIKiW3hp6tVqBi27uuWXn1vJo/Kt2c
X8u2lRF7xcQJVN4FXI9lvFmGUphswvDKYtK66tElBxebWfvH0CY1G/znCybts3wmVmwO/11rmqt+
CBg6Ja8I4E/O8GqezsxPVLCMPoQyEHNru29sY+MjDYCGC/nU0GaUc19sL2qjeA8XnAIk9HZh2mXF
CnQNJHkiezuNvcextAbAlPUU8qFntkzpGsezasv5tQC4zegJx2OKatQK9Y+0IZgXhHJtJbvy4OG+
jmVMS2p2oIStcPBlcI1gX8EKDzCHurtM9kv6lDQOiRMjWx1P/iCYyqoUhpK0lywbmInXqb0jS2gp
WM2ywLoCuoZ/ib8L+TExyalwdd43mWa3U9LuNnrf5Wz+KvXrVzsSKx4YKspWnKznjiAT5ksR/Ysp
tJmbuy1kIOR08PikzRewOhE7iS5xe/ittqXCpeYzaPsATcnrml0HXfRNnMLIkgT48Bq9MwgTdazu
Y7w6b1I2Hz6kMrWCaj0oFeaKIxwVlITOlPivo8+RmNa/ANC7aX+c1WkfVHvYZPaIviwWKUm2OJLj
HcvfVat1EACO8ft1N4vTHjc+DthEMQrP8lOYQWNFUeeaxLpB5Ahw5lXY88l0NZY5vyGNC/Vt5wh+
OGIx6HogU/9JkC+ilJMHbhdQgBWtkyzyXFcFon8QjnkUYHX47VUO8d4ugZnj98C9GnDqmMPZg5Fh
NwslEmIv5h5N49A4Y7ZCrF5rcd6qEkEd5noJs5JRDvL17mxLEwqT31bkSedfXPNjlO1/IaqyXHNf
W9avDLpwvgrXTVqcD8Aka3POzoXrCAAK4HbGTokLTquB+EEzZENe93HV1jtE8TxmskbgD3Is3twn
VRu/SLDkE2IdsKRt7+20fyN18gupmeoQzXQZzikI3yBiK07JFyNh84bVTHo0l5ClbiFSXWuv5M8g
0vPUDc+8pPlOsBnvCL809mnKxB8MnfZlRcN8FgUfj06MfA82TgkJ7m7veSlg7QaRprmxRgtSYIH9
7EBEuGVYIxTorjjX+Ahrb2KwFkztCjx7+5jF2E0wfEBv1xGu9MR3EuFR/kPXefMHv36fnCl1wN0r
IVNgNUME+6LAxTWJXFU4WvBD1F8FG3AREQrjqncA7vlNP1+U0A5VJXKCVn4GXJI5Phs2w9GUOtfV
oykbS9XFXZ7BpikISUYa2tPTmTEpvB1TDr7R6vlmTvqV3WOwtxBUSyF7vms0XOWlrsuY90dO1hYW
AhU44FVkYuwu1TDGGhOXxyNfc5y5DAJKCnhAIxSnad5ZukS+3muZTrpFvmtVht3ZOnaSIRBhoMAH
wITmAXbDRtNVSVKZ/OB6MSFdl1QoIVnvy7iSnlZFshoCsIg+Sb6u3LOaCGiNpUiGigDsazqwVzQS
/BL41Xme27OMDjQoxfnPxS3WhKP5v9HE10R4RnRzrGTVXTZXT6hkQ70iaLrsVfvDb8Jcw0EUswsk
iMCVEk+QTcl9kOaExeybpiHbVMxwZXu7E6k9tbjoktl7/Oci0Ac4/9/aBk6NRlNjI90bGg3PU2nh
tkrL3ESIpjLD/GeornShWW6jcD9R4ibJ5pmsyMuWws7kVf962Z3xQWtM7NZVRGPXNsJp5zhPUY57
Uj8XxFWm9kpcNq4kc3Ctqf4QRAYMXmO+DfI8aJJ5FZxGskcmAoiKph8epkC3m9jZsRXF0qz1GHDd
q+7c0gKLdXwbmftB9TpVCD4wCXwHthtyAYsR9MPoOZW0psXkLNun6fpPdxwQhJZuFso90rGgvfd2
40n141VsOADXIIKxhbxeAFzD5ZNa06PdWlUpRtmKMaNHgR7yZc0gWzxZNl7NJI5+GLCX2m8N3HyH
GVf5c5dWAK7nLhcHelzYZ4QjPXku9+fqp1OvgitOm6P7pB2LpdSBfz/mV250lzLnD0hT1Ks7w3XY
LnqrA4UfKR/nEy7e6X/ol4a38/E4VEWJm7wlRK0PuyqC90nd74cRZIXrOuoxe45MT0jmu9YYFF1x
AQ4HBhajpH6vLkDs95WnAMW1zd554qG7spnN8d8pwy4K7/c/WCAqb3mUKUX42Ulc1xGYawo9dZV0
geLLP7hwSSkjOa3TfeKgFTuIFGWATE+wBLi/hp052JAPCtjpOp8WFrFweMAMoMw4YHYTUl3PxNzR
h+VC21oqascm9wdLalVe8wdyNPHmMJqomaV+6GOqCa1Le/kl3ogBR/Qi1uoomu4s4hYyaJmiQJyj
HiAYtyle5EsVqI+1RbZ5lPrmPfPLXEh/dX7KjR8Jdq9ycBKFI3YUma8OfNPoGtZFGZHGkGf6I++7
8G7jxS51FIyoIg8Z3SxW9zTcsB35VkzbkILWGOxyPY6zA27vssXfHkuialLe4EAU31K/Xcd5VwTd
E2hKWb3n99KSXSb1uIouLV1GZBAiyvGuvFrDoPpyaJg8MAX+qGo+TqmYujAYP2MxU1l2pjU0j+m4
3uy6EG5zZ/ciCPxq5EvNGM4TtaTXu9N0LXfDxM2AgOZ4717XLEPLc3tYzooJBVAAGwQsYg2F8VUs
QLhpAXKoDN9UjrM+0HIcguWu10sUENSbzjXScWusb95FilpDxCLMps9/m8S7mDhowzhQsTjfqJ87
5/+n6yB9YqwF6r3Obn+EJ3DRmAtQ9d/uZFXR7zWqN6YWoK1hb5tmzs5nKqMkwpGxQmIvNC4/g7Zv
cPesd5+1bx1Ix1qZdQYBvVCCmp38s04GuTjz2W4OaLzXkGFNmU/i2llz4OEqQEw50nAnsPtyDNta
XZEpz8seqq9/kn267vmt9NxPQ/kmMDnoBj2xZyQv0ZX2mCIUE8JjnabeefLHSW9fKjFpxo9qyV+f
MtEo8MBcXdtmJk613TvnpXi2yYjvLOiAJMmT8sIme3kSz1j0h3xTf6uBt+eT6et9BaD7w/r84pEn
bJA96sOwQ/uLp0Z+jrqkay1lslWE55vOKDE6eRqHIZ7Ktveb7m5r+98kceRJL8wvU/iwjhaOolP2
javNrOqKVj4FxAv+GATa26CigEVVjT+frfRsat/7+xjTbPIFbG2ygNATcZIIfsLQY0NQFU9rF/nA
i0utue+peEPFS0862rkFKCbR8LEk7VKEOmx5vMKSB8dxXiqISHMGhvIMxTeZvhECBYAf3zuV4VjV
uXrKDFyH6bXtJfNnXcL3uggpLcIiofZ4UdWZTDghWUF8YEqszP+EUD9uftS6gCFTK225efXDmpiC
XyXy+3UoGghQtIeCiTUCoqVcd0vrmLvel84K/BdBMA0vhG2sU9Fd4ffqVKo6Cx5pA3araL7oHeXX
8R5ciVTDS4+dDTwFlyddscHb1S8jx26HX3FWU8KFCRlpwtWZis6JAlCkpch/n/HTNPXX2rzuCPD1
vx7/zC4ZQsaX/XItelnp7ph+DYNhc8YV9TlxQ9OhGVQtbXyfGPIu0TxEHQ8jjfrAq3MbKqB7btMV
5Zo3CLPbrve77Cc6bu+P++AokZGL8XA48S4g9PxX/CIR0abuQu+RpYhG0llaVbcXCPGn9j2zAIGQ
A8U92giFEhyxmiyciQPQ0dKmX5YWmsEyOr/76ER6mzBsXix5TsXpjYByWc0EYwF1m+zquOMsVJU+
QUK/N3m/GORHyCR1mBy1a9THVH33Iev5AZQ+nj+cbLDvTk7MnvqXJSrt8wntPaoz54e/F4ewqaQ+
mIlDG7zge7tkfopW6g48qOte81r0BojInAqdP8Fuo9NINr+QQcZnJ6FVLg80vilRRcI99mond63J
V22c0L1eIYCTvWzpj5SyoOg6qNRCf/nBuwfoTDMlIrc+eXlv5mpxxKUcAkHx7O4zqhkVFlG0hXHj
PjCfZ2xNOKswlHrDVMILvR0f2asKfByI9+lCvtN4ql/bzeJkcthzey0ihCT3p+5DwzPxoob/bSfO
isrxPc+oMKB8Q7PjRXn964/90Sz0lKvyv6uJC9Jt2pTltguMcj0jJ2n0GEb0pQavT5rYSvpEHBA2
QzxS8+LbFNrptDTTvYrt4sdfd1L5hdEHjDp4mdXk7CZMZVQrtHJDS+Wk7YsFTl3vY9hNB/26bvjj
BCGJtjT8JWFhgzB4Ly4Q34+M19y4KZ+7L+BJovv7im4PQEUvbW+aO17sPLP1vuHWwOHI+p2FFDkG
frdmzoxwNEEgBFZkO2hw08KuEiZmTzeb+LY+++kdqi1NN0leuW0LEEYGi6/8QX/YY8XBcCKIO/1W
UycE8B4RcohtbwgVnspG+c5wCfmb2LJbVUpBi8ZmyMR1vOAh6bOxG41GdcbC9pcN23HouM8qhJs7
YhyVhq+L2I7ArnlO/w0IcwweGULjMcPunoadzHsickUCmGTawRcxpc/CsiC4p+rZEJpdm4OWGlp7
FTjNycELqlFw2QPTPySESMZjqVWtAOFzuNcATL4z5fsloK5R6jZRmcD5fyyq49P3N0k+KwX9I8Kh
Gz1dugRhaI9lUWhcOI6omxC0I9ssDLokXdNI9ZtZZFxts8rcN/ZEYJhTEMUWG2CAmMLNeOlpZ9os
Fo93K3B+8AfeOuh3BszEdvBWQEAsKglltoV2QNRiB/GFF/8sAJOIV6OTyzQi+/QYecvNDvHZj+7u
iF6OPQom0UFF62M6bO1fe7RZR8i0VtXcquqtEC2fP7g0utRK4BX22HA0+S0Ws3Wzns0Fpg/Jzxea
FYioULyx5/OzHVIyZ+7UiOYmuhaMhuvbIJavBY7UoTsPY996k2Bo86GmeXkW5RY4GB8v3djl5xQK
Ff1vhtTm0VQ9miT4fVeJyDhON2HksBRHTd9wp29VUNMKuov51HjqmDwByUOe/OY/w5MnEg+bX8Eo
7/BkeUWhVWVIVjY469PMxSAZTfGF49UdYOZcc+zVgXqgZbcWAUa8KK3m60PAnhOiMyw2has6Lmim
HsabOdKSjRiaIv8QRVSgSCuiwOI2brpdmeuJn5f0vRnx05JWKdbvQ8+oeWau7bxWjXviquXXo3Yw
CvO9T76a4UmorahTMXNn748vAIr5SDsTl8PVWBDKe7DBhT70xHcxxxfP+m4UAGOGi/J8WonBH23C
Bo15kjzRvDxsja1IJCBSu7RpI7jUH/Cuh22At9SvEvL3evOW/AO5tkuoatzkgAb2oAsxJ2MsSo0C
OUJWI9abR1e6JO9edIHwPhFdvbhOwLm75trzMJX/aKu47FUc3c1QM53IbHLi4f/nsw73gWM+fsTd
tTZ/FYFroQa4GArat3Wo3QonjY3Y45J4IgUoVBk9YH8wk8NrXgtmZtqUqODFE44zzg4jLeyXN3xP
Ac14T4j41amzJAEkTC/gqxXdaeaJFt1kW2TNfTW4KG3oMy2UVhQDV+zQzSKviOFp9PrTmR+knrOU
bRXLi8KVBS+/EOgy88SxvcB6mD2wHbyoM7ZtveGC3tW6M0+TQDrRbAa6900ugPhpMTaZYL4BwVkh
y1fSkjysyST/WQCdvSQ9ePAJD8Y0bJEepvP5tFP6byv+0HHf+z5D0sqAr0fqLJNL/mODXal5zby7
9j+gnVzOWTqEZZauFEpdrDWkvWAyIj82czPK6lwPzdrQJSNWZCH6XCWWhgfOp6dK7AAZV97eAMsC
p4wFquld9kOpAw4/pQ/3nsmWcr6+vlno2V9w3Eh98ftkpYk66IPunZ7Z7oLuDnlxXEPJCG0v5n7I
EDCKABpMuc3HUrs8NOMeCwZM4Fw74UMB9N9RJ7KGDoMV2OZ4vqsTNig0XDZiz1aFtCj9VWWuFq0L
3r4e0Y2vwsIj6AAaZhbPBekxiTro7d6o18SzH77K2C5Nhh51x7TmyXOBXgSGLmftdZGPGLTLPlou
4oEYUjDgJFC4YMGjqZGcqa9uOZWnpuJFFbbUFXznA6risLrGXj1ei+rmqX384R7YGar3fJlJZ6RC
tYPWE+pHLSSTkvb3SU/4xzmclCbB6dzGasrnB/uLr+ihQV2gy2onNvIwdgLAX8tiz9j5Yr0ARZcc
szJKQaM7PW49/xQU5L/afjZ31wyiqIbCsRSWlRjlEw+wI3aV5FXDm8TS+WALDSxdnpW7vs0lqI9a
+UGXscYHf5Bt5+Ll3WAnx+diZmHrpkmYAGl6vxhTUyZXJ7AVgoH5CFFZmhoDmTTW02wJrMKMOKD0
xWVkw+3RJvRmM/gYs1olx2KFO5LhFrEIc2G9pIMv4fJQryFzFmKxfplnJP/R8AmtTp4HvyW4zK0O
/cUGSz38Ak8EoAv59qAYq7gufWuayAaROuASJ+uE9tArVSpaErCJ4tLMosrSTxrfWD/QxS3l96rR
PfnCRL1X0eqIgEJHiS0I6BDX1EKGHNrfeEeSO0I92J2GqGjryixevsJjVNGLNqWlOJwinHvwTqWh
hiuIu9Eo0jDXmYecr+Bi+CZ0mmZVF1oj4fMIfTIWWeD26iNtKmRGWQCXPGZet1F+YqYmOgxxV1Mj
pAFBgaaFTPR0fV/w5/xbrxt60TXuMBWhunncFUhhsW/4t9Z7Xej3RUhmzJpY83PmLy5SiQskqpPg
qcthqa3tpW+4gHCQQsl4gcfErrPSugMF1x+No0zP7QGBQDx43K66pbq9R1D3vQYnrbdUD3c47bdT
r87lqfKSqITKgiuEP2QU7c+ClzUYfI/9jdaRiD/ou89Auro9orHz7eEk7ugQCzMMFe+Hxl4iWVEH
CVxMpnvhuMIBv9LyguZ5nOJEX2O8kvQ+EzGCmVB3AhR0qtskfckzK2ffbO+F5MWJ+yxQN/qTCjnH
ikJLH7qh5qylBt3IpEViXfEUzh15D3+Sk0j4XdVnFbLLUfcPCobqq8nfcy2jFa5iwpbJwffVu4F+
OQ9F7J1i7Rq6cx7vLP+inVXXpO9Vgc1ciG+YXBCH39ue0qaKjDWvZL+9qz8PBvgV7TJvDJH/JKz4
hhocjn647Bxmw3DrvNnM75omzL7se6MV6FJ15eknXPW4FG9KlOGM8bvnRGeaejDUPw1rFoBzCwI2
FyHYcZgOdk1mXNMlgt7M80+pfYhGOwWwVO0dlGD/Pv3FPtwUtvK6n8DZMTHFMGEWclZAFy9ctfrY
PCC8/Eeun6MdKUfcFkbTISZKvMxPVN6W2BaGNN1SNYmoBA9iZigLTwVDj5dWKOYm/6Hr83jPnKDL
D5tsXUpYaO3w6/HU80GYJ9xJ/2kC9GAekGTW/XSBLssJWJLMopfunLykdjkysnEeo7GcwTHQn+LP
dVX85ermfCkTphtsYzoHieihDyiSpNfAxlsEAN88NiOnAIKu0SljJYsHW7MGIMG8RcFl0r1fjMr7
05hVHBv0lE+XhOy7uSiaoDudsToqPmkqbCmc84pca08NRB+uvTNI4aqPWphLi1Xi/hlwp9LyJqbz
9Dblfl5f4tKa0bHp3gXHKcPQ3239Owd4U1FQrIaMq3j0OHMT8wQ90agsJivdcc3yl6/2G/R3J1H6
yPvWMhofMd2plQ5VOwY65DGgJAfROAJJ/m92s+hUMH13y2UnNUoWad9yvXPf5pE22o6O6Cfp3g4y
0xW7/+kqRONP+KPX+Z9JMQz/ZkoHdQBF4fID+P4wQCk/sdtiMZKZJBx2tsWoHivCt8bFvKslOWQc
hlCJsQrN6sAhlaGF+JzZ7rP3jhTdCxC3t2SPLzwyJ2vrsKtwra2HxxgS8iT/+evHy5YZKz1cZES3
mRad1HVvkuEiYIGpsAPSOLfL17o9CeH8LAQvAQ7Z8pZzdzUa7cDpsRnH6esYZkyyLBxrkgYaDS35
MleT5optZiUBUHlMlHjonw+CGJ+uaviI3pcAv4OjqZwfa9pQxpUil/mMxlZI00egLjVt9an2wZiW
C2ENnAIneiSCYzsuqlA5EH83ZT9z7xDAqHnQTtF2KGxSeqIhWCT5/jv7q+ZSniAttPg80VTtHFXx
NJa1mTW2DgrLK5RlQmTws/C0yiJwgIbo2q7Bqsx7LBcRpvAcNAuq2TO1ycIcwD8/lWMpWJz3XPu5
otJVHwUoSZtNNVIkjwMBotrkxl1HKjfIzIsqHe0Mq69QxuB0U8OzBHc/bc+16NNaxHr4WNewOBgZ
f1hB/Oreh+z/m8CGa4ngsc1b/LbEtD11NuDNtw+F4CyRpUd+XmiUVZlIlQjiFFp+8eZB6qvxnXwG
wbR5S2uiQeaiS2LUbH24mn4q8sBRuIojUP12hncLqrHcRC4YbmE8mxjYw+/4E3sHG0jXSOI8Zg8d
xgQUO7w92HR9nzsLbDPTMRygA3qdWh37SHVDee0BoFUdL/LiAVtexPdzv4Q2dzgPutT4ATStiDyx
GYHQW/RYlvSfFB4GsfQ3w4aEfNeId5z7xzhcLLGNoksQeXqGV77Ud2eF1OVbTZvDPI6eqPAKwBY+
+oV5L59mtyKhpURyTumCck015lSNziD1ZDGLMrN+WLAvXTeFo0IRKqIkWTIFrmm68kla0whhE0tl
ogFQwJEa3PtJIKclJaZK47CX5GgmjUYiB5JQ2JJfGSme5qkYwh6phDPkIhaA+c0SVDi3JEjZPgb0
1V6COOZX4QAnO67xgZjg7CKpkB7sJYOWcN1VJlCW1Ddr+QEkHTSuiL8/hDIPwn8CObkNNnnh9swx
ufb0d68HTqJvu3/bARkhkaNOuw2aOr/LwgvjQTBLwAqVpy4aE2cKBqEOAyw2+Zhb0GRCZlxZiSTn
WKAYfDnKZgq0rJVW6YSP+JkqXni1ds1OEHRgL9+iqaO0l5SgtGP2aL3qTcPkV6Cmq3O6NFDU5SQc
popWOUvcZtclhIr1tpYIUp9zeq5Z2td0quXKqYiyKvIxN6u6YJ/YccT3pA18v97xrC5Y0qYNWiHN
SREe3enn9UQVaQQXbgA2CYkG08flrChUkzNS6AbhyI5TEiZ3YNoTwVV/Gb2ZZcrS5HDupEEieyE1
XKL7N8mVp/PEnXX+ZFDgMH3HmsBh3BBBRK0AtOLHadvE63+jDCD2bVOGq2iWCq/T9PRufTaPjX6x
txza+WwlGmSyUIxcVAs+pOtj9WpIuPIGPxuB2MAFLyzVIGuo3RpPlqxLYcO9WWPteYbxbj8Pr2nD
P2A85JBOmRzKGOG5964+HhY8MQPkBskQQr+yg2Jt2K9OOGAEZRWjYStAAIUlZYVM6uTXlid9MtWa
2mztrhfV6gFwmMNxSREXQ9A2NcYT/gxGJ8nZUTFNl1Ya4Y+lVMdYSJH80h83lMELi9moHFgNbN2v
PchFQWcea0x/aKQF5fNm2Ed9KlDpPMMKCc9ubEBE09xqPEqE4TeVcILAwSz9eTH1Vhevj0p0pFs0
EgZR5JsfnGRCO/PqXBbBRbmybyKvHMftrjOntv65iMJGUMMephWebb7NnjwK1nc76qXsDky9o45N
71TxdS5AVNaVHFn+i/Mp+RsSx4abyvP9FFCFpXVhdRRaizxNqCxLTN792Sd+ogsRqQMqQzrKrrkA
hKt55S9xuCVf46y100Mto7VeK/zzM4sloLZ+0lKVJH2PDmR6i7RidjQifDIld3JRQYRlrjUdbgHN
k+XQ7slvehACA9l8RiXgaVCD8e2/1ndIqB1u7nvvVKWB756wju/TKOVVXY9dwtcSLseBBVvXAE1n
Ge3FRc+TJHOlyHv5sQTbwFD6j50QTP/dM+lgrcq5ZS5oeMkEnSYlWdcqjbBwIKXdkcxrOCR6HtVf
7oXsoRzh84z3WrQ3MKH+/YIANKvig1jYAEbps7kssYvYNaN1MtZO6FlHAbgo+IP4dc6SlmdA0SGJ
Tjtr9AnIZuMQ2Q2cGcHf5h+YA8yf6zAghdsrvdGna8NYQGSOppvxmMunEOmSowBpmSG5oUrjDYhR
yoykuI9kNkeZdzqQW01Q+3g5sv0KI4Uyoasl5JcvLGTe8s+jUy9A63XH8BNY48vqqo4UXltnfwmc
/tdO7CJ52bwFHH0gwRvaQK8VSDlJMCE2pNCupSH8t1Ph59HIptDKTQU+lTN93D+1a3Om3RUIP61I
U2UaBxoBVXUjq+gsX4e2CuDAqWLRFcofSYFiHQs1ZDCUXsQZIioLgxGOQ68uYz++H16yx4tFnlUS
KvTMJ6f88vPTw/yRkQW1/yxgx9xUEwj3yMT4nZChciNGadpwx2uilx2BN445bfeVeUxzL91UM/U9
xC+Y4u8ljusPN8hcjVyquX0RFzFGEzoKq4Vk1MMRdu+LrbByqGbID5++BNcdgqRvtXkjKeUa2vyG
XMPWVut8aEVGHPDikxTBLX5fdC4X3LqYsBEGWq5v6vNtmJKSAgli7VGjdu+w8V1x9QXHMxbIblk5
ibO+hiYdoRMn4N4qQHbvOFhKP03WFoLSJGzyhXsZPc+6GLBV2MzqKpoYUcLMvCQd8Ysxo5VcgJwD
vMc/MfrRRMMyIVf2c66SIEo+UkkNgYG+Ba7FIo+37iod10qicFl/kymWhF0vicmSo6A2jjl01XB1
WNFY0t4zZuGihbUoTqr3xIlnPMrydLjqytz2JkYuJqI2ohHR0aptmOoVFvUzpjJlSoGBkyonR1Fn
5/WiUmw2dLPxHb0pZPr1WpBEBWYECWetq9drHhZjLCt0YJCkpAYW2bB0Yp5B852kEujgPbTCjauq
CCHSXo1oLkuk89zcFlYyd0N1Lx5/uV2QM7ZnkVN4PaOUK7DKK9C4tBse4bAjbFUOr4jHkBX0easg
YUJAwrwC7NKZU+SV09FJDm50KLR0c5mJDAnP07rJKGJtUQ2PWm0MqTJvAoDAQxCvw4Lj20RX7ih1
J5URhHYg8LXITF0V0JXKlPdlOlLBXeomRkUCn2ciC81Yi89rkE3YHHEDXouVCVA7kAqJ92zXhJbq
Lkdv5aY1KQRVrWJSGJMO4LuMkrquv0xesYsFH8+6R4Z7eIFIJ/+zVYk+ab9lYd22+MA2wfIkagsN
83PMJVW4qJ37g0cDE2a5mqMN+W5DvO8zjkrTXTF0ty0UloxhqeYRthMnpK6uT/6yr97DcmntTNAB
WfXnEtBZhNl8+4+ALcIgld/0eTZJw+ut0UvZuLYRU0SaWP4ZScTX0PdTyeHZeRFR5a7CBGKyFSjh
aGqZxbl9Cd43BQdZFOwOYDF0a6okZ5EZaGUSBpulUbHCDvzljd2nYLfPgATt+o7mZIzzYE7wdxe7
5fIMlzqIeZzfWX6BVXXUdTbCHSuwKp1iGWZJvWp3rVeqyL5+XgoPebFlT6oKgfi4KGMeZ0T2JQTS
29tUMANhtqrGLefchrSyEfssSnam/t/rHHzuph3VkGMzj85ORDBh0gNRz/nWpC8o58Mns4j6dOXO
GdQMb7QBpZDj4wclW1TLUW41zc4xnM1TYHkjAm+Ug1jNN3orh2Ta7TA5hkl0T1TntsydO9Qis8Q0
U2cbQl/b06nKFVZYvlz7Li7Jfu+BGzT0gmki4Ya2ChzpUfq/gY6TttpEo1hNKvvK4MTQoWhLP+BF
h8510+W8j310Ta2sNzvCpGTtXb3bqND6l1lBBGrBp/G2dVA+eVKbwisIpcjqnNiD71HN32gYX0pN
8iq7i0iKFvMgL6mgFH9Nk9FlUvoLXD1eWyon6PD0JZTdDWt+XECbRTOQICIKJB69e/OyvfFFHV0Q
ct/hCE77as/j50gmu6kXJUHRebP+r6xoPabsXjYSlbFlMwj+qev+EpRZHesP5tNjvAEP6yaqJ0lX
5W8BYSliOWXhJ91gyhWv+G+OaQexgQr+tZOnPCvtPJqreICpM8leqDhNo2JzX/aCdEE5bhRDGj3v
G7h6QNfi+kJLuInc/sdvKlatZQj2NysYy5hP3/X+Iugm8CLkl0X4CwF/ISyAcqBxM0bvEy1gHfEA
V5jVFhjxo7m20XuB2c87ZQUNh1YQ7YW5WJ6BxkLZTeVhm0k6EIJWoOpExJ0+HWJMnaXwWv+RYrGb
ZKlmsuMDx03SL43XUw2HLz340vYIXOES7Akv/gJAHVUNJLI0kadog4yHxg0omdN/rcX/I+/jKe1V
1bAAV3ZyurW1OrRAdGFw3LyKNHvtmaAgnP04I4JRLk77yPw3Pg6tNyJfJFmy+3o6asUwo3HFZQTk
g0WOc6KAhiQN27b3EVb+pmpIuKJQ0tRFUlHOz6ihwZgf4+m6fphl6IEkhdugXvI9b/kgRZRLC2xv
/djoC/ClkAdu32mOxGnDwcyWbgDkdS2b0gbEMMlrfnS8m3MvUIjmuUIFh6qc3h1M1xiqN+2x9GTS
PtTDg7Zwq1hxdLDo8wwEBm3rBbCz+iFDKb8elku73lvzrCwTBGF4v37c1zbhG/qxrjKmxroNorXp
hiQ/aMJfzRmvwihg7zNKappq0ctSQFDoSN6jDQA563I/wxpcOWMLXEudYpSJ7eHXpoSZ2f7vSuiz
tKK9g8aPP8oAEosb271NNDIHfklIGH6EjHTJmeDfMoosc7JuOL+1xp1GBD6eolQTwMHsQK0w11lB
EhMW4eSqquwgQ58yZxEWnlZ4/gxPhLfRZOWkmDcbeX/2VPO9LoqEvqQYuMFmnkfXk124tWRs0MaI
L3MCxjm2mcaXOL8BaMaaDHuiNbZxH1jpYQMBqd4dG15kQfPhxMK0UOWmTjHqyL6kHjJtD0tnP2oB
WvDbQ1Ejfvqsj7X5JN/GLN1CEB56s1ss4F6OhkVfglm8VNPbgttGaziYkqp8PQ8fuNlwCU0A4Jsa
NG01+cW2L18P6gnvN4OS8anBply3aw8lQIjepJxje53szdv7lmf0QKa8dPaG5FjyNESefI8A589X
DONyccux/UZaYxufIR6/YXuSZBkIIMV8mVyd3Yi1h4gn/RoDpv16Tm+RkyYNxUPko3eyDoE9iBIZ
MTDPxWf91NgHvxS263z6vVaJt5TAsSucfthbIX+3ZMMDoj+lzRNmtrVJQDzUyhheY71Qh1ICDk3e
cReW8WC+NmbbuQPOver9tRuwwsFLhyOrRqgf9IvTOx6ySNvLAg4dhw1SzYJ9XgXvqqpAfs0xN8tb
qM0jZ73TR7nEswkI07Wq9juC5Kkwq7evF1sDsHwEjvExyC9fq0JIQPGTravG4qzpas2MVEFwFUzT
feYb5E5r18Vx5Y/OJzneFYFgH34AqN+mk10AyPqeZTLS6I9LhtcYYxY0VE62YPpO53JUOG+MetGW
QK4f2y3cdICFmWheZsl17Xxt+0LNEnVti9sJO/Ez7rfMprjDKXepjLKcgvhJFZIjwyrPA+AIwNm9
T1K65fBHcmLqH2zYVfw7fh7QbHZnOyXN2lT4EMU7ArR+KV4GbFDa33/sKtqEJLlNbc4oWTvmWdwu
TnwjOO2OXWL+EUU3lF594gRb9BaXCnhCuwHgg6qukNxjxrtrN7sUEWRUHQwR5pQaeWDdA/LKiMWi
Y/hZG0TOeZ5wtABN5Nl+sE46OVLaZxYC/emS1GDFQdg7WTg60qHk/5V6ZpVoTGitpu9b1FSfGlK1
2blIh04nut0DCAazEkvUjEINi44X23wPOxIVGfHDemgH0VnISECI65XJeWZ33AoM2dSVHS3W//XX
LIL2l9OgqJQ2NCBIPLIMLZq4WRWi/9bzPtBDzDJH21G3Aucv25ipVQMgCIMC7E0NpiC9zu+1DTxk
5YOvwv7/KgVz6ZJbkmLkeI9ojzOGDAUm48tFIr3dIH6yMNz1cofkTLjTdAckNZAtesYVA2OmaAqD
Ee6FD/+6CLCMmSNCZxH1H+liFmqyO/4iCLx6aDJFqDVX+XcDMBKSZK1kafk+t5kEUdP2dKXG/vYY
+cmpgRfFZe+svAujn+1BjLTq2jsbv4DMLUDhbeuiSZ0+IFptBU3+f9KlpF4NaheMhuEbIhhhEElH
3NAPctT2x4bvgvCbiFW8LwPvBeVwTMSX8a2EVk9OF5aqrl+WaTg9usdoCHWwdNICVFdth5HeRTkl
+0EtsIbZ9yOPmIWa1T5cQw1ro9vs+wnMGO37TSeTiUHyK47v2WvvSiksZaRtu9kvPkWxt+lltu/a
ZHjCGu7+Xr46Q+UROJAARx1vNc8QQ86f26Ur4H00WJB0jxyogf+veZP15nyjjjJYlwYJjX4z5AvV
/R0QBV6fALRb3hYax6pArU9pfNaR0jnjEfM+CfSt5y8dllaTYM3A/qVEXO5ENS1OHyKbyq6SW37d
N/rB5x+cIpMpFSMoeQv4uu3h7DPgC5Fmo3GiIFXUHYDA1jOLygCOayYiC1x50f1ai8+RwHyUaVaK
Yf8JwyoXcQdSEpExpJlFGqBeK5ij8G+kqEYHCeIGE+L3Xdvd6clJV4Nrmk0XyVNokpazqkTuKIqu
BFAZp5EDGO2bFgLkBBpkt2pVxJc7Xw+uM/0aarV9QLPBkLikIjgC8H+Az9OVWAJ7nsF+ANA6ckqR
9iroI9DipVuxOhETtCavhmHheBLz7RbOvgmHzVrhQVG6ryr2FxMRtBGXCmbE0Z8QfdT2giVYnwfb
+ajN29Qv7t3nT+4TwiTTTMZdHROK2CU7ILNGwST6WhpO0WZcHK9VcN4J4OvYokG+LNY8eyVr2YQh
EuGOnEERvDTikUqBbuVS1OiXYM7dcd1Qk3sLW/tr1aK6y/icUCUinZhQUBFC3ExfSoCYTjdiyKq1
TegEm8ddO1Ef+J/uKwb58oAnTCkd9G583VB52nxw9nRhEPaNT8rXF8exJEhkLFcIKg9lbLzdNAhT
gdaEjzKXHyZNRHdjY0G6pdnUrx8hStuzLyZcG2l8kiTob5eCC9Y4iwZM57Z3bBwHTYFlYr8E+0X4
fVE1er2qg2D7dkfDV7aysGJQ3qYRN+mS5B53dkCc2jCqGdFcpIBoo2Yl/JTKK93JyJx+LvGjT3qK
CcY/iwfyYhIMgxpzCJ/KgcTSmfZ9qNcXfxOLlRjEcJzRK6wqEo2TEcVDaWB6pKr9bRb5Ycp4Vgar
tWaDr9yhdE+TtqsSSEA3FwpQ0YR4vI/V3bjgOa68jx70k8gTylu3yZhTxaa53GAfNrdmNwDNG9Ox
W3OnoXgz1CHkhDewK8CVxuo46sfF8HbPivmyd+0uf23FsIEh6lDsf4zAe4SwzEKluMO2NXqf7OnM
cucTMAxpEqWAIGge+/qCEkd12hjp/o+mhZEwknfBLIkrz0O9YeSxyCs6gma+szPjcpqicgYexk0Y
3K6F6Pd3tTFYkLOl66o2wje2vwACW2eF6WbH+Ks2RC03nMjdvhOpWvUtEVpdxBfJexp3flcH9F1e
7/IvQz5M6/pybCy7h/rBGQn4z9HAQtWPOjapnkxhWq33yY+jH1OQfrbZJau/TYYkiaYiBwfy4LtM
rWE6XWodCyoQ6x6KB0CiCzpbXHGrU3N8+amFyZdle43369y8z52Tgh84qIUThwR6AjaNaO4ncpeX
an/g5HPQQoDXUh+ixYf3IoFJ9BHkH7lvF4cOy4dTHm0UJX+iRrIHWfOQ5/6eYr0gD1tE/KaYTWeS
bydMTgq3jDr/kqg4Mecjwix7BXL55mg1SV8fGMwiNde94vJZGARGnawYi1m/pqKZBMlb0j+gVLCm
Tj46QXgqwEXB51qd3eru5iPqQiTb/gN0J55h8HujWu721z9FcPTWSNLqIM0Ie0BLIC7DTCv/hGy2
JJ0Ppr5O5oYywRe1HTNCMktB0JVN+YHy52R6WQt4Hyvcn3bx3A54yV7OH6IuseI00CMMxTocqpfl
8p39DazGFW+NG1U9f1fg19DCEtmgXQO7W1BG21ul/fk/BVaEHAQv5Lr0EHfQL8FHo9BSMCssSI1R
q4Q05gHkdDsmXqnofvaySU1p8ws+Q7hwu/da2hZy34Qb/2o50ea6ojI1MEDR22TGjgVvxVXOu2dE
HM/x+udrlYrfbPn7itLxzls68d2/zS4NdYmh3lfDbfEyFx5cALO3NX1nJrPaPBQkbrL/49cIuIAD
go2OCH/V2J8yXTl8KxT4xSPyi8f+qDOa/D0C+pXDZJn0q5P/b10QUNOvgRoMgibNL9S3n5bJccCC
tnkkOVgVH6lH+iJrtiqI+spwuvU0OSeJTQMsiXqrMozMMMWaCw5NsZMVvCqumqPbG4LBSFnBCu0D
7CAxpHlMcYtlOCvQ2ozpgcUbcqky9rjZRMZ2tdUa2cylkrFfdDFZM5zNM0EjHXItf897JygzQOvy
gMidp6G1QoV0Z3V2SL2cPbmcz/8rROatFutGXjDu8qvqS1eN1+yelfVeWKZH7RY34c4IInUTamOS
nfmEjG36CObU0XgXsdx/xcbgA75PFBtLNB2nlv1jztrhMblLx7IHltSs+7PToAu6cEpOWOjC6dpl
2wkg4qJctdGjPi6aD4wijGSI2PcKmTrA1aWZHkk8l9f/cEKQ88jXTEIlwXxM80T1eX99WmNYp6Ji
yd3k/WlinI4aeSGnT+LcB81ROjhU8+7Z+zGWVE8JQTWxj5kHhr3SXZSnngtetfev/5kfFqMu3H0K
IiLTuTfENoKViFM6c6CRTVtCMnnmbOwQRnlXLH9mtjODXHW/qqr5hCgT7JqjuTw/Yq3W/lBWTDxt
D3ja4CwAWWZufuFtZmLVdaP0XvphBvEo0j90YlqND+V9eLG8KMOi0EyW3UiiyJm8jERCUqv87H6v
NjoWP6cX0E6NstrdkZLnQ5JAQJbJ1X4JRNlSXHZoeBASkuzv/DhRAENgV4oE+7LkiHJdwOTAcADO
te1fyjFVcUM/OuJ3hxJm8DyAcvGw0Dpw7fTc1OMqn4j6tix3MCW7P9vOU1Pd94vGqqJVbrv4qX55
p/zmo68cNVAKSOEQ6R0bZdFMca46UUda0bdrZKQ1uZ4ZLKQ1hoZjfMVDq/PeRz+o9zipLYP7+2K/
97E8tt0fSwxF3g3DVRVLnwGfqy65fqoYf6glt0CueCpdJH8p/XCgIL7vfSf4aV0l10/wFw5DLUNI
Dogku6Y815Eiaxslv6lIzu+Owl3L0ywEj/vhEvj8R89OpOdGHz6kEhoysK2UFSGKVJvNA3vJJI6M
PqUe+gXm1wGnd3twAGrXv3rbaj+px3amlipcWF+n/zD5jRn/eDYnsXn2TFdpQCmg4vs8DH4ZnwNw
UzIIzTKKxOztnZI3RN87l/NOjDhft4wGINjVYlk3xP0DK/sASs5/1x6ZW+lkGLn/jdWZlLs7qF2H
u2cR0km2tDVymb+0i2f/uS4WmkKXXMoUfDLWm3ZyN0ZYojmh4abiMaNGb3xCJULzVMOieOTXDfx3
lwlGRhLE+fyC+GWZVvLENyE0R5zD409qJIzG6rd0Y/8gFJWXQkEPoZ/9s8CRVViTtt03op02pCpU
UitLjZUwnmp9EEIVEcdFos21MfXKZ1gF7eZO0+8z24XZzxAXTQqwf8YadKzhjUSooMsTj17t0KVC
an7L9jGBF6D9Npu5o0vuDfs8TsQ9aKeK2ef6G28Cz7EqKfs+fza8WzdnCOngIbneSf+VzYqo50Rl
GN0fD//LEJJaeeAmdEtWg3ope13KY/AzSI+9p9UODsqiuNkEPyneMhuBFE7ch8vmXD6Ej4EtTHm6
wFTSkq9VB6KUpv/aUrKo0WHsPas4wbdgkItBMkvNl5eMkAZ1LPWLQ6yo7Rg9XCElWtfMjcW0QKRM
jPJjzd4bjLYkQKy6rfeRowBj799HujDEmy7c9XLBZEWHeqhA2s6dz/Irs0/s8CWEjmR534GExXPk
w6wPyFFyymuoiwstacCacQduzS6d6vWVurmX/GYrNQi8AhpnBAGUpN1XQ1Xw6f662f8EA1Z5/wlv
m41i8VvFTeEWV6WQx7OOBxKDV41dF8sIKjNC81Sg3FF+AKLfABA69K5gpl2QrHnA0ha0sqz4L4cA
gPKC0yoejClDv3yuGzEMpU2vkEjPUG1rEekPV/MKVcCGx5YRJuBbNCVkA78xiSA8Gh6VlM4rbSNG
dVQo/eQv+u0aLIw2oTK3yGwf2nj1C1US9cqIMN7GJSPMEk/EdGZhoGM3zjwQj9yfk6ejZeVosi9O
4+t8Q5vXmkY14szvNdBcChlMGRC0G517EkY0ZC1TsyPB1UBcvGQRQMLR0g7+XznF0ORjeoCx6/M9
jsKyf7+NbidNmKWGZbiVgitkCPRAx2vR7wwChQOSV03iBZiU4Mk4iWX51RJO3qmAarDfRuIicxTv
fMcIrseUZH/jRG/DaimCfN9EmgLLYRfzU/mabCPajTRbBrViNX6yknPNO3JIHf1AyyR739qiO3U9
3pndsJsHidR+83iPtP9rwV2Zx3lFLnEQlNzcMC0ugX00OIAftSta084z9R1P9A/HA0d4JGqtnXDg
58REqMxQcrLCuMtkJhvA8lLbGIPn9mHfcMgKUKiU/dqbGZNqpjqMJU3iEZpwOhPLVH1+l6AzmETJ
+vmqf5rQwdJsjMPUg/DdYviqeaQZxyW9JutzIb9NUNnpPGEZUyi8k9KPXhVGpNCdeUebbrMOeh7B
CWe6/gKMLjulLyYmOpAdCfPWjWTZgktcIcPt9Kh9SNOl7RYw2jeNJuVSmgvyATGJiP8jaLCp4139
wjPGnBzPCxrS9rJQHemKEqIH/F+H5Q8ghc2P1pwjXJRdzCThim9p+nHISnHpOTKOk1w0THbbl3/O
HG8vjgd6poPstBai9nK5jaevZirROfqqGFLg49HzuqRaSglmDfmBven4g+rcjzo3Yl0rhz0eeCiN
0cesL0rVXoygmkK+lCSZoXms0AHitIfZ19GM8/aaMisLXAZqsw5C2dq0Ghjj696KdkGijDlJg9G2
4ml+/TWuXO8H6hfoHqjKyumJ4V3HHNkrunovka+izYzsO6wX5yZq3h9SmWpR39hepruR7kJE+aQq
yZ0Hk7oihZOTZ6Rexrq/QG2fac01tbcaa/1V709KlK30EwdSPum0M5D7uH2yGKcm4FnYuoEDkUUi
xi7/ML3usF5bl6OhV6EW++/4deTZr/1NWu0K9qmoOQQZl6aIkisQprbJVbKxKMwk0++306zYcrc1
aSLNGNOx2IKtnjnlneM7H/Gu7wEuzAQ2Fr6qg2qwSMG5XIp6s/YzWbn/Jy96ZD7i4XytSjm4WFj/
pySuZYJw+jlAxLXJYAfyXJumxvgIx9xopF0ZDJimEW4EM/gfgKWKeOTXLjG7PvT0vIicnOHgT68b
56neNJJRO3S3eVzAK/loCNizpe/yNGK711A6vtC82TY5Zjw8wf5xNPwwydmFUMKxXn4P+cgCSPLm
dgS9uvARAx2CAROSbnVEB+jz93RnMGlyGKRXjW+xG8g7enSyT2m0wwoGOjCxW1wxlTste337b5AH
ahV2qgvGXCOKQGYW4OMHxBZmuljZ3eoDXXezg3niWH8gT455zSf7Jtd6UHT1Fyi7FqkBVcEHqxdh
LwQ96hwjpLb3+kL+fA7sfNrrO5TxF5FV4yiG6QMiMEa+cY93A67TfD+pKBSl3+r49sHej4bFOYkW
zWQzYNQbxgIr4Lkxx7hFbXH1PFinBtivbcGkTr7lFagSthsl8+5jhxxj/zMLKzZEhWz+e2zbpMVI
I1sf87NphHcvctT49NRkSWTHLjpJIl6H+b+oFRfkUDhH9CLNf5KjPOR8FTcyu48KAMteI+xm34Iu
46xKIQG48BH14QPfZXGLPhE2Ytg4LVMTL44neYOhf9Gpunzverg8HYSaMQKCZrN1Oo3FS6DVen23
8hU1vJpSwlg7bK0BjZHfuGIMRGnoD3uqXSH8NFQ3tfRzHkRYwJTU+RQ3jbpGYyxHffcZ+E6/m30m
cWqr7rptswntIEpv2PmqHq6NBYQDnS7NAA2wn0XLMfPeIUgCsThZDmUDGyRBTiFf/HgkKVv1GNPV
Tfufa4RYlD3ayHgHchdhKhHtlCZDRU68Hnj6J2Kn5qzN68lD0q6syK336d3Ca+q7qgcjpTDV5B13
h9bdKkrigYP2nzBBYycBjDRyF9MAfwnWI8FPqSMf3YeVgZ4IPMA2c6IQLVG79rHRcBrqEKBjCyKS
v1G0WEq1y/ZazXh/4FTlTCSu/0s1QYqunqIbwKFMFlxGme2PKppwxAu4LFA8Z7go4CqnVNythWt9
TRfuLaLRA97lsj72rS7ZljDq4wQlvBKVqDc8EnQ9oLsaKanDvNfcLGOTWkS0SRiphEjMQlhWBK1y
AE9bQKnNBVBaiz60itOIKfXKRY3Zshy24oy+M5LwGSS6Bm0aNP0hq0M71SipxbUG7WOgJ5glmWOu
KZdiRL9Zqy7J4dHoaRSRHcvQ6xV8D7+j58kCk/QtJFQOTO25gBCDbxdSlgT/2QVyauH7YL5PWQha
i1/R0Fci8IuXYW/NQxD3oNqKB9/ZQFQoCVf1sV/5oWwj7n42QsnDDCn6tOYjBwuflNZhCxkj0Zl4
nxyYmaMyQuiZeXFDonQMURRvFpaf8kLWXxZsLUQipG03oqVJJHtGJC2Fv2mm4fGJ7oA0rGw3WDWW
oU1kdfrL+7eBosFpNCzExWGRCSxvcNO+kXIoZkPB8TWzUkVRSvTZbF3LyvmFTcAleuV46mscGvtQ
FaK6deeMHKPbnAxKYjfNwsNORpQBy5zcoP0hY7mm5xnlg878KykaXB/v8VRqr8oo+T6+5PNAaNiW
LIejOj4e9GD1XBrcCgvDZbkVj0QzpGw0qOD9aIod5AQ6SMpI3W1zq3MrGdVXuxBVcp9BLZDugTaA
ujVCPkxG18tKCt9d+q4+DfZpgaB2MBYXPoA1EdQJfxoRlSnBoHA//ugbTzPb1R0e9e+VHMCaaxff
XKzuoCiN6rZw1ODkk2qGqkTP1lsuTekf6x22pQIolOEexqy4ZleIrOJ20GSVh7NzQlqdnexPLvMk
s9HbaTlAH8P1n2y2/KMjF1UmT15SRWS66GD1V7bggKsfFsgAO5ZeXIE2S82H8E/TrSfrlEMz105I
5+8bkX09/TV7kSKcyQ5gda4FTjLwWth/9E+mUUP89ShwTHhgiIf9qZri+axTz5D+k2s/Ahm6y5cI
yy3koCrkgfPZ9UchoFwMzmwkNubMaxeU6YYDeU8Dn10Ypv2GW1P9bYNkpc6Kag4K69/p2ohbojkm
Uza/wbBqcHDSqNiMaeaeX/OMgS6ScpF6toVToD+v7bEW074zAeEuWJGRQ7QbJvD614GREmmSWI+j
aVK8FYRbc5TlgAjOvfhe5kewjnHsHTB4PNIhnEbQbhO/e8ly+0f32nAH1PenU4Jl2rsMp/+qOlPc
/OoTxn+VBISGVE8j71tKMvcgpaS7oYNfVx0tVSyiPVnxo7pXQ2HMEW2e+h/cnbPXI6UCGFobSbNh
88ZZvpu7CTBUuiRRdKwX4ocv9C9uAnaIZZUW2r9PSG37ocHfdjGaR8FxDoULvxlCHLGOWfF4YG96
sLgYccCSrrj19OJc+I5uMzSbRtW2KCsOHDrlltn+6VjyMwXyJ0Ai3x5TTzPLngMjz5GZOr7sKZ1U
jrHmmQ1EHbB3GOhsiE2y5oHmc04riKHsBp1KD4xJFLt6iVVzhAd+6Q/TqjnTw7Dflvaz7glhNlGc
JaFwkRA01xOT6e9upUlxhGqXA58YKKajNbhqwZBGtmr7x8XbWEtPayxHgUkdHYuciPyG5ZlOBPym
u4DGxMDR5pnUeJ/Aps62sadri6qvlva8nTiOfOApVT/Ysa6t2X8gsGuMfTlJquhxWZjhyJiMzvN4
cY0lyN4jhNLggD+AyJOTMVvB4vL0P+Jmamzu2LZJ+dQmyGFiv55baOQ0vJ5uBCTxTvh6Lm5OyCgd
UHoQUFTWmSzTtJn3TTaqgk/XVHLM7vixoXC8DUBYdY+t/sCyuFlBhdkFh2f3GjS/Po6hunaJdZf7
u4jVO3YmnlSAWOngzl7gbrBWCrsQ5kASIn5WjRGKejTq+5qJgmOd65lkxJqV99SC0DZ/hVsNFprb
SkyO9RKb7ewI+3QOa5IhiXPQP/mMuGpxDuhQM+tr31xzsIbhyRgGpt5pE6RcrlTLge6doN6gQ22t
9P/9W+zFT59d/uk//rld/msphpVFhVSAd9Iw1ccxh+PQKbrbzAd9VI16l3boYLTbldjcbHcXyeHV
uqWJEwnc07SFfFXsd4NMjYS8SxoJAK/2QvZIw9ICKaWJmgj/xqeMlGyOlPmxer26dJykyeR2F8EO
CglVfHavsZ2gk7oiktdAq8hY3zM0tVNgXIT0m0qZWUEeEfXl88oe17YuFbOPhnkatKO/dLFIsJzO
al49dLeUrCT/fEOJpct0AuRXZIgyESBFYUs7ALj80nbxP1kotso4YBjYy+N4+7mO4wlkqtAR7HBT
OGCZdSkxgOxLMLuY7m/IyNsOSvKzjoEwLT+JXw2HTMQ2xKnhPQgaOLOHjuQ+dhG9MYC3dM4RBKZB
ZIoYCGL1cayhQzTXzz9SZCuKtAk/2ZEd4AuO1zizIc5TdG7Be9YzLslpy5FL3aIpnr87RPcuuTaI
mJdE/5lE7jD/95EoyuQhUD9HGJPASgjsByV5AEMGk/HsKLCQkD3ekhHaezZVGbU5nzNJRU82AceR
p3kMMtO440cxrdgVZv6yvOWt6pWoAh2wb+FPEvWq9V3lFuMTEWoliRWsbW3OfaZuFYTBYcsF70Jt
jApK+z0bzg0+1gdpn/ai7hDjKddjmbC1q40Z7JKnxgjeyIBD/Nehv9ADUiQdMcRXXVUCCVergOkI
BarOgvuDPX8K25bUycFY2ZjY141n4lyiQNBhSA67zBIgqa6DXiPaPhDC/EwnFg6EToopT/xl5FNF
S9yN1vBJOaKXn9KsHbEPm8r2Mzey14cFSaak4l/8nBMiEyzkVqM9ZhQuI9ytKtIGvWdnI3NRvP7S
QeMwpbXS4UBEPm6gSAy5ZxZhecuau9CX7OLxzWGfq8Yu557WKbvD/PLQ9Cw7yCyK2lCgkBbUqdWn
n8oGaVGG+2iXFKjlJxn/VpnwIS8JWOkqmubA/l6rPW7V/3lVfrxsZ/LT/vjeNP5cs3JpYSaEUIOZ
ALAPa7iDtLRR1qQZ+hgXnLF4joR+Sa/99yleczli/htTHw/vzy+XBx/MZD5nGRUWRBi+nGJFSH+N
XCQoXNygMno5EtytU4H5Qpsq9LSI8cONViwP3XMWs4EEC6oZJjmla+PTwiPbR+Q4E2qZDa4ZYMIf
/phajGSb0AKG3iuFjMv2a4Cgznrip4vdsiuZIxrwtJbWuuVULMNWYHTb9FBjtHT16MmyJOvgGZ1k
igio8I9n2KYH3GIJMU/mrYHf2PZ438Rw7hcery0dvpmDLKova9tRfYvDnvVKVCfi0X6CtMGNSPfc
HUX41X0WINAwtaB3Q0+bKgscYDNFa1ZBhuPeKVm+t/XxZ7UPMVA48Dq2ZhS/gPuU+jqPvJQ3mN91
wKtUAfzVuHtNx7F47AslkX5UYBppGkFUU9qNwHmteu7Z0NAacwuQi/drbMt9L/eAamvj9Ro+nKZS
C9bz9bEmPixDS5W9Iy2/R8b37s6eBbvtwcOiAqb2aN6iFMXsbP4ePoUo8Bzbch3zGqkVtuYLociq
gMjfz+B2pfEt4NavOJW8AQQuVqxknANFzKH6/odPIsqpkon52U+0xlmwL2d84oIdG5vBPvIltzXQ
ku+lhvIymNXz997H9kL/wKaEJzwYLBrK5rjqOUzw+tELzRt/tsN2ldnzUn1jo92B1CCEtSlPAB3r
pxFh9SgvaVJa2DXpeK+gtCLCVAQkwVJkdVLwM4SucvfugJg7JOYKlD2ZApVmNEKPkqtNFmAAReYy
1ibNS/BnZm86lBqpCDU15G6eUPiFvEF1D+jPvTkgpkgXsTgAdecupUL72kTR6k+jNtkOF6pdd65K
4Im0kFX3IUPKbnQaVmtUTC3n7tcl+V+Odaoy979xZ3i8RzyGG09zF12eDQ3JYE4AFmF7xRmUAc/7
0yHRW7gpfZLdd1SgmAR5BG6bsv3cTlTln8/Q5aVNacYSk1lqdjbtByK9WWxUEQNn4VLZuTz3dlo7
fqn6tmogt3FVTW7kTtCfSoYvWo/ucApoMjED6soYhynMRAm+a/Hndwzgy37tR1MHfKSL8L77e40P
kyl5/oMUgwThqyXleEHv1R+7UWtVX0rB4eI+iDIwmlRkI28QMCYFguCzMCUrcVbCsL8ql5RaXOVV
76GPA51JwXg0LQIYZ4g7pNLxBGJX/FgZZ3wkl2AAVELMKlnprXUY71USaUEqcUGKYHypIVvWVrpW
l631QpaBU6QP2tiXB3bDSTCXFqM1p1DSdh+CavLLWLODT0fYPxpCtjP6SfPqZ64Z+yzhOR/vgE7O
5xGUnn8H4p+W8KaasPLuOm0rMEaLtoZrVuVgGo8oVWAjSiDLgHLINEpOiLWMyI+qGxAr3UDP3WRP
vdQzdyShrioYAckmT1cjl/kkGAmmHUPye/7rO/1pREQyC4zH4jg7dpM6si4DahjlTIZ1NHc7th+c
uoTHZpcPc4X19YbsPCaIi2/Co52/R5HurR/4fGovWbt8X4uD3ERQ9nfxDYxWyaNB8vxjF8EOG2ar
qPZoy+0QdWOHaCOMiJc1zcz98dr5yJg+w0innPN8tm84L0h0+4Ze/qXLKljwkJqph76QVayYudBp
uCojOCxYPHzFgkv8se0tf+XswQFBkZMYpVI4tpvQAd/VES1VeCgA+UAZ5x0ffGyDSF248x/ntvOz
iHc3LbxumX5K3JigQYN1rVnJkfU8s1v8wqq14Ls0dFFy13LIFUGQNsNIMQed8cgzHznzNQ5qmaM6
8mbCEtrZzGATXt5Z/POrBHok6H+i/I/G8TZCKUwIbeIn1UqN+JajD09omb4P4C3bvm+pOCjjmwMS
6y3frQyDNHLPPjoxajOEhlmHhJYicJ0Y4w5HB/cdDotlXeR87B5zMpsPO1aAbUOt/Jwrq2oluIon
KmY3FNnU8cT+Dtr3YCnsilJWRXtuyApkaXQNdL/v+6EiXpi7O0luN/BEDe/lmtkl30Z9LpxMtXHe
6aaW0+zES2FjvRbdl03MG138WGJI8p/Pa0o+u7fP3/w7i/N0CNIOcr9VNd+OZpvTmm2Bi9uUy/FU
QpXhkUZNxl4eS/31ZVllLnciNDtp5mV5ArvE/fegh7bebpChpBOSFYe8sVD3JYFE2wn5bZ652Do6
z7zsJJ2nFdmGv0obZzWyNT5BDMqYAboXLPU79Ln6xfrqei/ZVmzXxanrgKQ34eqHcaw2v889QMLi
lTMec30GhDaloP2wia6m68uQqJSEMxONOqaRC4dUxo3erVb5VqNyjE7E7bPZqmCurbOlmFJAwE2a
irmYHKi5+JgEk78SL0byhTbRTvBGLcx2s5al8/RXNMWD9L8rtbIlhPA0HZRavNetrCNa69X041F5
hxxPjiChUdPYZ6tYU0lsIr7O0GNbWz+7RSF2iZ0Frgml97+9dCnOdcfCEvFIgcQpuVAg4DaaLL2z
l3DcTOZmYIs2RxbyiCIM9wKC+reOTJjKC8rf1l0oUXLLDtcoSvufS3u/EY2YaMDbv4Avv1p4kO8q
JO3EEwGdznErEb+yMUhkarW9LJYarCFnyQqaq/eSleaWeiBRleFvE4tVHulGDlWcpva1+CNK2S62
mQhKNwfXjgfmzoBgU1zAXrCgnmAPJYWImtChdabFcPWrK4IQ4oCE4H17UVKldEtQO9XXVOi2/xV8
4c3hFYqumFy20LD+quUuBXaTAmPBiiAYk83qeeWmhZb02E1tYjUDhtrmcwi+r4GiI+7ZKEFivSKN
2baVSQv8IwQY+QUEPllhlRtoB3QVx4Zu8j8OOEKUKv2IM8mWriVHMwyU6MAzNkFWgVvfu3ApxPB3
mDOqZnGEx7PJHYl9chtQMH+BBoWE6nBu6w+RTCjxOissqzSdWnel+zHWyqTt7NMDtaCF6j777ad9
OIirsL7ENGTA2xGL2zgfgNLo1hT8EAp9s8/xgNPyT5Nn9fudrIzgZfaaloyNxNKg5LJkujXnxb3y
6urm/UJ0dI8MuLk6efJDQHQHu0I4vVIG8MwYqKkQYqIRgrj5cSccdcWBLYQr8qSzdWGDLKrOH+eS
IP36d7VA2nDYVIi6LKq00Do+7l3W6VzeaLqOjbCcpAYpY58GtFuGWDjfb86x1NS0QSA7+b1N7+Za
Y+ZwaFfHHhZwSU0YN1hlVIHR97pVkhTNheObzX6/kPb9jE4wG23OBc2fha8lvieUB4s2anTIYi32
Clvn9ob8Yu4+bKYOElFTD45eXNC/SILozmvU0RP/W08rExjb3bGnWZi9haS51eP55zO/72vd4DtW
9v0czlRAjEWzgv9ZlrtGAkvUxhmYm/AnjSypukX9CK+48bVFeEdfWOyaOmy7F2Xf4JpnoA6NhYYv
cT6aPXqFB5BRC9eLKEpA2u7wcqNpFJMZ55Y46+AJ8Fc5POrpFBSTF13zTxJnkgwNGFUwBa3ZUt8e
+KGkBJVRNu/tPQ+ba4en3OhCtnYsLgvV0M/XD7nGed7w/Uw6/xXabbVr4QI8lEGyx2QTMkqCUp6B
SlWL69mM/93yd5kFRmF33+vgu2nHzX/oSq1xjYD+N/89fajcY75d2u8fjC715jrzx/CygIfXW7Yn
YJg1fWIKwQMS5xTWeEWiIUH1nSNFcyH55pwnVpk+2hbdnXLb5EqBoAhf83yDnKv0vZn5ajY2ImZJ
AxM/DYal5JHPsq3BxM6iIuOHmCo1fwC2yaK2of+cjyVSUMJXXkjt3AiHnrJXeoLjAgkVdsFKCep0
jNnKWcLh26THQD/4Wtiyy3Zi8PP1oCSxJjY4tItduKQmC+ye9KUlC5z/z3UldoUFkSX01QLk6SxI
obpZi1yEkFDPelJ9kZdnTbSPe92kS9SN0b5pdGK33gP9pS7QOw0gk1CPu/kE/ydQ/RqKcfQN/LXp
ikMx0Gm+i5gz6I5npMfn6xTIc+hu44H+70uRD/pj89Rqn+wpW4gNJUzeVzxtbiKSd52trl3SqfTF
J9hOi3NW5vWTwEaMFgRuU6OCX5S8Mm74BMKz93nddLURsm/wbz7V30Bj17q+fG+F0gakSyVINB7z
GqJOpg0+CLfMi4wD7Rni+g6rrn33OBJ3u/vlZgnECG+DsTIF0I7LONZ5cUH8eyQmPxkvno8L5xpW
C2pjGzrSAAi0H98Nw4tRfEoLQYVsos6MH+Q8zsS8AyypTKprwRGdf6p9Hu9WeAo6fMZDt94/AB3Z
YgqsjdF4zhVoYehejowzS0MXT60VGOhetZBwDr+53kQUFVV/TP2An6McDQv81eVdXG4+b863uhDK
Qn1SvBj/m5yARoGHQDb6hJ2boHxcbyOyjs2xKniP8Xh9c96+c9IWFwpTuM0yAIbY/Gtnwq4OujZD
bSqx8sbprwar0HIDce8sourqJSwNxCnTH2nfNmpcWedfcKsq92JjCL3dNYA6eR6Kunvxz4eik2Zf
2mwUhE3wKCYDbc4oyU3+yz03SI79CyIArmgLd7/bFbO0woTstB0Oj3VKtIs01A2MHdEA5NXKPeFV
4aOsG9osfHKuLQ3BMpvuH/Zx4KQwR6hoTi/tjRdNJOhm9fk68Dvag4yHB6WJ8a1l8vKEgKWfcyaQ
I8GrEf+RJ5Eb4ezDsgr3ohzPBuDaZ9txjEQKsyvBrMB2a/Py0daBCioT0kajqLSQi+S6BZGfh0gm
jaP0gk0v3BxTUNzI1GfSe3sKG0lOqyiH2WrDx8AY4LhhXdmVbP6hki0eNbSW8PVRm++mi3iq3evI
NW6OSu7DfBfh2HPnHCH6Zhi96f1/lTJYn05METY3CY2kANKGUuQx/e2jJhNh53lDu5y0WWbu8rY4
HILE3O89y95MHRDGrdMQ9TbgyjYjZYG6mJN1Tu3bA4N1KKXSwlyJiyibpcMLauYa9EbvB8thljJW
8il7Sfn5UwxVUXpGyKMR7FdMVYQ9byl3f1D1AeqLluevCFYUBDOsUAyiHFOb+x+DnUNtpO7/17ii
MSYe62pR4+izl5WUuzSZAMVOq/L5EyUBKzvz9qIi8Jonm8z2sLI2zcL8dvJVN9AgiUbAh+VRVa3v
0jnopJjk+NvkpbUaaNyUupWstWUegp+e8otaCtkaxJGjQgwFASOHO7aMLkIMjVxIn/U6byjq6Fcu
T0HVEbgAL8J9x/Puj0WWm2OHaJf22vETejro+5uWQhVYq2x3hxiIaCugH3/k/udzu0B/KZ+77mRY
yxLa2FIkYzzT9uEjRyKywSE5BVCaQw7asQ9HstOVvi+SXENoxBYUqRoppfA4twqWBvSvfDAqsCX3
rDZgvjwx53tWY4JAm+nNSPpaoiM4+u3XrXTGKk2Ue8qjmwv81VPb7oinyg5t19b9zpb4KzeqcPFw
FmsI/abeTY/iNpEpqkTL42zYvKu5ObUmoIocazXtOALONypRTYJ98L8jwCZ/WOjqjt8zDH1+E622
4C6Ppy5hCL0DErA6yAhyfogXms2b72XSuBJAFKsEOzYzWeQ8ihfY8iWYcfn4DWiUyW173eBvwJ7D
F0Dv5J7B1eb8D8LH8pTP80Rpg0pw5dUJKFsyD0ueAadVN87j9sKnI3Cn25YbxZVbvYIRNEUE8Evf
26yLgrxMVnCle7COesxrUd4E0X+26yMH33XgBv0bHTCX1vIdIK6/ncuIT5Tn0Iqg39sPF0vHk1pI
e9FPtpttvdWwJR8uRzN6GT0+m43Rv5BQzv3O6yu94bBQ12IhwGfqXVUR6Yck3tJ1VV96Ad6qXUhw
rMSwba5EGTIGPPWacN/9+quxbPEI21psJHqPh7naR+fHVQj0n91//Xq/EEYVKv05u+jMHaK+uZId
mLSls+kDcOxX3kSG1mLZfpp1MXT5YdbZBQNv48YJ6bbpxfpzZTSlnJBWQemjtzrMIF6jDumly2oQ
Ex5gu1DxBjrSAToE3eYpxkdnbLK+8bQITGxFNo54V/szJ4crq14+6n1j0e2craBcw7buzBDLAPUC
G9i7YfEwSCrmHHs+jZSFHTkGTJUy6jH7AxbI4tKi1CwHBk5ux1+9rlq5F7DCYNovDSqE2v4sasNc
tCtpqgmtCuK1MkTwVUF6d5dOGibbKnjGB+yLL+3SlteeluP0Mq4FJwxek5IMMU3CYfM0iuKroloz
N7toNnzVlX2F1hEedBxdgJ63y0Jg/Kh3QTV9JFumQFJp7n1+8tDm7fgCyc2b4JciR5mRZ8y7onyc
kDHg5uqXehw9l0jMloaZLXh1zvJg6t1oBM2nmzRohpnk9Zf3Drs6KFd9g2j6Bt8QpbS/xqddmV1j
HRVzKKGAbXpRl0KNzWGno2C6y6OxCwozwWOB35oC7GZv7AOJvxuaaWLTaxvMDWlrC4a8mp1aIZcr
V4IqlszckJm1py4kDbFPHxOHb0GUg+GI2rIK8ap2G1Qe+izyp2zHxeGe2ArmpadjT/Kn/1CdwSYM
DGXTvgbE8USCXXR9TbDUi8kf+UlDw3z8Nf1pMquM0Rc7p8c1WldsjdpDaKgHS3hfdkfCxSylDKR7
EEEtu7fxu7KtxzxxwmLihETqXfZeLO+CtruTu9X7PmS86sulK/RLSHzXvtQ3KzQUT788ljHua2qq
0nm6oXvZ8Me7wCsBtI9RGTyielhS/DbNf7CetCqJhQJUDBxHYIi4s2simgbOhhTGos2W7tHUrL3p
P9YCcgPjf6WTTkUkKMXNC9sn0TbJ7hRvDhTzKPZRXvGzEVy3nd5R7p2mdLdsuH+333fu50dtMh81
RfMf/vQ+LTtNCoHorsY+c1HSjquYxKHnUnQhzlcRzgLAhhE39gMYJXPXQZfkUdNymMLyFSN2qu00
uWfHWtGuCJOmFcfYbhTGD02Z7Qui5QoeBmXDt7eoefGAUF9MxQnjY+e3f3XnYyODj9E6Twk0XQiu
pLWJm7bMiQMpPBTVW3ZaM6uadHMDtyzdph3v/GXE8k6HVlP739F2R90fRct+LFG3sne0FG6KZYYL
buAf1xmQJqOLlFrhRGO5kmiWPDET3jpNCpeSGUnsREgBNGfhX4mYcBhAv81ymXsNuWmtwRpBIp9m
QvmLi2Adp0A7JmpL7B3FK1KUvIf6EbtyRMkmw/oTvvcaZsVcFZ5Rxo+Ix1pWGBbOlU0nyr5PoEmH
q5JVQ7RKLW3eDmszqJV0k+SMw9EugofnSkZmNl5udDDA0+iSGW2+dirgM4RyvYv+MliJKpl1FFYM
ErReJdBuVs+m8oFRNbeaHLyibnajCXUyBE6sx1KLImUlLiz+3nEycmkoo6sidXiSHk+y1yAykdgN
J46L4v0uNMAT4WGhHf0B+DFjmemO+LZYncC/tLlsko+bs9JqFr0aQjdj2w6oEMdosiAPobiMxnOd
juZE3zTBo2Q9Uqylp/bUJMu1hlvREW9c/N+qPfcW3GDR+ZXbXcKhSmGT2amji4ltlJft/OYrGJq5
PyWFm+kJE9xg9HrLwyzd7MNtw6LTYJO7dB9FAyD44LWfSJBlmPrOsE+eJ3KY4en+ol4BOe7dWzAE
+4Dz0bliNsFzP0sGAFV+mydq41TGaIlnzZMt2QcGez7axyWE8IDSAiYfJgcUsF/rJD0wk2BsebQJ
d2LxJKdJKTwkeWD+ZXkDYaq1xsZGWFr6NqpNAT1Y7/yYaHGo+K3pwe1JRH3uBxEjmxdq99t+xjSj
LGEZIekfVWt41/IuDyL09GLBhXUaWH7/V48eolh7/42q2yqvOcy2cLYpo694IqJCn4g2kAqAkqeU
IhjpfRIdBP5R5ZQ9cxW33ddeAqfkBlrMCXDcuFbLLiQBQbaGeCV2yu10CZ8NsQK9JSDwviKw0y7G
id00KOC7afCTWQTsaU5UiTJB/To4+i1ZChETcwNbeqOIGNCM43Fsn2TXXsaHH2Y6ojHQgQDGWsQT
9/5FQx7xnOJF5hIe5pU7DekqMAAGPxXnm4KO6UDA9k2uo/CxmkhLKseeCXpMqDwgZmxxg76ieQKA
/68r/Z+2MTwtcU8Ke0K8jtmCDSz8rCZ3Bt6mcsD8iYkLILGXaZeIClAS7T9Wq1e7+2hVwYbdz/7i
sj2dtryLvtuuYrrfVWhQc3I3fgmiPcELHx5yWgPd5SppdvE3C9y3Nyy4NGS0oThMBLk7msYTGZRG
ua8MGLB5RmCpWHx1G72JW/kjGjyEE0bIP/09CbL0N/MXaG+S1v1RKOV9gs0p/qzOConn1kIqXgRK
p5MXxH7d80f5axc0kBSLVUdxJcCbbVF/+fkouJME6d1NxTVNA+vXYnANCUo/cXSdlMnraxQzjZjJ
s1CxmUSaRlfV0Mz78U9Eqt38ZVmrtzgNhewBp2vnXSraxduK1gCxGGyJFD0xFTiWPmmDrEIe0XFp
Dg82/zoaJ/EhCfFj8oYdXpe5fXCxWkHK8ko+oBpiOAr1W56wvU62iPljP2GKFxr0Ox4ctIjztIWo
jIAoSEilDlMmQxAlWdVqv085OR4FguGF5jlj3K14HxAuEpDnLMDyuiU8MXHIt6KH0Jl375elRaEx
07eT8AaUHsZ8pOLdiml/zuVHTvTlFAqnyKgxDmVi+w+wmAiIaTi0+9P9CSPnpCwk5vHjiypiFPzo
0flS6THLAXesCMz1mt7UZ/0kYw/UU25Jzr+ocmLTiYXnLlZnc+MVNA0hIh3hKZM2YbtyOn0JGeHW
v2fFrySM/ycF2clMKRngoHIVa8aUOgvweuVVWBrr7t8qe9neci4bbthFQqi3eANK0EtC+TOpYwG6
0vM1s5uOXBSmSPHpcH2SKV2l0oTqmmlu5iRhauPeuQoUBgfeHk4AlTFo6ZLnOyms/zor1fHtb5jK
LFLs6iK8NWFRMqESmdA4GBIY4phbHOvuam+DmWhg9NO6MBfYiR/noNM9ZUDWu/+iwQP1sM38owqw
4YzNpSnlXRUACXnwg5NjHtlxjHZx0vb5p71a/Ecqj+z1jgFzRO4ZwmJkp2t5zMEps7jAJ1Smw97c
h8HsCAUg0VTUUi4HgMLlenOq705/mxXOzDc7xVf9/s1X6j0/GAGXgWzMaWk4mSC3OYNk5ytZUvXM
Q9gT+SjMeKqR32BwRTfPLfFUzGjynNwQWjmLZOU9b8r87q1Z9Fw5juiv1jbRsI+jQZX1OW8lp2zR
UTALsbwJa+jmt9q+BawKYxgcfxbqIUFnK8P6TzjUgD9CBxpHLnFdRcKK/COMgGC0lGevGrckcG5Q
2YLSn+IjjvrsEUI8Kyh8ifpmo2Sog9KkNCsthSWzkFHdE8gCposiWt0PPDKVoribyVl4cVO/+W5H
wmaBAGENdTqRy6RWwuHewJLeMfKt21VY0YTzrQn2eXiujXc+EF8KXO1bYiVVMx680boMq5leDNDb
Y3joLWoMKUNsyuj0OWf1MOKyscYWU/2pv8G4qKycCJQRaOpt6oih9kzYk0q9NE2eJGMJ7JoO4zPK
ie8RT/36Z0fgVffMChG/dXQlYj6l+wFG7k7mUx+t8b1v3yUECDJb9NfBsiqjyaDsng6PO4Bp0BUB
gCZveDsSYvMk0AwP53Zg/VgR8yxzurGo9QxDL71BQd3Qp6QrA5mj5szlXjezEG5J0kz2bCnyv47U
R4JJLxjtG9t/h9j5gZJHutYnILFCK5DQdjUGEJK7Y5OcyZ1fcTYwgm5HxvWjauCMaKae+0AH/Kx4
PEj75JP4FjVwv8bo0b0TQwpWMcJ/qvklvl4j4YqSdolXZoorKVgRMqm+ImKQlbqU2VRYMdARtYrq
yCGDG5xuQgoaxYDCUNg5rU3oGuAG9qdNmnhHLN/8aCp/xDoJXtlRh0KxbQUppHCzQGQ7yLA5OOHV
q6+ICzP6xU1G+CByg4+msWqrLs/URKAjaxp317j/vHh03k5zjnXKRniqLjK0SMX64OpLnpF8jSaB
FeAtcvF+RVB5G7W8ArpWVeKDoJiDhMe0USQSHie0MYONlkzcz88EwUMIZ0aLo8urnK0PUtejoYhq
LFdIfGfN2LSaFjZrVXKv4w7Kp6uZUwyS/ZrBWoMhYZK+eEa99a12y69w1y+rGJjSTZ6+bWlSx/99
yjcG+GkKo38/VRBa+MJVtGsyPAE7k/hJetPAqB2fl0NjbxrWuqtARcpEDp9AAajdbtSr4uQ1yE9f
UNTJsr7PllR4MF14bknoDuDTPe+ff1J0P3qY0/g3KNiF5zcIOl1FhOi58LL9bNPzFii8cXofH3zQ
ANAnE2vUoBN3CsAn3S9gQ5Ga4n/Fmzmkv5ipLLa+yprWGTZMz3ZfNyTe/GoMEEEOJ/VYnH7431gc
hGOtsEgwY6yRF38XrKu/cW+jI9Lwf/I52IZ3vu2/wRVHvpcxF4pbYfILk7b12qgFTwPF1KJbFUBr
WWdl1SWgHcOjEHqzSv1J97v0FhC8zxA7G+Su9Kw3DCZgEp/G7USSZ5tMDQXxrp2X6dhrRnryGnL3
okmHJ5M1Bj0+QcilWDVQUEGL+PeqdLCXV/dQmN5KwR4YQwewBGEBcQqLeFkBDtHlRRejrVCl0KdZ
R/wGlMlfCI7rKobqHyriQr9mWQHqldxw8zWNGjq1KNmz/snlZyXmK2H0hu5wn3ukt2nzlyPxUgtE
mXaeYqJpJqTMG/lMZE3szSzAmxrhGC2djAfee5abBaRKLtvn4yvOXfc+hwliny2vn9+1uL+QMh8r
YLhsD9JPjjNah7UHphPX58nD4tzeUy0WHKzwfYFfH5cynDv1lG1f0oEM1Lcrj0MHqYFFNfq4iYxC
hyMY6hOYshEhHtZnd5443JboWQQeMjjOjdpPvkgupd3tqsYOF6/5wU4WYoTZGufIolWU41a+DEzw
bHkH5ZDeXb09mHRTGLeClD++NnOR241GIzUQCoZqz06oyY8ZsfFE11Ty7z9xE0xVo3TPQ9Wi5KBo
kpuzmIIrIk4oq2fmJ5/G3DNt9KmPcjaJHKiAezv6FErn9Xo1o6SmZMcDhD/7u0e30LjPd5ML5h3E
QDaldCW00eUtftO4g0Tay4Y8Tdxgvzza6wJ+AHVp2rmAZdOvE50YUTO3i1kFHGXRybm38ymq/2JK
vNcMIEUqVMWEbYie7T6vjJoCkHkJ8rvdrbrZNa71EOqBtMJi+16WlZU6OUHRK6uoRNuLJKGQ4Hjg
n5NaY3DcfMzYTYBubUZLNun+Hp63RkHVRQ6t/sn6MffPMZUjWDgCO76XVRAJ5x0E2VtzWMStDqKL
O18oc960bWo5bAbDM9SPtPHswAE4ZgGrJ0JlxckLYekN+6ZxN2+WWSXtMsFxy+8ZlcIlHkknO7hf
gQE5Pv8U3tKb5bfSWFXstHd5f46GTYfMp82ENpBh9pR2oBg0ovR+YPfq/lYxVaaRjanaBfBr5LFE
yry/tFaVhpJ7sjdj6D92Hzig1QsVPCwX/3G8CslJwHCUeDRnOTe++If4Anzdo7qMXQ7TwfI5pEVX
M6r7gEhrCrPBGzEU7SyraWHugniq9TieJ7q8rj27gXPZ73OYXKejjpPMCrOe0dxytBq1Fkhs/IGm
aLF7wKH3UARf7cvShhi+UmRYmL9qQUhZUV23/pNOM/OLGg6rFCQ84xi1uQZd2H5abfTdEGdAVfR5
3sirL7yNkF5Wq2lmqqzoVWwp0c6oozpEEBfyo9XU6hSDi8pNu0/mAXbx6HlBKdqxoYCsKqGxrWci
RPywzhwtO6vlYKie6L5fVNh7MZOU5EYOVWkVd2yAqOcbUZp0QSmgm/v2AhBT7Hg5pu3DQx/Ovia2
GDbn9Z4/iYVbuA+57x5P93I9HvrYazJlBACHqLEAdQZUY58jHg6xphQ/pegxg5ZI4TuKCvdbcT9M
+EMd805iuUbQ5lCjjTz1Ef4NGu9cmkE4B/yRCQzE5GRdB1ape3vJmvRLpRmPOmSv4VudAv32boU/
kstmpac1pSjI/4agUqZifZ0e8IJSOoNFYyfG1xWLJudO2vXrtvtSeNtRwTVb8/8Zu7hcXVuzx5ZY
eYpmatFdTDuha34zpWPEflmZBCn0bwtbspVSUtfC6Vys5dcNiztgO6+WMRMpsD75AvfcCd6beAqt
mAFVOaugt+mCVfsurkeTXUNPHNImB7jRss+bn3Wbc1PvMvgDdMu3xAi0+TxtOLtsnfC6AvhTM8Fn
mhQncIDwTBN7Vo09aNau+LPK07L4UXTQTbe+Nw7Bwq6sfF3pwDkIeBF8RfXB3uSXI/vJDtOk/FiH
dbiqVXSTyVN1Yyi9JKHj9ZDwAU0nx49yHrQiAJdwhWjUy0um52Zv8nzDPCrRu0A6JrH135B3dfKz
+Odv/Ur0fRvmNn7AWpQ6OiIiaSl5A8sySTxJ1yslcd9DikrAY+rRKEP55ubJQ0CSoqwOLaI7NHFj
e4rSSpDp8wfLVxMGfRD33FXKapeTVDlVWBXsw5+0vh9kK/6kCl9Gzt8/cKabidaUmvTYOaK/TZab
RSCOxH81yQgty57ksAtbEJgLfaH4z+zIwZIgJQ+juZGm6qYKz225DIEt8JG9QPjO+E4nt3GYla47
pgx63nCWhjJ81Xz3nZCZUg0jgK5agJQi1XyC0xN5MVlaY+vytC38ML+BPALHlZjoENZGxPH6Z5G8
XI230aVv54xmuZklvH5H2CDO4d+Ma/WPy36aNYrNERE8DIl6aRaSrqSUPruQnJxAKB+OXZzTuNME
7JEXcqjGIgVKXZamJYdq0i7F+ojn/KV8uKgwlWwZnf89G01V7MncPw1nEVdWtxIa6DqMLP9KkffJ
WMXZXptLcROtMTIBou+uQKOx7TqWEb/wFXAKLhGyZDhuBy6nZzWRqietn4WkCKpiH3G6KlQuUSnR
pULCTflA9KHbhx/y4KvpF+pcuXpx8yv028BfVKEeB5fIj3oucnki1qvngwh1erRTUa/DvcSUFnFn
F9JVPfeSXKIwv0Byevh7rDyHMaov+WLbDEzYDuH6gFU188N7kQS35HCyQ73T94Ze7wY16UH2LZ5g
PpmyXh295segiryY+gijak/87e1S1mVlL8kfR01B2du95CfLkoPP76tL7Or035h8SiaJ9v9zPnZq
jnNc/0zZVYr3DG+m9uhaBgakP1qO232wt0ZdMQ2xwl0PvE7iNIEvlZtqTzPDzF7bOjKdCkGM9hjg
K/lT339PSfiaE+5hhT3rgWV4tQ/exmsCZu8p1K9IEfp+Md9+9u6XlfdoV/O6pNTUo1d/1S8gkx+d
3r0hvPVaXO6i4BbEIqrMemfq/GY4NONpuGaC56po9H/mAizEaILwQ9S14zQJuJtvgcCTXH6e5jT0
WUzBaMHocejcP4HRPLGUkmlmhNpCmfduVrLwpmhvBkBMQFmT6Ljry5O0e3/QwBU0QJQt9XFBxTj5
8e6Nz9GDgvsi8atcHCPm9lsq5Pvzs+1ymoO40pyLpZYAXadqy3wMy54QbGkdElXO5xhK2R/6YRPC
AieeW06CTeJDVyFyJmDVvItjMcv+6AdYs6wyfC0wi26DgjZCFlolIQQzKRYWK8EUtOpLcBzeUU14
ZaRoSdpC8PGvm1NbsroWcGsDK5LgOMv13CgUIN/oSRbRDywgfDYaoPOORaFxXRftY+NVj++8mI2z
zQHCpVYtJVNcm0X/bditS40pxrvuxIO8Lrznvcq0Cr+XEDNReIum2UvSEUid8qvPnWvkgRCLnuy4
fn2WvvFh9ig2kbYyZdQZDnWAaldRrmE6QrXR1u4hUo2CsXueikrC8RRFtJYza07Jaer/6gVeuZOi
Vz+xDhvOGDKtLZIUgRiyFsQnc/XCOWM//UCDaIXETT6nCaNrc8QAO89ogiDcrnZKfX2/oxdMTNLp
or1DTacihrGLQTAY+MAgOlTgw10CezxwmajaLDLQaSftyljELSQJvQg7NozdjndQSzpHKWl4d3wV
rVIQVU/VpLsRyPedNldCsfts3ujw2pbzIxEloFMwgAkIhTHwhg+Nev/yTYctC0gUiGkmIe0GBo2S
4QpgkrCu1YbwMpqpYVmtDMKM8/0zXoVrPsXTl13JjosrnTOPbOIBJC70WZy8TFL4Uzd3V4P9HDeY
1KK7ng3fj9x2MbqDcLy3qQrM6SmanbJPY74jJpbmDmb23lgAjwIzhDUY4Qc7WMqXTqIlzPaF9ZUB
+4eR1QcBPzTuX5nBMzsnZUHPmB/cm3qH0RdilS6KFdNjZxLEXow0dZT+Lx5jarbeGILfypsCNXSR
F66mv3nDQaqhUauzh2h0dH4goPxkBzCTDz7ZuHzaFESu2DbVLwzofEcJdQEFqE2vd0q1Rj06pfJS
wgLUSK4P7h165PcPUokDsWDWG9V8lBdaiOTcAeqPeLHoilxvEvgGOF8W/7Nx5XWhePjAIiTSrNu4
vgR47nWR8VZ4qY7qeH2wF1OLQsIABFqiHGotOQjREzBFNcTMtSxgw7nPgOKz6SY0Txgc/biAhrAN
suZJNSDcxlQEPe94lXdY1RFhqkVMfk0/B1t3l+NcxSzrUZmfXZRyDLf28VscBfeyJzaUUfQsifRz
He2AgSlgtdk7zvGDLXNMxRfJlIWt8FUlvVBuTeCop7m8xEQZNlAzy7vj5A8SQe1TL5BeSBkIf+5U
crhKxpXqD6R/rp2l0AG4OeLE8eu4rNQxmYsXsajh963kVDGmwpCkCYhWLXJPQB5S6Xy69Z5thLDP
bOGc7XqLUMRlgLFqIl4PYS9TmQx0bkvGc9QO5vauXu+Mi0HkEfzjOf5SS8SwgtS17Vdj5nb4cRdX
e06sdFGrAt80vAPuSoCk2EdjJgEqxKYddu9iRVEhqctnWchT7Gg2skb+Ccj0akVH2cf9X6Z0bybt
nMlfHBVQ/hSnkvzIfdf02po7w+xhs1+cINPsnrUN3q9Zb2CgnqS4kmxseQFDjcn6OmCQLR5wG9Tc
URsMl3QLYYb78UE0GC3bQZFkySmHSfzZwcuz0APMOXtLTroTeKj3D+KQy4cm5E57w1x1+t02GRWk
K5kp7CYq14QIO7yboT+9TWT573zv4zOfA0FWPBHjesqXKFaJYeDjAK1IPYlVBgjOnFqWi9jkD5E3
ZpeoWylUu9mn4tn8s+7mtiS6x70xCfCsiCiJkPiWD65GgFoHVmxmas1NhZH3D0lVgvCgw5+E20dj
4QUaaWTKNRUlqLgTb0c7Qipmt0oxEOJznPfMAJ77cLZWR2MIF5ZOkOg8pmOSDd+HDUG5S3PDqTUH
DoSv/fAW/zxIm3kOTn0NL71EzNrzlUKg6y/pvTpvxK93BdSD094NAUxmqnd6yCzRqQOaFntQRhP8
kaKz5ldC4rjVdtyt8x9hvwsRi2T0bNd7iS0nqp83smEM36tNjvVsMZKRCq55gh4Kgh2zSnRss4PC
rqu5b+Bt9elAIOK7Ldef653MZAfgDhvh87loek/Zj/1Zy0dtnALYhO1ZiCXqQe/FGuenEd0quwEQ
9SESfmqQbGstfdo50lJ6iFfx0d2Pxd0UbhCLi7gqh3UF2YdYT7XOiH3bHt3PzDf5QjUapfH2ICTG
C0RXxH+tb9jRrDgTgyFgdjudmWUgIqiWIqx5rzTplKXJJJKal95t6I+4mrfqs7Y/kHwQJ96LMgVS
o0FKfPjoBYPdS4ACQBzKKKwRB4hBuBAdt/171wp/Z3NIU4L/rdg81NM+rzSuNYhxjnHH5+NfxV5Y
L0Mv5PYLta+AP7VN9WXkBx2ThyqQig+Ud0GkfWxHg7JAeWQhsxJ8Yx9nl35aufav7Wu//K6GdiMt
Zcp0jshZpx6ZyOFA1xMVMLv0S94e8DwnWCfRNZjaBlhTGTuS+e3gI9JThR5ZyFfTS2MRs/yJvh0V
n+Gam6eggApCO54Xaqvjym7fNmZ9ZN7eWRUKW0nyGMLpyTU+QbpCHgnrOreUcJdqJaLOcpwEKL+t
N6L+UwtMW4K5oDJ40nZ3eVz1z4yb2kTDWNIAnn7hMsof4tn/5pQZan9fJqhcXjSplPs3PC13QfD4
dxR01mPBHauFvFcDawvUOGf1b9iewxh/B8xZdvjui8dMbK4saRc9SeL2E/ikGn4PLiWR2YPyAZ5w
p0uVXywV3MaaIdnYTlJEkHS2lQBF8yRhHmwT3lszVj9Y6akcLWH1K208Y5I1tNZGbIEzf9z7jd47
7DUTJTjXypOYclc4BlZVvcj1lkNqLRmFdNVJUsmbN/Xp1uEgUN+h9Tj6kriPc6xCCTw88Dli5+/p
+3FvZb6eEgowsAnUW9QhDiuFHskBfyoS1GDUrUeG2YtbEqCqtqNNHeFtEqOs+p/ObuoCwqSkSAqY
VNmeM/YD7UjZDL1d/M4AVuYbhROtbFKvLkRlW8/tIx1Ws/Yk5wJAACXaoq2lXbcM1wSlXC+w/j30
RzYKqEIFAf0KF9jvRhCRFHSUPqOXo1mWdIPVGjN/LLQ72heqkR5yPM9khTJU0tXlno238/D9oPlo
tqOw6DP6t7pN4L0iKG7dYs3EeSlxyh+BNTCc0yIublYLK52pcTjykHT6qycum4iQ6ljekE+NzTtz
qCpIJ9urYTM5GNSlU64uBD0dBpAdS33tfA/SySrhJm9wAxyIMvHW62COZ6kwoLQesfXBVzgCv1WG
Pyg1h7YbeMNKn7l2l7SCtcVJiC780LB205L1w68VcMZByLbTYX11f/t6bO3jOHZETyzQn9412CKJ
1F5fhY6pnatVvrFK1Wn9+/Myk75GmEh3v0LUsJ99soaYRbdbL4Ql7qXHc05xcrM6P6p8wgIUviQg
imwkOaGFyIQbLPxH4mxOQ8sSfhoeUAbJwG1TF9LWhrk0zVQ25D7hrMhTs88hv55cd/JU4tFhbCke
AtTefCbo4pvTZzCjMu4M9e5ulqKafvIqMO1X8CZxHTm65BFnM0U0zUxIt7XvKLc3aXX8IArAlmsk
fYb/5XYu1iE/63lyAMgb+Pz9y8BEdqfSNOfL8FiW5WKTwGfkKaYRyIhM5FWBIAGEVH621buY51hb
t1t5DbNcQ4iaOHZoc6yTUP+L+FSH44+Dc8P+ZZSG1K4YuP7ZVgJS/0iSmWQTKMJcEgV+ZjH5GY8D
GJ6Jdr1MzhF+qRCW5IuudxTlE2VYFWmdRLsBBTq9hbUAR531ouXPyQobXY1aWyduBQfZEaNa0usC
XffzSZXuiTZ+/iKVD8K/N3K4VE4yPVPGfVW+mjdI+UVRk1Ms1ME/57ZsGRGsLlieP+TAxPcQi/WT
kRzg8hS1qsM1PQ/DJqvVOJLHmBYD3IW2kczdpbpvRmZ7gZHMIuz+Fc0MituXL5d1yfAZ4qV85clG
9WUREXPPN6TI1gQQ9eXRm57XG6aCnPJIZ06l26BuyogTF6ri0Ylic9FE3wK1AooFl5NPQ4t3A9ZB
oNnhj9vwWwVOi9PZj2KSzz+soQ/m/XQglTF6M5SrtdayBW5+RVkaJHBFM5klsM112C5KgkysNMTC
u/x94eLO+3J6cdSV3pGDDlLC6M7J2Gp/u80mG+3zm5Iu1ScOqLeCUuQdIFwWY7eeo+/PLqXi1/ul
OtrK9GuK5HuUlIZ7aGERm+ofgzff03XjapCQYcsjMfCb9KCzj8SFq43KQ4ynH5gVM0zEVmq4P3FT
9h/+GH8zuIDGpfdXaGr5FiG2i+yvt3/tbU/GJ1okhWHXBHZOSY6pH5C6B2oNhgyBRs9ouC4tYWcm
DAi+GznNulZ+sV0kpuIuwAZuQmtIoUY8LE/7X8QY1FNfj64vuJHK5O3uwl9jBOMibgiaIweOZGVB
TAUAFRxQsa5Gj5Rq8fQ+9dv3VgaEm6p7ZmDdnzVc3iPXC5CG9l3UU9vBaXURsxupfEyPGGYu1chN
HUrNFjht7wnTKGJXNzzmd9YrwQjK9lwNmJ4AUqRrLAkM7HJ1PQyfMTUoTvbsk3FqF8zd5gfAEFyS
acyDNftyagWEoMjbYHx9t5pW1nRpg56TldEi2wSwbIqent/Sj9UaJ1/KywKkqEv2QFHd7MPgmjYp
vpAQ47boHd3tY9tIHD6Wd5N/7MU0DP41B0HL0T9fs7tAJCrmuNM4l7DVdxdM1lXFeuAU1BqLcIYF
Jxux5MU+X2l7UCWqoCYpdXTU5ln3oDR1k4aI1SgjhJu3KRm/VyDHgYnjXWId5tcearA/9WNqJLyi
K8S3ihWulqpKQ38eS+vM3opWvbsBR6q1xr5cc7artuhqGl+7PCO4LRznMhGl4Fgf8cDAifI7ts+K
GYlRQdFpMCT2AM8yWCCjM1iDuMmyOuwqABNFUXgvYV6pnbF/jkZb+YTMkMDZsHIDtKgKGvX05bFP
IWgBUyYFAxLnhyGI4yeSBL6XBpPf0fbstkJvWhB5mHh+3IkvnpJeOap0WHpaEBBFAJIT3HqLd/SP
8v+u0YSR6FKPOkOf53z/EakCq2DKEg8dTmlnvmFu2+zKMybRWjKmL8Zxl7SfLFLGOQbUUxi7QmlG
tNc/muMa5iftk+2xyrg0+6ZfWqubkenHRlc02cScoOk9/ES2j7NshDL3wI+KqFp/hgiaysHOPJKn
k95XarFB2IWVma/AirBEGn/kffY+jZyWVW1oOeoZKF7y3hS5CIFkgd/wW+VTCs1j1wMefVNVIKWk
EjMVncBDYI/EHMsXiovMZ1Y9mYGZi9bNHXpixTW4pfaarO3+E8a2cyjaPetKjN/OsU+ze2Mdw9tw
ffefF1inAT9W3Gr3Y0uT9XqC+sBi1Z7FTpjku9NWSJBpqBnH+5MdLasDV7bsDFyvn07a60BBiDmO
FYVdMw4hknnnDWcBoFclgLhOFp0tsepQ+bZb0G0fgT6o9JA41aMu7fK4exx6ty6Fq3LgnqO5xXcG
a4CSekfdMxRRTlWRzZEw3SyZPLQUAKHVQ6j5mPLjwFNhzwIfxFyYF6Q1brWi0mTZY2T3RHP/IVJW
7HFdGAXOOOWCFS49aclThpTW2f17ll98J//0duuy6zY6H5p0BIy1nPHEf9EE+hJoe8L2hyb/QWt1
tbT7MfAw8ctAcvABYJdz2dQQvsEeGPy2QI/wVBo6Uch6luYgDYZ0gUEpWq+NBUhtAi2gqJKQi6BQ
FmbpHYoue8iMiMluV3QagBlAFZUovrSSugXLnkxXeV1L4zCeHh2s3HxOdpM0/IG+WxCp5PZv9sU6
Zy9ZyzjNaP74TNET99Y23L9PGsErJvzVpC/uBY+i31anY++AH3f9YZCe2ZYeDbfpJQsKo+UThF2f
hp7FqEwWpoGFVCX2TBUDvRqkCvrsScgTkYCibNyenuQyvt8RcdT4aK1dYVIQH0RhdhbpgF1ZctFk
dzvhx+YdPtD5si8shRky6aVUpRDZJRYlEhS29MRnFDVADuQmGlIwq8PmvMzRT4S5wYYBc1+3do9W
o6tEe6IoOu4dvvxD7FC3kQqgD3mC/N7uC67dpaUBFciigUUCW8G6Bom73x/7R1PNpW+rt8cM5B3u
mbyuA6Uh4g8/8ruylxmiOPiZ81UitNx7TwV8lSZq4QUySKgFscMjKM/XAHSl50KOXscboEYk8NMU
SMtxIw+CzD54HgaH9NEcD3tIgCWPG6NZ/3x5DOK7Xi94Q+hnxye2kmjfLnxAULhUWTwz9dbM3ZK1
y/5Y1DhiVqPl6jeYmasV293uEJRt7mc1pa0fTY4RQFQg48kH0c6eA7yNSxsOYWkAh2clInsCwvDt
g4LChintgYteisuo+OsSOYwZrgsZegBgYcrdrI/6fEY+l6u7+lqsU8FN4SChMFkiJI10MzV9FOw/
sjx2J32FstefmTpfWK+eyHUTVHKs0I0YcZx8djDP+1Y1fggAKSfJ3FfakkFpffgMIlCwjY5hmOek
4ZvYcf0OHAUwtZxFe6Eu/YCoKPtLofYjSCROpDEtCeSV9vJCfnoIU8/zEcBUyXlVCFqdjLh5YAGy
ZsNdimiH66Sk/udSF50NJw/jgZiftk9iSkoo7daomatr1cZ4BOCGXPWV5JYXWF6sWMTHqbBTnLZG
0lvlsaMPGDFtB0T/bcFQRuBJWscruDsqcoWPoGA59Kp1hPPjczanQFkgovSo6VOFxGKXcb+M4nFD
yPbPLWaGeEA+uwR+BXKGV2cvJshecJujxmV2owSAR4rUrKazqv8pXIVQZP/9ukvQ2K9jh2q3j728
WtteQqW1nbjJgsNEtVi5bAnp5SGwAdSPmn+NRmcacm5PDgnL0fmqmZUbBPfZk1DB8K3hceHTi/De
NiQvqsRkM+u4v9lnVW+5RQIDIOIf+4xp8Rr+zXPFVdQ1hipeDhw1gGVp8EN/5vlCLvfGs4eaQgjD
VfBR8rZMlDR+0cnVIPFF6CsUl8FExmCkjv7DrBd7i/43RUs+2Zhm1KMcvXhPiCHTVHvW/NWR20Wu
P2Dqem25+Pz5oJ2sznZKSen2SfmwMAvMdRMHcjTlzGScIeh/SCMjwxWQIyGt9A15g61L+HdPM6KX
HhPtHW1Y4u7k4FQEuQMJU3zMnJ5VbOOLkjkzzAk8run39DF49C2Noxzv/DSfsDVM1Wy/S0c3PusA
S19R0b1FT7lj0m3Pxjx2IJ2QGPXgg8kcoGrHpApPJELJJDY9tDlXgQsX4MQa8T+O5XvWGYU7Ie8B
kTg0QPSQvqR1o7oeIdVBvQShZIYcJ2aIE87LopzXY0DetaOC01rIOuC/rUT7r4T3mF0qaS5WpIXv
jnBzXIjpbN+nXynG1VN4KbMmTb98OqR/KNljVCYnUPdpktoNXlkAepmxnhkNOI/nVjqtxrYIryue
KvTeEx91L30FIgi357xVgzkBioFRx4RM+7drbuxBMA3i21zvGU0Fu4LF86q/QIFOssQJEQqz75ja
5n/o9AHwL7ERfL6evFrZSyTjWRR1OmReMGWbdYByCPKPyGawNVSMGN9HtJS7FO/+Kx1NyqdGoxFd
m6CL35etr9THFm4yK2VWO84ooIbUth6pvLkUktVBKtoAKyq1y0bLkZaN96eIKD2uO0kvMtxPOpna
5Y1ZRQaFuEcgCnjSRsDr9uyyDk4bt/6mloLHrF9kfqR/LUB0tRTCoS4CRfO052NuR+RfdCXtysnR
aZEX8hHdXGRPSjClVv+i1sVefi+geaWNQurdagr75GrrNmyCqXLwUnv/n1QWS5xwQat6NtuzIKJM
YQJoMOm6LPt7lKE1Ootr1jO6AlMTJG5QbwRo/JGFO4DA9aSNBw5W5gLPI2nzoQcBQisk0CIuVoHY
da+7uPsnuuRSWs6l9qS2xCB7RPKsIZj2Blp4a9fizmqeDh7Mzq2EAqcZurW3uUtISqG6zI7SMbxN
/4nlHcFMbFk2YzKTRlmyf45noN1y8ua4yFwbUp1hVhdkcHuOoaZYcFlQZAptybdWSHQ/OtysavC8
pC04Kyj3EU/TvaKSdePj9cd94NRpLkglJNcCUQrFBoRNsobgxkrCAmif0CGHH6yV+fFylcL23VTI
N0VZolk+ekqkZsmJ/Gv4RElB45GYLFKSMdUwFDfAwFLHca8bSd2K5MrltEsVreaD+yBv7Mu6v17s
TQsP08toR+ZTylGLurV/37npVrdk2hFv/7Pcn19yts1dSq6k1yvS8GkXEtxKyo/fAstCs/GCeKe4
ocFUzijCfrlv8dS6PTHnHcfLTdslGRMhhGwaDouePmlAV1eTOr1XFzoBwEgOpU0wIJVx0mZ7PCwE
IqDYNrLcGlXuDttASbRVVAzobkToYn2vGSUr31grYFSyDK9PrtRznQ2DD3cXwGQz1QesF1BK61DJ
qpmDof0Kn/u780fClhhd2kxZQ1Zdz0UKBv6Jw3/W5DVOCxJ9xjEq6VJsUnxj+L13uvMqCQljlE2w
zcJnNTSit3eyvJZ9+pxSHuVxPamsjuhl8Cd2M1I4/Ebem+ABvRySXP+rb7hnEQ6i6sQWZGVnGp/d
OAetAtyTW48UhDwaoEXvkJr295DLBQJenFzMGQs63BrCnzD/meuvmZncgB2Bn6nr/61VDpA0t/wk
zyBAVx/P7h2r3osD5gSW8Hwx7O09lHzuJqgcAwcyyDJPNdmG22KfC7CV3tZ4gtyS9NHQjl1G69R1
sDrUqkgo9P2Xb4Ynljk/2BF1cXhQz0Pp/2wZcQu0fmddY2oPK/e+4blJxZ1Ur8QSPNsd15eLPyDc
vTcUz7z0U8d+qVmXWOFaBhlOLhfaVSokkAxvrEv2EK74KvDN3c9/dmIBrnZh1L/BbQtNSNBqCnmN
jkncYUdHSv6OIT65YerJ6ImBQz0Yo1WIF/aICcNf1Rd/dcRUBk7Qy/WJwd+IIe6LHxokeM/4KOx9
LjOvTKwds2+KIPOsq+u4Y30a7yfWcVOqYPRSgr6TuiTjCUrhQbjPFgJh6Dw1VT0rtljccenYycAs
k0p9MeB74ovf3gJLvRZan+mpgta9AmEhuMXYCH4H5T2AxA8o4oxedg7dyQriB00lSloELXqOcY1/
L0ltCm9QZ7IpiKafjgJn2YJuNW2em5D4ZH8Ez1qiC2OEXlJSrOUNQBDplKpgPabB+rNwDPn4sDiy
zF7QHqzlGev23eqLX43wnZn5S9w7zlJbvC3NdQ6qzkAxvsN6VR5X8T2gxuOv/u1Kb36pRINnN6Go
10fShY/vqc9c22zFL3qBSqhDt9NmV/XMxGbBwtmJlrGk8tlQMniv3fc+K0w0ImmmtrDgcoOGFok+
HdI4S5x//XRTZvRZR+bEU+rBQXesJjyYsfo5Pl020GwA9NqbJch4HdMnZz059Z56zXtiuUh731xz
nd0PAlVsA5uAtouZc79QcTwY9xcE1FSJ91zDBkhPJtSQtsb3Te4EyQpuASvRjjDa8Kd8X9iFHl7i
lFs0cyUta+Cwdy7QVOkMrBNH7hbnxEWLhgN27jT6zFgBmtFMXLyydDxYU4qDUmh0jRkwGj6AeEMP
91bKFZQFYw6TYO77bBi87/QKFtLw2pu3N5xaRqb07jxMkhxBlxy946rpBrP7lbOggi/S57fhjzWi
PuVKlPnoG0ytyZQMpGvC+ROJq7tG7pcyLXpvENc+l0ZM/jEKWGQCW/SSv/m5CUoSl2zc6SGXoFkA
jUgYL3bR9K+71tRrR9mQodVf3kEjY+Y1Gts2RucZ4QXJyH2o9rIP8I85C4Lyr06E809aKeOw3sry
hdfyVEBeJTE92CG9Cb1mcEdIHJqnreS5DdgvDuIXKELj21JB2VbSbaazdtcmSnZ3sW0QTIhx1aid
XsQ/LHI7UVwJQLPBmeyd/TOlZ3coQvpD7/LH3bjljEgvFV/FHlNaKTbNJZxLbhA22aVnYmjckybr
mBrsV8+e51ie7JbuZeQG1tvzXx76JUkOvwmh3ElNCnWkTenRzTt6pQcgWGczsu/9TVppFBw8GSoy
X4KqBmegkWawUHryOlcdrwYn3Kcm6QcC5m3ImGs0LS4eO04hzXE7hjDsJrUI7KunSS6f2UuxyviD
E3iKWu5F0AbfLKxHqDYxheTttmQc8rEFuUK5e+1wKHN7vZEVW0kF85v3oKqFsAo+Gw+tL3o1wssT
p2pDHY3gw1B70Y+cH9oXwn3UgYeLEUrjRnNlVuZ0PjYDPoX7rahrhYo2J7ouNakeFbhlz/oDy9zL
UqRGIa7FS6fM/rZkTjFvYRgRUP1NBC/2WYADSSxuraVtYGmFOejfnwu7MzByPdNyoRPFU6CE+uhY
5dL+a3jjbaEYkMLYhJJFEuTf2pXKELnezZVU+3Eug57V2mYuEq5/Olf44kNHY+wH7IunhjugW37L
3ntgvF2hKzXcYI5SQ3BS9dMRLJWH2pWuHw+CvPesb1BZY6zGq/f9NA5zed+W59XsOK0jvDMXiYs2
Ce4MY1lS+Uuu0Zy7DzYlr8eh6UWTAo9o+sYacF+GLRMZr8UREpYB0KX2wnTVos4+9JSLRhMqr5HB
KGsJ8g7kgQhUJB9kg/bhxC/2NXtL/38+C2lObGdd+zNBw6PQuWth0JFbG4mV1LhCDG3SfNLtRMjz
JhHvjw3D6c2addTY607I+EgBcUm+h9LR96ubj746GeQHAz8fOvMfPWgAoaY9sfFHLGhJWvEujf4v
PBe1Em/VYVJBQ7LUsvoVaEKRBz7apG3MDCYQwLnscgvesZPszvrf0v1Aac3O6gjdUQ165vq7MBC8
NVyJOx1Nv/YEwo577/dChVc0/yK+K5usljhZJ9lotSNVpWsC+VYWjUlu07BwXQlxzSs0HoFeg3YU
WViYBjYraVGxkKo+dXRFZMpFI9spioy0BGTVjlvLDu6n85VQHaA0bvF3KPj6H9SXQ1FMfRvkpMZH
4GEzk/6pXQE0UI+Lkvk+XCCTQFbpPTWBmCqIp6mruxNeHxb6ett6sKW03SCckIpdkxM45GMWhsWQ
VrOTN7rQFMyJSyUeDbEO4qBVeQ7KcftvS7ZEvO4dZuV9GqZObzdD26UGG6TAO5XV9QCaghWGHaJv
RTpHy2ICCPkB6tyMxlrlyNBZQO8aywbD3/iAiJN9GG9WSdCUT8ArMuFL4EfgclsI+tz9yKURW6S8
pe8FA6ltmoJ+0Ag/YSFSkYHp79myM+Bg1yHBQ/ltg2o5LG54MDmd6243Zmm6Rs0mp0znjwdSJKK2
sc5PLJLGO35qbEH5Qjn+vT+hOeigH0Pmp833e5CE3XiM4TZD1QYQH45eFiycwIeK2H4hYixGGFL9
DaSIEh2G5+1ZR2DcJ5V2Z4Nwu4E32rEOcOGjsECOiD1GaIyuvh9bxpy8vewN4SPabfI4oBFcDOTl
t/SCK72D0SFvYYd9su2exJuuVpZZL+N10AP3EaCEV9P18DJnHHtHGovSewi4jJyeCVDX9sgPAZKo
0IWpR3riyMqfK1jq+6+S3Y5F0PUU0aBKk15g/SdnIOh0LvuhfddCvuQrgenOg1aljPWL9RtfOxYC
8gE4g3+rsRynvRLxrAnmLumHxdAxBDBhuOKjJ9ZZEgSMKOCTAgLsdcCFXBGD4E7lIR2se1ghUO+i
DR2sLrPiX71AYIFa5mWUedAcS04HFZE6W7lziHLxzrkoEeibdninhY3bxv0SwKePmwuQpBjCtOgs
j1WOdSVmbyXhfeQazKaJo04+BklK8v3b9RHoSJijOLshaJaFvWLU7QDeoEFKe3OwtGczVwxPde3+
COXf4WHZcB4kzggVk/xetQokBx7wHOW8qNBB8S6C0WH88sWuqRHbMMTTc5QbTSuIRzeaQm9bhxd1
DErxmOOWYhimZGyfBLnpNY/12h4W4ubrweKArlntk/s0FwVcFD+2Vz5eNwRuSUK21EtzW1TmIseW
vb+pXiFFOGOI85KxseNEFUU6dQOWh4JkgewFgzCevDLM1U5NfY/HbH58QDtvwxYQoGNR/IB8ZWnK
NXSsIYs44HQ6kQWOUS22Ynl6VkgdlmKTQM3+0n0mZTpE6nDf2t28SUBU7JbClp47+oDX7s0tsg8f
Kw0TD2OKFXW51nfF/lFpiA2WHIoPYeNLLBKoFNih+Zq5ny76os0ZSX2MGNILveZaI1YgMfZbgRn4
O7zBYKnWIvAR3yVTzNCNrdd42bDwkI2fHA1XxAzSl7fL4JY1L4lcIrCaHDr23b7imZnte6+AWfNe
E50uuHGXfhkhlW9D9pgCQzswummeyerb8JRGfR6xHunpApa9D1N2i9jq1ictIbaO7lpSDiWvjtOZ
bkmWyyeMuUOFho0BWD31pTq6gw/QEQ5xZYAt/FjZhT4IawPzobtMNXjXjlawSmgXLXUeUBcNvGVB
4yGrEVjs4Pkfsa/j8Rk+4KGQZ8lNPodHAGCv1ER6PPMquKAuFmuIdYrDkAhlOBMzWPqgSyv8w7Hj
m4bpzfHlk8qeApDTUgP0RaFtV2TLRORCZwspFcggsii26Kp1M/zjZHkZRdQAqHjRql4z67DNOQRD
5RRB3dxXa++kOGzYZoYVdA5KGPYoBNquYk0gUPAF41AlccB2RZgfPSVUorCJsdWzQgieLeBQnmpZ
9NtxNUPlcsU9HbRKG07OY1nwDpj560mFMUMTqqVs0YcCipqH/tK3Ymt+DLFiylUinqUZupf87ktW
Cy84THh3SvezO7aOAFxSZs3BWX2Ig8DvHq+1FOWalCvdCDZFtYB8NUS/q/b1bKdTLpth2Tg9wibG
IRBoADURtD5xTSE0/asGvRQYjbvxAvOnPfA//dRKoTDGJeH3THOT+5IQYrwBNFsfTEK1btkFV70r
CS7hTPxwIErw9N5UloEBRVnSZS7KFKH8WE8lncCJgOkpzhze2sCpY2D931chs350cFNvVkMVItil
pmONM/gcmTtQiyO2wgxhMHd1VuTePdXLvbfFoKA450pSNBg43Sb/5NM9ObiruuJib0ClGYxBHzQF
oT87OKHYMnlGwZTEhrQbMNyH+mbeVHZAdSBevXjv6HWDXaBMY0H7mzOQR2n4odnwIb9KbNMoOjfe
5n8/1FIQvaCrVYUElhvT3hLoKOS+FL1g7N6BhF9X55GpkHRcuhG5C1ZKN0le+EkaXYsS/ur0D7zY
cMLXfrG763R9+pI3W/arJw+BLJQRCyj6nU7Pl/TCqyYEIOGxFl/FegWvK2RKMIHMj3j2TP88s1f6
mZh5Nk5fnaMG76GCoG4jNZVbynMnHLRM9lFV6R/mIvpkTuBYBJ8KI1ZuH0THFcr5o3eOAwWud4aA
7Vt4sgkK/AvfFjqM0k7KJiBNNDguh8VNeVmcV/ibAoym0MBYDxoMXv5qlGxAsrgpNffj4PFjdrwb
bt/UPboZEGgmoqnchQVrK6gl0MR5lFeBFpwr/8rBRoJXdzOmB2zjMeYmPC0DClwkEVo+SCs3uF3M
2WwlpQw6sH44VV3uradZvl2/HsnUWRH5JnD9xKq+Q84g5+hXo1xJtPpyW8XjWI+zxrtyGGZGm2Uu
bKUg/BO5f140AVBWGUs0v8u5ccQV+J0jePoHMIt3Cs/vnU8mNYTir9evC64vcNQcApFC4cgpFVZ0
asQ39AuhXOIRHmbzrrsjqToMavoXi5SAqqXgzZ89BsDeYfjUT5Y2qZ0cYY5yLx2dZEgxkH0r4eWA
ZiVhfUVfgeHBonyQJZSd13nvJGRk6kBn0Jz9jW82EB9IUqkKdjIC5jvVv9qtCBfmUFwYGc1IJfKm
HzbFwomMDbD0hXzuRZrRGnlKuIvWBaGRB8zCrkcw9E+LVpYUPQGGAvnGm1AuFsVkGy5NjF1U5i4+
4p4egUNUrBzeB+M04Ui7u8ki4JLCrqTJhgb2oeqcT2w8iJP81SZOqD9x7F8tUr2MAjRNSTvTJzNR
7VZXnHp4jTKslnsm/YVR7ISo0xYVxpMMiBmk/O6xdOzLGWvvetbppJo0GWWucJpWkaM2sSGbb8KK
fwm6/H2FEVkjo/amugXjNa7l5cfKkVO5lJzk3QQxqa6XJQDngHDzCmtTg6a3BBv11cRwtEJ5oSEq
AMtJD/H9zW/hJza67iLfBPKa7u7b98D4mh2RC45k4l6FBSG3nEWCknCDMCA+qx9iZ+2AhzEschBJ
0qXgjkgnPYIWgahaxqdSNkaqxs17tE3aQuZ0C+RF27aTZb6r93IlgC6bYPUUx0iHUcr4sxjaezIJ
4+c/mSsaEyyF3mW5yFp2cXURNo8c06056F5YRmlZe1siKu5t2oBGG99oEJfbsddN7DoxQkW1b1Dq
uSDmSFjs5PO4u9aNQaSZlqhurtmMtJe5ahNsIveqKX+JxPADMze1krP33SbHm1qzOXC2BOhLzd+x
RvhbnyJUP8qzO2kQnN/bjYY031Uwc1kWObdLPKRMb3EpCs+PJZ35iQfsNUCmOy4lsjiQFsqUtkXE
gymP9OxGoXx9yde591UQT/TfTla58P4sPvq8FxWWl/fcp/Cb3Wmy9xCG31/jx+kkSTbDEcC5G78n
tstd+nb6MA+1qCN7kJPxYQYRGaUfTVj3mczmF2Ipn72ELuW7DiubF2yfjhZGG9QVys6W52X3sftI
CncNviACUL3cWanHT5U4WVTdpf9pJkMzbMY6jSO/lka8wm5zHJ0OxII0pllwMQ53SLYA5GhVpfKX
d2L07JYvvl5JxoMVbSrTwkajLT+YwJQqSldBp55NTlOZ5CzZyS9d+QXkTU5ELCAk3BrO5CohmZE/
P9TvExDKKF5aPk5G4rA3OaRWNqcmA0Ip8GIthny4iIqn/ws/hBbF6Zl+cBITYPhIhxOk+rut9ikN
NHa3oiX2Nojd3PCizA+xnbvOO9/W83QxxG0Z4hN5Ylh4JpPpKLaXUY2KqFRHNh0SCICZ5zFCiziy
Lw8i8RHP3NRRmgm9T7XidFv4Rd3Q5LkWKCsIyzm6ErFYtmnWR+mjMVFo3xW4/1/IBIvbWncKLwUi
skqjEilBX0t9WVDXypbH/wzV4udu7NVy3I7esvyl4skRcMgWXuagmCWxP7ew/zJbhrKLrY6NUctQ
Tx2OrxZ92uM4fh7RpnXDLLmJD8DhtBSQF87eMQChWlBLJdUGm2qdO6/P3wzHXZ/rn/TwdS1rvMcb
an4XR9wCqpQ2MeBiXC5bVCJ+Xcy8xOV/lx7M7Kt1IeL23rl1lF8yxtB2RE5ejCwjbEchm3FryNX6
sAUvEUU4lQ8XDajDMTYj8T5Fbm5VOVIJoa4H9p6DLH6AZuvLO7y06BpZqrudF1l6XH4tspTHeS3i
QDV4UWuiLp/XaNnMGRzRlrA9xlepiQ00NomRuEQz+4VoGx1fMIl8CP4YehyJw2hLsy4jV5JrxAHF
S1LhoFWtAdrMzZoibSkeibjE5miKgwQrkZVXj0IeojIjz/K+1BcG5ugnm8vh5i0nwjm/vYv83L+X
uQoI9ShUsYYyWtg+ZPD1KqPOTC2SuvZhRzUtRl8ccwF2FiXfpE5VycA4McZ75weyu4Zzy3FxCMnt
wYHmHBzDSB81ciShkIWWu2sGi1HNZdaSVk3IIdzawjhVFuM1yibgK6S3QPCsbIxu2zQjuQqsTxQE
Z1TitQ24zbj1PW1C3f3XfyboBZcShVJflmTa5eEoDnMOXfB9nufRLbvLArWhaB9nskWkmr8Do7sI
b5/S08/NTE8S+LfFoiS9R8PwnPYs5bGoanYSQmXegUfbHW/6TaGJjZhx8nP+J+aX+FSqIry7ZJ7a
JnDWDcY+4z++qIjUlbZxuRNguhK6YMkxrcarTCqOV/E9WdCelGqojy0ewHTpKYnJAwkKkINpYqbR
Z7X6PWfkwmNZzi2JMSR4TAJqO6zqS5SfEoXILVYuI1K83i2k65gtTL7PKqjPG/0NoLUYFLDVY1Tw
UuyDd9S/k3UxZP2ZhQP+xuvXakx4oyZPtyyu1VVXNh9onO9px2rE0G0nMopXhDYPfJWTfMkfbBa1
F+G9jfizyWnSy4Nn07XytRmXf1VEbnZ/2+SYIclTgE1tB17WYdSQumUhfUphWjO1f9WSrDtE8N1Q
u1IzvCElXmVc6t+U+hQ9/ibdw34HaqnzYyZpHOhG3Cd5VUIUHT5PMVZL4irk7V7f1F4qbBthtjFa
TIKhx4kuVqtN+FEPzC9u92xSmcwWJjvR6oh11sgeQ7TjBUHOgF73c45AFlqbAENFJVK9B9pW7tM/
hkx3k3lIgJgaNEhuY7X31Bzz1VtQ8Ef5hq8LtO+WhZmfasiuVe11jDwP8Drp5pqhbKTaP5X26W6O
5LChue1DjJhUP66CgMy024L61w/te3aMgrHsfHAC0z1zSWoPBJZMKF8fEayq6b4Jra4bFEcH8d4U
ivtae2ax8WRU94/62GB/GQKGvoDDJLgfHNncwsU2McRUg5iP7RLfiPiuX5VH9IA5uvji/rvLlzOX
hhGoddNjXi1v7s99e2TflxD8gWeFFbe5j7YkTMDCfeEArGr6BgpZERR4UkzNxC/lvN2VMYoZSJW+
5/sQuvvcIwnrcKb7lC0f76yUoRZdE8JfmNnK0ar/gA9pLAz/j70fr74qolnoq4PVjfniqmL8XgaD
KBcv1g77PDsrRkRCl03vJgliYONjmaGfnAI8JZJ5R7h0eCi10VmfL1fnzpzBRxuCU26osrsAy4Co
qK9XE8d6d+j3cfnNQxj6s3uoZ1YuKuKQbajyVePdNVNK26bVjLfq1gmj1WBuko3zpNWx48+BTD7j
ItdpymZzQdBYgZa+Hb/BY9yE/okG3TwQOV7GvNihV90WzVSZGiLeVUyW9K7wB2msTmCuY4O2EbwT
PqoSyJ04eAmMnEvPfwD9hT9DWt3eecBv9gz+pZAdAYdC3bcuT6rOPleQKtx74Xni+Zlt7x9G86kp
bZEU/g0ALjf3wyl/9EHbAFUj1y5sarTH8UeGBVieHE8bpVi4Kfo7ZTvyKw/+qxr1wsKybB8y/f2a
ikJ/t1zWM4NBjJV8OPzsdwMRIY1yYeii9vSSBdWmK+9VyxPUz5uyCi7GmnrFnK8uc58Es90s3FE/
w7yD41m7KzyJlt56rtY3/2AT8GxSBcEQ8XOOVGLct8DHsPGLRQkIl9bbirrU8c4Kjyz+/RkWF3rv
yNx1W2cqo8mzScUM9C4AcFYG8L8xQoVu1FhEsQMy6d+y4sWn4Hx95cu9u2B+30K+p1YNY1wWrX3y
wbcY82fglqqh/UIuWnSMv73bNV6obY1XB5XsVLYDEZJYTRsXn3k5MvxguocX0sReQSlGalA5fty5
eWkJS3scx6F7eblUxz3rx1TXkOgyIIbRawIwoFUNmV3jSGSjiCvpuA8+jE5Z/O1y0DJ9wFBW20yf
pckyPf8MDPgDLfB5YpWTEUZPAuiToL518apMtEudoC9jVeWdphKDaWNFMGYtonent8ePQabIxo5F
7Rtg+jHi5GfxV6nGOH0Wnaq6sCc0tt04Fs2akmvrtGfKN7aozoKu01hFl9xpEO/LmyZe6jMS/Ti/
IOBF1HPEP5Bio51Izpx5Yglj+OCvzomiPBM1N/Q6YAGJBy8qXohVS4KDAQKlkgLMio3et8S2NwE9
3nP9SGP2H6DB+xAB3qqRoDeCgo07p+NmTt31u1sOqYUqHKgWohmIRD/mZ+NDKKaS0arI8nOFb+yR
CX7B+Zqid21I7zy00+qVOyETB7VKyuHFL3NZQJ0OFvDU+wVD+5dcYRZtG1rkR9MdUOvUEiVkwntd
1yxGsbvqWrNQIzcDHxGDPj0OZfODRTnyCAJbKGO88wUgPeniLS6+GPhIT8OpnewCrFqCx7gtkEUT
znuJGiQoueJbsOUfaYcEz5HltCkAUGLMTWIwhWKEMy5hyJ/VOQcajEprsbs1KP/s8rxrsGIBwcP1
ob5q1da7ZYCy3y8cYC2Prlx8zV2fIeL6KR1TU4+Nafrfb+75UYhXpDHocQEv3IZXbPseEMAsbrf3
QxGBGfBanJNLQBK+KdyRlxjlJw8V72R05uQtNWYs59nclno6G5g0pihHzfWHb/u6X1Wugmf5ZtAX
t5CPtgzMIpoB4v8GFsOAtlEB76kfTb/ac3UwtELhvw27v8+B820D3FNMO6wlUM75jCHqIwbiLhLj
/mkWPyvrScAbTuCaKBJA+9CPxQxXkYzzjy3d8H7HKgdA4y83EuNblIgHv2OFIDoLflQZ1qEnEExm
MULCh9KyFa5lspqlg+5njvZ00ZI4ewyg9B9HcBf0CFHfwHoL8RxsVuviGWMD9u15gTKyRpS4CN9l
F4cNvkKagPSMszPmmKFk6Q43wC08Msv6KL87Zymdee2NiNRRmRay/KfxbM7JqghFEaqxcPqblSSn
c3mJdGkAsgztRwjUGnx2zOsJkZr9RujWTEJuO2wRmSiFaFOk9SAghiLw+yI06GK8izmgCYZSttfn
ECHXwZf2GQN31FjK0szXS0AC4y9ExaeTi4mfoWiTmHywjbe4ce3FFOyzLbQt0fMLfocJND1f3sVs
4TMfIqeGFj9wjsh08qqbDcRkxLl9hAhDJDu59OuurEGcYujQ2nCFjCZU96hHc8pvIn/hR4ctSVEu
zQZzy5jXN31iIEl4Iz1+xBBXYVEJqc3KwwGL5TkI5kYWAbsxwUE/qygYbcOoio8mb5IpJcRGioF9
flQXWk+wCEG7EGLeVrfI0Idi4ImUSQgb9qZ4ENCXlyKYW4NNq+l3WjvImSeS8ASHTnpfBbJf+FCS
dfVpQE/RiqxfWwzKjbLVTknL2/RPrm72DVmW3YFt05ImMsG8JNTh6anUoRraIp4tb4oYOOWI6xK9
emrRCNqIueJTQXBo0lqynOqYDjKdZWnW/c44bEkjqxrBlxMyJmVZDJf7+BJx+uf14Abw0LkbD1h9
UYkC+3eJrKwzCXfo5pjzPGup2mtPKLZpyWd7PU51SNbI6IgI8cMmqdahru4Y7HnjG0QwZiO35z0q
rvNLetARMBZjFyy2Qwwt+mqA7SBUkmoO+df7hS54bTWPScCyUQwK6Dp5RM2+sAmsdD+hpf+JJtYV
DwK58HHoUj0GZL52IVZzbr7UCjl3P1qAgJFcAwKcP7F7bOgS0ke7bkH0sknt3z8z6Lg8i1kt182P
MIqtVnD34F4pBFHYVpM3edk2sqsg3CLtjZciBEGQxx34zAetFYNslzM/rrcFkTkLhjF35IeQhktP
2ASI33Ith3hp5KCsMTm2Va+/8r59bDxZe4/gtqAP7fDQSot/K3bcwaJUwGBswuA8cuiGr1JwOU8/
Z+8KrH5UNyLFGVM+MGwsaNJBFu6vPbidTo6Wl/XyiGTJe3x25Qa5rX1BKpoD53/g2cs6nqGYIwmC
CZbnjULIwU/cFwXf1Ltw47xjkWL0QgnveMhW2nO2P7vLNbhhRyme1k/llFW/eCFtURvMT+1e4A1G
WTqe/AV4/u5rYMZdpoeT0jlW5q7C89i8WJfVUWTCS0urPxmGTKOLAnoIpuRj8npIQqWM10RxIT9P
zLHlc1AesV1+EeHoJiCgqMJ2dDriD3O7gwVYIw/3u9WlsPP9xZBuHMfwFvSyQfG1hp4nk/7Dtg8f
UHNYbHXcffPFLFklEEXElP9Q7HXGzlHux+cutYFZYBEZu+x9JK7nmpdhrBBtsKW+WSefJ3xJRKNN
zcTxI1eq4P9GULr80kRBkW5CJstszvhy1iqaRIYKhDl+LSZqOiFdUibMNlCPHArJOFjO7jLT0+6v
p4BM5NFTNx8mVB9oSqeR/25ub6Pl2L5Ovo2d3LrS4lvh5B0eHBHh3QKXhRsggZMemF2BRVZKtaTl
VC+dmPZB66ZzHzuB9ySRpvXPusV96pylcUy4KvCVRVWkggfSGJqhN5ory0bByp/F233e+YuUibIJ
1F0brPeMeU6NdZz+yDH3J5FI8NcL1ejEcH1TilKiGsEsWllbpDnKtB7Zqc3toE4Z3GskU4yZnN+S
TbRWEJ7AZJ0vyd/RIhvuGKG8YrHV4yfMy+EpDZNxkpiuVnJpTmziVmV8k/AnHVaCzLk8TRtxUSu5
09z6CaYJcCTuYsG/Cp0MSo1/itWNyqvIHcj9XrLWpiC5WdN6PH/mEU/QcEhD0okd6riY7mKTn+Nr
ud4OLT7OeKVAYOaWvxRIQ6aR5TRoIGCKYmOKxGxIPPBRLFQMgXCUETiZJ/so50plgEJBsKbu9ygM
WKmRsYTtUiKbMBYR64Y9zbK7GuGXIcFP0+09yybLuncNsSMYWCUMSiQwKEluq0+OtY+aXE3LZK10
pqqAH5AA48pxfy3ZcNxYsv3nNAlU44vO4BqV56ob9/LM8nQWAucLGq1CKrQfarydKKOwmZRLRAqm
L+pGk+pOyyiqV6qPBvTxVE3c/lecVH2AnCns73b2Dekjkh23a5/6NJrr9MlgNwvlO2YQ+LlGVNZz
EsPBKBFt6uP3aS4+ZcNiJPdkyfKZ4ewPZ1tdgn7B5YQNJlPAq8bNfzp3VoN66iLbh9482tFXX4kC
wu9rbraxETAQpJCeSYUJCqtDUKvo6hfzpsREbLVysuMxgGT7XB4vQC5L5EFV2WKwQA3DRR81eCMt
Pico11wVP72+6G2mbsZ4GZbnuU4R5/1Bw+wC8jJTco+O7JRdDdAeZHhcRN5DjW65WCotqF7dYCRZ
lNqfjV+MXdHt0uCiJsbusZlZea4BONbBnQK/DSg+wfg9Nc7XvNYXANGjj8wmk3y+QfBN145u02ft
EglmmYvYseJZF1a6a54iXDcBbwWcCcDXuhPHHxcwrytXvLRgo0+ktZ4oIcp5EhWTiuC2Qyy/gtyD
HIkbyqpnmMUq3KmYiu48QRFDp6fhL5zELlu1T6vdhCrv/cxzyx96i2WBNA9NT3+2b6LfmxoRs5r1
ot0bXvPPRuIHW/0XeUBxRgSiw1EFvI7SGIkVQ8Cr0WbZEfeSQ6m2ROnYtuAxYyEmXGHVhw+HiQU0
ILf1Uf4Ok3nmHuhfjhj4CkUPBnceFGqRN74oHzSJha41YgQW7Q4U8ISp+s8qMwFriN2ONY9NMezC
9AiOCBB/VF8NfYsNfXXIkPM6YVwXBw8AgJdTjf5f2T962DWFk6UmjX78auoR1I+GvxBK/Pzv2ATZ
Lx9SQ4KMjROjnZDhINe4G/f3I3Z9e0WZAEowtokPFCO1ipAYhNoV+/KPo9XO4S4myZPvG+zWJ+LC
79OtO9dKEKL2xMmy1HoUFYh3JPp7sedTGxNK40jVDd6UDMOLnJ+x6+L1iW8UCNgSYkTzl/gQYzIA
96B+Q3S8IU/VjOZ0ft7Rr5zTfLsSvaNxSqnI13+jvbf4XNMfrGBto9o3yz/aPEHpJd0o67H6otW7
Z5sL9q7yD7OpwxLVhW2o3RCklxKSKUxCm+58DAymqthGQqyRoiyI/o4lGpyfsHf76uG25fA+gQh5
viHQIyWSa1NEfsBJ9GedQ6QfEOyXEH7DirkRu9frttdGIl+l9wLqCWtCJgVVkhN87ZS0X47ul6tN
Ylogh5d3QBRFu0OhMCw3lL3ukvsv5pohbYco7VdLoGyN0AwQe4J+DzHz01W5D4iXVyGLMpD62HSC
LbDHycqoX1oNIICKSjokjGWGdoxyk9Pd+qh4r0rPHCru2LZNJLzRInMAsDpAEpyDwayhAPuqBFaB
PVoPc1asORnaUJphxJVX19Z5DSLrT8aokOZAuu96FQVsEFyu7PK/9gVq6+6yaTkeS29ARtm2LmAT
CHLctWgxsEJ0HGAZxRxyb8vtGklWC/yIA/ly4RCK7G68ZJS3aFHcv2rrLqdurGaUmSyVfYUITmvE
Fc2SH8hIGG6ex7mPoTyx8+Blwi6BHogbhRNSoDoOW/+5dtvypwhsgRi5WIRnWfmvq2m/xqWKc+se
mHyTe68DFQPjpeDh/uu2dCHB6GdVrgnGwptptXIoirAgbxNgTUT2EMXvlNzb0L8mHPa+qR0rqHzZ
vum/Px4vYcG4M8whVgR/Y9xrnaWZC4m6gRNRnb5FdOytHnP1Rn3vrQ7l7MUjol2VUqHd90MfkNqV
vdXOZIQ8YQDbFlqIkb2vEZXeh7cIH0vDpQoo0cA4SIA9XrfGxkkZR59TNBK13qa22WPl2E37Y7zn
zMtroHDCn7wHcu8MtjhkWxdbpT/m/BTc7BHDg5Nsu+S71MvlHrzW7kmf2F8p80zLC3QEPD50AbCg
+9kn3MTTXUndNJkZI0XCoJcBm6t4l8J1CzRvZmV65aqID3uREc8eOKrr+WFJyYo+pifDu1H4D/Q4
hOd0QS16yuLt6QNm/GKFNPl6uvHbcmyKpPp1Tro5UUbYBOjyt0mGkfUoW94IMITDf31Mp9ksUmJi
J8phPSx2ry66vFWLb+Wy/8D4egmq40hbAWotME58120SJZTtRmoRL5HK3KZrbuix5DAX4d9gGF8y
1T8n/99jRvhoPHeF5/erCYnLdezceGVR3+wEe6hGUe+sNJ2pDrbbd5XDNByP4H3782GJYiQqJH0u
YXRUbqABzbIg17pBizYFEdPsEzJN1sId0AlqiOaj1QCA710oG0BLpHorKoDxGRtSk245qR2Yv7VO
8MUo7i2EL2HzKFFTmMDW3g9Y96rNvRqHdaq3d1puth3j0FgchsvRLK09aN5s/4G4Xcigrgn/a5Al
myqLAzNz8Xt2I0410wVtuAPuN/cIAN+Jp/NA2aSUy71vJ6fOxx6m5hsnN4ymjOwxMjckqpmgSHFf
9V+nLEne5OrfxIVxCtGmpwlgwUnfs5R9evevu6mY12hAZ+G2OurCmT/bex7SXhhGwdhF4QlkcaYr
zvxF7s+f5W/ET+Rb7uicy9tYBPjr/5IClmUHRibiuPqs03NpaHvk/48gtjK47pqoQVb/Ym/vSa6/
Gy0ZgBRvSy5WXsJLtAAhGM8oKhIUW79HQvBw4tGv2qck7XPCnYEThcAZHCiruX8JAq23ye4oqtBc
sYJI3SA3H1gNOpWPcR0pIacl+IvLNkBZTirngzVyJUtZxlN3UL6MELVn4FoSG9DEdd/CdkhvaRQh
uhSDSjwxw4vMba48F6f4ikXUp2vw9Mg5XExT8557+LYF2DD/FYI51pQ1kXAVXh6FLqcH5xSGlzP5
pZpgvajT4njJKFy32cfYt2bYNI+e+y8F/o34nZL8RqXKOp98knbope/LZHRhftFPui7TCeIWu9BD
nDGlMEIcg3Guhkxp/uJozStVyRYeSstVuCPEtffKNtFWaT5AlLwbogbXw1ZnVyGQnD0uLwWOt1Kf
/DrlVY32CkK/O36b6WoIdiqojK6xZKPmFgT7ZSvquHJnsczJazemw9CvE3QwtobF3KQ7LYUhewp/
/Zce5ppxCrlzOHtzalBhDw6T1EqUQbeWH3MyFnSo/wLPesJOS5RUVT9bp96EiNKLeN0hidAoBKxE
KGkmsk/xhKqsLgY6USlnBgyWtXCoXUU6DY+mEwfB6KGlkAQGF6QwpsFUBdanBSiLgoOvqK+5H/sH
kRtui8C/HHre+vIAXFpofU19oRQ3gGyoQLeTUTmRRA+xkVbPCHh7oEoO4AlkEPcVomTcn04JwgJz
v6W3N/UKu9x4B78VCUmUrbi/yz0GVpMbZAioJz3asH/b1oblJe+cmwhsHz5nWRr0kypF2LirQSEG
4ZL0p22MIeTop8WLWtu9caX4Gdpx76ncpW9sBjVn24gJmQ98ggq+zhRWbJnHRZVyBg9pqVPiPQ4s
QcMHEc4jvYWHCWzwTuM8Y61aXpNx6InkwJSBQxDuwsIae2igqTxS97NfCO/5eBIsazxH0X1vDILX
2Q4ZNgHJ/TyIkKDBK+qy1zZu+ApbCj7Q6rqqUWMwlgD446gqj1xqFPjaRsDzXPFuTQDt7FNQLZ/F
gxb/4jBmyxg8cNPMhsY2dsUtr8EwPO0JF/D5KO/bvbD6Vzw5nqXBL1iGJC3IeHdyJsGYs/ppouQm
EDs5CjoSsGFdPPP4NXD1PkuvizaMIQ/W9Q0P+EinJdIr8/OQcBAgEqZwxbFxAeClNfN39EbJT0JL
ISh9BWaMAtSsECoqjl1KC1iRnvbiYi7+phX5viHxP9YyhCjUV0F0BeolYFk00wm6yfSL6U2tSqPA
5+G5EuFjkoqTSG8uWzCosKT1WSp27Pl2H6ryjO96Lq+3oLIt/G39ysK5gjBLnaqEQTo85hKPEazX
/m33z0+Pd97p8GydP2zWqQxVNqGZ0/fhAOXGP3BurNfT2gouLNBsQ22reGFzgJ+e/PIBp0C1HxCG
htsVPz3ouK/KbEzpfv659nbaYAgzX1BLQ7xEcBXWSrBuU3GA6x0FKeJb9sqPU0leMpmIEa6SoPH4
VUC9QlMkhvrMu0xGD3dh/35z/0wZuivzz8+l0hF2Rl1D2hpfU2OMqSKdVtTMNN0yjnW/Nxpom45s
HCY5uhCWyBMtXnClbpslQdYN0lIV+iWrek0OtQOayNr1gotwRM4UUxR5cRXtoYI6XSMxwrmhCS4v
Ndreah5ewkE7/ljw5ZsxUiLJH3bwzd+x5VFhiWkY0hMzkRdxQmsg3KiNEXsdMzyKiKEEuZJ5OB8y
LbrKK/jROsXcLZRWdumf8KXZ8McAquu8ogufl5XR0k4jVFSidwOVD8ogmRkmytUivl/1/m39jmRE
xwkOkq1pVKX9duU3s92dOtFNeA59LSgO10KCm3KEwBkmf5b237BnpAuSU6qy3SxnBuS1DdwrxTno
IIeXN7Jck6M36/4m2Qav3RO90BTdIJ2b/47ZQ8rFnASWLNlTS5besifLmxH9sLsnIVCNAQXkDH+n
HVFGl/AHDzJplH07whDYouSIGiU60pxazD5x+O9gS++UW0V92H5cgy1eYuAMF6w/zsyYHqM5tA86
qwAeysRUZ9vk8msuaySPpND+J/wEKN5LMNHOWLN2VADA5fbkE+hc9yhXZUAPgrx/pqCqssu1D+4c
XaLzbeU/nQ2jaDOOPe3M/hoKjMwQXowRok1VpEO3XhKAg+7ZSPSRebvyMFy2farVAoUZbrDfO1x6
hR6qyVwf2QL2YMXwTn7VCwV0aj7cnhPkMVK8o4HOpR2NjlWOCGS9P2tGNgONysrz6vpEavnA5eBU
bYrr9nGzuh6dM+IHFfWhHV3moH0c7+LG0JOmg8xxan3tWGsPA8Q5G6GuE2xyOC8EKzeD89YprQ/G
uG1FpSx9zHPUW9mAz3nGeBGj6qJYZB226J9CsYFPWXrRnAoHYCpBrtyMtgISwMfVXayQj5diXafN
5aMJ6rGyCEjsQCoZAQY8HqnXwX1kHJHY7T1nwjOWXM9u3wKVbtPwb9Y7X1ABkB6BgpqOPvzLASKF
ULx4loJh4NeBq66l2douHXE3DoWvPVtpeCXxZsWE5gOf57CSrD6aYooMXTevXb2YsgfB4pjx60+e
n3XMLadP7qKcncdhkc+ntgI0zNNUrkt37Es0ajKix9kuYoEd+XjgQZ3GgsiWm9VzAwRnsNqvk3zt
kd7g2w6RhRaN5boXxrW7zNPmmNNkute11ZaEqKSFzYMWSdPb7tRGVPRfOoE23pB8aWD2TBp5uLnD
rHhkxVsjCb/cr9I6xGPIdJdGm7DjeS2vvGAgP7ep4qZspdZ05NVLrAB7ZCyOzXL9pTrhfQiPGFat
AHFsXvgs5VnK8R2z/6UpccagIL5h9Z7FwOq6vubQWiL2z0kLqtJb+hEWD/QtaIfSNMbRo4mJsb5S
o+qmlE3foQ2LQe8Gn2/b3woOlQxZYL8nmwGz3Xl5gKT5CrzYpBINUvH7T5a9En+jcD9kXc1RxlJl
ZSVwz5uJyKJ+97eucPpC8dedWdWVL/yYr1ZUpMh7r3FrQGk309qllApQtszHY2GkuCZz1utJJDgB
cOY2rXlgAXFIhF0klEb7qI6A46EYRv5u4ONW5Pn5jJjuHBqdUDoCV73sKrw8h0SRj2UUFDH/c4L+
LV22vpEFHY4nNbiiUqjjlMkpWnTbdpQGhHw5XXOzrIkizGbgFaUTzzUCALUSIOtAm1RH+b3f3Ry0
dZKzlKZv5bRGAwWgrXnx+7gTLk1xPCKW2UINdJXviCnR4e6t0I3/DjZXD03x7zaqeU/Cy6YTnqap
UV34I45tApCe5PaQq3m3WGtQitMQ0Fz6GmCel3351KBM7PkbUGmY9OtlabvBA/0bDxgVJkKsRlOc
Ln49tsiK92KuAelLDmXZUm2L+7r+PkQMQtJdrvrNYE/wGEHNiwBMYExMzPYLXp8TQiLuc7pZuT4c
t5Exw5TirU1Vbus6DwsVWqV2E26xSkzyB80eTQo41o+3/lEwba1lmSowkBGtG5/jIycWwlYk4w9r
gfczbpFZbvOlFkHJm4DN5TKW5+sc54VoAQ3UNFj7a2Caxx2bpt9ZxRGBWiSrPAgnM1II4JT0V6T3
pHQniR5T9ScD/Jid7vbc7W7j08I3YK8v6haiBEZSMX++4xh86yAlN3BgqXHu0Ql9/VvdKMFbLa0W
uoDDKP86hXAQulyhs8vDMdTZGIJWOJTmo7V93Z/HF5wrjuJij7ufayesLTrJWtZTrpGlSh4T3XbK
+g5BYEdiCw2Hyx4yCorU+F7dFCvxHttpz41Bx4q2AO8O6gDcyatK1OLWmwz+UdTitELT8P1zJqvV
s0KQNeRL/YIfSQpR7Ezn9HXcaLpkhqKNrsb6fTFrSWCWktQ8p/+PBKT1gZK7hllNIr4QgTAxOEr5
gvPWshI/uSJisZ4BanatJcfOSVk9gZjPD+rb9bzSiZ9rA3CvCe7zZ9OtU7rcKe7ZT6tJAQ4yGByl
giMwzfM1gZEN/vZXp9bmEtWJNdL9spjMLPrM+U+VAZihmsN2Y3pVocWZuXxGK1gc/BRx9WJuJvtH
JCQPwpfzoD1oiOpk2xaTI5nLvDG0RRnDeS4k9sYYPYOIVXTiwZV8UmTa8OP5kudf8Wf1QWSaFDgY
uCJK76I2PVG9b9rxeV2duzc3OZpoq1gT2MjAw3FBHl728E3UPd4Qz7Pl6pInS5Mhx4ojxk6FwkGI
ZHt7DuqQKhY7xAPgVBYzuixo5RhnHu/fgccRcW1bejDX1uVIgIrS4hDKev+vqZkLA+wHeUDNNIQX
nZRP641Cs79sYWuuz/SjkyeSqS4xdBoM+Wz4t/sisnrgzHqN847yRBHsONg6DT6YtoThJwW+ytL6
vh+szqaQXJAqgmWSM5pzxT38ZOf11Tqw61XKm4c6incVw5j4CCBqh5mT5Qqmm6+N56hhlFaTZO6N
8OJOkz/CGZyWCetCI/s8qGsY7RY58GeF/N+uUx5Cf96ZYTQg9vqmcax5bGXoHPOWHVSJV3ZuNoH/
9mBnBmZfTiQhrKmXgVwzt0vqDCki1tE5jO1YPuYqdG+6hU9lvxMqdTBXaIP6Q2AJdNSwIIEoenDw
S05Ze/4yho62oHEZGfF/+UqcpNgyQTDDiqQ+l5Tmdd286OchHd6s4LjsofywJxwlcQs4X4+2yFLq
i3rCpBmZQwtDj1HR7+U9MJCbYxBKvl9pwPMEXnJN1lqqBNisJdCvxBsFQH6j6UKZOFvEVhAaTROz
KMv2L0mu/ZfFjbW6NWWutWaGFScpCuBR5/degGeSBWAa0FioAmSa8IMChlK6jh4++i70R09BBvkW
FvGeFfCFjLes0YOOSZBhFsM3qgIBUCDGAPwd7DRMnbn5MAyw8n7IVs8RubNZbWmst8tYVsTrstz+
eh0zNCIiUzknnwsLQ7NnZqvr+kKi9mfrszgFNvqCzJD56CD3rhoz/Ldo+JnpNL5Ip/c3RV8ZNwG5
L7pl3zpkLddO7/dN+a2OMALe/Xnm9Wc54YVZkJjlN5vIbeeaRia0bDQ0lCU9JBEm9z3sYxR4aXq6
z7Ih6ftXmhPU1HL5xlqYs2DKaoAY+Q8p4nZ98THO0mbyPHK2qDegaHM9ssY9WT63fbbHdus+Ncoq
/6K/pSQVWRDj3D5Ire64FWmAeDSqEB1pACVIgGtlk20dwu5AIy8IyPHpphZfp5dQnBRIvZNUggpx
4cxEX6li2MSxUcgtaHveqpPNHNl6YsJQI8+woQaUpwveMczezFvFwnvlGpB/cpOnq16Kk4Z5eu3k
xMzgPXB6Nu5TI0SUbdP9eI/1nLHYLKZU5zAGZ14ifbMQOlZuPHQgpfNEaHkdGCdJsrNfWXyiWBGs
wnqfXzsPcAXZ01q+Z7Oeinp2HslycKpcoMYoq//3AJ8n1wNwb+dNPfH2GiVXUagkeD++u2rvCF/z
eCjDRtWZOD4caF4kxOoAkbjNOeHuJEpduScP6vIg/tLhHKNQ3whVoCMEek7odDi+cs9HYbEgJ6xP
I1u8BlOqC6gzSgeuhqW6mLgRjHBsEbtkyryEvTq5nvjnZK3vgo5IvgPeMdnvuyEU9zk3WRL2jLxi
oKmleGYvKQ+qoigxCxNnqtIKcjGR7hgLczRCajwg096dVWH7XCqgVliE2mHLCUlm8aJTuREkHmfW
8+qEeFKySR6iZiup2TugrFqVZYZzjDzrAbz7+R9/6XnHwJjoQnu/wNVhyeFr0zPTw5jR5KhkyXnx
Ww1BTNlF6IQAicnETU/ERN5supRtYJr6DpJQVB3cr/vVkjT/318Li3n/S15n5sprvGDS7Ko70nNK
e5ar70GeEGmeE7G2yssoBn1RhRnpZN4rHsm66Y1OSMWsNhIPdJPz43TWt6q5PXS/sGmIj5z2/zL+
dot2WWC9JUYO2V5ggAOy7jrZSoTm+VficKLvYKVFWzE7VJUZqK6lp1K3q9GW1D+gRUrON3WgNrZc
NnegvW8HjaTo64GM35TInK7z6OAABwd4XW4fYLx/MmXRe0sIZKeruahBtICUTXviWqv5KWDZvZ6e
E+QlAawG3CbESAaOke4JlW3sVGNml3srxelVevjof1FsCZYpT15V9JFTldB4Y5L3Yd92IOHHKbMI
uhMRiPAz2KQOlWoG7BsL+UNGzjI2gFEv1+tt5MCKdbWlBoKb5yKUollpl7hI/de6S63LTL7WySkT
sAgw6FtXzBXcM8FImEwF6PDufneAhAqfQtm2I4obF1sG/UEWx75zw6Z+BOjKLeRdsuik1PYyylgO
DuM5rl6rJZNbpIW+tM4z1c5JHEUqM6/fQtlZQk0ILG+lCHNLt9O2051v+iRdsOYDnnAbyfjebb/L
eRcNdd/hS7ae6+WAfJRFbWh9L23FhC4nVxcYb537blyCLx0kkjXEcxJ440ciDxxmUUga4fDJyn+O
sTF3Evi8P5hmrQVSY6jF3pAFgIS/b5IHU1Fm2sis4Bq8+DV0715L3ArZbcww2N5E5iAzZOA4tR9L
Orh42nINBzDGy6o6P50KGOWqA+wo0oACknH4Ai9JWSzv9vv3UARwMbx5Y4x4ACK30kBqfLr1Wtnm
xUWrfTJ95Q9PQ6vjKMwT0oJwQcAwNeHdfVrxm/6TVzK7BCFPukM5xDhkHUJuk4mPlYjEnSluJUV+
crFTFgfa5HIFGjvlZJ0Th/CFbR54//fytowaP/r++y8xmyT8+Airp7hb9T7mRYlu9L00K1mwT0yo
oksmuHueSnkS3M25GpNOTWZjuBZIJJveJWlqh8CIcOnDN8JOjVMCfziFqdIXdTAOEurAePY0tbTJ
tfhgwiJURkca3ja5ZzfILBYqyOdj/YdTgNM27eB7DVuT4RKHsA0eqLTnFwUDFDZAfIy+R1PJWtji
xpZ5u3dEX1fVY1toIcL9rpkcjJfJJgXNSo7ZNAcN2P4wHt4Ggx+TFAWUFvWllnkxySlKMpMVgJ0U
TbGe6uY0qUNAamZIcMip6HEmqTwe9Ne+ehOSPPV18MiwaOaFVtN2JMqKCO9sE3YS89+k9rnBdcGD
zWBzI7LNa0P+MIqGDqpZqPYFeM20oLhscYS3J6v5wWxxgX3Hs/z99B4591UevwlU8wcXCrYr0WmL
vRqsYh5AJ/yiXBKGAdtC0haVFLYxlJtjGRi1NGljpgzWqwUzvdOQtUGjQSyn15bqLMByX5QrlZdw
hekAeFuhBNeYfJBwfZ/4Yig5akcclW3H7gz2bDN5pXrmpGAmICKfn2dRa4iYkOQK0OVbTuWbvY0j
999JAo3c3qXdPJXyODZd3OY/QM/aFeVw/gDO+p4BfjNKmwgX3DcIZHo7Ya83+HgDh+4h1kQSQ8z5
86lem0DTdYCz+kBe/GP4o+dbOpGuWPtx83AfAhwC2e7PgF66RxqcgAw6Zh8mL5MUuCkm3qCInDQs
fOigRXxPH5wq8uKHsCby12nI/vtTUc0pt68vZ4zBfoqFrFZkvaM4bpAulsN4GZqnaSJCsM5OP1hg
yORo5sr8p2lmyoGeRAxGr/9D1icYBxoa6DZVd0TerpugvFUyLUKkcZdvTrN7Cde2R9jh6TBxa8/b
VMpFrDdMoRUMEZFqOLqdpeCfYp9EgnXbY5mgWtCVNtuZaMXmFzOgkUur/6keHtGaQoSocf1P3gLV
3Ls/jrHN1SjDQFCq0yIzSSKpNSHOqrdgb4pEB+6sQG4SuuEmTb497ze5LljXZ0OXE9z07AdfQVLa
aqjY1oVwtPlUPnZirhWfWRDxA3WdS6avHK+0uhMxYLnUoc/G8pYMXjFU1uLh7dJ9toQMq1oWSapg
dDEoyPpGWblZaLdR8qexvkCaCu2TVMrXCcyqXdcae85Jd577wAGfp80MiU6aHsNLzE2jo/miq03A
80hUWcMVPJ4UMbc6gptgCYZA9pDT7M33PFZ5KXd0n7KGf3iiQRzuU84yCt3B48dPe5dcdm0IxPq9
WwsdpZSz+axeqzBshaq/o8RKlN/l5nPQ/EoGHwfwYVvgA4jmR+jTdmvFc/lqkjOefS8CPiUOlWxX
DSckUfpKKBK6p/wDS9WrDRPi8AznkAbWWxphDkMEOHGiiYIelM0RnJ73/Y11RwwrN9IB9E2+Creh
Vqpp6wiY5RkgnhE3elab0RWszGPECClbkxWQffqAgxJiP4VQhWDR3GqJRY+P1aIiU5Y6NjdH4kwj
aY9gNCuW7nx6nBRg99Qo//IO4oKwzUF5jL8kB7F59C62qG3eoURVcceqAFFQUkAeohSCSLWzd7uj
0g3f302jPkBHE+3LRTU5a5xL8g5LDkuhNfXa4YqCA19Le/lEAnE4170Fcgc/hQ9Wcl896rs+S/b+
b/hVYG154zTUUErwNPhQeQTI+XocvD0gmBkW4oq7a3vu1VxROzqbmsS10lTR2JqbmJZ9BumivSGC
hz/9XaG0D16HwuUZhGs0xDyQWzNH9JDjgivaImdIdQRGNVMVc1NBkuKExqYL6qMhZpx5r8BrGMm3
5vE/nXyqCoy50U2IKvU9HNJRM/RVQvtSFGzG2mff+Gk+jaHygK6iEZrehAs2Mf98DriLhgxFICdn
tDh+OMsPxR4TfgIaMWW4oKCO/K877tzVQ+YtxN2x6k3dCwn//zqi5WZUds20uj8uBMAmzRmbncxF
KzQSckaRC6LKNoVh4SIxAwMi4Hk1tFxvFawnZmfmXWiHM6YmNFrjIcjDayfY1CDXb91MKZp88KmH
PkKxuhcPwjvnqDo5xxGaJUugfHGPqjTa2+1myZTRwfDjQS97phOkeZWJtingqtteslGzVrU+BVic
modL3AvZcQPYD5Gp+4R15Cn68SFY6hVZxHUJVT+Ah993iDlbbkKk+UpVI9Eb8Anbp7Pm7py6dh5Z
Ah8le4svf5bmpzrmiQ6ct8HRez3+xlM37hM6GedVyUjZGgpldo4ClEx6rsHJooPLA2VoEglWE/91
55CIMDK9iIbYUn7slKqegrBmImuErvn5bPdDBPmp8bDBOAM9CCFxjy1YgYdtqjZgR1bli2yTPHZv
1KW31b8NtT6ynqJmIg3mJgTzI6/63vSEcUSliqJjcStxIiu7DB/q6gmYw4XCwlqTeGiEmOPIZRJg
3wTRuAh/wqmdHnn3/tEJpxD9MALlyBxhw2V9OMHarUtRu7Y/8lJwitU9PCGSw+p25ZNWFvqkvKy8
uERQjEqQzvoYyr+J5QrJ6Vrnd6WE5VoxEQp739SU82mzyBv8wBXFGvrxlCxM/lqC7+7MRzjR42hi
8N0XBfiTV3u5WKT3wP6RkFQm1dOaIcjqa9YNBYRl3jLmHAA8wU5Opi2wsmvJbW5SaL6urd4D0hnx
XN2tLhkE7pG2f4GNn6gLWWChHXvS7YeesFUYhhetNm7CmTXr7PWGj2p17xEUNMPg1Dwrh30vS4I6
romPB+OK8F282mPlqBVUOCfYfToD0hmUQ43j8xD6rvFly3T6E/1gei5LThr2srWyeGzKxfA5RBdQ
+wK9kAoKG5vv/5IwYbkDMWTLf1Q+HgegxXMlY9pFjFtp37/HzYB0nMm7BuB86r0C7/mttgMnPFGZ
8xvr2NPMo/1g1pQ9ScK37JGHApZAeDrKBA7SUHy9ghFiCfJehH7/4wS8lGU16x4T/rurZ1EryfK0
G6GkYqRbATTEqbK5CoQRqcm/NJG34YARtViItDuosOMBmWBkJ1uXTF2e4o1zqEk50kYb7CWJOtSd
WkIDKdD2eaC5Hq3KX1lKR5/mFZaf+VlW/UeaVVZLMCCOCv7nWJBplC637sUkwp34ZQOrKqaIw3NF
Q4UrigxKPj9M4jddtVmg4SffELuYVKfzcaFGv1x6w4RmWMHJ8IWdetTJN3jbh6sRGCwiRHxunAUM
inObjO4wtv4LexQPSpg8Pj5pbthAXS3+rhjq+HStwCj6IkEPUN/VUDv3oNyH+4BThujg1gP+tP+5
QrW4rfxOdQJtmL1DdMMNDPTOdOiZTdGVe/t4J4zd7cQDrn+zDBIVCjgxli9wVroUwCl3nvjE9Niu
r0LvZOlhQYylbEXf2FvaLaCifM6HA+EQ/TZnKwy525H6SgWwqijvh0w1OeOedOnS7h4wMovv6hK0
QOxKh15Luoc/BjA33DTwqZx6F6BDu/1o8Qsdf5qzzxwspdLrF+0gaVPnXtr5u5/WwDGyHTinhdQE
BLMqKO5ybAGxO6tFD6o7U0we6A03xoxNuu7E1xzNgadZipduu+TF8ESVbHoLJVT6XvUHGNM43MRj
YaK80xUVe6zFhQZq164LiN35zJZSEVEs4yhM3c0C/91edpXYD4eC8Sr1LIX8YcqvRaHYze8u1w5+
sTQ9Xv1ZO6we5pdumOGdpOXebMOLSyXi4smUD1qb2Bbf7xB7kTOsjcJL7BcTIocufj2hkjGLuJW4
mu/KtKAoP+tG79gQYek+eXSYkAllER84SIeJQJpKaR5Y0Qrrs4NZFia06F3IMl8qSeDX89ImJrbU
cIsT+8g7OHzy5keG9aOa6lLf0qt3foGCGmFR0/ua5nVx9D7v8d9993u4Vz6fBQ8a/R+SnUFGFeBm
RzvDh+A1jl6//sSPiytDeiXbmxvisIDLu0Lp989UfetbZYsqb1/ULq9Mm2255+r1C/zPQBR/hQz3
6nVuOIMKWFsXYDdtey/hoq1yFezRfpicfpZxyjg8AmEha8dnn/ytbu1MLwbwQmhTsd9lrZ2uBkzo
BygQgn+Wn7yMwTu31NLGpvPFweABdBHULsjZvtEjCRBzlcPaX3UgOXhsoALuFZUlsf+nmieXRItX
BZVPLgv99Qx4QHDnovonluH2VVgTKluWWpWSZuqrnDFv84k89cjNmKh1+ZwNEknMYPQcQE+6ttDd
b/hY/YAJcrJafKcLsx8N/wBDxzLviAoq1ifhXrmd8vnZbxPJNLBSimjkO01ZFHlk7dOkd/00RA3b
MLyMOGmiESdLC+AJ4DNCM2dMjPi7AK2fyfSN51m+h2fRj0pjPctziLCFGdBOQ39FEJsCkopmx4om
lm80xDj06gY4LMwBqguvyRWt4jAY890yz2ZmAFscdcGZ3Dg8/JutdiBw9QTlJ70xjrupiiIc6z5d
TTy6G7xoQh+d8p/A3aHQ1AmeFbHeZr3SLJGejWOhQ8D7+HJJStexFDnv9VtCFJHNj08lugUFgXrl
TAiUyiM5Jwio7nS0PORJ73vzLT//AXWgyZtJOt6Tq4/Dyk2Np1/NJGD6+HL6x6KvzE8o99DV9Qto
/ZgTm8VNcEDUpyhXpfw/qvAeOqEiA2IBQ4ivqSYdqIUb63b/kcE3j/+v+Ub/C3CUb5FH+9KGxJFS
gXvnvD5jVpw/aUOVYyBEv5GxCFBPmISx/l3xzXnU8xVD9y7JLt2Y84PbzLk53wk68Rt1OF07QW9p
J8THbpNrWUZruKgPP/8DNKD0GrHF+qLVhp+AD/KV2RWbsi8JR4aalh/Ge9Js60pnYxGe47LoqbWr
PvYPruGpbPlmZjOFk90K6YlqUWrNi+bwSxNZCYTlQ8q4Dwbxp6oBQjIb2p2MBDPJ5Y+liAEyJb3R
RKPy3IIeV2j0Ht1rr2us2Z5Fk0jWtyTX7WPuvuKuTywAC5JnWALVb8Rs9YmzSOv9k/gr+Se5miMu
Nb94bKLqqQ44GhgXZXz5R0Rbv/kuQESn3bdRqxaFVC4EaWXefMhIRcmRlB2xy6k7TWa1MSgS76RI
/zEZ7u/1INZUaADX0t1yXp2qtqRzhjZElNrcg/oL14tTBvc10xGTRT8Ri+ywdCqUQe0TumMaLyWb
9zgH+3q4Rg0w09IHo/EPxlNh5XooKflbZA7r06bxxSHxo2jEr3pI4cNm2OZrCv1oxc79m9HmIXSl
6/P0a/A4M1uZf7GIGaN/M7lgvv3kRWChUUIIkp09/Pp0ynDA4Xcn5vHF7tlVd0spLAdxZg1MKaBH
oRLeCiOcoGNJwnF82ydLKnH/iTsg+kgmwUoS1glq5jMnd4xo6mFAdwAw4kb/QS78KxbJLcISpgSH
Bftu2jVRusgkUYvfBr6kbg1tEqEUfpT+xCOKK2EdhY/6dxO10WKLew6bZSbz0n+ON3o31+R3S3oU
GKMnYhBH+KlJxdBi3UQmOCpOC5/JzP/XKXIn1BkMJ4LNUvGyyGXQmBsEem5PNhVg6pPOGX3C1soU
mYx+EDdvzBPPWlm5lgUGEh5f+wT1M8VsfUYZI4JMEdpfm4eJDx/qoZGufMR0o7Vow06na16UND1E
hTwxCwc9kbaiJSNOCHUKCCOXv4N4TC1whlOO892CHVR4bT5hKQczy1WF6jNjRwSD5WRWmzvl4SuC
8pCUtj894iByLgJNq9Ji/sYWRGSTaKpefZV8ErjcpCAVp72wve1hEgwFaxKbUO3Q61gg+Rr2Kg2f
V5JWx+ngSp9KbbkXlnDAlxZ+EwjTux8XJQiWC6xaAJjXP12EWmmpu6nMjToLuuMwr4bnzaMTos1i
KBGk7ecMcblGQH6QUEZn20R/W/vZpQZqjyOK8lroXeitAqO5b+IOajH3uuzAzxu3l8ZFhHraXnRS
3ogq/g+cNho1EnJy94PCBAujQyQfkL1SkoYg8r/0XcA8Di7pXF8U1WrZkfInvENwUF8K+nDOUmDr
9GrkVflAlXvr8lyrB+WUvQFWL60rThvXF4bWQVAm6FvZ7Bot1Oz4AT58zFm0VJwM3Nj/UP4bYswl
qBEPaE73uZk9sHArS6LGmHaAcLDJsykABmcapcs2cI97bk2YIhevnxc4upvx9zzI9XP18AweS26J
NCW1bR3sCGZtzTfIT29BL0Qt9JStPA6FMsxMmvfKfiYcZGMDxyuS59dHcpJJzMQ8ncODUbjT+Fav
j5CFu7RmvAI8i6uk4GjODtu/NRsvhLE5aTvKYX4Vcd1TMVnkRiqGO2L4kDtH2aQRDOyhbM/LIa9p
fK6h3tG+qYL76sCt3sET1zEsOSbcNqF/W+g4a+ZIgYbpZHD3WUjqPnx0Xydj8kZua5uPAVdttPSz
EmdIPGno32FhmtCQ9Kc4nsE3ns40HNyNmysfwxYvC5Rutam1Jkdo80g9Q3hPVdmXtBL7R//8f1nu
FueqN8FJu1o4d4EwN7FI4AKQgQTSD8JSeB9QTBOq+jNJJKGYrY1ho7wEw7as66rCDWnBU3CIGRbv
CTLsIcJ5MzgfWY3VzM3gLKlRuKZ+xEck6SkSuEgEafxoUHVkaTMY8+EgjM84S11YDA+xc1ef9f1A
sE9XiwHENoFQXS4bf1mBDi4bYgWmRPMaLQikZR6kfykfXnQK2VfuPK0rWTKDryz1JiIY+9yCt7Nk
1+zDjegJmwVVaJ+Il32+5WyGUZpU799r9Y6FQOanyFF41EzPZRml9kCj7PtGuEsrjIl+rrZ/8h37
ZuR/BM0MRq5PkiYmM6SpjOUnoqRl165w7oHVs729rpl8cbkciKKQGp0YSnkOx3WtgzJw4AsCF1ne
1z/bXi1Whc+B03kz4Q6/1a4KZ+FwUglf5HmWxTEKCsa+fDIaao931wWelMNCYrnT2WTStEtYp2gQ
cvZaJmbTkl6w88aMOggFfxpx5dcT9551Zx7OI7fzMeSrJczEHV6XqHJpn3frcNa+jsLtfzDefMXq
ajycvA6RAQoLqLd5PTmqQSDZW6StwsRNNDcuLdZYcKGDGK+M+vP60NgNx/cVqWFg5odYbDqNnWje
CiSXq6W4XoBhj/rFCa6DqEXH/yyrmPKq2x/pXA8d6LY8eB0JGk2o3lc0hywUcut/24YvR9x3HgBr
/24xIOvnl3CMp4L8nAVn/YOxGv0R6T3f0yuPmQMVmG4t334WKbh8yQCAVgUX+Ah6hULJDogbK7RR
cmyIWane2pC6NRtN2zvAW691Gy5SXPYxqOUPTG4TrXZmhjTK/m7Kqfl5PMGfV+aKaDZgZWy4DOca
8JQV+JTsrHOrXAW6VZmB/u6PFK+pclsfblw2EiNJm6Uyn0lB1N5dG3TiLTYWJLA8IpIjoKwA0f/i
5JpAjMes/CVJMBFVLGOTGvKvaBFKz4KMxm3StdnMeWOczJAtnwXRXmcT1Ory+jiJDqP2kpkWv72r
8NnA9I7tOTGl6R4QsPxjxCPObfxpNCv3+vkkP5O4unQVQPE5P/C8Ixv+eVo7d3bw0CCGyy75YlIp
6THlzjDjkbKh6BB6m9lURMHZwlX1vdb/+/nRgd0RcVF94JUw0syP9+4opdFeIksAyff6iXdGtEHi
4AAqhvJgIFCAhgUDqfLcOghF22UfnIiYOqZgSwCHBKIxgiqNQ1weN+x1eZyTNb+niQnR817eGYqp
F/Ng3DF5wPEpKEh6+ufbDxXbx8nEuzABd+uQJbckTpQ08nSlUuvEGp5/HMdUp+apEFePlWyXbtVv
+ou/NXHKaLM4n6xqQWP/eWYU5HQck895RgsPaZKRl11/5PFXOiAM5BXDOSiT0QgFiYQRTJBbNQob
UbwMPY/mrtb2g4EIMqNE6uwlhyZ70vFk6GDXtQKpsQAznjLlAQ4JhSOm6vcx36vEftZStaPjvnKL
RPee3alRtUmNs5F7tCDD8DyhjKPC9dixM33pKwXYUBmENEbPWyPd9m83QgEpxALegMk7/AFoDEu3
0j7quUILYDa6oX5vCaHgdgtvdLyh1tZ8QSeVhWJfrjGIsGcLJR4eBKsu9LREslBT87gk5y+pZh1d
z1zCKm2GFWlRsr8YJ76++/xES8rnp6Ts7MulAcxW9DmRzc/0bEfh34LYRtOcqd2DGbPbvHXcbUsn
wrlk0nlK7tVN1TrnLojpdj1HGGxXyVcsXxVfCh+ZO2oj4+EKEKtplfAbl8r0SCbt3RQ2uvxJocAM
Ls9XHEtHo1iKcwsgsTRNF7/gKBZ6Zqn/FdublbFlKj8gVbo0v2qvYP+tw6lc+4G5aN030WdhgIsJ
VeF0rmKrgDIrWfrDGLYDzCvehfGG9sDAqI2FaUaWOS9OPQpAiuj4LVpV0CInBgx0yQ9D9gvTEGoT
UiRHSqxLeY+mEyE3lsdv+CXbmj1vnLxrwfbUt4T7hz+iiDKdSinlgvGxdn4Ll/0olhfMWz8sEebp
TCzMudS5JIiBzs0x841UyHo9ybJhMx0NgN8snSE76u71WhZ7SeCAgOAs7+zu5prjF4iwBenBaUs0
sTdAhaSDsEojMj3g8HPdW4VBGpVVdYBH05JxLqSn2V+Pl/xXflI/mjp+Who+/c9c0TZdv7qrkXDN
y3/a8TMekFgon5mhk7XVJ88v47eBQyd7fCjFC48gjeMBMtmwLAp0mY14eTVgX3P1O25sbCsMuAa1
ZgeM1jkIX01NzZw+TrtNS6PoeyI4zVTwq3+pWaeS+PlHXOFHkf+vT3CONg7oUUdWpDNfumbQQTWC
NIOOZnRq67cd98wfxivBYLvGOPR9Z1RwP8w0+onNVxZ5ea6THC/Ul4pVWxDv7z93gLFQivuKg85m
qApQ4ifjIGaKqvVYOah8wVpq00HVOg9GnlM6hXSdwJNd20SKAy9XlIVgrlZ1IHvL6v5OZ0B31YoP
TrE3wd9dMXzDk/UP4kwMK7j3HlRQ/QuhfdSde1JseFxkeMu+q+wkhxeNKXbyOb91046zxZF2Xsag
d/RFpdsqjQLnblGwtdfkK/PmHBYhXFjO2+wLJF2QjC6zzRLkCbTFzoRFFNEReVcK8Bh/kMane+5+
2o2SnDiGP8/NWyMgSglopMGlvbWgxWMqB9MEknvqPMhaXpN1hqFkhtGwidDN3tS4o0EiSLXEYmoV
17QyYMHBg9viBYtM7kugFXzdcAoQkx7FfX65IkJSLPHvp5iIzN5WgijbeoocPUdPyUkSE4lFqzZU
uNJLSWfzpGR2xFsJHGCtxbSgnqtFW9gXeRGW8SnysdAf+tFwgVxTWNpbfgDHcaYQ69ZtH12B7xeU
HzEh8fRVlDhbWexerlzR+EG0RELsyZpWtfLo7jeM6Byh8ihRClwlrSs4sgtQkHqku/bpduSq7wGr
M38eeaXHTDE5exVIOlsLPuZr9uzXJoqn85nfF/mAH/NGSBD3I29RfLxaWRfVmyMAxEu6jwVCPaH1
7pv9noIXQfs3a0Fe1uRRrRK6pEGYgSFO8+3iPbV1JI7l58llLNziavod1vc/YUrcoCKJ0W+xtCHn
ShVkbim/s2+ZTlMe9+6zc/EJry4R/HyY+JqWbVGRNn/dksfbT2a3A3LHnN/Mzzd965PCQLV3+OcD
8xFUx/xirl5OdE3Z7vRoh8+2+HoDNw1AdgS1ALI7OSRhSvnlCQ483haWVCH5T+LQyVyw3xyfbP9C
Ao2utY2108zBSe5fKLnaZIDWbsqpM1/dv5PiRyAwdsSGXsUCNwjrWzlSvuoCJIi2Zl+VLOB3Xt64
s1PgMxmxz2L5lmTJ4gbl5k3CdvdwsZn/PpJY8GRXllwQsjYemLNoalEzPI83jQI9joDgoFvRV+u4
y4tb+zJ7H6g3UdTaGidthMeIVQhlc2/0jxV2gLXSljhSq0h+9f93fxx2FmY13A0MqumqhBxpyjN8
8LLKU1cG/so8k09ajc7646Z+eX9dnYycmzDgcJ8VBF8tG/OGMWGwbUsO5kR0a1fZ/g7yBI/cICRS
GYLmB6P+tSs/O75rz4TMQ8SeGnbCIxBZkTDDcRtpNorq440FTFl6MtmgFPDErSSM34N/o0+NpjoJ
jRbCdBrS9+dzqyXQmUPQG9eWh1A77ttXPUe6XYAcN2uqQM4JxNaid5QV4wMlCuBhCiA4iTiPeihk
L4HzUlFBu5Jm8aDZjGme6X1Kn3c15q2kc94LoFOXcbMgxLH68qLwA1S2oIUX7tI5WAQQbYtUIgeE
lCDN4pv/VayI2NX1HCr9yeiaxPi0hP/p+8a+giPPmNEvAx7n2Vrda91+U+wTlnLScD/qb0Vw2+XA
tU/x8nkT2344JX1SvIJfzSLQqQwYi6x3/2JBjYbSe/xYtmqkEQunXXJWFYa+EEP6eeIS6vslL7NI
rYWn9a7mORLm7DUHi/ehbmgFDCOVuv1uqj/f/9RDsl+uQ+bMI88XrA09xbmNG8oYbdbadfmEjCp9
7qZY6AjiRUhW5Wi7Dq4g6VBk+RjlkBInaAzGuu3FVpqqppC8mFYBgd6h9pVpiVcto7qnoiJyHR/1
WMWW6Dp3iy4Qt1kRk7eYepXMhG6c9JBp7RLqM225UYyDsh+kTX1YdAxTgkGJNagF3lwng78gaqsT
bB2hqUwqhHy2aFaZnao3nPg11KiBR45ep4MflWS3HetDEbErZe4sLOXycYVCxP7EgeoltEUaknQ2
dxhHOxaMMZE+I/z1C7i4l3XG/S6C56pm8okzbF3Rpv7Dr920iyfXfuKH6+zSx4tAe6h63R1h/Ztr
nfT7VUzCgGeCPAtsSehLF8x7NnN1IfqvuB8aaz3EbNhCc0J2Icf7amgY5SwEISBCXWQzQpnApUdy
lF7SrvzGLRtUQEtV/t+6my0UROs5MzTO+xUa0530iTXc/tY7vxT/X8gEaSiUbnSViBtlnE85pNHS
9WLFWmtKS4L2tuiG78II9+BYySpxhzsfadeciG3PXZRARmm7XW8eQCDiV+QOVsoteytuK7jG/QMr
uTB5sleJMJVcmIoK/ZUuLNYTHrtNWooO/Qp8+h/+DpN8qavpCRVZEj9txincqrjlZlUuPHulZd79
C0yAhwmQ7KVVdoQ5dEN2GvDkdkN1+uwtxEAfmHwmH8sI0Sd2OrVL1IdMZ69TH3yQVfnEZJGrF1PA
hxQzVsNPaW8fMwxywn5qdtXKCC2F0rQ4wmDZgby1O3rVkdYuL1JQQltMyg9o/mUfW3GWOyx8yQo2
FXZDppWSmclvfYxyO+TRiPXvMQVJaJGCsBpCqBMM4qLDYtxNfdQyZ5SK8oBw178AmZw8zV0Yp4I0
XuyIfBsdCemvQykLn0N7cZ5uHBSZ/FmRin3npI0AuYKTfoxQEbe4OhE0g4PE82n3K6diwWJIac7s
QAYSWdIkYSXdloMAU997qAUTU7RHBRLIkmLnoZq1hD7pvKGEofeZdicHzOQATeYaUnLAbKKSovNl
le9YGMRARy5S0QwOe9cd45+0AjQsVAWMCBlVQr6dQ5ZN3UGXXv5eUnD5VQQ63Zt36Ct9+BnXNyyG
y29ikE4OCiBpqk60Im1QX04ZIKDz4HQHCioQJoDnAynzERyIfgijY+Rk0o050EqZOV/Q28JnmO5T
92DSS884nD0YH45ZXA407ZG2VSP9X0iJmUWMcgs9ntzfyMH/64xynfufdgcmlvU34fxLtjLSKgh2
cyI2BUgvhk9Q7VjRCV5z/ef+hELERM/JecpYnhEdvVoeRwc0oIvVFWpNUPkjscSyI9Vc3PyJFFJM
EVkj7Tb40qs8KX0ZcgsjaUBbGU94fu+9i5D3ph51EqDjkMUvDkds4a4B2SmQ2qBG/xfYNEb6pKSp
7fSDCiBBbGL/9bwc1t9GGrGcARgOLS+SDz30XRXaHRgsxXX4UtKo2LzhYjnNQCzDVDplznCgkcbk
quiClljypeA2gOqDk56iTmMVPxgauqLw5ZPwOh9OBLmER/Nm1/0/BMGRbsw+QkvQ0npf/SE12RNk
Y4FBi/W0pEwd1L8YDx+UPaULtsNbuKnUE+O/rlUlMYhl1FWVVdewNyd45uQxImTjeMKoaO543deM
18KEEw+hk47xrP59UQV7dfedj6P3vHIsF06GPoOZFydWLJnsQSsE2tU50rDiWBH3HPr/VVRxcNzu
Xxe8ucfXPf0btwl1TTCP1MTKY4QMBnhQox+ELVGzbnoXavUWM/+HG5pbuKGqc0OPj87F0O/KIsnm
cd8Qs6YDXGJNG3KBC7EA2Udmj7urQ+t8Jnm6vOrHRRKB3aogPlWF+vVv5RAoGlU/Qz1AcrcipTpo
zDuMGhIhegp7HZHEtfJCqXlP27aCFKc0jGr3D6s6igP/wy+WszUjOM+QPQWJt7uGjsdsI4MQ/o3p
H9HmgiTXZofmV0Kdy/rYST10SCk4gKASZTbttcCNjUPwtHJmzGQodmi/L2+F+rtk8YnWV8tgXkdH
sXrv+fAW+csNGNACoogD6sC8zRCgQjmo7sS26o8SwgBRpShjTw0waJr2TyC5nex5H3QdQ6OCzQn8
csh+ICcXJpqTe4oqWKos6zqS4d2RrZkZnFUxI5kcYHjWXKtg0DcHG/6jpIknFVyKI0pyP/CVgWFN
9IGWwime+5seg07TjdQETXzMcLvr38NtVMWajRPcTtuJUk3w/faY1jwJL7kGUu33yXtAtHyBYU7O
Dp4g8nZL6kEVbU7QaEd9PvBNg4WMV6Bhi5cQrgpt/ko4/oBLNu7gxw5Gr4xIYTdTVE+q1d73Q3DT
jg+l1mesJZ4+LnOEhXpCQx2CxckTKZa8l+k03PztlsQqYlp3ovbCvdPGKntabCrozV4HU9NQZjLQ
el2f/agqLSRGwhiUkc2ILC5hQYmEjfFCft5KAjflq6Sojtb3b8ZMqBDRCPoFopOCK1Ry0mzd322J
cBwWMx5UHl94tGK4ErbopOwJUX1mkJixNjPi6yYgFjyn9uwW4lQG0+7uiES5qxkHntbJgpjn62Ii
PAYRDQ34jOJo6CtqpPlitefXAEJ1ZdWz+wEve5VBoE3Bzv7G8kTTRYDTbqlvhjNS1pJ1hof//hQB
KpZtHVgIk+xKq4IMsgfru+/FY8+6ZgvXuc8wvQ8cE3BRSWoO/COjMNrAGGBJsHwXup3ApbCwEyd8
B8+f5iV9dywE6AMcWgnzo8onRDVfSkR9nGHAvzPntlkqgXl4aM8p8ymHX8Vd2GIRHTQeoky8a13Y
uyUhyD4lBZcf5ZKtT3iUOkZ+vVndPaOEKaPhZ+VtZW0SuQpAzpgPICbIkC94jh6zuQ8P0LToLyn0
VjON5xRNjnDEuEgvwxJsEpNOB5uBChjYAtEz3OkEQxuqTCLEkXZwhUAfh+k4FjRcrTJYceuvFm23
6l/8919SARAE6Bo2vbgN48xqr+n77aYh6pUPOSiqSjh/uH9BGGDIcTnqnJrpITjkQVIXIopbUOtv
7EJvVCkAFCgTkhaV6KN9k+7uH0at6KwguhzIn6GrSxou661pJESLNu+zrsD2FMVCySjxejyTiSX4
AH7N8J3+hqepNbiza6bNHP3AM9qtLZPXPXLpDyR123tkuOK5slaLCmXY1/5Yq8diBDw+41ZlNl8e
6JiyJCdT2HQ4gGr39TwToTkfQhhkffrYJO4D8pk/EIVx7x3qGFtymUhECVh/mMYQOdZmfbPSKZhQ
/KzNLXpxDCC6X1kHja10NdYUtZIbOOmVbNwj8zvS4sv+3yUBQdLaLGDeN9RcPi0weMZNmO36ieOH
Xak7ecxWrn/j8n9M6+vzRTIN1VaMaxyPoNuNaPnwl2rhD/Sru23nlo5Okwe7WGX0BOa3nCaadBa3
arf7WZBrOLHS7eHt9gvdQRssPzcSuOznHWEt0hCoRsv/WOSzWO4eAzQRjTU35/vDpp8cHEDv+Q4d
74d4lkZpMK2u/YYKEFDtvgoGL3DZc2wlatcpn5AKDs4ITU/49pijHAy6g0G9qIe5VYyJyJDTdAYV
oHnkanJaGphTODEzGRcSVlTouRMSfZL+cGRYAxjdPXRJyKDMYr/4OpokrcFuiSBU67ya4QVnNxmn
O4PtL1PiTHVj7XqOG6pQbKBI4MPXOG9/4so/Z49Ckb0n1jB0s1XYLvy+Y3nQ7JF/yJDMYd4TM/Sp
zVpBrEHYPg80vE4cUzEeFDrKTD9zD79swObtDk+qvgIjhewsYpEyRrLDRbk9/G7vV4NlgSXefU36
BopAGGlLL7n7UxCbzUU7PPQplQ6IaaDKJf8/+DBdiMVyE6FikoV15F85WCUIO253IXcJElAbuSnV
eOHFwFV2kyb1NdQGSBR9aby8NbUWGt8W0kTu/yBjaLRfpbHTV6ORBsR0QmUcRgzfaNABr+Td92wk
TxUkDjj+vhC82eIOvfqSEQrSOZInifk8fnOMZ59QwKcYJOGG4hR1SPTZg3NQlbLaMns7DhOT7tZr
XGjwCc3k6bkqlp376DyP2umL0S4JkDw/CuwUGBwzqDEPcyVw/y5xF3GWTGUEt57otCoAQOi335BG
Ybx37SaT1MCF/xcRZ+zgslQO4/KMdlut7OnUUZuHT1Y2TI3VMFBD7eXYYxEst2ALyZdh+AS0LA5i
xflkWobF7rdwqIWaUnDT0HA8yYHvqnX1uUTG0F5XbfLJIRZnyoKQY/DoZ0M34/3IwdJUoxmFlivN
zCkpbHGdvPFOujAW8ELeQB0GL7tMAHD/8xBpThuTPKzMO9rVQUlcBxnfUYnLhrcKiAXnJGyF6AEb
YcHBRuPm84WaLtmrst+L74UT+EgOPHDYz+zW78nTWOJBLr/QB4kpfsvNgD8oy0xLWWAHAH/NfMXN
eDZN7kS5bvAlJKK8j6dXW3UuARhM7eQrzRlVQ983o3+eUiT+V9MaDYrF7n1fGjL6d+EqrkVZwYdP
1ZTToGIFWNTI3L+kXGXjGqZdZppJRFkHEGVdVDyE9MCwJbIa4m1+Q94++FfX6dw57EOM3M6T9ZKb
OQsiNcUZwxdY3rsSDBmhdpH70aoHZoI1pEONWssRdqkhQZTM54CiiKdCxbzDapikaQqFFmi7K3PM
7VtDz0jabvTEwGlVpHY93MJFI1vpzrYkf3pScuJhhPkercJ+4h7oH4qN/Yk9NoiP4NQSqM4CgHa9
1nCWvh5gcaRONdzip9AK7RStiCxlcdT8it9opIqkyA+8tHJsx6sI1nnEb2CiBrTWBYeljbLJvxNy
XJBoQ82+xzizpqoh5tSkTVCx7dS+PEr98Ugv7XliyRQ61il7uBxnuDQNRTRm7ncUEXWZQernH/KR
K/9SJJIXS0GtCRT/oXsNz/nA+/Qw8ARIF7PBpjqEdXNc49rSZXr3gk8W2Tg2sVzJY+4gHnZsZp57
USME3PwBqQwXwobbACEnHxLRJltCeJu1xRSCQf5W9DkhNLoDg8SczSupfFVtuWzIWmlEqMx4DIyN
WAaszeRlh7DUYLxUlKW2BIG2ycZZerH+7rJyG0YozWrBLp2wW+/rJ1dQtQ1+rpGoC+alfP5NIkoK
V1olUnpHkNZhi2YRR9pObcVSWcaSH0oRmmw6Q3mbKipyznHm9dRZm0RkZ4AUDM9Aj60+WLgooW35
WOEIityZUOsUuB2JP4Jqcs+fLIUzDjOfb56JVU3/60GQkiIZfdZgKs3bV0n+s7OSaojRM9Oyw6fn
yZR0MLYTjE15/ey3cPqtrZ2wF5EvfV0baUiGpZJejWZHZIVr1zcVp85r7nRcveWpuHtXKTZT5q+l
6AyG8oPaJh1IeFTEOBDDWj8IOfzw2EOllIIaRqNCXCCKHOuIS04eFF8E+lYG9SwaO/Po7q+m4bK9
1urc/09HObzYPyHGdRB+ndPbJFHiSrvI9+m64ZJ2bKGB/9hLL6xTscp9t4RfVrQBbhAMNs9Tn6BN
s+ylKN8ypQU3ZahsKbyD7hP0wxTA4AGurzPt5aKCK6UGvqa1g3b7VxBMjh19x+MgEf2bJ4EMqgoa
V9SkNbuvPykife01szfsApVu7y6FFfrx3DVzIZjObfh29u2koQlR9pcj+NjQ6BOEEwWwl0j0D/Ev
5CNGrHLUQ6IUFBWv5zf15JfLxZhco6tXt8nuM83WOm0HY/66t/8q6kewPjTYbNYxhvKQYtvgZe64
87lF3xEiVr6qSROoysTg6UsjpM40pN9Xw/ghyPaGUUhbTRwK62hFyVm2AURHeI52qg9Bylb6LFCk
4Pd8Obi3BICcmQpmNXbBM+jZPBY1/x18KEtk/PE2Fm6lRIP8AXwuGdgavYcy8UlFITNUDVuC7nap
xgQeRpAMtf04SNKMkNi1+qD+iHRzKZTqHlp7yPULcEtKHBfFR3KaLhUmrtshGBce04TSiJwHQ5J9
xc+KTOT4oKT/IsqfQRGJ41FAKSpBLV03vJrSlyRhMvbYCcF/3oU6cyYeLSF4ML5WBp5KfDMsTDqe
hnzqeu+arm/fShf/eUecpFpabt0IlmivrMX6e85b5edr0xl2XzOIX8xERACUve2gDseZ+YANsE9M
fmZ9mz0hcgAPSFWY7sX+y5toq2h7tNQqiP07sgyAxTU2t+vgoHq5YlIXnSrGFRnHJJA0FBWn4Mgx
6BsH648fgaeCxTPzHyoLKFQ0eZPhGHzd7J1Zj0tkZZ91hOTOiJ7O4Nwzwk9fVaDiDPiI6u16qv7A
o33hkMqQjh0Wv7AyB3Mgv5G/KLk6EFO94kcTo/eOsUfA9gW8qDJNIdRhYyNtVeVlv/x8XSlpli/X
YNVtOEFaLl2WOy6XbHFmCBYWvcY5f20VHbWTj9o//f+VbC56XVgBZ3NlW0o4Iisgra6fvmfGDj4j
XX7/tdsXWXuovjoQV0nt3kG2k5feEELK5Bw7zKPxT7tO9eNefzqjY27jGo51Qb/Hm8iCplLe5Sb7
ZtVuMitwfg7V5Ud4HXya0QvhtVpQnytf5MWjLLSfXOdr64FE5QWhpGYScispf7elORAv4oDTs2La
F0UD6HRvA6Ly1mc6ATTYXxWtUxZPJfXQiIFR7mAXHFafDTRnpoE+/6cnfXFJRTjpKkeeYh/AXWSF
qwE31XqnVmDCJWpASBJrDv8AYzP9SyFo31PrwgV8wlq8OPU2nTjKcYzK6lER/zSW6gLzvvgteB5x
RB2iwB2wqKpQH+MrXs5OHIj9fLPDcod/n7t2Fq2GtKXTSjX/tg1vzmRQfKJqyaWlgXm6KKBk7U47
eaFWHGo+YiqHYgyOgbF+FUs6i9yGCTo4nMztT2M+YKE9uSiDM55RbCZrGsbLhPR4RLrc9oTVqd2D
zyJkxoBaA9g0z6ubWCKKzdqPSx9SajS6luOP/kvmxYrkY0q3z/D5IBUGSCWaoBdSKTQCW+9ullTo
i29S8mtqkZECyfrg9Aoyief51gnfPNt+W3bQ27vDbvZ7JDOgxEQXz80xJmBBm2ze38rqTBL5dLar
+v4mpdhNKfs2+hcBzQi/sne4vzQOxUYjpzE4hacD4l4gcnN/C72HU7wduk7haFDA92aWHkLMmrqp
PrRuB/0ZEH3Ec/z5iK/5bia8J76uuNtknRRjRoIg1DstJph174Ws5fC8cSA5fitg6+pBC15ecmYn
eqyj7eK0imSZNtxmBuK3LqwRcUVpQ8bWLfzE/CC+gohRz/f4/c3UxrLU5yju963SxPVigK1jDjRL
K+x+zxTYnF9Wc8EJjpdM8nGSH7UBZiJIWBTCOlfpvqI0UpemqjvoH0jE+2IK6FNRmh7s1Dw2feAK
BNIJUjXza7uI4TSjAfS7vhcfWjTfsyPY3zIluMdd0h2Edku3C8aEd497V995kSX8bWEusrhNnz8J
4YmBfr7VPXpknJC+UnosAZS+XkbN2Iz9ulXTPmaXohPDK/ebPdj0ph+hR9oWtNftmflCMSPaCliv
cdfzDaSATg3wbuwTfvBcC4huEvWWsjgu6lBwQ+1PMl2g4rExjAtkFFnmfwx2FF41z+mUxop/0xoi
2X2n6L74n/yrm8na2wbs0us4tQqGRxaPK49hjTfdyF7TQSM8vNGxLBZxtqMqvQraL0oURa+wOXwG
0rlZ2yf/lK1KCW0SorUwLILaQ1Q4oROdQMRsp7UsySwOitq+CGZXUrs/p9+wP4iZNk0TdU9E9NlJ
474nkk1UnNdXcWyVD/m2vJjW1alY854t6wCF3vjjYk+hXjsk8gLvmVDWx5X2kaHudLhENk9Yr5kz
lEOyXz2HerJnzzIzY0Nkfy66m3C8TOzYu7GHG8oYBccwpe2i+xb8NmExc8PtIcYS+ez6NS+4fNSI
c3n+n5vhgONL9WIUmKu3wrsnyA0GW6j2F09NIpscg7gxeOBTduTbC973FEsP2wBuNnqZdP3DNfdA
ErxpK0uUzfOtAMTQ0MJCMH9kEkuDl9aueoZp0CqER62DW5tVity6U+bF4wswcrC0AorZeFyN1hBi
dTL4oyvJs0V3OxMJgbWdSHPG4Lc1RBUmWlWQxdN54+KLTt06AelTFx1LhUOtLzVAQh/7keG1LSC3
DdHwNrnMyxzf6T5VwTU2dEACdsj4c0x24SJGedNYm6siRqfLJHM6ZHxJxFYHtsT+8sZRK6LdK4cS
XY5Z5Bdte4KMe5V6Y6mnYMrJF6cVkY9zj44Lpm4sJbpocdAQq7W3y/az7NkS24zBxDoVMBQV69Xc
tmkqm0Wuq8eAepG2KdrNz3XRPF/KFgU0P9Mor43K/LVdFONMTLd52HvOdmkyhMcVBDxLaasupifa
UVo5+o3Ksy5JeGrUhCN3tpGt7vcRPiZR5xKb29o9uS4eH3CedJK8+zyAMpDcWcsglNUUJo0qSr4b
zImpcGdwpYXshH7AleI/qlrNsAfy9xoWIeJ869Oy9yualpmp9C4I/Iv+SyYxGpUw2MtXccj82Phi
E1IUVJxihfB7sZUiczJJ4MbWHLmfVUv523cTL8LGI41hl5ioJ1ej/C+Uw0dP+LAiMwx0SDTc5dk0
UmM4rLOgW7Ue41ZzUtpXlLNWobihHwNeZKQAm/uKebFbFg3p6G+uWJJD7+nxX/lRau3srcWlVcy0
UzwYUYwJW7nb8BYNu9A+6ircOaLTePDyLl1F/SF3DZCjm8ZbQRIjuPPzBfY4I1nu8a2aH5aSGZlE
TI8DCJkK9ojFwjuNZmrptopywrd6/kpZuMhtWqyVkC5BD9rGPZ4BlS6gVXKYyAbL9b/Uh9PY6XOi
fFhqAaf2S0C3sK8bgLiDfbqsSWJPGuofjRacBcVsU1a2a9GgItXjPGDlD89O8uA1834MZ6uicorx
o5pG4LuaLvQOBizL9uIDcOaymNBtaTmzFx55Dk/7sAOwow3w3wvI1q567BRcm/gwdJ25rDbHHoQH
zIXs1J1eQ/zsFuPiLaq0T3IgX2+XsgNV/a05vY7pG/xjQdgTybY7JltT5Dsbvwc0TNuFshzn4Nct
+XvwVrVikFjIMni+s9pCMGswcBQxRbFtDCeG2SlVdEOWBwHWTMzGdXrkFVld+eCQSCNA/S+3Bfka
stJOqyJWu+CNxT3VdBfOiq5Pmj+Q5HGgckYDXMcZXtm04Nl42LYHaFVRCQ37YperGNrhTKcpTT1B
k3Wi89kbBWIGvBw2KRSIzM1DQw9sRresyD30vLkb8c8L9XWYJucSNR8QxWYkUDH8bGVltNQhAQvJ
WU2ArRTOVl2Qk4VGBHzFsRvzuXruz3WDqIo5uuEGQYkReOggQPay7Jdrr8Ne+x0JfouBLo2V/A7s
mZgbeJH0SLUx6QjW7EtEtpva7lryGmJIcWj7wphOzeWqZb9THKp5WpeooOPmFIDweT0GQ0mkytU7
9kh95NrhhXvtY5YyuOqap7i+h+YancS0z5nWwguTsfwvkf8Hx6hwqACY0bA4ECCR/oMXAGYkm866
wf3RBjZndaOU4tod68/58bBBgupx209aE/7Nrct+fIPGdT67A7bQ1raDuoGbD/gSMsZ3vuzIHsvi
WF9DK1aFnVGh28nGdYX9pNDT9LDemhDevTLQoIzycLQJ0G/qsaEyF/WfjHYWO1isunUHTGQDaPdy
dj2SaxTMHR82JbxyVzT3ueCnvU5QT+jTtmiMrM/kDm2g7N4t/zdSshxtgkv1sbs2mjleW6qH1Vdr
hdfv/04S6lgVlmJYN04hyHD94oXhlp7SAVQhWfrlVjSPxL1IP7/BD/MDhvvcnz+wqoo9lup/9Hez
RSM2+PdhRyMwwnhm8OGyxy8m1gpnq2eGPyTmAIkH/cy+SJvYLYQ/DiETdsFb4S6p5tL1N3poQPwP
OL8GxJqu0EFA1CH4Lfp3C9m/MAQiLvUv7IzzRiiJXo160OLxEiwKnNSbxV52twhz53ePbm/SQ8mR
NsSyKQVKeB3r+TiAYC14uD4dJgiMn+d/Wl7OIa9c+u5LtxKGhrv+XAU+0QiQzVFMwm/5Wb+suO9D
/2tYZ66xi8yfuPl0g9UsCYUbPltV38T9S1sRZfVa6kWGEkrtT/h/pvj18cZyfq6kxLaJPNHnYFEr
9BT43thprNUPpccd89W3ThhO/25AjbkBP0ZpP21kiX2H3TblaQr+K7kEhnUt5/A8XiNQQwChkaqo
UlrIILJCBQGhBrnIXH12kG+ru2KbrGpIIx9hXwokQFKf3zLDN0g7LSXTWV7AWu0FbcelBgAOlgXz
gXpUsa8iM3RVrQEoPyDjZ/JrXEwKBUIVB+K9IyJNHkNx6QjBXN7bYZ9X8Uq4bMP5i7Sgw5yg2/ix
28BYeHf6zLh7kMzxCWh/CkqVuNB1sHmgutgZHrIRrr2w13br9vrrf7kwtXLloQNkdnabVVRUERGL
dJLcqn2IuparVntculJCIHrFnZY9ELkpGBwfG9NAH385moTwaBrphR9Mfai/b/AnB9xBQMduTKeL
2wdhvLRX8qnhZ8GIZ6nhxzpZjiTJvZACrubfW0KUmI62xFgXmmNLmtjwieNar/KVq5i4k21omeOh
/MdxbkN+AQ80SZCXA6eV4IF2Os+AuQp7Xwhue6p9ZSgf6wPuDPwqkS4wz9e/26CtCbnHmNhKVw8X
7SmKYO7lj9mEfZHe6LQWJi9qNV2YG35I/V3GcUfW03uQWZlKNarf22hzCOLDXd21vJwVyYwkHO+3
6O2SgERRkw7zV9avanmwMTKW8UO+DbbAu0wHYq/+A17+pwGKGVZFHSfMVIPws9kkvRBj1EmD7z+w
v5N5EK0Ab9xNX5kekfPcWWnjixjK658Xb6jv7HM6WCHhdeFWUhmJ/3oxInR5UROQFOEwKiaKcDNs
wsMvBv/He+ThToXp68gSmR38YKnJ3Al27b8H+R3irkgqMN7LRiETkEUnnyO9p6nT2ELokeEi8niR
oa9ueluETQMQYUuaQrONzLcUwgB6kMA41wtowf5MtIzTu8SmSY+nuo3MBkkl0yx7rlA83Yr7Ku6H
5CnfGFlWpOaF2ZFcha4jkNdTzpsvwwV6zgQ5FjJ2pRfR6F0Pm4R1g7q/cQLWz5AW4D/u7GUdK5Qo
pIDrITZWv1YjQX0dy+9iE6ddYdLByFU8Gj+tHVQ5XowrZjbnwNTiCYKXwenMYmJXEtKBMVRvBZ7s
l7CQF6nNd0yqZ1388u7WSc7cLsNkRT6gxVZxsgV0aAH+4RAr1WJUfCNIU0auIqzgOCEN4moniyti
vuagJqfWPLEa+fRxGfc2D394srgi9F77mcw2D4OJVbHvhcbnZq+MQ15RXk45HSANgYH/suiSn4dM
r6piEo2ALBxU2ldC/kghlmCCu5OX519uHuwVOKlY/kPxTUwuv02sbOYfL6X3TPZ7gvOl/VFIv8rw
2kO0LdCfvPBkOZLgYsLt0ns4bRAg+EEhO9j0747hfO5AojfeDdyBVrGNxzqDHLGavRKtyiLoqF/1
5dDqgWBw2ShpOhh4j1gkbj/IvC0WAJNk/U8plbDGOAoX62eokfBkDETX2XzCaHdGrSOOFrmkGlCP
Py5WwiHfYpD4f700ZlLl5A4Evv+E0qvLUdIniteLrJICMaNecFXwmQ/U+qOI7KKSLs5FBotPfD6R
5jfQdtTErwKOgGClCsusq93sHpoIvWt2vzs6+N3eYWID1bbmoVrCnnPOEM400Mp+scOV2ueDQGeA
uRSXvwb/OBLtGJXnf+a9l88xvkT/FUlPbKi2XzEBed2MLqs+Cp+8mycG3e3+5XERBmR1LQ/nzuSG
erG8sKqmswX/4YrGxc0ZRjqR1e6j+6Zi+LZzxJNa0j1Ra38IEGdHztCyH7MuFlh9auG8F/YODCfJ
ZEp8dXyL+sjtdzlPDgDBbPVEY8ezU2SpmshPQfEWmrz7L8KdWS/oTw+EMAt6AFZarFtRhS1DUyRa
JOP7vtEJ1xN3rxVn0BApFPS544qPGHXXQnKCpSxQ+D7ivsRGYmdeIoTRjkBPMgSVc2MUnbkz55Zl
58bUbtOANTRy2Jtrz8M4VE8QGF0/LZrZInYfrjjLGc5Tiuppb5cEbHmcub6oJFkCFu+Xjynv+Q3o
3Jm/jTSpMiw63h1+pK49/Js/gypIaJq4s+bTNLZNe5BoyfDQ8/w33XLujDNbuVExK8LsaybNkEkX
yVLd1NGtnpEwNstDHdXyzAtslALaocnBtvkRtKGBiJTT5eXvfLZwKroTIjQQG8OEfWmloAyXFbRO
RDq8X32ncl0eOCBGr7bRmxEQqpcnn64EirJWUDIQPDe9P9dDQfiH9KQPnZeNchXFSm0MNyfB9Kza
4PF7SZa0A0jjeyjMwUeOTkmUXpPUeQGL661KrV2srQ8Mr68cpHbXZ4zgk3z6REOL1pI5I7Fe7+wH
6h8P6Y3jBBenIkle157u+oVG3N+hDAdV045z4s2UqQwLlePQ/ZEyqTSrmU4mIMVR3sB75Mn7q/D0
dOjE5fYHdmjbV4RedkYd5bOSTNqQrjPTPMX/V8tuZZ5FeIXp44zju5yahCBhVG834lxzx3i4nwbB
mkSP6umqNkScFAGmdYNs0cbBieeDcHFWqZMuq70zUe65/r5Ak0KeT8mVzmXS7tmgF1LlWXVrOxd9
BJUqKasFx4DimqqCOmkDbyQe5cV+3xN6YhzUQWLL3GBD1av7fG4m/kQ6ISo5MtxYwzr9PP1MoNFz
Wk3tgB4Sa5jj1vJjHZsfKMt12kz7cgwp8qL+6mEa1b6/BUTjpLkMh99sKRfsif66m/pBoB8SDvEI
+QKAbOFcgKsoJhLDGcjkpauwcTuundZIPDeJyq/9FH5VwV5mCaEXiEWVnjpuxWnnXj9CYqbvEIgu
4BT5gCxpyozzL4PC12NWundMMavkJkQw1tnwq6IlH5NXQccIDJOc1wbAfDunzJ+ZdWzjYsxfLz+Q
mNjdlN3F439BDpWOCO92FKw3liqP+CBDbJCKvfK/xjg6X+15KYKNc/e3kOsD0OhcEVyVofQx6Y1x
swHRvZ5VPAR3CWVr7p4S1mU7fm2OOC6qxbfkd+ScXgimiOR/uma4dkGqAHiKRGlzUcPfbgHJsj/H
l+EvpYYHSbvZKgZSzDrgJnCMeygqezSAeObb9sKmNe2euharlb/6zpyT/SQtgG4enXz4ZC9wnF8s
SiMSyh7r5twJnZCqiQZDqqlN5Hpos+x0trngH3wkrq2AuzwmKLFIwCEohp9ZQ1ZdXfvfLeP9WbCA
BVNtNA/ev4NeW+8HmsmqOJpTD/M5OSBVJxrruiz3MdkJYZJCWsMpDHG2ddG3tea4L94Oe86Erk8E
1TxXr81Se5QyJM0wQ/TMVxekk6TuslX98o+E9EpJA+GHYaGp5P4ZPh6D3YklGxcq57rTEvizjyzA
/LGYO9QmeHVANbhwbaI5jFK5mMni0wzYbtLxAXARjiTWM8nknuwMf2cXa4G2R2FLBpdSpGLekKzm
EneT41cvzYKtUSNmu9qazjZYQf9btDhYIza5Uup6WkDZ9v29csDjtREILXvKhl/6aIuMCx4AAf+d
+wauT9VoAgmahDcrUDdNyGyQmuBBlW4U8IA6vWvUe74RlaAob3p99CjpMR8WXOXqSLDWLmUolW0k
oLhl5fLuRQEMtYYUllNLzXCjOGJBsZd0QcB6azCJCpvA7MkcZfPTJaJj58j1IylMPRNLQu7SaQbI
q41IzMpyZfdnHEqYP6A5pEk1wrH8jqgAVA1PJOXvOz6yxygtRZkhDqj0vA/eQu0FvWA9pqc0ocQ1
unxdqkyx/FVS0DZmwIGN5bj36mOqipZTjhU5qGydI76yjSjTouiWx6dxsZy3EN4iF7dltgh1vymQ
rMc2iTOO76Elvgf+1mRk8OBxYPxs2VrOJFd1jlKCWuZiKOuk8hwgGa8/5JmSoIrSDoJs5YGGP2xo
J8DNf9Bxq9AwlnHOec48Wj5TOVLGbRb7qW4PUzqxTW7br62lmkBolnjIZ50xRg7E/EHHkoDpoUTM
x8mXXC9YJKnYKOgTmN6SCmUO66ggtZWCnM0Vd2S8uB96jVGRjmvPqKcCu/YHwrPfi79pUuzcIqx2
JH952ZRx0C/J+ucapM7em5KCKmELvBil7JQnep3xVsXa93nlviPzf3H4E9B24g3Mrw8IEthk2kBO
VVab5/UP+4pRrJLitggckNyTMAYP3ntqdL8cXM6cvPjqygRBjjOHBF4l8gQJgh5sbHqIMdYX/bL7
u0Jz8e4S7Gp1dZrv4TiiNBghHvUSDMCYnGIcJdyPUCHUwoa6K7tg2GDiceihr0dUNzwhTE6GMPv4
2R+eL5JhmrBAMAWwfmBIyFGV/14v0TVPH7Pr0wB60qyCmVMfID0BYFHMIVO6NoGSzSztt3Q1z7DM
bS0Nl1R5brlaEgxe0OxhjS7U45flc77EmiOnIeLmqK0UqRwSDx5zlBPK9WTfVgviwDjo5Y3zy8Tz
qFFcYUiPVckHfOC+gFVXEdbFCpcSQSwKoHWzo1EOZguzbEWkhczZ/y4iH6BNGGZGrh7ugyV0ZV8S
SDfc87LuM+9vDqRuy7LOdViwhZkrLoQYBsXDCZeCZPJLJIgC2Z0MnmRjDJCF6FGNhBgIT6c79wMv
b88Wd7gaBhvG56xQfEH83zHgywRKcNvBEUxqpYK8Q711z2x3IZbilZQUEZN5APb/3iB93Db1Dugx
zYgrGUr339zwiLrwq3cxcQ7nLkZomxZEF9CFNQR7H2eLPy29L9DCKhGR9YKLvPlAalKxwZLO3F+2
AOzLQ2fyUcp6LDuidBPCrDVTytb3ukux32KCSLoeiDRBURMH3V7mPUlFc8AQ9zr/e9eA7OrZVGPZ
iYUfJ1wMOkK1dZnWmh/SoT7KRgmRfnh2yFTpCocK/BH9qfePALpHtQui1tuvfaKxGwc+3hfQSZqK
aPjRWbLmSmRx/dWJKAitv0yw3VRO9T2vAzd7Ma4DUcvTpvqeYDbJtwTjqQBfWhIE1TNPlcOpcNh1
1y8FpVZ2f9t5enRhe5ZWI61euyLnBJmhDLuPxQjp1PXnfb6DqwESik0Vxfq6euSSppQd2VTQ9rkw
iOSrWJahYltw0PTOROCXC1EXJt075q8nZfB6wgmltidMWAmqVyoz3wVBLwSud/89Jdn2CMX0ZhAq
QMJAE6F54CzgMMXt5X/gKu2CHUtv/Sehu0FcR9nTBIxvwY52o8MUAOOWrLN+KMecjiWBvhUrIdmW
R3SxsjuLzI2xhMe6eWnl2VtPEyYiLoRBMgA2dPhAybYpcT23beUBD3HB+dcxtPZHksO4aQ4FPl6i
IH+ja15QOuR+gyBk2safo9M3XLLy+kFGzQzT1LtGaZG07GqN95fHWnAA1pSjxtj5ba86PXE+9pWI
BfXfEbhahgMozuXSDgXcAckSAFupaCYmr2yjIio6PUmJaY/f18utGNgu7HCWq1SHY9JQJl2MI5dy
TyrKqCUCEElIZb1iTKNF8Cofl6h0fbiWd9cwheu2iLgZvUXEjGVM1MmQllX1LOyZefzd4N89t7lq
stbM6ECXD9zyXqPp/qlFajvZQu9t5V/1oUv9zl4axYrlC71aqrMDOOb9NaqSFft+YuLCHNyp/+D+
VyIzdC4JfihM1ND05Ag5m7wHczyMO1RhZfmdn9+ufgdWm4blTPo/drt6rytT4SgorH5yeFl/LFZN
65JsTPbg9pr9iWaOLk6cYhZA+5naHJ5d17MGsQvJ9CYGMq9zM1vBjh1ugjOp/CgOoYQJl/XbYQks
RPrfJoskQf6MhosNXzuKN/GyGgk5KnDlnBsKE3IJ066ZDMQlmuf4ZfIP6DfSbvpz1646OoUCnAO2
zyfcmUidYTljhgUfKooFbKuM8zhpuelHyvMldoe0UPWESMSnToaj9T2/Ha5tkyQicPsR783bTmTP
SK2C/qV76PkFQomSlDW/WoCuOjAeUs8Oi+2nEPokHQYwGD2xvw7sJt6sNuLM8VDfelHYGCjaIolX
BGjr/ice7P2ycSeSDG2tkWjUmwn/0lyGHfAcE05a1nYfjFMa4hPBai/HKsJHjq3croOjWdG3Wcr5
8Q1nNp2MC4gLqbOGlDi9rGl3dUTSCazrzJUyZp+b/EEz1kAEadmcMr6OuGZTjfI7MIgCv55zwC+U
lFkAajTLPV5p/20nWjxmk74M9eMdyOUHkB44Xjh3mre5dS0QK+mG1gWF2ADv0IRuEiVcWCItepTt
saeUKs6UeK8JZpSh8HEuJ2Ppl3A/XURssXLJdkhQ5JbwLkj7HgbnP6yIQvlS3Qgc6LnFS/uDlxyp
VG7h43daLOuG9oezU4kIYLz61Slb92COwF1/eHpLuReXPC1c01ndFCNUmL3aJx8IQlkm06bLRiDd
jvJ1j1vI//R7r47DhJEtsYrRK26Zl8uPFn9vfLMpcDYxFtAR3dwJdg964KenMpaIFJWDnL1tH4Iz
fuwN50NVoL49XEhhaaXfgTfbBZs7uvsLwZ1Pc0gCD04h9uESJ0GMMX7kxPbf8TZlCiEWYkFPK1q3
VfOv5lEWgf5fvMCogVyTXK1FoZz9oQbtvp4ZYE464nnpiSoTH4sKTswz0e8vDG236N0dcj49RBCk
Hag04qTrMvW23JfhODGt5Y0rZAbY7It7Fdq35wP+ooRR6+YfNBP2aReiv28Dt+AfL5d0Y6uFNyYW
7BsE8AuyZjxXwfe7dgI+OYQshscKnX+ZprkzPAx7bj9bTokDapwyceJvyVRbrqK5xEutVVm+xDiQ
HrWp+8XZlIQfg7Kizmek0/wHogEuLvotUpiMqeRwsacL/JqI34fKSDWBTrQZMqVv5xPJzpArkM+F
HhKxP7S+QR0UGuHZTbN2VFwOP/QZyf7dHuk3SVBSMqkFP900ohkAsRa5D26hA/8aonI+1YD/JPNO
SsdOuTxs96W6b7mn5hpwjSmggWLlDwWekg4ESfQJixj2uic7eJSmK+5clBJsHlH3QNrpSl1Ad1vy
sm4wMAAwSR2TQmshwBCr9J+O69ohKdwA+LO/6itF1ftodEa3jHB/CP3zEa6DuGrMQKdfxVYfMWf+
w+5ikvYkabS3zX3NLtOxqI+esc0K4WCTiyHmN0267U0Qrmfsf7RlwoT3H94L3jmwyVsYO0iqgTQn
NJVosR7aTali/4TyK9ISbyPP+JAB7xBKe9unpxFZdiSqt/uhAMlfmiZ2m/VOsBwyFzZSWIU+1GaW
8DoNjTPBzyb4UMtV5p9bXy7d36S/xLY91DCm+L20/IQUFbr0WofWz0k92D3oSdoXmf7YskE5YJEW
+nJKC7238baKsSa6YLV4jzhLSvgqTGZbpqTs7qAm4Hr7KZSwSL91/Sk6+uHo/fzhYHcC/labCN0E
onrrOijLjXl+G3aMsSorVE7yscsMBR5CVumNBatWDxXJX2PsTsPVnQmAzPwNxkvKdeapMD9SnQED
uUsP7wyUUZfUgHIqDDQBCzG6l4BsGBsqU1Mc2k763bMDV5oZZm5Zh6Z0QKWMQeFsGFsacRJbXweC
61cQ9MpbZado+3hGDfe0G05Ri/IUo9UdAKxKpeYp0Doqt6C63WQbJy/iLMH9/T3Gn21/d/M2wain
PZUgf16oGbp/FHdczVISocHoW+IJ5Ccz7qbU5TrkXD7YwG9Y32KRwxNVF122I3FnNsu7wrQNYvoO
zWAW8mzNKQhfX2OfpBjJaxOzYyYtZ3UAIQUtN7H1GUxs8q7LZATAWETgIrDg0mI04Sfm+w46g3R+
egp+6Sj7WtMiNnvB1uSZyfJGYNXtGnQUpnuF0K8evNe6QfOfy8OSH1fhEx+Nmu+cGcOG0xJSwgnd
S9gH8qV+zV6FbGdlJK3I3zTAm9YjPE8MI0tCUSa0mphgOiwh6F6noICO5eX2Cihoa+8+3RjIr1pB
f2bFYZJFHZv4QjXZtUQgD4vPYmR7SAD7s3Tz7CL1YPh9oe7p9xv/1WFx/dLxVQrq3u84vHQpPULU
CnngLmA1Vi3Z4dGM7TuTOHnAlP0PVesILtm11bcjCgr2cEeV6igYADY0p2ZkzzeefzlOfto3zp5L
vhAySSktwepfBkozywODfY9lIxX8bzyHmSDRWNkbVjijx4mHGNROwbZCHkO5zSHU4NWOEAIGykWS
AeQZJ5VXh12gVrKURnVghHVLIqxgRdIaJzu96MuIOynvNaurN1D+OmDeA/C/+/dizsG+Pmk6DJA3
sJAHLxP/FzQ01QO55a9nwFAh1Zeghsriaq57vhvbgSPtcQGH+G7vkbopPNICw0CW0awl0sjRNrty
tgb8wH7bq2e5DOUAc3IQB5cb5mBBO6kQxtW1WT1SR5jKim2OeA5HSa4GGjc6xbnsodbXr4ZA9dZr
6w0P3RXm+21mpuakirCHnKnAvxya4Ub6Y1n8X5Nt6kFbjy4xC98cH1QopYKRrN6J/at9x1Ii4DEP
mCQB/UxohRLvgm/+msfIznGmhbxgeP5FOp0afMYSH3NOWaFRoxngKcDy+jJ5Aw+fYcX7lshGBRAQ
1LW/iJojtQ748K3wedHeMOb3w9CLXE8gvWATBOHvVuxV1OsAYtC16P4FOdACWUoevKd/8DP272uD
pF/vhBQMGRZckJnW9tLBTjAYdVw2sY9ocPGGCgdymTFvIWb5bSVnFSt/rgr/My8hadHH7kVeLTZ9
p9T9BJresT28SlgaojbkTm8Mb3GkHFsgmMvgliGufzpOQAmNl2Nw1R0upYftsy44HOHh+WEjMgZQ
fVoqj/Pe+z/zlMWoevIrDRojygRjkdF2sFYHCcENeEh2SBlX+35/sw3DHcPcWpcYhmqgfFNjJAPQ
acSzhXlR7WOnQ4fhgI9dLRLLoxiXf1jRTK1gxVpHJqeCRETDtNQ19AnQjRI2LZcB7lRsin4n2avA
Xg+sSY+RqPbF3XTCh3hRtGZNj9hJZO3+WVkuzgRAsNh7qpKYR6KoN3kQ7+DqcmFg+seXjST8Cj1P
1nlkewYPVHH22Sjd8p7efrxD2a4ieADKFG6ksxCk/312Bg8j1x+QfcUcorQwDBPSR0RU6fKL1ACa
zyk6pHokhd9d66p2yfkgqAAtKitHDV4pYTBo+VJ27k+P50v/LQw10jDUyPiA/b7NX94y330i/AP3
k4S1KkJi5PSwd2ViY5utVpftCYMnML0Qp9umJ8oruuHce7mP6Gs8yu22fOa+cN4pjbPn5yx93bKE
fc3UsUi7cGzmZ9302GTPtJXFTtM8fM0PvJWxwpWt6y6tNrX4ViNQtWnceNBCsH6LDB7vIxz4Ph1E
XAAZmd96QfdtLw8Y6LvkE0aSObEhQwN/aUeki/ZVGTzw3TfORl3xGHAunVMVjuUw5HvJAOM1eIpE
0ObiuPp+nX744uhRQb9mrUb/E09uuLCU2/hyeeOCx9o9/mwfJXZrZU1M6Krh4SxX9MuufUdVufX/
phDQiFEd6ndBQubuaWrnNvydA/uLSfrnwL2xmJxSz1bEZz/20o511Nxez2KjOD9a9klmDKDZ4YK1
nZShNqJDY99hnQrilsJmtDkonsNR+Y53J4mKRhzOmDdAK/1gzuarJk+mktMAzmAoPXqns0gFRkVd
pREVIfcsTyOP8L84+uC6/jc07imUbRhHvrMhBBILz8h/ncdQnvhd1GBDicpLk60YNne/t6UTsMJC
PRDt6lYqtLgG9poqnWAdSCeF1Keuu6+fAzKSOroh1iuBaYGbkRmTMdisFmNCK6XhLX6WH9VtBWIh
h9ck8EqDJWI58n0jWsFVo3oys4P3JCPa60RJ3WVUh8pfCPryOzBTiqgZQkMRVmWDBqsT5IUIEg+A
kvLkPTZgMKMhh0o7+I03EfzbQJMKoLYruAmEuvAhPA0dOAOp8+A6u27IwHNKuTMP9LPcLNCSTi/L
80fC8bHgtt2FUabqddr3dm/UC0iO0ZcvdgS/n9F/lVyhhgB/IgEMif/fa88wNztM6hvBUCjicFSn
9wzYUHiY86GSdOds4EQiPZ8zL5Ln2bD+zBTMVdezEJetIm5hu/lnvfXYK/71ugf7v+ijaLAqbImx
epV6kWgsJjMvT4KnaiZavo76klMs0WEACnYtmwcp0WeGflPjlr2ghkPCshrYDKsAP6Bl5dsP6afQ
DYDEb/UkHv8rBYVDdGDyJq/zkMhEoSPZee9iepcu71Q3U05GN36GX8qbxixrBeS4ZqiaSX2ZiMix
JBKCX+tV1Pj/qI8PJEXCtq/tJ2woK+z9mOBgNk8dTxo+WLyPh7V10A86gKV4FN2zM2jKzvXz8vuQ
5Cz2vL9jiJP7ekf5TAjBzP3VznpAcHsQBK+XywfWlL/niaLyY/un4M44zEffy/afmzyphdpgzCA+
oR2qC1IYXNlNjFiO+iWhvKZJq98pGau0fQe6XfSaP8lomnrAu2TrtjRfyu4YZLlmcwen8aV62Aqt
++DKwU2Xyfn+Bk7QnjBnV+XrVjx6Lg6tkPrm6pzyQRXaff/S0e5skcSJVcEeyLGaFEPyOS7btwBi
jNe8iOfKBLR/XvzJvVJD9j2Xjz7rhSQcERAcoAXFlLQhQNj/N+Vle6em74gyfogCcjmRLakDDv2x
GSP4WhNXN521gfdthsrrtakij842rES/+L3BqxzYYRxTwBvRHc+P4jRhqioTi66GJYU/MG914yDR
p+/ReggLX24mnBAyt+kRcklfrpcfkY54ak73jLXizGsI/RJfAFOmuAiXz9Xo0gAAzfeHS1ldQy5G
rAqIfF07U3WapxGQqoyxtfcdihq8OpwnaX3n/QUjHpNrdFW0lv//V0BoAOBDmiwGPTXUyljF7yui
r33rx2xQZguoiLWUpPDfxDhhKAicivK+fDCG80Qgcvq9/Kp/DncX+zcY0sFe+2mAa8dTMC/2NOz5
+rghN3Z0nrtdXnGUMNIpeMq3hMXYhN9+hx04SGsjUVeOyTNfPaYIZjMkFWRt/I3Pwa3bG4nIZCq6
4RWbB9wIyDDpWwcnOxuvfDyjihD8ugPvVBM8Xv7ewmoa37qI40W23ndsxVLYSvB5hM4n6SArzipH
1OhUNTuKMJ2VL/iuVHEJ0gDKoTili4CbgFNo8ZAarxp1CqaZ65OJAFE4IMk6T4axWrkx1yp9lnv2
4gwh+LDe0jaqfVBxy6yImIdHkvtLjeeBCJuVQAV5HfFAqz+KuM5DAzp+8rWvOo/1abYubcVQ9Rfn
BkjA1n/tfYf9k5gWDuSZ8qbaajx91w2suLdmxXlfHfl3ARiLNWgAtsIVI0gAJ+lDEale8EFMUGH9
6DOvwdQLdQwjubp20p40FIcq5tI1oP1FcKtdbnSRDnTQI3mqE370cBmXMRKEADXyTcn5l/m3AIyT
anAm/MOjWuhX2GOrFeshkGar/In4kg3TIhNod5BJ8NHs1eAVnyfE+wboGc5oGKfq75mCu/+W8Q8J
gigX0bDFIA8gK21hssryz81Z1Ncj8cAIgRJOmQyi4ST9gYsgstVYFtI4a8V4tbs7jx+5GeyDKD2o
N46DVbE3MbZMX/BzoPy9w5KxgpIk5bSKFLdH+zsvVySImfNcBOyImAMgnVGuH8psQrDegBqqL1iR
/v7d9G0Khce3iGrx6wQ3D91j9qV7qzqDNHkLk+EGp+46L4rAFv3iguYpLa8Fyaz+nYEvp91H7ER0
lTdMoKIjq+zhoI/Ohl7c3P235b8RozSlEoEt2u0Va8h6is+4CUDXgvT+EN+dOOviTBUTlTZxkBez
B44G8tM8ydutVu6lDI00Lz1rHGQxx0pTjrz+y6Ta4LPx8sTZbpr4HbhaEjTNdexkiIiCUrCPHCX/
/2lMu6gYiSgiRnnUV1f9KhZAQ2zsGLjpVgzAK9kL2f8kBxLvgf98yg/6D6SUWyfJ003eHgX54a03
40XFncdmCcxEFkpTQJqH7xtcYGrUAG5ZVx7snJNm4TXNF2GhKlhI+k16k4ktALkrQ2bg4vrpFj8T
yWG+f+wbkbZOXQ8hGPht1api/UhIFK27rZv6Hr/yKqVFJKHNiaiJZOgjhKHSE67Tbs/m3OtSmHh2
KUC8l6k3QGVqU0hdMeFyWaRDAhAICdfk0M0iCjn3D4JX8BPiXeJ3ZHcp1Uuork4dRgtNlf30dqd8
/OhulR/geoZhipZxQU8TV4qa0AU3+0F8FG7Y8RQSJCdtW9VeaD6vYiwYr3NQTw4bgdoKHhU2zWDV
MTnMowwilswobQCymttkJswu9VxAE1Y+Ix9XXXH/ZfxecBqZdmwcQpLp39cQrYeLo+ra212u1w18
YrKmDJm/FNq4QQSIuTSjSr//tfh67FDYBnuHKIKeLaPIvqtAmRTwNXq4tBJkTk/k8GELnpeZ02HE
oxNTkl30LFpFlg2voPUGA1bKN8TqlUHvbOhBUkeMNBAhucY0oFDpYEcICXL642eTH3+dzGZpbukk
aw2GcI296W2URSxZSQUHhGeYCmzNjKVcuVPwN5IuwJjJFJYfijHqPqQois8TIi3CmzDbpyysBoiM
cVw1Yyj+rlFhLwch2BvbHrfhgSuG8xL/kEmygxTjR69DIzdHb1gyUK37r1jXjO694znooRZQwmik
XOhlqVvjnLMSzHA6UHIM30KdpHs2xf/HVWxQ+cP/nmetU68fjK/Dwn8M4ZaDHczw2a3JlREj/Teq
nKAaEA251hztcRWY8X6YZurbnaYCqo6nnVc6nBHa9zVyvrGxBwJZE8rmTa0AIw1ZEJ6Lu/kgj7eF
/a0SHfWlBzzJ/Mu9h9KXj0FoOGt6k3ZcSeoCSRxceK8WfbB6OmWnptaBDlwNbdSNueh2veAU5Jbn
h0sUeLXSrFmXdg59VKuRg1Zj+7d8l74+3INqbDaPA4ZPUqm5czQ8PoUBXgiy6IyVdQSr67qLT1u1
ZM0PE3Y6eEXtJTu9c498pMXZQO//flZPb3YoWfG+nio2WauxN1Mrj4mr0YgK5BHfV5noZmpt/sDO
8WhHjsmf8d6pUMQ2GxhxnOA/wjUmNLiB2gDEHw9LY8ZYXGPz+18bk3Dn4HaPh2VVSERiCZaIJhW/
cwVFQfeIjqUBIvWZr06jO83L4wiNFF6XGu2k4EbKqbJZ7TIu4PDTT12y4I6QDkuyiPtcnMpW8INR
OGVtU9XZ2HgKVlEjqFhJbJ+OyXtknJbxX4SgHLj2TiyPpd36Wy8UgLHd9ogOA7EDvyrvoOQG29K1
NaSWyCA+9uUf9Hj/AZcrznb7PZl0+SeadQYoNq1XDjDJg1vKlntIyW/Zdi7MHKqyKiLUmnVuPUC1
hAONBW2ham5BeDtJj32jn/KlTPm7ih8RfD24m2YK6MXIO9EnJNroNLn/7kxMwjmaXlgAkleeTtbc
86KXQCXCMJevbB3WrrZ8hAXSkXIb51JY8JdmXiBCp6G9z/PENb96XKK9R+h1eT7xo/qd+gZJClWX
FHpBxc/sm42e4NqDAoz5lGNfilQBgg0D+vVDM27l0iUIxjlG+uY8kJXg2EGhc+7ObvVdNp9dupgZ
R6YgXXQm8UhtaKxSV6C5NrOmkA0oCba63VPTFvZ0G2UPXMBhWdk7O8pLF8l8nhDLi923CHD+n6Jk
mo0EguG/zdxqe6IZugozYyPulsvR5ifxVjtHz92T3Sy45euWGtZvJzvpRFrH8jCymwFClsq08JzG
pFeKY12eYmViqkY2Qju583Vg39vtq/RSj9/ZwohmWRhMXeQU3RgVg5ijH4bABrzZFlYAxtjPUbRp
iu7Ywo7IkFg/V7zMMXZ/TjgpM+FmBt+n+R74C9j43eGVn4VOh5/uZWIvsyR/7ZS5GAIXzTnDwQZc
m7uWYjYy1dULcv5a0AQbZch5Qwfj3RNC2Texloeba0XOBx7Hjs8keaEMT/FXxwYOtDe4HvkHH1r8
13384iyCEIRiAeLxRojTzgegan1yDfOEPEYFgiPnaStvtOSBA87bvlvdynYNa0CxCUJU04v0usPL
Z1WmFY2oN74v9zaMLDZBVzmvthXy7CR+nVyVk7UyRXo/2ADAiJngH9zMb2Si6D3RQvBSopZx4wHo
X3nFLGwlmcVQTc93zn7XBAK05kWCVQhHjJR4v2zfCxLoD777zNnIgwNLBbU7IwxC1jbijyePrzSr
IkYue/sJ4SzaZxpNd/Ndcqr9ow7d7pW8DsVfp057PtFyg5MyYIX1t6iEOa9qEuJ+HBZZ/9zfNVgM
UIkgFLWn8GeZlpbx/HajVwWP0UUQFR9PSF3xgOlzd53DwJ4K2OqOKOSii9h4HLJF+/lQbP/D3hJb
8eo4krFZUGhgMzQzUR+3LbKnDIZ1tsONf0MP/UfE8L8ovip+15X3YFvBorkpxHLOF+wF5p/rI4Fw
V6c5EToBx/mVmYw7sGJIhWQ02GxO3v1pQ9y7kNpx/G6dw1SAL4Vte20JDLqw3AYchc5Eg0ZUEEy6
Cz70bjDb+nC5ULGHgPXMOeiORyRXcTcf5llF35P/KDcB1PoGp0Owzwid6coaV/tOX03L9Zmyolfn
UPbuqB3PFgx2O4gSC0GPdafWyx+dXg0KG3f4+m1fcXhXfy/lnP1d2sKmPD7FgJ3g+QVcswTB/g7J
+Rb97VOZvOj6lshV4POdsdMpktT+d1ndrDGp5BrEnhmFVQtLSFodWsgw1K9B6/mbwm4cagYh170e
sscJ26jrtdqlrVWhQU38LpdC7OlCiCB4mpMdskTIwh3HsxLar5dbPJ/TlTq3y+NJBE7/yH96N2EX
wEXM6NOMxlP6dqtMPLyHxCIBLxXxvGpxo/a7HG3PBXKk13dPjYOIIycSeVmkP8TYHb8ncHfHJjTz
hmGIgqVHCO8djf0KY6Imsas6d2VO+7FAF7rR5LC2Oo0MzRWzdAc35pSIibLCwgc3oHuhl3wJXvD2
MOz2dxvK0+QiNi+qh0RUt9g0XD3ceXcKeYOP6mhH98wL2MxkAT+KhIho7UmfhrHO9qAcPsetuuxr
idpZmfHsDaNJS2VYQv2+miR6XBGKk2XIAhRx9aEdEvwf9jJ58I9bLTYP7PPwgqvd0dE3qoWPtdgs
lK62z2Dk7i8demdfZHY5HvIANZBZ7D5m40LN6I/+e486Wt8MfyNQhSUF1FESNraVwUN6rpdjUv7c
hnom3cGnrP2MvBi1NyH1Z0lAwQ5PkB7BwSml0zH+l8L6hOVGnCeRxZsGy5BltceJpgeHe0gdFTIr
9JLYouzc4JEBWi4JKSqMqzyMvsn4b1Vxn0SFGvtTUctLTH0WA6wLXX3P5TgNW909II/i0zXrmKux
62WKnW0yhbMDDvRDTN2AVQQIYnm8qa2WL5371z/FmfQQVqwtYLebLPmGZMKQxaM//cuyQmyb32NP
jpJ9zBXRZne8sUR0kGyCnA2mKvcKuNSHrIQYvk/Bvx/2u5LOU2afr1qXHPGLKs4AOUGz9QFph5Hb
VnjEc39UNyPVU4yZFlDQZKzU25/n8ZLRDsTnOLzdYcavXUAQZEKsyfLceVE7PQOs1yt8W+ERfbQ7
QiDaMI3TqN9oFYeE4jyHSrl3dWCNs3tm3hLK1NZJaz3Ho2OeOrJUMRCkFmFj2oVX4ydIIGXjIkFa
XEq8BqD5kGGVBFGV57O4KwtTruQfKAAkrUetZYveaz5HVTT6y+zs+VG5pDvKmr4m0O7P4WNOHR6r
boiYzI+yFQChssXClBYg0Te7jlBZH4/RLNVP7wOr+CvdZcG20WP23Y3DMCMhDDuKCXs4uR3jxHG1
jL3hWWgFzaSonLuuWNep1sDqsH6Jxjy613bK3reAWrc7YQYxil6F8skSlTQ1V1/M6+TcYX0kF6ta
XsW5Y5+sh9LaZOQvmt8vc3OyAYEby/7M98vNlmBuqdzpLyeFhBymPnbJqDcgWkHuwuUoKxvE5l5B
9G7RGijrLH2J26zCBZ8lYifN01llsyIudOwLIQhHw+GKDtN5yYUvkt/JF8a3Q/CpJRdUTDIOeoUz
E4M2QndViv/6+2NoVhhHpHjpV6BHE9hm+vRA10DUjEJd0gemnQU9uDLszt5jEfZqKzk1husvc7Q2
xzJ3NF+e4ZOxkXej2u6ISjfUpNCc1bCNcLYLNtUzd+GJU0kTylV+6VSxNXnZL5twPky9RDEEtkRs
g6gzBfGSiZu72e4p0rzT0ZbUuMi4zjpZkQNAtv+673UxG/agmdADPG+5AGCEmPanHauaLJpDsHc4
IiV3Xhb4DY+ohlklxAwKUC0G/1FUKq3ZqdQZ5r7tkvjQfgbbzddPsV2VhHcn5CnDXNNQC3xR/xHE
OdGNeDr5UyyiZ2DnJOe5dkWuKv23b8dh/jU0G4Teu8DCJr/28xNJ1Zu3vglQr7264OMtOlRIs+9o
KNxtfyelWPv+uG1roZQm2j0+ePDvIapN9gIiMCuUSIfcddcXku26AgYRx5tsO/a7ToEAtaVfnN4E
ObIllR5vHc8VqU+X5WpOGBEFkWPeR471QOzVooso3B/xrYj+nnymu/+I57TIpoPNzLCcoep5n30v
8DDZygFm9JzXgInI/QTI4YBNUPAec4mOHm7x976hgMwtxIjaTnV2mfQQowCxNDadzzkKmKEFrNY8
rtr4V7ilTIrOtBbmKqrDmOY7HwgzLfVrPxpOXPh/yAtGEbu8MoCUIOVjG8fpdKajM92Mu+EPIME7
Hh61adqT+F6VgHEeLD8uEH1sLAyEAs3jznQWDATCqpqkKglevP34bpwo24MBAvtMWfAS5og+trKe
r9DvDK4KpOMcl/n+1Rkp0qApQX2KEFKh8BlWN3LFtnXa7p+ayTOXtLI1jKegX2ZUM2oKUfHVAE0K
dIDbNVNAkyDNepl1X3QAlhet9OU3T8on8z0xZ7oWpZW3jMCaxujn8vN0faLI2vXFLiSYN0/n7tuH
ZElLrQQNJ5obRaEzEy1Wmn+LRpM0AJj6YsD96q6eJuXfEVjr3KpsBXJXaUrp8yEw9p8Rip+OBkRP
vRaEzHHQ70eZiyx6NjGk/3c/W6FWJOIsOkyy3uFyD1Q5Z0z8H7pNfqsFcnKZXmM5Lm+5OwYXYpzn
g8xkqMOiWYgmW7r3f9Kxy5eps/B1X+q0uBk4aDxiIXjSOVnjMPvxRwNBTAVblNIMEIhL98Nn/ISF
fdu/qqMZhdaRYpD72X7sAA/ZI89hPt0SNq9/qXvHDN8KJmDMC0EQeRABU+WMjtn7YE5GKggRUbX7
YbpiVegTWnC5F08brcw+vpKIQegrhGHZHTagfO3TP/rArqAWyVVCc5i2jPQJe7oLmR+rbrRn+a1O
M911qnLXcxRO6Q/SneI3stKkLg9oC8g5aTfPIUIHZClheIzLiO2SIm3i3uZrtIBJL8ipvOR49teJ
+thCY6IWjEyiejP5zcvSpB7anoKXRmEFTchmjZ8eG2hWDiy8XJ5N5HyiMrVLrQhAaKzH74vUlDJy
wF87v0TyqDrIqF0zYg4GPA3mQcwHMoCbWOcv6UEm3zqmGpH77BKpKMN5u767EHjGGbzDaXEKztAG
MzcLnrp31BdT/GZ7UddMOUEyDHCHklfnUDq59MgAkHEUQ8wHjBMpLIgKiC/d0g/QG3rTQfEkiDSl
s4BZYcUluIRJhEGNM9Jn0vk7FGS5HLjAl/3ZFH6d2n4fCMabxOz0Sq1c7QOSDfCljQyTtztdV0Ef
eVp+QOeMA5hH5nCGX5qlFbrG/2R/h4705P9sLNPHS95kRG0hTDf03FxZY8V5FqBgomvpj5TUcPx/
b+e/96cXZ8IBP8+j+Y+V0mgsTpy5DqlPwQWiGM9zCXGPGQqCR77kDK9WQyh6lMGwjCNKvZMicH/3
Tce8jiFtSJey77ve+9BU3SevXOnNNsA9U97qYfygUnT/j3LVL37zzxOnpuT1MB4Kda85NU24SL24
ZSOE71P7BiPUDYYzHgvvZx3g5LMg3hpskTVhN2i9wGfNPRGvBVO1GcOI1Phkb6yIVZTvstWSgKYm
VzHnPj+9ZbhRrghdPkvGXVsUPBBPS3sMuac2Chww4N7IUPch5BsUPFTbo3oZk0ydCEnFFc+jYMUi
LWxpHxaGJ+tjo6MW/WS4+j35pUo2ezwnc9S0VOYbGSjKiis/NdHyi5d4Q0ccY6EBIgHE3KZNUkTP
Qcrq9+TvFRrni8fNCxq24myzLB0XOGAq6RUhgqIbPm7VyQ8ucDRHOBQ0WPwucoM9u05xWl4DiD59
+a5vI8e63IZoUJTGaKRq2SVB7s65yRJn/JnkO7PeiwEaMxe1SabaMoxlnEME1wn9Dpk4/zmtab3k
fS25tmHt69zsHOpyYCHafaLT9YEYl9ait0rA6erX+SNPskfiJtCGhpXldDHruiDM4Pncq7d45o4Y
BFtyVu864mQIR0Trn2sLU5LR7RmAbUBKPu8/d7quCrC5rzAPTT5PlVZp33bwTLhutfFtfKa//QOy
3MAvpApvQ9sLsrzXNdBX4rf01OHyXb3RU7pv0kxu+5umSaI4t6sKgp2HxQxSiJVjymWrkOL5HJ0l
OHlSJOizqKL6W2aFoJHSgovIVKxgE+hb/9hiINxqeswZKaOWx0e3WcbqNjxQpD+BaoxKnZ3ckyrX
hNGIr/2JMc9pUuZISbuFf+QHJGoN5/DU+/8b3BkKFGd+j4A7LWfBMOThPL43t+0ePl7+4hDoaCnK
7SZfemlwJib0sz6vpHGqPwQBRoFBYF9g9o6yJOwoNLuV+YDEiUb3KWWUlTtEAqVwhcRPN/QLF+0w
53hQmMAQ9GzNTY4nDPBcGzhhtmQ+jCxwZ6sYQDYDIjIY/EFVd27Bg/IE6bUdvPzE9OeDJ0cI0VlB
xV4PGzGC7eR2eQ+2M7Srdk3Fs6ybT7uTfdE27JtSsC0tiK5R6Z54tF1kHfvzq+OoUef9PmfEt0Ck
cAvE8StzytBu/U2RODQJgOr8YIKU/ipSjXavxDdnjWDzImXOVXMef/R1D7wghknSe9wiRJ/SNH4r
oFj3jYQlC6nlnpZadFHZPWtvTAA5AJjQiira5NTNGUZLUBVNSaK/i3AuzR9pTHFC0cbWEGlGMSXw
zzNGJZ9HP5zURq3qdM6bHtr/cJzm2H3yIQQcCR9MShlnZ/B8krSHC4uWrjwkt/CdIF2iy9f2JdVO
UkH1Uc0Lmo4eIUZIrDyt22g8SBPP/PfKxZhcpzumiHZCJM2Ijdg/pI5VBr7X+VyHb07K1JUpNFzQ
6kYkAn0+/29A9BH5sA7GvjV4IDoYeYHt/+65HiXJScMU+wdWjYhi8JaaSpubzvmokhgzr/TWc4+S
l2VZjPqQmRgmngHmn42i+x9McKmA9EDxfvXQMWMDWIVqUNTEjJ8BYBWKi7nbb43Y+qq5ps1RGZrG
mQBHMlpA+SN/vs0m5xWCKi/qeuIPPZDmH2w3RPujZa1SxQ7f/Hk+duwto3O6Vit8CNemJ4otlPDM
MaNkoioulZuYdBuwfp2M5KVQ6zuPUIB9SVuQpBGJAGdSBcEGDsfLd7O5Uott0CXxC0+aLbrDDzOT
HmXAYPEDkuINQ1ZMtPyu+0MwM40BQItkGePg0bVvv+lpgTqxQ4g/leyv78tfffntsGI/SykzEfSr
SzXWC2+AIussURDJczgRgQuNmgKXtufRi17rRNiwivxG2vY+RQEiAhAH/rzubcXXHlRdk4hsKJw/
htcglE4cenJ/AifswV///Rfppcf/2PiDy72Sl+FG4Je8N8faxEG7G1Qqy43yFo42nFqZ9ZTQlGWG
U9RRQmT5l+s6RkWiKxuQGLaSF37YwVMpPoEemvypgDzqQ1hltJWNJK+PGww5d52cH+l1i15fS+CE
4ENWnGyamT7kZ00PfbYyjH5JzicUvZAM9aR7xstp4WJkiNhB3hhvLqWnVsA5E2zpZkqW7LPl/IIM
KpTdNYFMlfkvspvNhRkkZSblCWlSp6f9XFjCpqZ6hflu8LgTBPnknjSLc2ipybgATFwEuFDmKVx4
EbGrDpybcz0StskP4smsSRa4qfaVOahQSLZZtyecfwxTwZgRU+5uNsLHZDGOqCAC8M2wccqgTz/Z
sO9jLGgZRVqd/5Su/l0eVPxbhKv6A5x25tV6hl8saD749s/jn1mT/EkhQzZlCfbRf/2C2oT6l3rn
RevtfOv59UE/3sT3N/AtQwnPEPjee5We6OAEukktK8XXu0TK0CLX8r8tggyRlX3qNN725CMlgbh1
UBEladnpQF9dgKRMxdNbx3laIBniQzDR6kOCNZ8qI5QUUibBoGIXoZccTFfXeWXKjRvzd91nNsK8
49/edm1YQe87EXV6HP37FzgAT1SrE41dvygSHYyaEgmWqAP21bfdHXLHap68jDfOtQmtb95iLF05
PTmIuTkUxGUsstddxwMcvNFUlT55XboIke0yCQRwqHgUHYIrT7w8cLZ0TUrwYZAFTeLWD8Vm2T3Y
Us6CHL4/WSs76x9JfCyxnVf2J80oVzpaVPwY24hjYxCGhrr8brp64/1TemojOJxN4UDmoHtXVmlk
ZdfbwxO9AtHOO0OVibd2PqIZwpA5egq799JwIpXL8ivLWNukSoe3xVaPASO79MBRd4I0LFuif6z4
zT4oucouU5aTzVgul8P40F80SH1PM8vxOSCBDbV5fOaaMUGQ2KT8QQkhxUeXwPWQYprmgh/oCNgP
hk9xmkGgEn07OR4lmEADe6Ux6uXPUcr70KlwwpbBjBrbmzKYXWqs4yRbhWrvIwdU/Wf+sIzVFCN5
tIPyaSSRkrdrcj2A1ttFFxDR3P/A2Dum7ZP2qRXLh2xQQelfZ0qx6CHEpxI8JjTaCA+K1Y57OCB2
ZU2NUR5MiCGSEx6JxKje/cTcfw4D8J+cps00JECeMN6edFUqBnor+7xcFzPQKC31Eq/3kDv4yrUO
0NHHK7+oGJ16O0y/4qJ7JHHg+Mvo9IbIGX5Tj/2wqmD1H9sbiPS6wDjBOD4cBHMz0r+fUtNbMpZT
KOdawLe/hzbSyEzIbuDcMkse0kFoWf/iJMgsSA+NjBFMfWEwfrUaxDerAwMPVvje2Nnd4rSY2XJv
+iIezcTKTK0Y5Z1SqeztuaukIZu0IV7m1KKxDvuIphle3czgWLaxqIahNhLeuSiBlmbsY9dKZMAN
gFsIfe4yMMsBGdpaT4EUQhalNI4wIu+R5EbzE8qev2Y6WUtR9+huyWgsegKrJQWJIBpm/8ebTtaP
Jl/E5VFRN72E7YultItzGYtTbQD1IjcQoFlTXxYlgeatemyuVfA2y2SPjzY1BN4t5JqE7xeEsCgO
7u7GwXnnmM5o1vz+glMrTif/ngouTNSioTAZ86//Ul6YGnNFerNrAA7DKkAsdMSNRmRBvKZyz1CA
J9DFh+SNgOhZg5D563JZxW9vYjCZ/IJ83tEUPB8ntkBeW/aPb1bvJ1Xpt0xoUe0BqfDV/FrThEk0
MO/Ji9CmarqTujemH9jaNk4btyRVFDLcFKSxagyuCLAV+Df8ViNJGXQsDdUEHiMCYdbiM2RK52A0
JqMrTvqoBZ4KSOfdUibS0Mr31pbmPdjbUvK9NVYsoFECRFrJznouzD6XalE8jbnbj7S2a8qbEEEy
WIGEViy1qp8UK31MXxZWK5YZ8u97zlASeD+aVXGghO1aFrxWnks3BezReqgqFUBvrZ2mpBNFvCZL
JI15ln8F3wEkjB2FcN3kngN3in7aBpxJvLyLBvqyH7/AkawP4by7uzu9C+Ft+cQmHgdDsQOZ2dpm
xV+Vr3NwrODWDGRfvL+Hbqe9ZukhObaeNBM9fWhpkOcGAkolbiUWvQLwOZhs+zM3wb/MmhjFqW3S
ODrcwb6ZoM0SQCaGDKlBCbeGHw7WP2MS84vd6gp2vEEgC4VbLYZgzvOlYsU3hWHZqDsZwuEhsA9L
gIuqsiujSDltQ4AR6GHQhPsy5dPUEWNz4ntpZKmjTuCUKFQwUmZcSk9IKp2Ml4tcb3ky8oUMHChm
YT5gbmQDTQBZ9tKxjz0CIRmISn8bO6VV3HfQm0c/HrSmcJtPMlorE9zxNlhNKSdYMVGqVweesqJ/
eDxeCxiR+o8p0CPdmm7xr5kPqntZRg+RowZZyLS9l2lgJfbmXVw3rsW7BeAl1NBnE/wdZXzXU37e
Xat36UN6omVx7zcEs9g4lIeybkO1zRvyEhDQeAXQ/iK3QH/iLVrYJ5SnQHN+OT8h28VbDP/3xo9D
rOXdyDYpCFN5KVp0GDfzhTrIuqeBW/4ZDs1pQTmXtseqAWe5AuSMY5sHzZ/pswBsP9H7cfxYENpi
Xs2dQPrkP7ErMxB0WCwkLVnXyIf+27dIaWT6I4cYaDUGThEn6K9SAmQVAicG+BymVdH1im10xBJ4
WM26NaYFrSPwieP15dmFaxVTAYW/jb5K7NsBhUAvUa8NpF9noSzbZlV3X95+T5utW9RLtbg80O0X
+Z+vhN6dE4zRZwMi11s0R+3pI38e4j3A8arUG9Zpi+1gbKH0EVA3j+WQH97SQ/Uhcskxa99Coaev
Sxu8T4+qGLP2dLAZbS5/Gmd67yaMU8bn3TV35m81WzWEHpvDX18T6pbvotbajHl0pg5pdHkX7Jyz
ZzDG6WTmRRxdaV+J/pA2F0K9tlGrZrf1zo3iEUnmfZ65HKZk4JB+QgTUbpnGQxxYMeDCJagWQgmo
ADp6MChT6z9STGaHe8fcHpkrVbokG+BJwuhgxMrW2AsqCsvqTq9a2W6SiN55lEeEq/XBb38bl+QU
2WgCOOfTv7hKFWiQ8FW9Nsy+w51avT8TIZ5W6G7aDfsIXJwA6F0dqZVM51a8Wzm1CgW0zATAqNkb
JanUfsQJjXBVXL22TsrDO1M9R90G2LBR4FATrDOMo27SS+ugLHN4p4k12L6FOrWnthEIO+OwqK9Z
F8LOCI2iXIJ8ejKSrS+Lt/VugoTHcAIuXYTA2J/ZwxQO1dW/ZbbAYIOntYaDg6q1rNI0wo4XtzTq
qcMKpM/RnrLNEGnxKJTCZf9Fd1yzhGHTz+MmXbgqjXfXDHQW8hrAGqCaosM17kF5ptWoRhLti6VT
TvFEDV9O+fzwqwgxmfOZ5Gk97JRi0HsnJXRFXZ2prcs6izYk2AS4rNpEJaywLmsoKYaJLtuE1RHU
kuU+0RJfxCaGf9vMIgV7LkGkr5DR6sWoc5qHh29HfICqQ+JEL48c3kWfXmHPOrC0tDvqa68u5MVG
67qo8KoYYxJHYaejMqfAa7xHtBdDHMJCndsXDvkSNXSgspFMnlLWGHN9fO4shnq6l+aeSIvCt0ai
DVkBtHUj+fu+65AVTfFVWTGyhtIpjDH6vkG3AE6zsJC1JWIw5+5DLHI4lv73ihYQn6d8RmiW0xGn
+/fmMdQQLY/fzhbEt59L8tVps/Q6eP5ljQ/y/42HomQUBgteqb/euGqkJwF7juXwS1yS9h278jFj
56fs2ugSWhqI8W3cMWkAo6FQK/nqybkuxgxB3iMGSkDaOElKvNZZOUWBUK0Wh1W31NgWmfStdOQk
mzS7u+SDNpHDJS73uuVkCgmKStzFmAFjbNmj6/Owt0ukP6Y8p9Pl8M4N86vgx/8trUBlW3QPq5aX
qSKD3RLBpJoOoRnwjc27C41O2Z8q4TOXENz2tB4m5FDNracUu8+H4OVXoox5SOqAKJJTGmlJkzJ8
L6pub2tGnV9xdkc9WPkBGhS7aKBJm42IPYVYKVEs2WzqjDLCZFgprVuZPYEeSAc3Amt2dtvrp0dH
k0W26xsVtu3Rba33u4cgMlxUDR0+3c124sJi9P5WVraJjxDcdwuFVo4GZ5oKF0V8atP7fu2qllMt
j4tX5zWC1HTuOfABuKmtVM8A2Fhjj7OFjGsAabo6+jWW4v9TuWy2Tdf86kTfzF7Zb6m3eagfDmxA
nYFskaUyPIgVENAkoKW0SRKfboxUdBQ7J+VhI4+JR2RUn50O6yFYpAvyWJ2Dr1RkqYyO3YIMT7+6
NW0o5lPVMBzioGBqUGC+35H8Ryp0EEdaylbZOvHUWXnQlITTnxr+uV0hrLR1Lhr1MZZ1UaMCrXKz
+VpAixrrdxVMxVwBKFFlU4xCZGqliz/yLq9R0L+93bnwIQyhoO3G/MVF1taVJD9Zq5ot4Zl45C8E
wVojUPkJ4ip0nOSbxMXTX3kMF46H8SRQ0pcIlRnWK0kf3hsL3PfuMKs5k8sFsXe6CZ3i66GBhiBO
3FrBFYGEhh+TayWsJhefnICaLNJx3tF0swzT9kaZvyIUmWcqayKHRy7vGpZte6iR23dikfSBx27D
/vxWhiDC9zyLkXs60Q3CmJQs/Yuvpj28WXpaGf+e7VKyKYdSaowvg5T5P8DsesWoY9Y3XFOF+EX9
MzoM4gtcgdM1LNwbEQJcZDuKNg6dSM7dmPG3xrYZC3OvrQuswwTE2F3ve6WzNQTLn4pMMVY8g3X9
mDkx7/nh6LgO6rX8B8bumq7VReSMNq0GYXQ6GNqG8E04xazFi2Wbex2HHyzZFeD+pTBkEgleP/yP
JQKff+E+9pZ+zkS0777XLNhwd6UR26hkkfMLt9U6pMf7dK5LMbm0+SOKKT90gn6v3wm4yEGJwSAS
OghQjaqpAAXfkdBu/zPsscNz8nZgOwxnm7yeo3UzqC1EJusxUDfwQTXitqfbI61jIMfoRQauBw0x
O8+uSDeYMtVeGp/BekOy0cRpC/uMcGJKhXjUiKZHe8581LhmpYzy5BdwgBv1Iyqrlqy4hOcCmg/8
ceT5KiM5wpkjEyhrcQ+hkqZBlqp5rR9CRvc3K5b78SOkF+ekSjFOn9iTX5E8cinpn7AJPywgeVsM
4sZ6/vg0IdJi5lozFw9TF8SqGiv1BWrei9H7x8JTjBZD+3Z11EXh6Pad3Yq1bqa6Xa17kQVYykEn
zHGlVGg4iBiwl4obbtQqpl9osaozPFuCYmP3PtLtsF4PyZFC/G1GhsIXrtIQZoQEFON7xeeCwWBK
wS8ubW51dlP8TEoycIbJqOHFl/uFLq7wimek+Uyof7LHm031yh9uqsuSbJxn/H6WZUObUNNrym+W
jHZ+mlL4h1ePfIThU7cp9WpOYk+H3xtys38xvIKkFaKMS1jV7VxpVul37CvvW5SVmaRXtYNtUzbv
+q0MBdP77IWBRPnwjPqhJX6DrGvM1nb6tBBR7J6BV9tC/aXcmqVW5gwvwHjXpqbSfBUNoP/YVCGS
jlN6qBlIGe6eYaYWTO1MDivrlVdGV/emsD+Tkc9tMyCmpv7mXfQ311yWG2kyytWomRhIRVpFjbI6
+2JObEccthJxkqhQ3+OgolQ9XQWpNzpbcGCI9CAUvBScmFPJwNay5EsRj+OVURagc0fD918a8dHc
PH9ZT4a2wlhkDYbvRbdont5lT3+4pG9zthlJg21sI+iHk9jWLN/TuruQtk8z/fYbiGj7tKtZVXzK
uNr6TrNaOTosD7H0bhWo9KQKJnaGzSf6LHZzb+E5FpspRhduuMg4VbSmqVlhOD5IhCaOqzgoQH/w
eYIWGeRClYJnSp2fQJiM7TtOI1lyW0mYs27QKirariCvPTNqMNLenPuPseN/41cIMouovzBjPPES
qHL+MBMnyTSdJ0u3kGYmW3Fd6RwaW/KAuWOc+27D38L+9q+JoymNq8X8wqr8YFZ7/hBgflEBlXio
DRxaZfVgX8CplnYBp848ja01Ib2L6b/i0N4Z6nfVdeQV87oEQduUPhyHcvYPvwRaMDMbJTSaTwoU
v56DXBnhRroPzRGLvFTpCbobzSKu3iwhGr+X65CBnkAfE95iVqea1Qv5/2wEWpZ+kk679KKn3dzv
EjFJ5Ca7itfRVLHC7Ikr6koFIUJRP+5sNLAK7MOAZTfCDEQFIzd51fEPB/ypLrnQeU1AK2ERcqiT
d+wMW5o9zAeMuB70BAnEWmB56QKTHoAncL1WWH2PiglamPGb9mm9Atk7mRovzS/1mQug+TPbwJQJ
9p26F89n9GNi6UAPAWV08BvpLE2GqRvdr065nyWS616tDtgOxqKHagnXKic707XLBCRJnXEUbnZO
3dmCRPNtfncdXqzqZPkapyyHQevClanC8UM97u7W6V0Ugk9o9i2hAGOZOSk+4/mBdMamkT/ro0VM
GOMr34RHzUoC44roSKiqaDAdiMHjC9IM302TyzCFqZ7ZVevnqJIoqHnBoqBu2zY6KNfn9IeXSxQx
dEYsOps9zjhQHQp10dG6mgrfxVcNQR0I0UIPViZ/V1Hq62RPjC/L7goWEa3/udspw8veGW/w4DVH
5szLcN6CMrWEL+J0fFQ31G7GbE54hT/xSLE2cSDnl0I6FoQKhObo5CcOKgHP7KxFHfmCIldyEpfV
RMwib9i5E6WV1A4JwLtAm3B6HgBy3fcuaN9KcaOzQoNogDEEa2evoy6xEJdDuf0WlUeES8BctxPX
NvNM8u3602p/Vm2qm+pb5VTMvFfAQ/vdWFXiZeS1TtPipVG+ytc1m9G0OIxPt88NREiBociLLTPv
5mWePyUv27x94RQTXZ/kO2btkGKBY4AC2HI65ORhiq1Mr0k5Ndpv7+RNmnllHTJ5gpuN7k9XAKeV
GVIzWbOXYYn84bYQwyoC+anElIpV96bgznk2FHzqYCqXYTPlV3+sFsFvVfYvyHoIK+OBWg+9WgVu
Q8nrk0l5+OM+OgEakCI0uV5gCHyqGfI9YwzJy/XmK6Oqa84P1FhPdurFugATAN6JxZFF3eL6PpCj
pBiObAvVYqMI87n2vGGKwMdgw4To36KGT1WuGp9nNTAbe/CrChc7/VhVeTP0Ncall8ejdgBnFyD5
hgjL6m79cmJTtafmnYF3E21vp2Ts1UnNvdk//2P7U4DXxZF5tvySq1KYLVThamwsmIYXczV8W04l
GeQ6s0r/winMPwMFNqMDrmLzYIu0hCa0fSy4CDu6KHN+iLtJBqfKJWLl2mUV7lxCHiZxVFl7uhTO
hsdYlXtDb/DhWrgIreXcVte+ZQU3r4LAXQ6AtgXImgHWB58N/Yc0Fj+cXcNMPsLD2Li5I2k5KTSr
s37zX2fJgw1sZleR4z0z2KnxAOqCk7sS7PiobI4GJja0cXNgsW/2JAA8aXes4ymowIA6zp8ZctE0
P8ugnMd3UBdzNXW1TERp6of8Ezm+GHmQg2xHLzrUVNuwLQf4jOubf7r/iKzijvbmR3Z9wZUK174A
Rqd163OAMrK6AFtbpcxBBolfU7moHwnSV0Hs1ncnzfJ0z2UD1P5sHbo+SbNYMKxK2YTIQP0Yd0Ou
qXo1kL/BqgrwgiDpfcjrWaWyZpc1PtWXyrTYodVV18umy1jfw3A2GdkSQVtXAXUIRJPZ7o0xYC5J
d6Y7Mk8qBJ32dJp6SgT3BXFTNxhWQfGwX39PKYYBDjL4xuAx8bsuOxYprfXXn1/HGngfThOZJl2N
50ggCXLCGv+cxssOVjuG+t4Qoo4VYfsggsjs0XJYosHkxsLZuN+6tNSX1hnxshWSnnnoDuPGytVx
Gm0dPOgZDRgXv4KkxbgvW81/CsZ7Fxzqu47bdwpReX5HtoRY2dSqiTEupGv1tCjrvAeoN1eVjSU1
UYwDv8P9QX2TlIKkDiaYc0mvHAasinbgj7AXQPpzmC81TD4kA2F3F3GgcfjAg9vlY7mRfLkhM833
w2+207/MoEdqEdTnHN4Vx96RjnXCcB2l3n86b2rcFoWU8/T7ohM+230gRRXXG3pa/8c5kHR0GHfy
5jr4RuYFNbSrso0c5au61W/AdawZk9wLnUeYnUJ/+eq0cibQWW/8NVCC1V2x4pPpKII7qtOW8W8o
l9TadMxD9aINC7OAi2vzN2Gr0XueRr9VoQPABp0VsK90A6BE4fFMHQb6IqIwnyiUKosy33ZkLgm6
xEo2H6oWw+mSVRmp3ZX3hq/ASBP0OaElzTXhf6eY0ezPJeTbNh/fnJd8V2iv3rBqyPe6qQmY63Fx
byVUF3X8bGrWOIxKpuHJkGRg4nahImRZiy/e7bjXed6zZx+X/QWWK81HGzlvMD2al56+H0PlohzM
h509HWjq9gTzqZgQgRCuOdwajHpwpdCXH3Ts/QgIqmjvEu8l/UBTtf3Fa2JrWe2ttlHVxoZU4djr
pPlv6WlKd3SZUARfryl9liZe1V00vadbwTvsi3PWV9ZWmKSghVFWhif6kCswelk0xKofxSeCa8D1
8hEYzbqqb26ftrvLGB/2IdOFasrOgvl6/5moEMjRRg5hdd+HxAek6Qi6U5HAB+14zzquT4CLSTca
gz0Xtd0e+RvhR/SKBtoRr9DXBMvifNggzBdvbbW+H6NmJMFvM2ofgYgGUKLywDMZMhMKzZU1Sv4I
lXEYoXltz/O0E7LNjDj665j5w63qTSXbh2k9xdlOgYg355N/wwnswqYQ387drQkWykMRJ6vC/BNB
Mh44n13Por+Iz0OcvFGOBVab3D3CjHegXqBkea2Np0nw1m4FT1EoIqEnBr9nDQIXbuxRq4h0pef3
Tv1fKjIAHudxPB3WfXnSsnldUvMp55KtGM6ibPZSiaAESGe6qJRaLkipE4QD/Oa7sF3B6LENmCb1
zX+5li2NpeXo53QRGvZvwwqpY0wpIJK6nYmRCS8Ctu7PRKDNjjIPWS32cgJBLCbQZ5qrLY4zndGz
h00PlFVf/8AMQvfpPjidXwRit+9YHnPm4oCIfBBapD8pOJ5a22c3vTjHmnA/YKtLKZO0YG75Neey
asP9O6gctX+F+75w0zl/HbCEbQwZr13EnFT8q/r4MPRE2zo6OhSSKaiZBF7wWIzqypb4gfnspDR5
McTnhOCqvojb1zdStHmAy9WdrfxXZGgBDrnON/YbyWHB/vRl4kTWY3qYLrLjsRY8K9ekrAOn5zSB
exb0SKYADTjx68B0/c1G2mQYMXBt76W3ctglnlHh1/RZnBeLykDhekk1Sq8KVyCqKBSDPzbfrxP8
mSmY5VZhm2BkmXbO3oXsr93fuJWRz7lmMAyL41hukH+V0z+Oz/Vt27SW1tpwOpWWkAL51oy4AmXp
QHg031YKdg0O20n8ucYZO3xOv50JwVb/GKKl9njUAxMYWm9tyoV3PV2u6LvrncVplrDRctonrCpX
klepRI+UUdCGYdJCcFDlTt0Qh+vhF/Z/tl6E9VIxNbg03CV+pjE/hW5sH0KjihpBeGlH0qeKK03f
fwPWCkSIra/c7jJuYIlgY+C5vXuWsTVMrDcb7Z6NRYwEX1k4WGD83cA4UQrshUo5LDnE9sqlweNR
0b1d19UFe8I00eCacrbVf9/t/E3Uq3YbiJzeHDw0bp8rARl72ltBmE298lE648EnOK47/UrYXOrG
F+lZf12fudLgcuhJXz0L0pjleFpegKaetOYRhQdoNXt7RZ/VXJJ5IqkQFhmGEWxf+CpN5UMuJPQQ
aeMypZK7yYOWuj5cqfbs0yLyFIuovUQ8ssQYMEZidpucVShooOofSJiC5CAp1LKGvdBGzoY+z42y
GOXrPy4qSn3T+FWhdsUxg0t7qhntqxJbKBZUNCpjX+OQCXalgpXDsgrjLtbnkgQ+dTco1nsyEMnH
IVnCv9sOduWDNYqe3K7TSP8usj2SGh/RfXE2XAHO0uswVfGmDYdtS9P8ej5WliK6REw5dm9hQt7N
bHTdHr5gEBaw5kRQk+JTydnZokh0DRC4RwZUG7cvOahcFlY+6hObMAJ/VCTgybJ+kvcS4nU8AHud
jHhsNhK0Gs8IpleudTpqCrAWN00nhX4KmCXOkcsJll9qp4bDzD8LW0Rr7FbFxUNbXjdiuV/aVEOI
lQzxlDqkalycKNiA/YbUtcMTrmvUSbLfN/kifyeDtuASoxfAiT9kvf/76J/HH1UzGSYsfYgTOteS
kAf6tFFWoOQBjpbWZLbHzbCAKs0MQ9GBlBSwppg/rktD+minudVlV5CJCwT7XiSoVnEprXgIHG5x
j/2kZUvL32nu3sA84AfFAO018fGdg5co3E5H50U7mjya77dn6IZgjC4p4k3ui+PK0vseZZVt3F4q
FgTdwfVyBw84B9Be3PbGVNbX86WuMvXNww+jSl1vC77hHIa7f31eG8SI3QMlyv31sTSszzDhCyZN
5iVND4W0tGVZy4dAtP3nqIWKt0r49Ib9oUji8g6xGkYC9Z42gsmmgaQMXrw3lvR6k+7nrlahdyjx
pdAoRDT/6ilYuS153OWrJZMaFwFMPy6qprBZdndfGY2N0GVGXHgxatB+buLEkST5DWUFlVOvkRw3
feKVsZOvp5Fsed9n2JQAWcSRzHgP3i3FJJyHJqqbBouNObXFv8ZiJuW8vK/x6T9JGkSFfCU+UGwt
2tmrCuW/bb/i7nEL/sIjRtpOOX8WeKHRkSIUnOgsrRMAlo5g/SgLnf1BlVJchFY90eW1MaEcmh4F
sWn8hQc4yFec2UjmcD1TawxfS2+AWSfM2ISGoUDwNsm9DnTwFw0iRV0Lu0pd6d18OehgJ279sq1T
5ikxkmKRQ5p1cduY6kR48QdHj2gZ0GnookW9lC0nqGbH2peYGINnn/dGPLPInMBlgx05qoyf55Ps
WxsnUOK88R8TWNgP5V8QhdpnAD1W6eMzItVJOwXerigiZt5DSun8h0r0/WXcEGZKvBUOcnJgK3/w
b5CW7UofFW3DOaVDxAKe267FjvFn6t79RJBCRxjqo9GwHN0YYzR/j3LjCE0rfzqKTMf6SO3FXpZh
UkcapoS5nuEo99eYd0kyG/8mXbIUHdUv7hHVyVuVlRlJ29eHIMW7SxgjDoeMLHkuQGwPhX+9d4FA
BYXg+bJLz8a0cVi/IOJv5Zo3CtSIIh+GWrN3R10D1mci2GGxI9IoRQEkWwrA5lBvUkeo4JOhdoyk
GPTs8hLZjfbHW4LRDsiEJQzDfk9a409PHBlIx4a2dmLrPIroGM58xpAT8vb2vgDu8+eGCxfVSsHZ
tCgbQzRtRSvtFldg/l4aUgYG+vveHg4nsw1MF/ZbEZrcsl88D7sjrLt/PxQfq032Y9VkUebemzyL
nDEssCkgPfdLfknGXVTQkxt6HxwSLIcW30o7mrQj1fooWZO/T6easlaHK+TnxxgNJlwKwNOB8PO3
r/He0lPm2FL0kzZOy3cW+g0bBYvucQLE6C/szxb3sfP2Auqp4frrvDCr0LBF0ga1bg+8wNlEhX19
4pGXySyoExnBCdPywx8DyEVcnvg31GMZdukn2J38anDIqU+aVuBr/5IPbjnCC+rxfLbLvG3M22EU
eG+CNcsX+6w4G9dksKUGSBODMsnNDJeHLVFUAE85kEkhRcnXnXzWqCa+me1Z0oc/8eNlH+E5EthZ
fZnDeJ/EVU4p7c7hvyAhwxcmtB/8MXuZS1gbRTlhY8dZ2I5RzRcTANYbrW/U/ACcoebwP/EOASiG
6JQT3EsXCQ2JVMKW+eVjCP8j61GnsjmX6T4RbCtt316hHnDvLy0uwHbgtiUg8e+y7rqQeVWhN48a
/adptfBt3pllglpOyNcsEcIeFNCzQRa4d0x2d/UqurIYky3JYSt1NLE3VhdxVHQffSWHwnv63Vsi
3/Lp6KtBR/t1ePp0nBkkhKKSLpljNINp3nJZdk/WqtElQeOmCd5zLOXXOOFmFo+kmidYyKUmA3MS
yeDCjS1TKfB28WHpJq4OYJ7IDMJmngVG3dfejLWKIgrOCRplDAELzc7cBBUZzCC6k3r6otSwAXRn
Q6M3+2NpbCEUA7r4aNZwodYQRM0H0RrthxkTHYgn48i7uoUCIoDbfEd+Io4jzcQMojYgVQwXVchb
HZeH8AJLM1ceiSGkr638GUi4i46seJXbSUVGc+arFFLfWLo56wO+T2/dqdRzclbkEdeSh94yuVuB
PEYMge5dyWtcwcDyI+E3FwtEJdm3JRRFGs54jffpdhWq4tC79Q7m+q11C8xNSkW4Az9sW+2NZVWw
DUPZd0tU009dAF0gyfeudHR8KIjZ+oRLdypHuY+4DcTLhMkvCkRH5524yh0BnIEw9cdIGLi76UJ6
k9+4n2Oj4rUU+YZQ/ax52/d2sP6wvjW+oQC8BhOCrMqxYvF4sqoiqmEeW5aHxcTNgjLA6bB+kaGN
/KFowZ1nImXa+t8zxrhTiSvskuTrKVWgeAARiyvtL9XhzCoWD4sgwsX3SNp/EMwa2x7XWKhjc8tm
JExQrBsAkww16T3kfZeCcoTuxeYBZHid97gis0R+iXmmxAFX1QDQ2CbCmpdSK6Naj8zM1cHSKS66
JRc+eepxHXhoUhi8j5N3oKFFBYiXx32YZkJrzSoHI5UUF71X4lLbvYxx6lhGx21+QO0pi5mDFnxQ
UWX4FdSbz4sfn542K2RqUbVYMg8/JwOo5YKeIuRNgUKj1Ay+pfyEiF/cC0giFjKsqoHQIE+vsspJ
yMvKGwqqwNQbkPULJPornlEHbOwW4RVlVLU/LQxnTkS1CEv3wfIGBkwxoiU53Hmd2J6FdnKdpSQD
OOnkYCfybqtdo+eC2CmHQHOGMa/OvtZ4HrburOZJCeH+1b85UsdGoCtOa6txKatDMeVOlH1g0f8M
G+G0yupnAwzxb+fpaI9y8XmDqMLgRB6aAMUnmFYYn6jIYTMj7iiIUu3TuYK0S8f9HOPv5XN7mtd8
JL5BG2j3jB69CRbZAdYK2MXufx3KWa2WAviCQEjWqtEDSiWNNC3kBomrAd614oClSYKbZI4k1380
Rwps0+QJUZqbwftPGaR0f8Drb91n/OeFepEjj6Z+D9wjO1RX2UYAodh/JSQguMCNiS7Sp8fRo4Wq
TkB810IdgHKKASWp6uyIIOsaUSHFaXb4F2Nw67PG2knUCk4PNFpowAz5xhx32F5fB0q2dbpL6lGj
eKF50WdT4JMsFHFdOupDOe9ZetpzhXt90m1b5EBdbzstW24Fc+WOju6jrg08dzCvWlYqBiy1iDVB
wYJt1WzRcdWHb8eq26j1bO+fLxH5+hOQD8B0oY146mC63LZ7h10/0ByevctHGDMVrE/dijWDwsh7
/UpvdmZ7duB8XZlrDRxm1BycdsZTi8yqmpkxoVOOrQJ4SrcjXG8ELfmtQIaN/fYsx3u2tdF6aA76
NqG6Qs1OMV+rHoGpZLcI6AfjrOJ1X3Nnl1uyfNa5Ou1/HvPc8TI6cWB7HAltlbCcaKh3Z+wwGeXu
AbrdG8msybhbNYbDUrLnH9xQfZlwebPr7n3pjeoS4oBo05RDAtrPfD9wuSX23OPZXadhtqnxWH7g
5hThAYeaHTcPgNX7f6lu/glH7T4Ud2ZY9+EGgFTLaUiI7iFV9V2UxzNJ4KOv3Ah3TsOpGvhn9aLg
6iKcg6aGN1Usej1zCvWDbZP3DY/Ni6lq+PZSwlPcN5sbR7svgfUbHN6KSrwJLvXUiM3aJXBmVgcb
HOGRbrcDkf3zmcXurdoWd83fC+ZTZhjYTrr9AUk1LkebDVa1x2PhzAiCJuiQbf1tgT/K+3EsfQ6V
/tzNXK+OkmOmSTTaPnT524MRnHaObTN0F3pClSXIQdIqi5FOplC7iOyTHLgAmsad9soo5fvDayrK
ijFfkyBY+I8F78PU8q0Qb+WrjMrj/NHyIn4WDC4VAEx2DJy1MaM0FgaNkpBVJ1Dh45el8/6IBkP9
oIg97/GsPSAI1mAoiCP4Uq1/GyYYcCuMcfHwRKMVAMutKXHt3IED0aJhbKw+jApE1Fle1EcNi07V
8bo4b8H8HcFS9cYdVtegr9h7L9Hjl7I0PpdZyTNrOlBgj8ASkKs4zcta6vTCe/qnyfkdBMQscFqZ
kc+e8Y/e6oIKdnyu3OFWD+7PMF9YKCD8uc81hd4AIakuQfKG006nqooqso8YfFenIjZS2d6Gf8+5
AHQwBhyxp6L8oHvYH59S0e4TpNQnQ8GCOMtRRP7P3plZVMbfmB57oP4IeUlLunMcR9VxNOT4Qogx
6FqkI3Po96zXkfQPYqNfNak4edza20QwaxP9dHZ7qJ26NvTCDfb5TWIq4bR0eZ52k6RTn7j8OuM+
wdJV8tLhs5gR2ywN9d5lp7w5va60F96ADfHypSz2Q09/Fo0+sDG8Snj5EHBLeDgMcIyFV+Yl8f5Z
l9d8VPszH94EjQg3OOV3x5r5DL6wtAT4WUTQjKd928di92MZe9808W9js1WFlW7O0fePaGFCW7g7
yWMzCYlADyOTI954+J0aQHGQvXNDB1+N7Hz10QvhBd25FqcmLzyF26esQ+XS7Tz0arStU23aVnLv
92e0rRNuOaol6EyLB/vEkAHoo3N1YgC6PgyZiFZofcSUnzuT+6Y7d7l9K6vDIktVjx4zIlQ4+ql8
okHfL70Sl6PdxViXPDyyOMUOZbtoEyoMcfDcYGCUKIMpqJUEw6isT/0X/lwK17a4VDI0qEGeLJhE
WcBpcqwlEG2GZuZRkmcwo2zfcugEqrMjF5b/3kJUq90Vrkl3PWLnEanOGeQf6+331zfgZ+7NXj+J
6x75DCLRf4X2GGaUOoV7Fa5uEqPHLcp45i2UM3DYmOyHcqgfHwMX7X/wnS8PLFIXiv/+MKtKr1y9
GvofV4TqG9CAeAAH150nhUNF5Xvivk+qi3LYOfPMgF5+bnYGkslOJfRL6l0qhIsC1pkzPLt41SiV
xG/rdHm7TdV4TnUIIOUy61GIa8tcnLdUKMAQ7Gp3168Z0D0AlALx7JmO3QMIf3XMYqOwYcdvGM3k
ljl0G5T2uFGie1phfrsqUzdd/MmxJYrYys4Kgf0LeKTofEaaGBCJ/ibEU1LPUlyAQBO7B0JgxKEu
+Cf1bt+Q6ywCBz/YUDQykSSyFlfTrv92mVUTeILYP1jm+XzirNFeFu0OasBfG02+PXGnRRqw+nHO
g5PnYY4qT7K6hfws2mcw7SVBVkD8sSd3uJOpYh3UBCTrog4ngGU4poJqV9ex3D2Kdo+DzAVrTbVZ
dqb9MidZ2wNAhIpe27d65pZ36N1mzXdkQIxuKvZAvT44RA6i8KJpS3iSEIjzeK9jfVTNHxBrNjDp
iJJd++BVQTf046UHO9b3md+5Ln3ASbp9bb3tbqcMjq0eWlyd8vjTi6ufpViQtxknz4OnAJ5dwLlz
ueD3ABPtAJKYF6x1IwIUEweXWi3T856MMzgGLQsWGViJciX7jEYj9ifKrqHftUdBxIKFUdWSLw2L
GdmCZWWOuJn9iKAasau++SA1ekNgSI+yD0aW7EfRtzRr/OojlzhvW5LnEgRIngGIB2b2bpsDjMGB
mW8gmWXdzAshgNof4zYfc2Kklm/+jFajiaYjSPpE/yw6/7VlAPQH/DWlev4MVdb93V8ZEeZaN1l1
zcGUVdxvaxdluTstEmIbR3lGhBT5kiRQX2R8oyJGqSlKhX3044+eqpRjkLu5yTbSv3a/3mfKwbkC
/C3pu9VDQ0M7aCb8MZ8NpFl1USdw+h9EwYLJgOsfJMriBoO+ntaG3iosAOfwMDCN5JgeguGh/s9H
r4huOf893OAUji1NccM3VgMvvDgCrVIRqqgQAdqayb2UwO9XHWO+VljM1WIWq7u23lSaByPMzAnq
tkXHLXHUd/DVjlY1sudhL3b6QEYbFNE350Hs+V/w4KNj/vCR4Dsj6bZalGc/90H6cqBi1Axl1qjl
Pi1gbGfe3f51Xd9DwQ6ckAgPjE4pPV6vwU/XNEM+jWcmDG06zCWzJ7mKt5+2ixV6I/x3IlNTQ6YZ
n/BVjpvtTDCaGBSQJ7ZpOLj/+6t5SOciJNOY+01Z3yMAuve6DgZIbDxOxNb0kOVjd79C2KlMW8br
KAfYamPZG1CIitzq0K/sNSlVVvl6gSPN2NtZQAUNcqj73jYBlN5HE86U3iLUxam0q0EJkq6HUlFu
db+EtQy9VQ4MCCBfZ5Ej/TZoq03uk9rxt46fXqMWXbvcaf6R8kgfRdqnTWhSew1clbpcB5H8TrgP
KwfPsb/LMKBWajYV4FEsAOOURTGapjkXt3czhphlz/RnchOBLfg1IwhT5nPuD5/uRGef3uVokZW/
6tbPhXN/Q4ZDud0qJemhZm3tCgKEK5HYep77zve9tJT4vGG4XOWTBHJ7/wmRhRfQTsGoCLnGFKT7
YJPtouhXiBEE9tP9ndoULihYU6JlGdMz3/Va1sY4S3I3CMy5Bvd6molwRcoF4gtmshrBJ1iP8gjt
GRtOeytyvi7Pd4YqB8jUqFTFnejEiYaPCCtCvH3BNPT/1q8asiKQHpkLaF9LM0HE2rPvMGdoQXK4
6QvQeLrsRvjVsnQz51bN9dB5xuJySPQBbBgTwrgNYWJe/Ni4ghmMltq+80HyYj3FCO5VIw5I7fRX
MB9CW/+SXRQMkJDC5ZJ5PEht8dmHLYWACdvN7tupEnEIXfsbv7YU/HTxiIB7jk1mOTcBt2Bm3DrV
oAtXN4qoWoITHdjhi2sGhNUfsZVdw58Z3jfbpQdTf8oI7kxSE1WATZ+3peiwQTaRvrT+xLBUxrjt
b2Sc0I9crVz5KZwcEdKCqdgyGBvxulshS7PSQftwDNgit251WfwTgXIoYsDbZChmCRB9DNCP4ZAR
DocLKC9hTAb2XCfAhSDax/x4MU00b/cxQyrU1g5cPSq9KCflOhLRteR5HxRD8pK1T6zzL3B5nQ7r
FtQRQ1A5xXKBVO4Xi+Et/2ifOt2EEsVmoEKWIBJHkwYZseAdxPcdXwU+uYHc4Z+j1p1YrNFIE2ra
5IB4v1/BlYomjeJ1NrQYtUi1cDud+scLis02sD1ZVMdDC27jWVpGYqCUQwqgxbQWHfwLuFUgOrf2
/d5YYzfl1Hj3BrCMvFhyeUU1So0NmjKNGG5qtcLi1UImm2d4En7rB1RT//xYNaK+X6a4rdJe13WG
r3Bgh6A663eKehSRNuYvFurOcfMcIyHvofHE/RPt9FO1B0MzXxKc3k4EOjq9/507nS7PdfOaZ2xU
JMquiJjSsVY2AiwiUtWIJuIr7Syg5qzUSj/2u1IeEx5gQszDxE0vGu26Ca7y2OhUezrMoxQI0ezE
ibGMVEr+1BhRhrXQWx/qDfkOxu4Uqp8nvVsh/CZxN5RQYDDlE6svYw2GIkoNRtLUxH9qAcFDprlr
rOCeL5OncpMXJJz3GSZslNrbh4538mhp8oV9q/utTh+fzs1N4puL130JWGuFtovdfZdZWaQ+hkPC
bLjmhK9y16TkcnSSOe+/+7y3wJn4L6l9lXCOGzI5T2kLp35Ib1QFtDLvPTx7H73luSh6iwsqQjkJ
9R91O1xk13kdriz3nPzP20iR6sMTvA+YjjF20uOd/vIbWKP4w1bs0k9gyrlF4kJvg4A2wtn/pHQQ
zkKWpiuN5Bozopq1A2Y/DNZ/Kt/s2ezQDF4/IH6tjlMpNMkszwtb+icu1kXKhBNNCJK6wePtbREN
o6dNmbpk3h9/YgMVl4L75xld3q2fmy/QxuLt4ngiI588ppLyW7mhLtiW2eeGM5P0xYa+C67fks1u
Uk+7krGyt/bLG66XYDJdo0XlCB5Y3qKirxKpu1tIb5arwOL/8oVL79ZIjB53qt3aVxvnpIC4Pwcx
ZUN607xpfS3FXVGlPEzU/esL7NiBJ0lnt9IsbaRw1hurnw5Ndkl0iqPY5pi9JUvWkFZwWWaAQ3IU
vw8de8q3o87W+yre5bp9YqgvuqfCi87/jeSie7yyV7WL0ZKINLN1SsD1dp0rRMVHCeMtBpMfBfKY
6YNWOIFpKONj2deUxiQYUr+xPw8zXCmqzTyH3OAsQMnK934Q9/u8UOYXOYyaXaCFqMRrd+sx4Yyb
+vVEpeke4kgm4yFeaRvCIL04rGiMSG0evBByuyIk0fRCbS9l2kJLZci0UsIo7Kck2g4Wb9pJaD8A
blmC+EkWmrBcWVoMnnz+D5FIQV/JbQWj6ZRB/GL7B2yplJE9F9NMNakpzXkeRbA3KmMPUUWShiVS
KyElwduXVZ0S0i/x77lSplERd4nWX0INQDLx8dIHgJ/UiHJXVc85+U7M6DnlymVO4DvfodknkAh1
xtalTfNbaBheLOGyCPhu0VvNoqBKHNurYKDlQuinLvCl6//mTidGLI9i0VxKCca51Ye2wlGRFluL
OKkkvaGEaUmD6jMLGwb8nwCTuLKZyV0HcZSfcBewrL5vwJPbBS1lNIJy0o1GfrxdoqCvhTsxFqSI
JtXVF95fjgx1WQuccRzaz+QnNNcwk2/JdWrDmxG3x1qUZhOHkYJOrAN1AX0orTqBMTSqx9Zs9vDu
yHp08V/7+2Dib685fcNZsU3dPF3mfSXzwaox2nGjGYi/JcVXLLx5XQZ8HRumAm5idt+o0eT6O6Sy
6v1q9e006QeLaS84/C/BKHa5cWifTaBlvUzp9ztAKtouPw0q+OkiyZHFVMeEYkbdHg2mxsrD+S8C
Gwui/BgdSIqoeDwCMa0Kxgj9y9PUT/x+Z3mLWsVXIj5h+1aj9NBE6nm9kfRILKsosOAGOsfyI8FY
kWP8+cCF/o6Vrxr9LB6E28h9IAbUTRn3dJYaXOjphi5IukGIqLBfECwnPMVwecrJyuPlx2F00Gbc
pICzdOmcyTFnMotLLMNqJeJlfgEmnhBgiwKgsp77SxHCI8LSX0CGuEHwncqY98RRZXGz5J09Y7rS
6FSAKtstJzfpBS9LoKlavwC49rmUFjtT4LlfIRuwJ93wGyrDOYnOMAk+El8LwGtzKxoqnEE50J0N
7+w7PoqJYmSezuL/BAUIlAHKScT0BoUw5pW5Ko/w8F7Mc0MB2CWBD4Rof7LEKBSO4lsg8zQcgXrF
2zvVpkzFf8Mi1mX2qYTS+tX67cVM/3UEBtiqDJ2YtM8gwgxEgAg+Ct0hYQEAVbEauB0aGT4MRirW
yVysk+G2UteI38JWY7lCp3ANyfxPYZYopsUkqIkAH+K4bXH/xRhCsYNnMTws0qBVkfOwNU434IVe
rp2W3DfClBQr1uVUXMYwMJMj4VPROc3H2lLzugRiH0CKKwLMp+aSQrDiAOv54ZcsGjehFZqxmIFo
izKET4caTPTvODAQL8Y9dI4ARbtW5VrBmiMKSL3n+AQ/n0DFW2VMorHqhKOqdlF8HNEgzr3hxYb/
PQ6mnIuAGM80Hje5Bkdahmzm3jsk1y4ba2W0hGjRfT3ynoMiEZPe8oj7j3F8eyBAx6v8Eg6NmJOy
VJx0qr4gLt4A6L4XUQW++OgAfukhudW4PKm9hidl37hgpWtOodMnuNKq1OZLa9kcGCzrYe2RohTO
vR+g9uF8NEVeTamAAezyP8wnxOYTNLGlxmLk/MrWQs83rncSm+ClPXZSMlpRG5J2l/Hi1WEHLmTG
KwRDowQkbRGhwaOYCKC+/tNO/JdKJWLGp6MMW3LQuFHJmOoEZOtzryCmIMcrZvpxdgVhpvyLulls
9vaEO/OXndJUYVMwMdOz3NYogt32bR6DbLsV1CPRMrZEp1QH8JES462tOAPl0mcf4XLjlmsmW+mK
DpctFOFTYfVdWdciRJfHrMQK0JMlPXWO1B++sQSilOBcJ0C/xfIQqDHaagZO/ingA51mqt4yNYgF
sgMQiRap5dvURwV//1z2Y3BqXWdSpEi9R6Q3+QqJsswPVuiBDlQoeAY2a/G54EAEuB/NbPOdPcgS
o6sOkSIASnovWLwVrXwsi/DvM4tSkASMCUU7RoYopi439aDsfKKE2ECM7HMNCR9fh/r90sMLiw1m
cloLhQJ1joSYH4FvF9IlUesNMHLkvSJwaa49H4Cnv/C9PCJ80QWY48w5odHyC7msGo7o7YgRwee9
MCOBQdPrqFq1GNcusioqeAE63zphFtyx1EvxG3b1Ia0oYvZw41vGQKPUH0ACRfXZ/DjKiU/kRUyE
VHa4c1p1YYKVzU8V08p8zQnugE2n0Jrv9VSmiKKM53x/5MTmQWs2noHIboDpcg32EuydJRXCS6d+
XH90CGdYKATEt0cQ4B9EYMxvHyHOiWZmz2QpdzQOL5svEmMYgJhY0ahAOZFaGJ+AMesiMrca7wd0
xzc9xq1gXs7M30hhLNE2wGueJ2rNbJqYfW7BDsZYSptsmy/ytB2yp8m4r7f0c8rI/F2FK9BYm8e1
Iaz/Pqrxiq3xhnGjU6e75hoCcR5cI9mFrg10SYkpn/SsQbvyZ8KqbnK3LNjnel1EJ2mybA4XmWxz
BcvUiEUZWtQukiXRFU/ajhVe2YhKnF1tQ06LGfe1gbEduPZC8oLn4gA6pTNmnIJGA2G/5gFQvzJA
kXrv/x2a7ZN9oLDO6lHY7RuiqzlSYEpCR5k3l6tnrr1VNhyJsGN35qARrpX1ssyaOANVbHAc72Wh
pWXiiKl19/EtgC8bwK+pEYL+XJhZOs4wSEyFKb0MDNfVubAVTxcPBZ1M4q7g//JAVhbDbg4XJ3KB
VXo7idcDgNlGh2tsw3LPDkIQhLaR6ave8lrvNc72XekZnwp2HcH42dIzT/kKcYNZW7wewMMbfRbf
smjQ3M5BwL7n8DYmUXMXRUHrTwvXSw8Il6EMOfPk4jeA3nFl5zPqKrIyY0sbRjbcNLAIK2nC97G0
FMgGvHSQrpzH7L2wugW+K+Az0YL5ZIgHbrOWsjfqyIW5bJbdIV6uKreb7bcsBg4z0Z7HJ6n4VZRW
xH/mdEDo711t08igR6l2eFN/YCX/SGBkqtoe5HGoRDr0d/kuLIh8mAkhFVgB8ewJ1WnVEp3WyKV/
lhpDXfVQ8dXJf+aKvx1EkpOyC8G5XERDpveMf4a6nAQ4UGjdcCA29XnA2vDTehm/qArao5yiUQmY
Z83JHQmnmOceL8L/vUBHLnBCNsJS8w8BkoIePUiqQRo/X6rutuqRkhNJ98sd4a+Ad9BylvQwD/jH
Di9fyAg5FCbcD/kHwhq0m7HPWVzoPonTiufemwbc4g6xcRnU+HqRoC+UpEWT6RMEPrbbsXB1RljU
vT5Eb7uRZyjL/IcqtqhVnAt73DB75BLH0T5li2jshkUsDNC9WwoUHTfAKVR5Wc4gqklKSx0IYKNz
pwKuByPSXS2HQXPM1ploaBhW1cmTjwFnwtcxhtsQq1oXvlvd2pb1jjLGrOgCzzZuIOvXClfHKOSc
EmFtU19cWJPxLtUUor4qAED5iPAaJZRe+PO5KzvuTH5rPs1nFIMjdOj3rmQf8i5XJA8SU+2XA6Ag
4spE4R1pEvBdzFDheGgmRjeajavHZPG1QUJPUrH0FLx16OER77roO8I/p1vlC2k4FlxjAhMJvgjH
0vwu93BtfS9MCRPnSoGWZrWyISea+PqAGSQpypt1fxFo7XC8KyhgsNkorFMC7zXfsAHps3RNtQpW
LBPOHCweGHGR8y5yOJ3aqAIptKBybB23CBmA64L56H3m0ZM8dplBZrrQk+wBY9wqzbhptTA6mqxv
RXirQcDgR4wScUkR7wcf+fG6L0xYiZyLFZIb3Jpq/hetB1wBd5Z8fXUWETgkIn/xh7txbzXQjddI
ycKznup5s/5Ld9yBhUZHT56lDCJFM8s2feyiB2JRwIKa2wJTH59Da5LKOYAWg/Z3kd5UBCqkdwSf
8Qq0xtNOluJ75/PwCkbWeYMDTwZt5XlUDqMW1nocqzGVJvW6ZnkJtqY/ysZGAKZiu6H4E8nebG1e
pHMyGAkdctwvdRVAdZyXh0hZjQltOG32B4QVds0NoV+p0MNjXQoAodIujHQDccIQBHUnOkqkgJ4A
5mTjMZX4f7mX1c7XmorxuVNmRhlQrbekcs71MBk4vHUpC3ALxIGzI/rGlRpcvzSdef3dJTzsqXa0
5apiSL7nf+roJm6c9E3Sd6iRpV5AMNwl0izkaXj4ty/appM+j4vHgO6p1a40aVDJN+HtO43afXc/
8tso1TpsHPBJepzPG8wP8cfxpdWCoWHrdQU6V4UX2Jv0F6whs21t9LOrtCyvMbADbETw252nHYde
2IaIdGQv4qbEEs/rc0digMnq6MMtpk9rI8yAoQFwZ2ZJiHZFRQtKZJsH1uBr64OXN30QZ9PiYLVQ
aXSv3r7W+swuM6CGUeRJ0c3n5N6bnBlEkVzsoeixyikBNnhC6onZ9ljrKFK49KPFKkjGfG+0cN5x
UiSlinjIhYjyie0juWtKmScbJuQEEjizva/etiO3MURhTOvAoDfPoT35NCXAARWln5lvxomUjwsY
bIv64Im6nBf7CMOtooKKyAgVpf89EHn8pvab+nQ5ukVQnjvOQgr5xRljrN1rG5K9RGQB1yP8LueE
CVGfJc5nZn2wMC3zNoiL32z8uXROCoaSx4asZze2xXOf69C5fgAfdHQQ16m3rEs23puu3U1f1HiO
SuYZ9kDCK/PBEN7lRph0ZefQUiixuvz2IeNfSX90j723lVLj+8arUrYRc286K41gWhuSi2Z/7LL3
gqi8eneqXywj5a2tOMORGQVw7CIAbHMHZZcX8Pc3elQW0bLceVhvjSN2A9kvyYxoLs1pM27D74tu
vraZ/7a7E8GHXpNHU7Yx727sHD9SZLvqQ23hj/zpk/Xpgg3f7mW1a6/oATxKV5Gmm6spJoUZLTWC
ntruYVZRyqdIy+QUxG3S0CTV8kQixk6UWYnHBpKVV4zRB6ZsXsEwt7tiEiYC1y+EgZM1mmBLsBoI
ozjNZL+FPy7XbA0Mdj7wHijoRSPUQ+qK5T9eQsiLIF4ZDrqkYbMCe1t/QZwJaSjonGLY4uSz4tD9
uY4TzB7Fult8QS6CrsJ/EUeTvfs9A2pL5oIv9F21B7kHKqx5gZxR/M96t2pMepIBIMq8PRx8u06y
dzl40PBflqLg37mGN50tAou5IBHrVbyAvmWVXiFtJajQO//0+r8/c73ikKZutsTittY/fpQzWlgn
4wMkBOaxXXllGRqBk/ZnCs70Z2Vo7bSneP1awmog/AiRt7YE0GMLiGkL8BWi/TTHUT6OhpiSKuJ3
Ksz4V0DphVY75K46rcW/YcH35lrQH7gQWVmb+fNo2K4AevwB9zeOyOhX7Ay0APbK5H3aL4GIgTYo
M+NK2xTWD+jdj3LjJgGPP5kJiqUfftSmZGDOhnK1iBKvTi0lt6S5fdeRBZPVUPfhSRrzofMNX6nR
dPGepBghvH/vZsd9nsDdtWKEp94mCu5p0tBxExCfonLvtYkyXcefRGzMDRq0wsyoAqs44MPPl6am
bZlaWgC5++5yRYO9uVrf0NZqu5pTLso2KNbzzsm/dHaI3Qx9cy0S8ZGHZT4zXXldRvMxUDeMZRWt
LaBCnRJZOUcu4hFaix3IbtanF81AtCPh4Bm+5RnarizxJzMIrSHQmAU3IVwe70Q=
`protect end_protected




`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
a2ftgqajmSYIzeiBCMjbtSWb2ZukNWEEPjvLnQw/DLFxSgbJC8r5H98uDEQwHqGwJN5xCIO0UExg
LszWFMGeEA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Zq3N1k4JZvjrx7Xu2joAPH3kQDTqSvp3VEDaqxYJ6LqbFUIsEZeCHDtByv+oQ/vSRjQ+7nIhl20J
uvxbz3NSAAvYvmGj3uSgHota4YR+QMGHqT+ZvH4drU0pYI0TRA4LOj6d2oJyIlSZzUs6lWxaWVlD
12TdxBpgumzh0PFkG7c=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UwqwZTIbhKNl9nN+ejl5LH8cGwFMEFaQKrCe78+aTH0JCWqG50xzKWaCFkUPNMfsDtOnXc0yaxTw
xaZI9J15ipTUWfdXCHTZl72EdBBWB4S3j7KoegnpTWYu0Eux/ThKLixN2T+60EvnaZC44cinlxNM
S5l6QEUQWrfpWdQvsBuWY0OH0BC+Rvro8rHLV8bI5OshoWaQfyvU2w52H2GVMmgTBLPAK+0VQ0KP
0EJgr/yqu3rQ6LG2tcxLAYRdLY5AqaHCJoAcK+TIY7JGeaKsQ4Vdn/OUCfmXVV99bF2siFnUg71m
oAY8VvsapYi+AN28yQkG2xT03q+nWjdMPxIhsA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
E2j12MXp+3Av8LyHKSnG87aj12jUIEkfcdq+wkxq0pgrVwZ+/pI2AeUe/Hebq0Ul6YCdUwssIzr0
l94rca6swHlg89p1I1sOyBouluzr0VCNMhljhrM5icWcyYp4ag1iQ9r84ZpgKS1hLq+3wKoEV4A5
StGOTWUyjP5VTR0+0Eo/6DWHxDAXW4DnhexsjuC11T/8rHNbHAjEWKuyy2jQumJgRe5H3MKfZ6rx
VbsmSgcZYco4EM9J+ph5VctCnJZQQjNFuo8I/Hw9qrnyejyctejiwuLVe7HN+yItJdT+mVevYxax
Ydhi3zOgKCaC0IlpfmqWVn5GzfA3D4n1dC4kjQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
P8++xF8rTJF/8YyO18RBPdEMCCxQpz82CetG/Njfi/V3YUvBrMBgGGtFl7MSWv2TD2M7sx0Ylqam
58phLx+xjIPg1qMMBr0l4zunH5RA6BjbW3zN7HBD0b+3hFjaO2ofgadaXe9CjOSz2BsYXKpqoOQ2
+e66gjHUvePkocfpjxWx5jujSqOdzrf4jahvP5Cca+8YZCoJaBmnkBX0SZhbtZTjTWVuOwnobMJ0
oAqsFv1IL14mEn72QTLUKvJL5/1ANHOq0ACKffeChKCfl7e6Z0pH81Ei6uxTM/eUiBjNcamfy9fs
nVzhAFovC7sj/C6/vB70VbA2sijr8WMsGxofUQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jOm0Yj27UmyyaAn3FE4yl6hZCrPKtbvH6qosvQpRyXEkK/d81Hct/erveBPP2H+7z6VgMu8AjV+A
g/N+wQsKeKAck+5SJmTLGvI/g/1+l7ez3kNpJrd8uj7HqCv07rirdzXtdbldLjn4D0vdyRtIS8+Y
9dOCDhMkc5z6wambwSo=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
C0d1SauKtm5LwuU5kPVt2s/uk5XEbvkzs/hABVTkFw+5opCmrARaGMFX4tQJYRW4GJxERkezgJqp
8bDuBjZEVx9euqZNNCxik4MmTMn4YSi41GLCWPWUu436gEYtFUkUA2HmTCx4ebXXvXIcKWtcg3ux
m1ECsrPaNDa00iSpGsbwEYXB0xds/oYJqspnGql0trwOPir7GTvDTcNCIRU/Tw0yVeU4GSdmspb6
hVS1aTnszmXR7QZIbMWSInToOvlMCGtEBTVaT/QXohs+wH+VlHDnwkNV3nrZFjofLFGJbfjqurdk
/qGhwk8vOoRk9bo5SHC0kHc5X3LHtl12BJrPuA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 921440)
`protect data_block
wPtPpPahuelhWBphJfvRG+sNZF7dLZN4kADiWTqgFpBdkdd0LgdMfnAYyj43PVeista6tc2Fyldm
O4LtLM3LqA3KwWu4xAjNIMjAYpmCUEaGqUUj5JfVkk3soqSuLL8Yjbl8JgpjMbqg5IZURvONVh7r
hvdKR358Lt+9YK9cRhp5fqLf4y0jqq+N2L/FH94/UPSbE+rwvyADeDik1XQPbqqAwAxkFgH8tf0S
2e+XPrwNg6dRUpd42GO9Z3EQoJNnxSazT7J6z+wIK5J7cKVDSuwnhrK1ubXoRrtbygmnZhGQX0el
aZvxFoFMTfSro1Ohog0a3lSlPgo2LgD4PKz8tjmZA4PuXK0Vp/p5pMMhKBH3Rj6zS0OqlORNMPBE
hzzEiAJvCPzLuFqhuS0KaEuYybbqGVCNjHTU1VLf+SWqvnM7dVUCJJzIQDBL95A2KmTZHVU7exUr
QtP+Lk6CTRLwHzMY5Ib4W0wsFhOSNaL6uBiIfUjbWIL1qGDPCpnR71GZM7es5KOtZDLqNrM04oPa
ish1rLXpNzMQVXw3gyBObefQBXmJKdMfM57A9Otvf7XLCY2bxO/jPo0AEtUL3GXI19VCrvC3n2KM
QcQDQJEmmRtNSktKgwJ37moKSIDxWwM+vbBtOBYKaWZmX/R+ZETunb37RJEnAMmdVV9ItrvJxh5x
GZn3lm5NqD6EyfYUs7sbiF+U3F1pYzd3SSbNanPT+hBZNsD0Q5FCs4JdosJ6FXMyRILDJcJRm0aA
tZMOEFYo8zsRwjxW/pfanEvPCMgci9G4yzr+rIpvboIT/uIB2c7cqjgN8GvddksvPJ5xBWFa294d
XONqKDMssx2ELfmvcgPpZ0Pv6KNU1adfrJ+USol086evXu4eNOkFkt1wgb0Ab/0pEGXCy7YWjxce
p/cgfoWV+X9H/bwliY1ybmppLQNyn7SXqqkxCCW7ala1CetARxjdcceC3j8jC51KGFWYijFM0jtl
lFwaCQP2RU/CUpDTdrt0MI2nD0xD516GVrtir8pR19X4PMHxudSN8xmVhkWyDME0PTK93AAM19+A
crDcXr+lbArk2vetgKuH+PdBZ2BJzr5cJKmr5PuXs4lxgh2DvIsNJ8Y83IROwTttPsjlqdjpsJAo
WZnoQXNOlSdgkWfh5LM+D+HVEeprx3oOB1wrDhhOcIk8tQM2UuywclNCq+9Gr01txVD2OEsFXwPV
xkYAQ6+9QfH5aMcSyqo0D2OXVzw4A3Hyw6eLdfXGIiZ/8LlWTaauOkbR39AnbijCLwMcdaoumQ68
9BhUS+GaFLPoOYQGZltQR/hd0SbZTHTO1KmBvQgwwq5+Tlewg2Z9bHUw6+yXCPsLJHPPlfeHlK/n
U5cTrqByrh2VecCdSaB/EsyQB5IuEKniGiYj8XaJGfJ2GSkjKaFSiEj6BSTZ15FKEETohy6/2TKr
9sNm9w3ymoKdaGRcpYnjIBWyNw6dIacSo65WMlwvlsso21W+Jlt7g/pAinXtxGuMESXPNEzVKOby
0w+MJkZ1rDeCYUSQh8pt0JTl+T/jwG78PGdqzZEumayyeFZOLFqD2Jj6SgVY0k7ESpmpORr7cnKt
MQBJMbQ3jdcfmAauthxkpw8JAjG2utnpD6aDGaeCj/uBQ1yLvNnZzt75eSg47kzH7PZsCUzaiJh4
6r5ec7XxkH3dbwVyhUcVc0N2/a4ERwVNst/yXAyuJboqifxx98A2RSAyKWc3FqXz8CenZnBvMhMW
Vjuao/5jFkJMcJ307sSX3UK6W9ghgPN5F/2Ns+kkn1srzcfJMq866lhhvBppH/DM19fqEw6ewBUA
OJhM1cCt1EPVkO3wrE/JfVpoir9iAV491YOjcpo336V1ZIFBbUun0l+/lAQqrb3/BGEUHO3YzvGD
HzO13wxSYjw8P6o12/5YVArRPxGaobjFEu/P/+Mj0LgweEM+szAeGewTeDJeVWUc0Mw+WA5ZreDq
RXXpXWeUD16QBuvGx8nz67oPHjuE7rsbPSH67oNvD7eVEHkBrM9hp29cQkAwOIcGIgkjUxOXpHXi
hR+6zDLbHA0JGo1sd5fLvuCKi/NGO+aI9Ep4t+rrrsRYla9j0TV/2Y5a7TWMcj99GL8LMPNrRZtR
x5ZVLiV5Kh48sVy20tquMvaaTxhfAbjmhCgIk80sAghF4mcVhqH5r1rJVBH33XeN943v3uim3CUp
5LXwkwFeB3kQyUGs2QXhQTd1t6H6cutYmH7IbmzOIctJaYVZSmsqSwiCVY49Ocmnm0Fs/pRMbdTF
fM7+s/35O0Smrvv6yPY+An1BTPeKs9zNLvFc89eXSR29R7Buw7rJwGWLfirEUy7G/hvwCttUD82h
ElG2LRpUCj54ka1NpbM+4GvEH13Vay/RyB3IsKHgs9nghb2THn3rtDx+TYUVXPnA8BHs7qM5FT6q
5IB7eTLxqSZdDn8Hi/V/2oFQjeMUmXEJP8HfkF8UO5Tso9B8K0rWNyTxPlqg31zZhLGDpp6nrBhe
ANTdvHb2fhaYabkFRyiW8kkXV/bPebUPtmqsCxJ8tAPm80VgFvHvA53dpN+yO4UkhjFi7yJQ2cqj
sFFB+b3SVi/TvlvRdjl5IwuYo1t3mWD6LmMIXkZ3vNuwTGWqPph2tU+nHnN1BeuJMHdkjFh8Sv2x
XnUh9UF3cWb3q0jFNaFgHuPxSYsyjgQCeN8SeiYDZST6mAkNa35fV8Ofc0R+9NQRa6j5r4vGAB26
FOAXgxd0NM1ZV2WLL+IDN76KX74sDw4nQmXuSoCRpwl5uMf4AlnHByIdWogseL9WZRB38L1GoHnA
LuqIivAkWbPGVkxNjLolM6wfsPm0/bFe+AnSHiuawfWFfz8g2KFOipCFvoozaW/Pb7Il/v22YFQp
Vpbib40D1C2rGRighlHIcgQ/s2dxUkX2hepZwBxdUOuvy4JqpnfQc9/WIOCv6TNjPeNzDAEM1eZq
niKkaF3RUNHen03i2Ti6PM/5H0WkoB2TyeX/WOpGNucY/QWofNCG+Yl2oaH4QbZeATYAov6e5DPF
FY5LCvG1axiNJiwUC4ipvKj5krUeELQUeBxTH+0hXH6omzXHXqwMmy4+ZTRzYxjs05gOX+J0xTrZ
djKI9TW4Uj8iffHzJ4gMdnz+Pyxxk12rKFUMGFlP/R0DNYViGpyLZ5JPHQbLlqjkpuTmIOASQ7jQ
l00ra1IdFg2s+wzG9YwXigdsWfY7CuyYAwiWX2FGqVWjatnCQ9PfD9JZZZ+ZfkU6d0QJftoryL+r
sDV1uHdgqcd1xX3l8OGx+xKLoKMgDj2b+EECmdETtYmZCOEiuz8GC20kyK0lmil5bMGQIFuVoo6i
VfOUMbUtRtYGOYd4Wf7Jh1NJwvKXobueo0HRUTydorTkDqBeJBVsR7zsgoLYWAOVzXlO7azun13C
zyLbUnWAS/MrcyC8CncyS6S/n5DCZNrJdeHwfE7TQ4TtUzCktljbD1y9Tdm2cQ8r5LjVRWwlzSH6
nRYF/9uAl6dJ4SdLESBnyp8c5hAizi05m0tin4hnJ7+cwOPrk00NcbK6MWzpUaLgDj1Xn/Z7sxxH
6F7INgYZB9fAUVhpsaA6Z6hZOUq5gT++Sh6VU5Pzwo3PH7xiWhLfZ4Xkd4R3wN/h8q0as0VzcsY3
zGubMYx8PNpR3HakSBSu+kSv4kYIuWD2iAoSkDAldO4X31dyyMwc+1sh1etqYDDdgmAKCDciBjnf
40XEmmcI6OJPAqcx1H1mAkVW/PaGLl7wYfRSbPvRGDrvjSj9IPr3XV2ctKQkCnSU02QXuIOlMU7j
7g7NS3OAb5Io/1gzp4qmHZM8ByhdQM4c+NkJqSmz+a/Tss5OxzUIANb3Z0ji8lFeRP0Hnr/i5Ev1
j6mZkAlycyLV9TdK9Z9Mslr/mP9VKvkNmW8gGEmec7d3RMgRp/AVgll8X69vV3wUvMCJt+xFwYBf
h1qKGGhd3AZszgFs3xmt1+WzmVgSTP6zh7BGuYUrwzAbYsaO4a6NtjiycHzzQlBXon/sWb1Tyb4/
vVuCogUiT3eIglK34WtLVZwBnwhftJvcSYVN9VLt1vcdqhZTnaqYGU6G0hGOGSd1yS7HRaACHr1U
UZDzKtf2RLD0FvP97AretqLt+85pIml/gHbGwsZ5ACcimvFBfNZavUuxon67718u8gMNyXJj/uMy
GGG+GulhS2AqLALpIvL7dyeAfz3XjMzUmIcB/6P94J+JcQHIZZJhTtb5O2+GBbQVQPfO3W3bBmZN
/Pdrwa/PEezdOvWjqpCmZX/njJN+dz7KUyT+g8cZeblzcYHD9GZwrhBcgbo6xT4Mu2fYZZPefkTa
1+pTIvoXpJpBmM2ds7W1mesv0jyfJOwyddlx6wxTGu6x16qhZkHzRqry9J5xLs3408ExoP/+8JVR
rtoLicOGcw4ElRjdOssf+FGt3QB55IdF1Be/PXVAenfkTs0GnU6Gd1xsoxzIqtU0qFc7wIQxkzfN
hFUTu47Q64mVCKdDx9ch8tBnfj5U/mYwbeczdZ2hBFLx2GgIZMToFceBEZNtbtlVDmiCkTuqAnsM
jENI/eH0HmfE1x4XfjQVOBbZ2iwK8ws6ALUq0ZJ4LAgxWUqMelIMKa+/mcINRN9+oFLL4nI/PYmq
Rrz/TzDslRkPUgLDJ4EBs3ITKkrTaUmFaah/aN0fpesJcVXDUytHk0Gxz+gKAwyqxNSmjYPKRrRw
IEWLAOJLxoDX9jkiUWuIZE+xlisenAw6xnCXWSdSpxCoIEvwHG4b011D5ZQNwHisEB0DDStcN6Qd
VreM+pvMkaP2cywHC94NrbQmPX0fb5bUUEuUmnr60+yHix4SnSqWmdQkXWOoi2gYRNHDE45kb49t
Er5VwY0foMPcqDQ/hcLN75T2wbFlAlgmAfeBbXGvBXP6fdkfcNQdbDUAWBlCHJmDbO7NcDLty1Y2
S/bCCioFeyNJM4LsPiXrew8/eWL6olzcjvZad8GN8EFvCCgJV8h2yZnS146OPjZg6cxFy5fFCmhi
pkyFBYSu+V6H3b9XduF5xsc71Uo9TzxOFr9mCk52c63v7GPkKleQkp4KlHE/qJokXJWEq82RMd7z
AdquJRaJVs3SJmRYssI2iO23Hgm+XJMHCl0Kk+SJ30iOG28OI0y228EGcTUYo948V78T1WoAAZs8
V9cm9pC/88DMYokHptOekxMNlaMJLJcuIbET8LXkCzZQ8t+oXbI//BSp1aK2QjCnBPw0LU8sPSDC
UG8KHEdA5EZVY2jbnlqtywWih51Mkrnxc67KUqLNw4e25NIkreTBbiONMo9T9d5GTMlPh9p7Bm4e
wUcVeyjcOFf5n6wHyBCOgxAAgzWzF2q8FqAeFq+4c/tiRt+ySmJA4U2dUh5DHkxEtNU5+DbPO7Ot
/IXyzZhUC8kHkECB0+Sf9wVv59GLX8/3vQvjHLYG025ERsEELjdFfibGJWfzbEgFhvF7ke7nZ9gU
bx0YTo+yXBDSsNZCWuyTF+acrTaQxf+ZszV4D6fMJYnQROFX/prlcxHHBU538S/kWejNTLgiXX4q
ZJmSwJK88MLHFHtg+RZglSJnJdbMQ376CeHMo+i5rvDUWDwWDgeXrqcEcGyXP1PoS5vWI3YR2T1Y
xcqGQZV1Mw0eaWxW7jkA8TnLOeBtdswuyUOTbm43MaFnoXiTephTJ3Pn6FHdyCNwbrVuJrAa9gsC
OArTHZDFRyuijVEhfIsLFfB3oPXS5al+YUBqY4Ou61mrk2lOPBcG8HmS3F/yUp+li3Kh+q9z30lC
+kQzGOvDmOYxurjREZANF+eojNmnyQr7zGWsEu4rCBVZzSgloAv+TLrXc5FBEUfjwgD7M4/WLQw5
5rSfR8Hmg58xGdcmyJ3eXkYlpzuU22n1p7eRlcNl4RkAGab5SPbtVYcNECFUpAZsHhQevPyM/N+B
N/u7OloTmmbDoGnSHJmlaQT7f7urgQCspZ8X7m+6LZGnb5vWcK/2lXFj0mLkwziPODZnqKjB9RVf
Q7cEEUjlz5laD9V7wG9CbxFq0tkEofwEFvqBCYzaK1VX6kIVKZreBQqHx3iszwCOD8kcrtICoWC0
ARvDmpW4Shc4VGU0p93Zoxh9W/LdG9Zq+997WHMh+oUnuYv374GhaXM4UeWnQ60ZEJbBGky0odM/
F6LG9YhOnge8auJ/zeKZCgT24Yaeadyt+xTu6rxaEOcDvGPnWU3SBTPQ79LmH13o4jE6s4ZlSj/3
Zpya9PCfHmAcu8ZUNyU+vwOc1karGLMqAnVDZEVvKEgBFx/9JhPnN7qXhxbLdVGcMsqMIKVexk8m
rWuWgugxpx1jdAmA+Yys7bHFwqJRZeFe9Efj8dmyl5uGUIIm8mNrX7QPpvnhjMuStLfzdb2IwWDu
Kb1/kD2HjvpKTDKgEJI+lGjABVr/guXn50nLTWMkXh+/PgMSKeeMfuyCkFJtO4UbQKYYTzSYp+L5
plSf6QYu/fv2y5IYgFhaqDM/UvG26y8UpD+t99qVUnmmOGcrPNge6RKnp/y5IqWLC6zzp1UKViEl
7ONs66vFjoqA7B5bAcVcOUAirFFfBphfMWmpcV7S2IpJEvvpz50uURnFri/B+SHBfUvgFe3JNMjK
Uia5BopjkSJtS4J3raIWMRwtNw54NdKF7zJ0ptkVRBxteIQ+fxyKVqSprX+B80bFKZens4/iniFS
9Otj6Yos3nlrodF9F6cq0BQVQsDGXyZdgkRejYKdvHqD9Lw2FG7XqXI7+3aKWj3oM5HpU5jiCu8h
uryKo4Xx5g/qspxabGV9oGb5VCJkw5Ol4yohkQtKCenUCwlLlcs1R22o6Do5t96znXPD0kPV1SYi
AGbqgJ0cFDR+mEaB8B3hervnouZLmE9rxmab1t7/uWSqRm2l7Bn8YVH+u5LaQ7Uw9CfwHHjajHcA
GmitBW1qwaWpvrlqbXQHRnZJMGjhxYULH2SOeRNIRphuTXbKzxL9eDB93RArnMlPrfT18UNRyzfX
lh9CjiBepqkM0TvRQlFWYp+03licv39U50cZjs9Fef3Wjb1e+0WnRM1ATQbYMMVSCY4RO7g5JpqH
YnexzalgaL6HGk7URRZUz4hUQFhfgQPgOQnEmYblh1Otoa1N13TOxLYeazohwUpMqiZfOj3XbK/l
FuIkoeSfn0fPN4X4U+kRnlrpyka3AP6A1mai9M7gr6APF0pp5pTm31S+Qzzrc5rZVJ1h+toeEjAr
QHpRfSt97P/8Duk25zXvprXnN9d16WnSH7eOFFitluUIE8ZpcGdQsjcFaUL9AOqMcUZUrE6/YNbu
71byO/8LBY1loXlbLKaXD1QnBHgpFrOk03fQ4i0uG88DuGAJyxgYhozjE7xdEEIvP7SkZJoNT39D
wPFTPavU6BwY1t4+V8PQA08L+fJpGGJcop4s7tr78iMm6JY+JLT6h2HOQCOzk950VUvXn3ykeKHi
PRklf8jOdR2h8pB/RriiQz7o0BpJFwfnMIZHCm2g2I5dr2UZw8jZuORJWk2zxpu8CaLm+C5Ylo+f
xZeFtKctSvKVQ1VqdU3KTd0FLAPs3wLa8cMdSf1UUDruCRALuCpdxbaFSSJeYdH0UUA+q+qxIX5O
zD+avy+9Qf70FiwQskJvhUpx9pGULl9QU1VJn8yNXbk8QvoFN8PyuTARlonmhlVuuP2NmEt79rGG
7TT7+LoeizIOV3JB0KuDqfNJ8XM4wkJCwdGyOeLNsc6n5jiPuTGagRRgdP3mAqqqz3dP/hlbMWgc
YxqLXrABrPdn1RyGPd2QNFWlRw8GDjvza0lccr/lBjfgaMQYsBMrhMCi3aUAu/VvsuUj/Bi1sRQI
Txc+/aZhJKb5XPAMHHZGe8riW/CBq2okeGsktYvE/ve6ZfhiJHF444+VbcPchhe2cnL1xmk/eWIR
PNvhPT1uvxhAYjJUuRbWTtuOHS99ksWR/fG/2DfKvCCPua1HETqkMXVkLizhRa+bJ1hStq7kNAQz
DzrTZ30/Kr9Ft0WQ7PrxNXaStNi3+cp+WQ1sinexjSP/XTFlL2PH5CdmE7TDbT5Bu/Pv7LztQPRf
7cvAJ/QtEPRT226qQkD1yN1FsbE1CIVTKc+hI2EZzneQId4UriqOkxxyNe5IcMlp7OKkA6nCee1R
SYe5PukwcwAEX6Mi2Tc23bVWOs/j5/dITMro8JMYtzD1f8a5dBCome2FD9wXQdKzCvLCAm8XIY7Z
9M8VnN3oLXt0hXgvl7PwHzHz2jWOGrTwawfbM7xN25p65HeqjouaP4kVPjpB8HiMdTtjZqbdyUAu
igzGNBKAnaFSRDbOR3VUpep3Gruo25RsQbBypIK7CcpkMDnzRb1a5XagRBPLaPPyZPUCsLElsZ+R
UIecLJrcCwH/gt2SUKI+D0W0+f5ybeEcA9Dlgyro19XFrbjGTr6N6HvPC8j7X+sWqSQGER7GGol3
X0NL7tgjWO8nceh0OYhRNH0I+PLPD9o5zHLeo13xcnl/Yz9COdwyRSyF5zDF2u9tafAD1PuSGYqZ
0h+rL59f5wSTg3CLiRwnEMSCk33VzWRnFn/Yq5fUcwBQFdc9anfM0a6NI39e4BaPbzftLBJsLH/n
plwTFAX/8g766t+k2RwVuWqNgZ8+EVq3iNHZNaZHuI3ex0lXQVROtevlioiNjUKoUTCH09ba23C0
hVH1uChGQAD1l5ufXrrWXEF4PHji+qr8SIPRXQAxBSLDdEg6NfYw+wSuSQHrVL9sgDreZTJnt+xk
y4eTa8A0CRmUzgi7k/RaPs6JXQQmeBdVod02Z5VyWLdCN+cUEOIlSj+2GvrkBBVP6qkFd/aGjrep
TCVOZpXnxtXuFEhr5MYT1LI2WQYjoIVjhNQOPjjuyH1w9grk4MVbLVNCOnO8W78FFkCgQhqZRD2E
TW+jQJuTxvZ8diKbNk4FiCQuP1BsFfmw3Tj4DLlynzRrJPK2DulAhQFAakNvJaaI5cERGvAkEhXq
orlvkthqgUs+cf+lUObBs5wKcNvgsBYdW5rtrWSGAuew5JqEZaG+W0XjKgltG1X3XuIjBspTaFOB
DK0B7bj3I0C0b2ioWH/E6ky2mFg0vtaWYPJ2ZNvGS3nqfjqwEAvAnuOtWFDSxW2T5wQxSuV30BEE
8Be6mg90p4COfCuXcJZT19CQVu7JRXwST21GAstRb/AN8OWbqPwlAn17H0LMD7SAh/EKBG+jUrG6
u5mvZm8JjDOBhpWuUag3D7PjdCMSdNKaVnO38TXlQ72VQH5OFyMNTw1jFKRbQ3uxBQIfMNo5IBOX
gzvfmpdwasihlHUtwYQv6SGIPolvtKZupUGgfHRF0kDnW9aTEdfa0vz9aP5RqcX0fMg6PLpWRjWl
yqD7TexgUVMVqsKDUd5iFMSmfX5YlSQi4NvTN5GY6nu4CLTpWHo8PUcIXQZEoBIGoBEUU2mERXom
A+1oyQayp7MUYXED+j8ACjduIWTdDw2f9hFIWh4UTBkjUVuenqM27JNiUJ5TQklvKRmH/KX4438i
Bwy4K9FT0LQo1fb1W5kzNbZVhFFhXD+4Go8XhIFQQkCOrZzxmAeDbZtbQcwK6har39rHpob+mY0n
c1f+BoCIBz0UZrpnwb/bweNnX4vXG5glf08gzYVnmtG7CIwkGm0mWkPM6wngEf/++gL54n8+0Ld0
6scjhwofocE7UzvggpTeabtsgfLQ6KEeRbPfJx2/AYk5kI4Lc0VjL12oSh7P9+pyBicdQ7hOVy5a
SdHER06k0R/gXT6znBWJ5/WEJ5GN81BW36ZIzUtohV0izzN5xg+47XiKNuZuIbA8oBEqG8b2oE5Z
5NfojYMVXM1/UJb9jw7VPACSkxO35ecWYncgAa+lNUiLp4RbfimW9zY3Z74tkjnkv0oNzjekTLub
9Naj+zN5GRTzaOA4bRGyrctsrD5YZKDfF0A6VyM+kiG3jnmdeUOMOj6alZiCeohHFL0sLivv2Eow
tJqsBt4MZWm3/TnBcF3P1hbJ4YnoDbd+OgJl5gBSYKXV4cYUMAHsGHpv4rY90AVZtzs1LIpHmoIr
ayMePkQELxTKwUXwIfrQ9SdH1CQFq2SZMjEwiup6Kf1WROgxKRHKbu25yF8blORw1VXoTzBJadwC
5hypCxwMx37uxWFjkH263Wo+3IwIeTEW7HS6tnVIK51lgOlNsBrU9adAnvmh+AZKBepB0+nC+7UG
FdzYa/np4KVMAKlixA7ZDH11229KB+McBxYl9aBGKwsHZVX1UF/pqb0030wZzV3F6k3UgLxt2IDj
tXEM9uPv88n6mWZc+krs0h0jc2ymAw9eMmHVwZceN0VtcFmZsbVWETKJgyJb/ZehOuwf0ASa/ohA
JB711MyVIzzhMfaskfFMecaqNYpkpcx3LubYan1LG3s3fb5cvHwkk+vchWmZf8vC/B8l3T7PcLQq
G+GprNv6iw095fWW1Hi7y32XKZyNSDysJjrMg5epUhbF+o85SQx96g3eGJ4kBgZ0XzfenW74YY5N
3dnM613rPoKZBIKFRbuDhhFAuKRTC12YQQJt0nndn4ZxSBrOx7sJjuChUUQCMK3zt80vSgfUQKxj
uofomM2cd1uwqD7m+1J7bJbw+CoJkTx0ag7sfYrBjoH6H6HRceE0bAvuZ39AUv/jkgZS2AiJbMmY
WzzVeffmom5rq1bU35Zm60Q/RmE4myrjGVyow68AOnNWmmZy4nr6u4BcdiJmRGuesPkLRAAjyV92
Jlx/zQjRQf49T1YEsXoICwVC5GOUw46l4HZe5vmmjm7EvLhNjoGs9EuG1MucsInzkQe5WTTxlkOv
NVs4ZOVZzkzpk17QeLMEa+sgSbLuyQp4aG3WuoI3/i5c6qas7XQRX18gOPBB2BRm5Pl6jBTnPVde
L/YqV1sk97KvDIcnlRu13Dr6f0CLz20WbcJYvZGJyj7PJJtfDNJTW45UU5Vmu7nqhpRW4seyEsSj
Uc380J9WhW+WBUHh6wj0MklXCpwx/d+6tVwQ3F3DjG5xF4LvHZtPSFrRwXWu2HgsW4hghCDMiw7O
sG077e14DF8O0eegyJ3PHF9Zbd+wjmIqKuBgXD27tylnOIz4s+gqS8HFyKP2Nn8J5ktT68pjDp3A
CqHpDzpyrWG0UGj/8fzpeZfgRS7xdWSDzTA28y23gbo5dFeHlj3Ve8kv7evLQ9ELbBOiwzBw+Ooz
gAwie6dXiQirxNIamMEwy6Q+wNVnXotU8iuXeu46tXVuQ2ZQ/tkb9SuQKOdOD7JLgpgZOoxe+Bqs
/gPX3sACjdGLlM8zoEMhglbf1psL1Po8THqxjz78ytbrExPXXr20U2kdvJ5Ym/VCcmVOyWLLcRKl
s2/6ttKBK8Ste0bw5FAR2TTJGEpGEbeLPN1z1YLgps4+NErbN5Ny3nkBdhF1PjPlRLkwg5BnvwJw
2MExxaCluw8PIjdEzuU47ojCeXNEPZgqWNCOmPM2d+RkXEReJSCf8sBoJKtKL0kA06sNzDqp5JJ/
OWxPkEKVIeqESiw/N26zovr6yPtycKx17auQBunixT7ltnjM1+1i5thm0WRmznhYkP7Eqvv3IvoD
0VfL52ZyoDaS9WE3Spfy9CMg3xuocph5gwjTx3FrJOyjRPAm2DYrCjonq9yviaJdUPX19ljpB8Wp
5+/hEoFIsK3xsmWg0XVR314ndHYd35QNK/pTbmdWEPtYPiRzcxjPUp3tlLHk3jVQW+5Z7tnADHNp
IhX0jRg7uSQiHKB88C+JGz9App7NqDDRPzQuIcydg9qaTc+Eg3qA+8lBbdVivpeXkt72UP5sRsg7
P8etszx3Ec0EyisrQIU2KR2Vv83fsRZOvuYy5ljdJNNmGo22xY6KMGRuAw37oeXJHc9XRjJmUBJY
2P4PssQksEW+a3CmgrjlLqwjcqN/EWDZE6jfamDC3G6ORohx0pCPJaV2A/41KcoOrrCjGGvdtUJe
U14UT3IS4KuiKEFm5g6NErP2S0fxslOdS9ZedM83vohDe2aOUZCGv47jT0VskNDg2fYCIPNMkZNF
IKbN/87chpjyFjj/rmOi91Y5fXHjk7+Cpar0m6e+TUHCzV4upbtIvfN57RWkWrUu5eqxeLEg7Y4p
7GfJhC3FZPWr7VgCEenIZU4jrQ5+7jH+tmywg0L/NrgR8zOEtlC1NWDeQRwtG68+Rr0BGjbVKpOi
fa85sPnZ9GhUNMlwh2Tw6RqBO+Alp9XNQZ2X/UXkOBq3h1aQABxF52EAIxeVb4dfoXsXrr4kQs5A
1JDeIKQZW2N65sP/ku1HqbXMQtoz5v+38HX3fO1AMWvQoC4H2MlTdTqEloCn+Dop9i9lmUkXKTtr
ovZoHhfCQ7WYfg62TTj4xhn8bDMXa3+41zOYubGUiMfgUxNK3lfUds+NAN0OsIF4fOcXAy9kGlvR
LrMVqvKG3g4Yj2B9o3OlC09cGbT+wWw7Et9jEchUb4VTrM0HJqlKZM/9/0h16tMHV2nofpuEw8N5
l9Xli0I/GLUNE0xC3uuz35AtenAwjKHULUKCof/OEvGZiZDi/I0kpFUKtaZcgIX1p9KzwrdNrv8b
V6fWPasLVZ+2U6IZfBfixwAfURroyl/ABHVqIinP3CdOqtTrByhUidi4n+Pg2zjjo0UxrAJHaAvv
L9X6sAkXankPorwTfDbUdfLizSOoAoC+8XENepV+lDdLPOr90zOWDMOcYcI8XpY9zIJ6SQkhagY9
uPzATmyXziLfRQuiJ1boH95LhFk7qZoFts/s/znDmwh8SniDL0Hmqi1/B2jCXYEYFx9kojA5gZuT
jesAS6jZy7TQnpyDOxbysetv+VUxy0H3JPxe/uaXPBdHiMRj70cqDYOicnhTXs8oJ0pAE+p+i44Q
7kp4s/rfjg6Vy3U1BfHExpnUnTW01ztslVhniBFlbAzwnXbyUtvuSNjLyYREPbDk2I03Zo2GFFGe
rnIcyTv1l3SeRMWdjgrkpsHCBN8LvM7kfrwxi//JkJ4nY5yAOuhRwBx4rdIhtqhXYgqMpicVQ6nO
5fg6EXXMK7cLPlH9R8gQxZN4FRcWzq0NaHZQBZwTgwVhGFjttbMGFkOwGklYLOO/HivVYgiC4cm9
qPHv7gsTP+hDXRLFbVo+rd10+Q//LesrO9mw1OfUd8pT7ws+Ru3/mzotP4jpgpTXI7rVCb8Qyp4f
capzFuHRZGrUx2cpo3fXfulTNZrcMWT+Dtvn4LA4dy7axHqLXCW6LP3c5nMBrYtYx82QrB87vaRQ
OPwEazRBRrbFS0cAafLzKeH+Psrl+fTEkaUDB+F6pwXsygYQpYZlWxAWrpmIjidzIPmVTFfcCm2Z
+vQd8jgs8K4pWS55gzjn5+lSH+HIT4HLeMs7quU+BirQmQsZ2wcZwAP2g6kFtmtjjqZrPWbLZdgb
S65TMqfj7iKxNnhmzB9UUPwm3+0kjqhX4gHpwpFkVhDfe8Lw7TM0K1sHLFRir27rP14j0VrGesgA
g6F4nuMnrTpEvP0U5ZOlUW8pSdEVqfyhrwzVHhLuD/GTglPFld8XCxQuRNKseT/wslGOlSTDG+CB
w+Lu9BnXOgaU2qHsk33+0bch0pYkj9EfatRAD4Y+NQ/e99CM+gCaJ2G+nJxrShqzWkO+59gqu197
+EmwdtMERmtHaNcv+G/uKvezMVU5KAnnpBAUPMVtBQR/X6g87D90hQFMMUKmqPo9fCo1Qq3K6XOB
7Qj02GlJqGJsGmxtb7RfboMAxe/n2hRjR8WqyZ+flBXS+BSrdXJGoV/xNe9Wgzu65Z7dCoYXWz8W
OlpNKHJ3ha0oI5rtk7EVpw/0S14UpQA6gUso6VjPIN8pOlAE0yiviTI5HpT5CChkLTtqNMBZB6IL
+gaLICAnlDryOYdMyj5/EakxELwdNtrSQRIV9zouq7+KX8v0SRAZK5tyGlAKe4gAIGBAoMX0VKkI
Aub8DfQ6FEtbyR5g40o2mjsQoUFHKSUV6o3rcwllgueOZ2C12xQeHWUIM8EkHO213COZvRX6wXz2
VvuQGdaU28XmD0PW+t5nH7hjmOrQ+oK98IaSfKmKe9tCUSCl9gc5CU5cxwQzIIi4FiuKu7z5lYb8
PTWxLuPyPDOkgjgscu40vyYKaL+KHy7Re9o+i3UI79uO6cf1fbkyk5G1JLvM8ScYVwmy0DSUXttk
wWBrAZcOSysZo5QfuQUVEYbwvM9sXYuy8FvCgshs8K5TxgYsekyB2ZjOLRSt3mrVgoJD12X2KOC9
nt3HsmHYRwVf6oSEA9KkzTMnfRocpXZjfGCqPncJjD4XQnCAzcbq+q0xQmMl2CPaLzMEP2Gz24nm
eeadA+iyJgdnHpL4QvQbCsV6Rl1xu3T5gpY2xZim1uBvDHXHQ9f7+QhoL2DzYg3NjhLVD6R2flSU
Ld2qb4BAjMuGFpagLl27Bo8tkkycNcpg0plYQUhTwb8aWuEYZ0lYwC72ACvRqFGdxQHAHPMeCXYj
aJYUZVapkNu2ekuwDcU5iIsVYcA1smecMIoAue8x8ehkviyUkIeFJntyh0DNEKeKaYI5meqkYHsp
CNnK5iwKte9oXU2gHOuIdgr9FKj8ovf147qXpOTo6zgzn0GEYNOhPt3gJrSX4+Ym4rAzK/M2IsP3
UVEekuzZYKRbcOCf4guHhgXBnca2pLsEPbQJ8cvf4DDWA7ytMOO5IfQ9+BeOmqGBUjsK9z3/Pldh
O95hC/lrLHEcueb7Km1IjxjoqdiLPSMOYMb8RSsvRccZ/xQ3kJrk5A/Bz7luBvd2bh5x09PGPO5P
iL34iuwnHAFj3ktiXYBnRwJ5+oqDkSsPFtcAZEaXuNHWI6m646xzbOUGNPMXgfcmCeCQg1lwiJqW
0GqoTZc0/ibyCPnLKDaYXzR72yxmRarkVf2xrx2We02qo7HJSaJiFLg/zOHKqmivqY+LKh39iiqQ
ezJYbNFXDD4qDLijFLARX8t0By8uz34yyGSz+YBTgycs/Py4Rx7v8d9JrY5DRIlUkKM4TLvWeyD5
XnEbA2Yl434M+SGg4Qz8PSGQdKm/N4aoxEE9OOnq0t6VUwOntv8pzXwwWSowEc8539Z+31aPSDsp
fGlyksrovpZB/XGqy0LN/YST5bILPngsB1bmSwmoIh5RCgiLUCv772vVJfnV/Zqqu4HA6kRf6cp6
tXNwrYcORuf2ZXARjn3pYpdsmruHF9SpnoJNhjlA3JOMU+zR46R3b22bSX0UZrv5P3/NXGyRh6IK
cHeWvyzkQghrkkDNEgXl0w266yKb9uL19cmfNtx/r/gR/yrMFt341APpFqK4HSmv9zIqSicJZ525
E7xpBedBsgTsUk7IS67x2tmlN1H8rwDchSbMtpvidMWUzZ2mKKHxyGJdiNC955SiV9luy3548DC1
LSkXllK2pYddELuyCrvStqNbp0yfV2HZdWPmEXf3eS9frwVoSTdosZcRJB5uRp/giDf6CKtbQyBW
sJYEVBDCETjUjqY1ZuOxGIZlZAsiGfCK7GWM51kOyePfG1cuA1MIaeAfo2FG+CYrIW1mjbvybWds
gkIMuC8qm78fWgjBIhNqoojMGWgy90hMn0DcALaytQnu7b84N/wKgWGAl0oaNqCsaQ9hTaL74G/8
rkEtZdhcFUvzfWS5LcM0MwGiQPmPNhhoLfkMW1aYqH8c+9fv4fynJLW8JIThzYms2taMLjbZXutY
Jdz11RLe/LsVgc43URttKrCd2KIDcuQkWWIv7MTPAwz7Tguw52UnLZFSbQMNZc+m1aO2zOBrr4LZ
39be6uZqcBteWi5tOwhe4y2Zcj/UXmlNfAuSq/hCF0a4DkjVESZSTuurWamS8Z13HVyEkna0tXCL
iASJYLeK7gEhj6Oc4JMKZRooAJga9GgfmyY21He/S7XSBGC9lJRafA3JHvxqe8ViOK4NbC14+x3M
FgueJ5G0dHnOBlMfb+lDe9y0QMie66EbmqPDGr+KZPY04RTiv7jZ0pE4/Dxjhbs9+JFxW7wckEXW
ifRFddO2PGY6U3Iihd/0SknPsi8gWCmgbrLMxvpYjNy42MiSlIAdaaURhIR+ZUSHNtymcADhxxhF
aTedp5d6DzyJQ1jbGFBxEGI8w80mNa73hWD0sSCZLHxrh35Dog8wpq/0+OSyLYmEMdV3bZb/wHNN
uj02Q/Mv2DRc04uBbEzFHPAo6FJToDY2snFF/5fT/7bCPzrMog0GHS7lP8xx534ip4G+ovKxrhRl
XXBgS8nQNH7TbxJ0PuYrT2k7SP+97owtKGnpRpiPxroWAs7Cmwl6hfpaKiqOYeu/mabDwZhGmrWd
XLIjcPXwrRNoiyahkxOnCi9mrGJRKXzRrUBfz1XiTelMK/CjlC6hjd9eb1llBfBVrnzcSI37qwqg
Ej0im/ti5bdrxszcsPsyHG4Mkdq3qzjRG2rL9MfEmmikpSrlfxFbNORs10CMI+LEifNb9RSCPtsA
rjRLVSJotnQCYBjmOzn5EVkdxxQKuLJv2yOn4a5vQAPEswEE9zBxmIscHO3vwwsVENukTWdObZUJ
uQlUdSSCHJVOn1ivybCtMm243VIrSRmHxk8ZO5L/0HzbD4MdduisumsgxPYNP72FiEmlEairnyFg
vXxK7gKxk/16/FrP84nZ/byQuSxk5XTe2QPRGP3+1YIHJ/kqQ/ucgt9GPdt65JHnLwvUb0+nDxo9
wFYZi/3K8iygaylYG8G+LKoFhrVCI16Iuk5Tkm8DQ1AyBEgkNy2TmUknPz4BnCVvIx74xzh2vwsi
tYooMYSopZShttYYTGEKgL6WzPAzK2/F6aq7RfXtpCGPGbcilrafsxy+IYABWbHlzllKCfOUVmXs
ok7PFn1HjHX7ixIyIed9rV1/5P0MEKnZdlLV3MJcaRFBqkakRXi3IOIEjyb8dY7hpfTgynmkZFjW
hojA8LdJ7rkWm8ma28HFBvUm+Iw0801xUQO5IIUsUvwyUpW2iiwyz52SOmWlL3NqqnQxBnuRBJ3S
rUuMwjvUNx+i0pzJ8L9NymhDN06DqJuQjC3DlmmnD7ELkxVwxE6ILwqMcKg6d46H2UAw4DZSEk7G
R+O+zsS20wsFSKH9gnpEdJ/neidQkzH2bxmMgkLqBhbz6KN1Vo4H8G2iLrQwD2ZoxmwqljsvnRON
T8fcdBwZsjeQJ0qhUyV4a+B8yzqjaIFC2THjpVnD2zu5vfV689OySmoqRljEZORN2B+4wBfzcqvL
YP//v5b0ioCvwySw2M+QIttWQ64yCQbNddAyv1lFV3pq1DnU90PmslgsQ60PKKjWImESeMo15IOv
zNofmBQCJzj9JdepQ9BSn65R3sD8/H97b9nvbniCawwYhQH62j+DX48RYfyNe+NbMOSHQYiLCDc6
3WZDgE52aXCyLPSDA+3Sku68KLhlWr+eAkYrEaNl/MY8R1l1puE7RZJNr9JYBDwodThKBQqxVP9p
pR/nBKSWampl83GXO1kr1WJgeMH/VpDcxfVGE4gHN6Q0YZ7L3lbG10VAok6dVMIzZrLTt+lUym1m
7c4hhNNInE7EAx341Y7LzX2rz/pomjiAOFF3fmgep9yumU13KXNgKLX0/vv+j7QrvxiksE/4salR
WyAZxV/xbBfVaGS2XO4VURU/EtfxFIwL3L2vjiEbOXmhNMdSVuDKkoBo4tG/Waye6Ef0WdQhYz4z
FC2IO80V7m6QXIffIFX6jMw3yBgaF2QpMBZNa4B706QmEV8XpQj/c/EYVdrHS9TidtEON64IU9Bt
kGxxiXr0v3ygdNtbAySyEQ58e8yoCseM6FVIPbRuFWXXC5FLgdvXCUAruT3VdCnGCKaj61y2wTd+
3iwkKRI4O1QP90eJ1FxcRFZXhD208pbaozBISDm1SwnKMvrT+5MpjH9SLcC1z4sJM3sROfM9mPOU
+pjEXg6ruLwJWmjR2EtMzMRjQmNj+BHQwWBNJj58y7B/e6W/qzaHOoXczHAO0ZBw1+hbyKAvrEqN
axjnhQzHU2IaOPMMJDV9WXybdZlxUKwvDPrsXFDIcXDEw3REGZ3dN7/KcRMg3D/oVsFXL2wZVVXb
fdbpyp4AOemRILVGC+fiB2emzH5Err80ztBCMgoLuz50vsmW2xjfgj27O5emiSc5AxbB513SHBFS
clS1qFd3BXMZckS4s2YPK2xq09gCdnu3O58zPdx8S/ykxWY/lVJBTtlORxPz4BiYROpLBqY8/t7O
MZlOV7b1fQmRu0py0/3DnEjFG6NgxjXxELtIwYtv0dJ+2Xibtm7qBh+YnrFZ4y9Xqp6gFSRVrjXT
EklqcUAGpCwPy7QRzIM90y7C4eDqhn4lCApKU/6Dbn8QqejRlbi2S7fPjdg+OO32dxTQmu7yGkmB
9TTqrVsuDYdjCLoWqelTmpM3VAYDDuxguD4AjG9d2pLsxv7b3DDQelLDwbdzU/5KSLurg5QfojoR
3/1cUCfFX9iPLiRYc4kVBf/emGTJssTFaUSUwIVe6IgOx8wHIb2ihOxVUNpTMUSfgPYxMuLR/UPl
uJNc67B3XDfZnxs9EAw5RFKwqV87PoyHyD67iaBukdjHPcv55BJ3audAOuPASk3atGfPPc3osKl3
g1lqsvgNLsd96Nc3RyPJhwp8JNHkctb1pp1AfkQOYCLDoW6UAFn+9kfLluMPa/A0/dFKvV/OxH16
MH7vOA+4+y8Ta/XgUOBdEmI500vjFs8G/DmWA9AlfNEpkcijDDiFYXmUkNnehaKtwYM8XL4U9fPm
0CSdn3OWkxawJJ3eHv4bwTLzsKTAFFe/14gKWEqszITNp+wolzuke/rGi0W4inv3kPnxBbEBLmpF
bgUxra+Lcpc+ofhzxn/8lwiDgyqhs+ttNWvgvK7fXZBS7nrjvwosPFbte0r34Tl8L4wTi5lVy6Yf
XujSYUrGkWS4YUTRzE5nbtWLI0aUaBYusw16s3MGCN120+OY5+KPcB6eURW2b5/IVirsxXegcEnr
Obrkkn7Gnz4sGDX9eLG60xHoA3hFCtitKkB4lkCqNZrNH+v9Kfm019XSFFfO7ZYWRlsU8DIPfsHg
2V+HAVnowznUmyuDjJAjBqZbVf6Z2AaIzfiGqnHB6h7Dc722yVbeoyelxjuBtTqdjYEitw/aEUs6
iUnb5hKiJTa8w1DwWvKuJvuQ5KZgMtXThBaYeDu4oPoOnBlT3CmMak1pFZ8TBBiAGXr2sZW4+sEf
liRNklX0ov/uXXBvchj7dnWRvKv1UdpduW2Q9U/DvHO5EnjZYZURIOIMSaqmt2HCr53Y3ZMZOjh1
TQ7QvqkR3rqocGowvvPJ9FvSym+sspDn6oaP4rK+/qbOmnF5GTf0a1n9iEDiEPYnW9AAFkwjv07Z
dKE9KbRsa3WE3CnXNbI3/94ZEmHUXumSEeGsa7qVU+CFCCXlwyavm5zLODSmtrPmdomhrO2sbGbF
comHZZiw6QOd4Ay9lQ2XownwgAfFjq6rVzFzxeAxiYw6n7Bt5AbAhfSpGgyr/p7TPAzCPvg3cBFc
b2cExp+7dQ/V1djeMnNdKmW633ZhOZJqTKG+6YwCfZA4/GfHLFpvGlSVzi9at4J5Ux15L5l5i9eU
jQfuhvQzpyPV9AwEjbJKnKUXJHKoW4EEVlYciOmfTVd6upqYiUWMAftp9FOqAew847dLKUQbr/ot
gzxFfwgdEu6+Qrbo9AoOsOZxcMx8FYxFzZ2NhWAoUSJ5bXT1qlL5SzACnwgmCxVbuIaGJgjyf5OJ
/uapzzUhMSNzROqwOKYYZF0j+pOaQleI2yQuacsNBigcVFsb/nrtLDJ7P24J6vzSib6tWcuXT7Z/
UPFPOfdfzGuQq19TvsfOHm4bhjgm6p8wfgoZk9QQl76LS6r9j3JL7tD/L5JVRO5yc1+Lk3xWJXxE
Hd/NHMUFba4j4lcCgHWapwXl1qblSzQ2tO4vNcuCmrp2O9a9W90f2b8xMKl37E1mJ6myUyCyZ9M6
iQqNabBcIOIjYVLVo/5UFLpyGUzbx/VLUFzcDG/iJtrpOekc9TR0HA47OPmxUHPQ04ojfaPnpWfw
zTVmRqnXLADN5eaurruIoWXYHk5n1VnzNSe+Q83mroPMKQ9aTx7sqxNoE1f56EfiAdhCPmTa7n+Y
dznmOnqvDQTHvA3aQxFIb97v9NoBaydwytLz7ZapOuLXl3WETwD4ZmVZc2gbSxsI7QE7qbS9vVcV
xaaKuoRxgVOVIKMMVwll1ieuKUx0kt9DoV1AgAOg4sUUjZ3uPltEbEgaeMxhTn8LdxpSB0SetilW
Uxw8MD0s0lNlldINVe2i02aHGluCW3CO5nJdFHg21xu8j34yr15474V2FYKck2YntAFbeHm0q4hz
4dfhJhMaadRzhHEOY8QtCjckFAYp3zM6GsM4FWFH/ZIB5tIsZ5ZpzBNlPS2w6gEeu1bk5VH2WUk/
fHdB0Q+Xa9a3aQ7zcmByKson72CDKB4+jOPOKCdpUpzsmH2tQYWBQzOarqkP3Cxc3xq0DJ951TED
UDnvLEsBzUeXzGu5rGwRECrXYqO1Vlah3luiclkNy7DPn3TFyW56QzOoX4SYC0yTYxE4agkSRrah
QdF7f5xrAt3htHfBbYZMCVm/sHnZJ5vIsCc9wnEjixKmfzUnU1wz+tXhdSZuQD7TyS3kuhL1HJ1h
wAkvKaEfQILXMV2eNCKHv0naFNklnxHS1CDJtzlLIn3Wi/ewEHD3iSu3jwkiZODpi2q9YGPBduTK
yWzw8pD7PxYhr+BJxCv7oLfoCh+1r0ibccy+qnQspzMXvhQ2xopAw6o4mz3YT9G652iI1uhG/NNX
F65REU2yaV/SF9JyhKzfH2EC3jC1kDLqg4B6SHUCmRRTMzWESvPz6lnjS+obJxO4jVkq+bDZ/y3G
vRoN1prWJcyTP17cqk9rXHQPzjXoaoKXM16Zv2JkFudzLVb0/OI5tWqLOJ0jj8Wvdifn/IuPSCRB
sJB2RVuHher4PJddXa5iibA9T0YvCwc/tolD9MCuI5RVMrEfTgEn+C7xLaxk7Ws6HAd8uXRmkCmo
BiSqugm/BKTLI+/D89OmGQ/uLi6JcSiduMVnKATc9e9bQ7lIeQpx9Ued7Pk3vtRlypUdFvq2IvOK
iWvVQoGMBFyDknH2OrCl26Bv4Xa7UvJPVUtWXzi3ckdAdbRzeTndkkDLwfqKLPanq6TMomIY+lMU
CBCopvVbKKe8b3ySKG4ZuDbh8tM30Zzngu4qU6SVnHtDXQf7gDqnbN3FVux5tSqBhAoD7etFIDdl
FxMcUWh0euDjZCh0NQQKxiyh11dmBmCGb/OritqM3D2ZYjxv/rIBeEALClWIw3agAq4b12NKzMJ0
lzn4RJHXGnlxyrv6ju0WYqfObPia5PrhQ0wGIKtJ9BigLuk5A5z3c4/EgjamJepX5GQwJeL+XIvl
NLlMZAbI0stdHKYyLRjJ3mY2B6U8cZOGoRHvCUs4ygukt6I0HANkLn4aU8rwT95pfDbCt8iErHMl
7gqt2IadBUPgAg/Bgo2/jyF5jWZVLWx6xvxtDNgCATgbX0oJ5ag32pedQ4PkTsv/sFefM9iw4GWh
ms0CmOHloUGgo+O8ddNSg5h/NCkVZ9v8haQEYvXCtb4k1XPSJxq4KVD3w/o3qC/A+NqR9RsdTPMu
EhzDSGiuIWCa9pEI2Zb4nGQO2fSJHfbMUQPRw9ikav6h9dr8nbLnd/4MYl1JGfwkZ3ItT7iiOfbn
OpwZxKuleQLXxQKTjoBH3u6uXwhuXpqdQZ5i4QmzO9lSPqgez0FRqqM1kNmY5PI5Sun1WV4XkrLI
R/MqoMhOWXSSpYm5L9DpFk5ZCImiBZuGEjwqeV87ep70b6HiyInUamgt45sa1hCs24xAnlKgGvyI
Toi3IdxsZxIw2bUXk3W7so0euHmZN9yquDVkb2T7bpzJwLry4mMfYUg6iW94A/ZoVKUUcxj/SR9r
h3v/tCSyi8rktpt8SAoOlZNU3bryUyOmRtGJd2z+C/6ZnUECapg3ne2U86/NempC+zufaBCG6Ku9
ibRJweWu56kBthgG0IBsIXyz4cViaJ/i7rv/Zy+lU2cfVQvxhBidAlB6jIDu7TjIaH/rTbd4wZ4D
FeV50UQNWniFQxfgk9fvwjuDIbw7TnykTgV4R9/Rd1KIIngGDrprqDyeGEUTXURc4errA5cTpk9K
drqptxwA3psxT743vmbE7XhBTaof5u9A2bFVRfoX9MpbjKUWhXLTeN9yb8jC6XQ9ycIVISH4Fjs/
ODblkIyEXI5NBfVOa1fJMwb1wjJF57DlGiYpHkNNbISbqueuX12NOVwn+4OmsRe7ZyjTfvIdCuy0
fN47jX7vwx0eTveBILZKxYW04lgd0izpeeHKtLSVolBIJyp5tLfABqKvsucCoSrllxUSnLw4Dhq3
1vTqijsqPrMn9R2F7GuVmJJIJOZAgG0tMMyeNkTBhoigahwBDAls973MpGEoHTHlAwXEh9h3MsyM
nDvh6/m76goWSKmwXnGIYbEHUcvDqesBDg+p+dtWQxrj28BUH7gCwTLDtNXQlX3xxB4/ErV3BhEJ
slkZ2IrMaixillAf/s8kKiyTQFc5hqm3j6riiu0spjmRg4yXJ4tj0uKZIIIGoMIzZ9CfZA1qghJd
tNVfOKWfLwYDIYotHRV0V1CCO16yu8GmTGvyCeLyh5U9C3BXTA5kudCExgP6bid/SnmAzMarurqx
8u8oKjLsCij3dqlpPLIbuuuC0E6TmMSGFwUnXCTB1SOgfS6CeZHh5+ONL/V7XLH/NM5dPjI9VlEa
76CxfdSrZWn3b1skRcsEh03iPQ2gelwMZ717hPA9J7mhENdVp+5J4AggssE6FfOzq/9HaUvx0CBc
dFkG7zHTE+JSl2ZCM06VEEZzfbgQ8xbZ1K0sgOULXeeuofJ8xn/C+Vj0OvUkYOWH460APCzjA5Ad
3qkWLkhJXR9c0de/ygvpAX1f+ODd82sHYkB9pf6y0aC00c3qiH5cye/AapaRud1ChQvGSMbSTdUe
fhgJfsQjE7cw3RdK1fwwmUjCDg7i8CVis3dfbzIaqSVNAwD5QKgdVMQilKWjvOkcg5SOE6K3T7RX
+y1P5HJK/6sjNDhUuU65fUmg9LizjpPYl2XQaA0MI6Gm5Cfiw1mG4IV0rm91zCaKTtpbjUuH6a1A
8cm9+kdL0vhplQG87/IBFMpHbndLTgIsuZ1K1H+52hZZNyyLKE14fmpXVDrrizbRtSN/JLHuOMIm
ZyEZ+laZ3zzibzWV1W6uaoKr1s9sEFsOmx3O1QQx5aXANfEL7pElxyVJF/Ufsl7pnDeG8cgJo3SN
qipvQ9KJGuwlF3/44bpANXSBSoEC3vLkjK9Yz8XkYtegew/f13i/c9U7DYf/YZExZ+dF6RVqival
CFwhqynLM3qvj2D4JleTQBwbV1eXMeo6oyqzv67nlCql+wtcbpGcXBkPXwvjXepbL8Twcw+nmZyM
ARusR4Gy7Vmr0ZtgtLlzQXdcmW3ytAyefSee1vJeKuZZEdmrZL7ytIoeoQCoBAFw4mdcCiB7RFpb
S1AwstktxkP21O9tC7yebbRSUt82PSMXoGDHhOUwUQdF3rvdovWkIvtXR1gtscvqAkk7dTomm1fm
Y3tRVkjtALVfUuWXmkcKkXIworcPiB2BEQtKMI491IBpFMQ3AXnnsfabHzoJ5Ui8WA5QX+FQJY6H
rkCv5aOfBBNyt/uSejWzfeR1F+qcFFRg3KSFc0m5YZFDBNXCtWEtYWcQjPoohxSOwU2TkO0/ekfI
+i0RwpNp7LvvEt+UtNQ9yuEf09frs1eIv9IK9V4X10xCL7i7zzHduetvKJMw0IUOCXq3MmNZP96D
sP/2rxsWDiN4SmwJEFJOLVIFu06+X/xaKp/jr9lHdzEn8xZCWy5Og54aSIpX+rpgz0N28wFbyKB6
sfnmYCAFcBRYZrvgIKZ3rV0TXv8gHO8zFS6os49RTUT5XRBnhFmdluXTFaXhrTIORZ7jacmPOVQ3
gNvTN9FrQlldE422ELeABZV4inhT59IgTMY8T6hTcGDTmtjN/BEgcLXAlnshJ+fTphA5xOyC5Jfh
CV/EZXOoVU2YU2DezxgM00k1OJgh7MTHhRTVq4YqIF9DX2KHymR9yoCfjK5Q7/W5lTrr7QGYhd/E
qRJPuDbxIz+xLuq8RR1Z4OTmFU9bYbkxauxjxDdyYhpwK7I3thNDf0mOtyP0a6HpXUv0EXFWDV5B
FyMxOK3aFjHv1xGFh8dWiVmIIc7YIJHFb4qP1AMJ+AYvLIjaJ11Q4G5GFdrJx8bHCA4GNnpTbbRQ
3k9974q23/lon1+ypPtAmRcNGOKycnwZFnGg5eo+L6Hv2y53MkuUSD4PYeaAuasTPrh5XKIyHblR
6y4GiWYLLBAiLo6DQCIH4jKSM33DdrS48PV05bfT97Pz0Dv/EAWGAG0U3XDxkhiKRSMNSbEZAmED
xJhbpSV5QA3VqX5pfObGvqRDpa/5LJo0xh8JDAUf50Cy9RDx9SCLuE7UVVmidTkAPwOwnFtNckLb
phsIN9hHMCT5+DMQSNJGTFfMSFbKGJJqv9TnWySTP2T2pF7zsMU5FSx7SmKJK941GGezzYgWyte4
ZlTx6MYaIW/ctPHMVnuayeOKTG3JLHoj9Z1pYdLtGq2WixsuyEHHRft5TsgFPpZqWncfE922KcbC
3TIPvklPgTXeZzVTUK4b+ffh8T5Qu8LqPkom79qFE11ZL43zol87CyJzsiJ2HAbnyAJloGfyspYM
52bSaLrslP9yMVdGho6Ru2mTfp/S6zlru3pMUwFmVpmwEUvlG+qUB8L5J2u+JTTn0ts9nom7DNgH
o3WNZnilo9TLY3U26Ko4IvwN7JU/USGCJnKSHyO72f4MJrz5hSKmhvLeFp+Uj7pPXahEWH7ejDaq
+qpfOyDPjEAncL2S5VLMBJiHeqIqDumIkuAI2kZxX+sW+tV606/jVvfh/ifP+bzNbzGl8MV927Pv
dSzzWrjZQudcq2eMTofmUgyXA2GeoY1v5+OH/9laG1kUgeUUJQHFoqWuv/pXlrSrO0GmLXe4pUgO
lFOrtgBguCo91vx4eq6aOEp0Mk66gS7tmGX4IEpLsNtN8yckxfzZ08xH7nXWNpvomQyzqREiAnh/
wYzENJgAn91y8FAMqualN9JiySOul+rCEkgHd9Lg22dnTWOJDUuuTm9X6b2pMeefjsYGhx2elyTL
3MiLFyVdx2FvMGHIRk/W4eqe3RjFHjjUJJAIbnq3Q2EI5ltJVNOcp9AQP1gFoFcU2GvE0TqGHWAU
ufr4mb+x6vZ1FuE57icKfsUDsW44dOC8TfU5hZrfXffMvMiSRsNT6ms/zl9KNjDWv6yNx+n+Erc+
emAKppmhN2hFNIROZMdljtk7h40ts496tU899yCn/cXo5m8uhmyON6jkFzblNBRcc8D4+4ca+KbL
SAo9mHg99ZHOpVzXhMBE2HOU6wmxpNmJ7J+E/577CsThkQ1aWWA76ve+WvQoQT6loSy2g0hSBDsp
FQk85ujBZ8SWJdu3tzqI2zOhq3l1LOeVX2hpkCj4wb8n7lXcbgSzEfATz8DQWZL8oIJKTADnWZEP
1YA0ZGsKZfjMbF52kQvW5ZRViT52XiBllWTxK70H//Q9EPLMliuVkfvPTjiikmRdwLh4KT5d4qj0
u6qTFJhMiM0rJG8NvO2jjd9ezKPAs1CKz1GNc0wZB4Y3KnnnrjiRM1m2Kv8IyfWB54iBUPs6yBrE
jxeE+D4PNtJXcctQffcarAEraqYIgpw2cBrDQ99dGBmxdisobBUFSvgj8prRTcUgQbXE2gzbomHy
FV+M7+5Vmbyo2vnK9hTOUANq0z+TcSmpKZpVMyfPG1t6BxHHII+3RsWhcKqGn2U9eUJYLMaPQGCP
TbVc3N7YdUc8sXifQR8AdVXGZ7yTt023WlOoT4ms7MRMZOg1h3hCqiZgmLSl2DYev9Uw+6EQQP6X
Zo6LttsGiTbzYjJfLLixtOJglOckbtUOOseJSNOi7BEDAW7SOz3FGeojWsNQFrOejyVLfF0Xu2N5
5B7HmQijKPSAgC+I9tAGC47STXU4SL5vU9TgvheKAlxAzo8Sa02FLEicPL2Xlfhf6YsOiNm9k6G3
JVZ+ivmlvHK/E1mSxGuiz3t5wUDPJRLCOT76wDHeYTja976w+tKoUQajIDApXR+YmZQehG71a2A4
yGxjms+25y/RK9XKYD5SI7sDdXHQh/5bcNhG+bZCsJCNrA6AaJZUJai+SnYqROFW7SPzRYQgLA5Y
Y1Au9Ydvo7z5sB/UGZFV6fRtKVsVBfzGg9nLrfOE6pEDcT1qNFKopoc21r3BYg4hYR2wq1BApvzK
ZMdMzNXtyzD2GpWKfeeXjroSHR+kC0FiioZqJnaG8BZEpWyRcobRvNlykTs6lleGX51vn7JU/Ms9
DzQ6kTf0zacFFP150IgINwJDyeKI9yaldQYeySIm20IsDzXkKr03/bXq36kFLwzA9dLHKDV747xU
BaLAGKOUTIovJuxgv0vAwt5Eo3kFSeGsknQVcmp0oXv1mHPGCXdBVUrgt4PY2or70JR2E0Jjmr2B
iO97luXRg/TkJRGRgIUrYNEq/rytpRQJZkY5MHB3B4SR0XDsXoLufSVMNYH+YilNsnGYKFjdaorF
iPhalqbJJircoc095tCMkoyzRPl3rlTaY8ftp2A7ZWIWWxo1PZvegGlp3zsIkI3o0Xk8Alm8vsaS
52mGoGuVE5EmiwmvQbWPWpyulmR22O43jllQCAul+huMCb5r4ROJiqhEgbrfPdrTJA8NaTz7coEh
Q5XF68oYWRmeY9Jb5RNfmBIm4/+fCgRs2KQvovkKrLVJVIClStcZOiEEqKq2QrBiU77siZKuRBAW
A+p98HTi6v/oMRTMsNsv22YDCUv+Fh6/o9CMzg9TkY9Xx5QgZhZR95T6Fvg27hND0pr15TD3J9cF
eiq3RWQWrsadsURUWPtFvn08wMqFdT8mLy52+50yHGd4w3H2E5kP3LGtnOpjUw2SR+ANmrDyHChv
Ayg2f3Ur3AS5UsfnfnMAetoHTNUhHNs0e7NgBuWcPr2gMMV+fF8tMzr05vRud5qn8DseN7VCdFl4
Sj0bvN4d7/xPxbu5qXKqMPhrBgspPqSZVn5jaFzMBu4Gk+NcljDD+USYeQQnx/mZ6eGvYdFYOmgF
pat6ApVOW23TFDVOKUHLRhO0w9NWPvrQUY2zCyHJn3gQshNp3vUE7zRnNVEibm2tNVXPW+XOl61s
mSMauRJR9RMwOFJ0Jp9sA7u++aHtI7Jfk1x1R6UzI11mgEf6D4GrslqRkWgjPeDUnFizXY1509ay
mwn8yGXo6l+UxqE9UW/FkE66kP/GFfqrVvgrLngXUWVtLAsDcOIItVzXpGk1gbdsMfuqbc68WepI
+ozf3dJbccD8zOGXF9Gwn+Az7UHkXEOtu4Ntp0b9LeAIN6bhVPH5WrKNAfNS3CNK56seavwhfTPi
/pm9by9yL7vU0BUu20oCE9OgfXeA9PSlVORpZlg0xgdy5wkFxyRJTDQgfkptk9/CMTzvC/75dqh5
KwrVM1jgZeci90kSjkV0b8Y3paUIMmdoQK+8peAfjMdLGiUbA8/q3D6V0Q7LIw7wbgill59lUkzQ
FiBx1NPA0ycqJSWCqpELGb5WL3pyr1sJvlriQapBwe6/gY82LpQkDjlCvExL/mD5CzLqoCIONBlF
0Bm2TehnRRlRqn/VwMjAFOKIGgLt2p0J40tDxVyEMsGQJJ+1Zi5QYoRq4jzpKpVbDQBCj+osUTu9
eKAKKZ3XXGeAND2fOiG7zbV1aOyJcE3O3DndLY5pVfrOaboVV6YN39vqOW3JoMMrwYow0bhWlIh5
KMlxIy0Yzp4GNoYaW4Ad9G+5Et3FVmfPU+bKajf++Hvz7PjHxKdYNxZgJiVWATmD8Rj5FRjyanix
GYTAewBVKUiWu0EP/MQ+2eQ9mFQ+oU6/Jsw2wzZ8c0BLrOpwbLXHMoIxCzgtn2Viz0JMylkrocmH
iVtennM/HR7CUty7tftZQj8CPX1t5Jbt9oZmCXRZOAY4bp0aWjohhhjqN49H9Ff04N5DyubD4UEw
S1s2DIPkD0iyijcMGA1xqY8S3oopLQ7uviX1vtLkN6ZS7B9150dTRpiMZOJJ5kCRqiaBgEWp/dHR
Ei5D5nmy2WuwqVIEHhGXQu0wAtk5ESwoaT7migxChKd1tx3DAz4OCq05WZHv0CeTJAaiF8bQAkxN
zNN8yZHoIXUxQkO8GD+7MJpWqMY0Chrt2gfX9WZCygetlMc6UNzXLmD7bnVvKvrCiDgwse4ZHykc
89J4oyANMXT57GIDpY39ZcNgI+6fqVbAi5vA43tTV2hJUoEdmUPORJDT80ACThiE80Yt6H7zEZID
E4g6/eX4OTNE7brGiej9tTBTADBhMx3wgSZHENxCPq3bariWO/9RAAwYvVgkhCnIUDVtqMAbk6jp
an7rFp7WWIxlJ92aKkU3Lht0NUbK2DY+vXykhdzEKhox4zBGXEu4agZzYKwxi4l+Yef9GXz/cjpx
Rcy+aXRiX9sSCiIgjhsmyti9fN8XpZs0YX66veE6RsyIjUxfgb+7qSPWSk/45oJe0MEliNSd5kG8
sY6ghovS0g2QgQThUsQZGiwJSc96BpbMj2dnsgkJPQZ2WU0V7wOvpyiCr86F2Y4KFddP+gcoKiQt
tjYjJonPeo5ZUS5wr2zgr7e9JrvMGio+LRpZQIafGTlwWrgJ3meFV//ZZ6IoJL2jvetwoCTxeXRm
BtFmWAYgUfYUmAuHxu9VVKba1nZnZK2fAb1aRTiBmXYKBIvLQtURfg29nNmoMwhb9poQfXQV/nDW
1rUIG90I9BI5qxIQoWzCCHy2O4hNdto8bCi66kMfC/IPCWoka49tculiPRWdS/zYlv0leig2osOM
NTdJNvnFShDLd6Qx1nwybVk4KaqwA8LKJyzs8+92YYgVww8UO2ibhaJR2148eo0FmFC/ecITA6Tr
rV7blF8LvUPN5sU9QAH+k03GoL78uopgUh0LnZlLKjHWAA/60nVjGJW9b6G2T5XvmsIFPcTR79Tl
Lq9Pua0TiulyCcDEwqa7v/t4uLK+u6+zVjMp1DfmmrN28lipZUtWp9mNhYpUq9ipddTuEIPzP4pm
kw/U90OGzv68YEs/MzgcSE3GyeAdZlHhoG+x+bjzXjpe+mu75Y2fSZfXaseE+uCZBgSdaWpQA2d0
ReGLB5dPs4tlZErTkD4zqBrlagz9b7R0O01vScy6YQ5n/x9xmJ7FDVN0Bn10WpzfTyvS9m+G0yXA
vhIdWntBUfjKfMGWcaDiPkL/XYaWMazmwlTCx6/VkIb/PNzxYQKpDV17gshD7NchhBEu7dRdAdvx
1Hs5Z4VvVoC8Y0jjPTCGXs0MDbhdCwxWELmbCNb5iMkl9YdgCpor1GZnCJ1SjRnt+OaWx+ElBHiE
+QVgGr3xy7IaHO41fsO4e4rzRPKx+Qj/8HfjojLCTntGscEWkmftKdTZQfPMLcW6joQyBF9VrO60
jXxVWDuubpgGQ4hq4jwZjcoLAiRDY806F6D5EBoOhVmCoSSUEYRJ4t3dLtFJTlAyPQo1qkHZl0Xq
enoy6qLdUN99oFUCkx7OVajdMRexW9BbpqnCb/Cp1pxKNnXzeQhZ0T3S55qUptYIZHHGfQTQl9pW
s1d8lm4TtikX0BsWGWCv61lW6HoneLlxlenvKXT2Jr/TIJDJfmRQy3pw4QI+yHYbEN9UAVKX8BGE
a1ELwknbaiUFJKfH3mCwLTT3OO/LOC12H/rZ6CCF0YhPLPsKVRQa9GNeYLCHv9f5TySHXWI6ZMLi
hTjziv4p9FOtWC/gpU5XO5nJPMbkkkugBWDIgsFokyhfEPTPOCF7r1S5i4pXD4hE9gCcUxlBNkjO
viBs/EmD6ETUqKPOo1FyoKWVJnnbLEZ/21nFUcqUZnW0uZUxoZ+laLUsuqWDJcIfl6SCfKWixWNv
+k+zw7UmQyxIfLUBmaUASdiSwH6CH7snRAYfe3nC2zo8Lp3rMtbXn3eWpHXd6eMOXRMuao51COCw
K65PF/XzqkrD5UhjFUvAQAwm6jAfbtv2bxEeuYCHpVUIMvt2Y/mNCJz0mn68jm/poBKX5KnIkm7Y
67sHRYAQ3Sa5cj1sKiN6a5uzIorIv7dtV5HWXyOC/I54LNr73qKWKVNXxYkl5/f7PXyZ/C6/zjkL
ulS+DMWUumh/FefV98DP4q/EblwXMT6qBdIzmamiNSxMO9JOKfMhAhTXxYwVo1tnpLTwNuPFlXty
reuEnGSkvmsrNrY7qm16Qb37UEZ22X1pIIXdTqSCa7ybJj31cPWlMhIh/xwRBMEnDj6aWRnNNEe8
pGEH64rXccZfvWa/QjdWybxWjD1u3JprJRfKFDDjsQk0DotXwG/tgJObOvnXh6qnm86D2ploPzQK
U4r44cEVO8OtH2byKPQU5QkxH0cezsCDIy8jfS0wSHAYjMN4vLfPd48aGX85Cc3w2m3Xv4Dd3E5H
0p4H5kSnTtI7gAvht4eVMvq41Nfy3S5gz4hRvRwm68uWeH1fmj06GZN1IWcc+1sQf6xv7jqaZJHn
9qEla92PTku9BTkUGlI36y+EXjm0RG1TIfjvurkvuRj0G42rQF7CsV0ZdgNW81xKQA8bMWKkKLyT
dcxXnxF+1MFhkTW1H/dKVOIvm1ZDfS7NRfp5//W/+b3Rl+JmNN7DVsG9vmRv/VhgzpBwGkDMHqbc
YiRuukV+M5UZuUeWPlN6534WYmk0n2Dp0XC7psaUqbtDdm05Ob7XFHNflUJL0bx1bV2QtGrBpAzp
dI0+R4T9ao+ynV7sVCbeMAbo8ZMCu4mDDTM5LmOg8tGArzGAl48IacFVQA88BL0hJPwZmKg2WNuC
bX2/Dx02GTvZLS02yawQRGh3bfb/RXOlyX++DOjIMthJcluOy+tt9VQCI98NPNd8kYwoZWIOdRkx
h/HbnqGphn+jcblCEnseyn/B9Qf//rLTAEFNRsnMU9kGnxB6+ny+akBBRaUjsGH2KaMl/MLJU9CX
j+CJS47uEMEZcIq44gPS1pjSoz6Z3PMrQiBsWCK+pTZZOFXGkwPuxWyxRcPWbpD54ok0kk/j1uGd
DvX8qaxv9Dlf8LZkIiiPY8o2Vtb5m8YOgilqb7nYwwl3TDuc4ZsW2JEWJZSM0UcVIrz9X1oncPk6
BfSfdj+L8dUkwoIv2h2is0Fh7Bx7dQtU6X3Fw8id8vzRVxVFmPh2o5X/lhYo/FM9YXo/D2cYucUm
/H4w8HjxtY29+32eRT9DclGP45g+o7h0g0G6/3l+CmWl9IKz9q9bC1VAQWGDwTxraAOJ9HB3hCJy
5FcBBM6Tgl7FPbxjQGPRBjV8zUt7wFZNrmhlkgXoSkkcKeenDtZlIUJljT0ac7nNlpqiminlh6yA
3m6Nwx//qD+l8DrlfZyFpSs/l20jvk3D+SR+bmivRsM2Eb15mrpBU5qlkYLSoV/DLV/3dN+7nYuA
ZW+5jh5yeN2ovvj5ad6GIvRVDJ25a8pvtgWQQW//ANTvK+JzmjweDFSwvlYkjFV3BJM5koa7tOxq
bXuSMIhPnoZt+qaWJNXQMa3NTnnuoONunYM4jwQZ3fEgmDz3OlhX60vsHwrKNK2kIuQEwcbU7HgR
M12BwQo5tZ7WfgI5jO9WurpYz7UqqWorQFMu6H/Exh7o9ud/yBd2dgkv6U08Q3pqrsvUC09Kxsqi
+42I5Jpv1AM6MXen9i6w0oTDmyXbfI6vhnawvYel7zNCOzVoy2Pt+7M5WqJTNkzhov2eO6nGIZed
7jChAZUtdwD6PgKS+cAdEagLu2eXRtppYwgiliSn5rADsKPrd48QWN30mJAmeKDanYfg5Nq672t2
lpXiU1j4A0FjIqBhcTvUg62oIqbl7BdREtLOMl2iChPIVReoIMSOk04btc5YN1Zl+6jZqywZYTil
hjHFicbaWbDKzbEzSCz9Zk5SQmckWXX3nLl0wvMG0mf25iShxtvW5iXfFwXEk5KVtY8DATvHbrRA
I5F2EzcUCC67otwr9zIiEWVmhniOMnD0RqhzOnAOfoOeTYdYoJsrjIqXLKrXVbOCsgNGVjWWSLEK
ao2QqcF20AnB21yAIbCzQFQ6xNnjFKF0VwmiGNn/FdR/r7fRPBhtUO+cvwA8Xc3eMvmQzh37saX+
f+UAdwG8bLpwPUNgjHbO/ks6K1LgW/VAJq4mILA9q+13ZVb+FdPFqtmyvsNG0fQZBC9voCgajGVF
AY+tJlaHwnAiueA02rQhp4427eH1K9Rh6/EpQtJ47nGWNk6FtJCztlM+Kjb9AmbPc35RqykEBriG
fH/7lVXfK0va592Koqs34wbrAbT4/vWtCxE/NqC2TFNZgoaVOgbCsOclrEirdSYJP4u+0V1dcTZ3
0iLdforv/F041zHJ+ajZjfToGnzEXGW+mB2W0Q7f6GBs6wAtpt/qKWtcv4alIqOeYWkDL1X3Irgs
fE58Vlmb/8cdBlFC1hvG7s6l3AhKBIPI+lVe8RVjhU6OcVGhh6wg4vZL+EyNYksV73QfSxJlztHg
nuFcFbyE8qgqFP/onKGykO4i1DitqFy1zqjOeuebz3jLkug0z+etyIK34IFLGfqvyC8JHkBnZ+NY
OSo4+JBtMJKqV1FYX9URZ9JqUYz9WflSbikRP1vJmJmWIIQe59BNU8iLYRuypyoVCcH6wb+xKWzP
kfr7AbrphZLvLdkXUSy4V/dHezzPxgFTurZUUKJFwd3ziksC8WIws48IkPozvsdOZwEC59VWMP1y
16R1pvO83EvHRb2tCyAfexbotp+ZNFBMADVtYS4q/182Bk7iP5I99qYO10mqitoH+2qXtvnHf/+Y
iEPzEJdyIKJZzUPCvmm6sR0vCa1YsLaBKYuXngcQtqtTTg05SckHFWBgADa8T2GHYMDY/rNivNE2
z6u1ZzE0bIzvNcERa0xVNv3mvXarx+l4QcFzO33jzvMtOfrrpwxH8XFmG6ffdgPG0XjVkqgZQU6y
/DsanEQ0f+QhdF1D9+XenSDltdTvtV6oFNn9AcdUPf1+qbgPuP7In3JyWotc58Ik6u/SJ0koBwFk
QTp/EM49IbxLfz3q9uWg1yNJvQxfDZKk0FQjAO0NiEV44kkHbxIAPnvXeyVw6QH5sHCYpUDlnD+f
IIh9MFizPHEWuTEtZp6IF0rfcatfSnlLApcNc7lbZ/aSjyfd6b29Aurqn2TrWkrFv1tmZh3OQUo9
0WdpUuOJgB/4+HWKwrJ7toh/4EAmEcQvHWmUplBIDBCQqm97/1L+IhU9x+FluZX8WhkHI5BZZL7G
CkeXBnMIWz/nu0eM5TrYCF/pCAkaK7mQH3GkOh4Vd2ZfVPIvRqQY/6nJ9SBfVguwayCiuwlebwOd
NvQH1OeWn2Nz7vjIOFHMn3l2on596oAw9wyNshiznqKn3xzerIFDcyOM71/mhOw5qY1rOgg7AALv
Wt94ITnQ+zVVAZq6OASTyf+J/jYFnz9ODqjtBXNjRxlunnmQYQHaCugfsRWk/3gVmiOPx7BKqFAf
EKIy7vUekXah0yduuFFS++cNkdtK9CfTfve/9Xm1TDxDCJldNaa1OFElV6nJASG+Mud7Gf/jOefu
XL/nkWTaPGcZWKWub4EhLanErxBDBNSWWSfzvqZ656wI5Vz//3Grc+YHVRmohcea1KigK0B1MH3c
gquCdheVGWiVhtmbWClpl3G2SCOJ4fD4ocXPgXta8OghkQO3VrKGPc39uWzifdbc0DH5vlgsxjM0
pzxt4umESKpMj4KRmIvGWIQaThoiH5LQdwOgGFOe8mGzgpg7qNBY/Iu3U+xHYiWhXXZaaug5Xgnc
nsC6NdNpBkApqtKb7QfNNtBNS2oKOuN+XJJuEqa6C8SLgSM58ATF02mLEMI3WgAFFY0jAaJp4IPG
SetGp4iVTYUaqF/HHh0SvS6GXVLcPMB4hATvZ2m/mf37Kvc5sLg9cmhlh9YWiaYWSkgBaANxL0pT
3Jcg/xKUFT538N71puPUU17JsqGW6n+9X3G9Fo/6OzeZrZEmlw/+jJfdKoEMWLVulogargw4Cbd1
qBI9SY10f3Pgv/EK/oCyV3ZaZOOtGor5UNJpaMJas+7xn9kT1RMx/sV/elViLbd2ZE8XJmp0jlnw
owKuKBe1/Kv1XJXCeeCosNw0UppG+piTMG8nnn8e7ZdH3XF+h9o9UMvPS+TjV2C8MzpQpSfCTjmt
Md3kvGwsMTbGIhxtUfvFstUJ9wFlCNTMzD+EfnnvuJ06Moj73IvVaQEJFaB2wEJ36stPfY4UN5fW
jzVHwzzkFvQh5Tm2uR3cYzxF/oFyL2NJc7dWYngWEHXIED8L26dnSCPcgLPQ6mbaqrWDcB4Hqm+E
mI7Wv+Svm//7zRCHM45eYOwgKeM+zZ+OBjs04x1O7TQf6ALUeAQucZ4VjQerRY/lRiHopU+4zZNm
EoQPVtwe1YcOb33YRzOFopRutNuQbPw0J2Oqy9wryU+s9om4wsGxhCQ5tHk+ZP2TITThdv5UG61o
CQUH0OUH++fwE318EZ2ogh6poLYHwpf5l4KETYRfG6xyj9qme4ZZQxY2kGyz87xGodPc7rAIAVOM
GN0tceiaJCv2NGOzdZd/Ax4XhwLTe6TOqk1R/SA8FRccOkVRTc/kNQ/yPRNGbDytqBCGi22KK5iM
eOaPbIs6gGB7KgiZfOwDiTQjNr0iksBs5glDSMOeUeoG9BU42M8pCZqAxVd3Y1h6MaTmPwsjsdf8
6PAHPyyZKLQ3Rx9g0wLLYALs/kueMpCwuh0DroANliSRWnZeegEWet7auI516fhVN+thy7xkALRM
WVCpKx5/xIiDF9KMtQCduyONi8OZ384GMDvHgKAgY9rKXmrwLL6Ke9ApoMKTH8UjjyDA6NIvXpnA
jd6L531x3AxnFJmjdqphd9GQG6BYtx9vkPZ3OKO9IYax9i9dIMdwyaOx0MOfGd6Zw0vKIlZh1S40
s/bpI7xYAoNzNdLLsv2bxJkZIEEAGIa13IBaprp2DD8h2ligYDhutJo6wAka59S/thpHUvFSx51a
tFsDDoZVvHwsqmJwgMYOEVpapR16Q8AhCYBXRNVEcgMxXRvJO6BO6A++c0/tEz6gT6Kr/PGjSgRp
hk74aY5+gggA/X4eWRZI3EQ4N4yLk+UAoHhsQjS2slTqb4xjQv1IVmImYfiLG6mlBVc46eny+qdh
UXYpL0tC7YNpmS8VdQhlX5KfkupKpIqBOsNTeXYrl+g045OBnZGgwRPbYrTujC5pIYo28xjBdlb+
XBXMIIFeUfDnkdbUe8i9343DQ46RDEJcBnRvylfe73J6gtVmOD33qVjWMt8bIrrPeFWpYBo9IeLP
ETJkDm+tVINr1OOw/kGUQFIjsAz7Wg17Cet8s2EZGyJjjVPb5r0kQYaioeeMvHYRQufbU0Okq3sQ
c2w67ZtHENm5pb2bJFsukObEuLWpwAHSGKqAz4gkqmBh157WPs8rGqa/Z9Y1dkfF9Ly2dlPUoFii
ufFSR5geqyZVi+abIqxxrE2bPrOsbJJ/ujl87GOTWR+kWTRtWmzRco04OKtb9hc815rtfl+xB56m
xtQynyQfWVR74DQ353/MYebQInPjLG8nD91vvu/q+6sPhoHBuG1NrDExRqjF+XT6b0tZMqAPjLiA
XqocBToGV1PbLEY3alXJXxYVj92Oio4ct7Kwf0K4VrQf5XpbvMOqmt9zpWsAkibSi5ARzuDp7i3O
14v408Ilbwrq0OTAJziOUok/s27N0fiNtI3V1TSCQi4LefVnVwe25/dQN/ZbAd7aGG0gOsxvHtdL
IzU6RBF7qIS2FhwyrRvZCwTBGsXmSiy7KMSTEU7D+7IvEufiqX+az+5UbcpYPoznMjpeg9UJ/Kls
tUFV0MK530EI7b1nRqV0KZPk+eYQFOp5FdThkIIRhLgc7HK+jAnrilpI0+2B1Gg1DpisqblrZ13l
WZiKz9Ms2je+u1uhUY5WQtD9b+MFrE+3xkOoLdlh1P8+Png5z031BF5+w0MR+dNhGvpIWYLRnwEw
LhuSF1H4LG/vL+3b2t4jcgFpXcJQYECB5217p54TO5gUx1J3mC6iT8WhGUjVai8AZAYXccmpk8XN
FbXiyZwbFmYzuVgi9bTwGyA7ZNE2c86mIGv/GWNmCSyTh2Jc2ndLAUPPP2kMf+/C5EKNh33OC4+F
1+7UZ9P9kHufZmW8yJX9kuMRxKKhvyg7AARtGVGDu8vI2Ei3KOGqRTCzyV9NeEggCFQB83vvtnFr
p125/vBOWZ9FFE1t1oc4+dpP7fEQzE9g81LmvodfC3smPpjpv1rNhPlKeX6nwQW5VYkjl0yK4URO
+FP+P9kk9nZRiq/MCVo0zKyDyFlvGvlvDir2UpVrof6eotjpzezQCfU9ZLPQu8kYnDuOfW/7BrDj
e5FKqVIvCpkQqUWrdH+svJyuVtrZNx77jPcOKM9Cl3X1k1AEcWLZSBH82aq3VaGPX+yYAcgVCMCF
etKG1Zs+RoXO74fxQXlLmbIkcvaruL6nABBRPTcp4nlCQP8rpYYneqqLWJ5cpk0Adb1N3kX7Sswd
RZD35MtK65MuTK78jCJx9C/faBD0fp8y8wnPOm4qETyVDvIqZYNYaTYXjiPnWB5Mt5bimIyjsNtd
ta5kLW0w5/awU8HMEdp/Z6nPXd1IKHC2pSbP0+3ZglJv0VbubvdPrUs/Wa2oZxOyH8i+OfkQsLSX
C57ae2gfz2MK7koDyKwxZEJhrP3PMDoZkraz+5Hx7FjWmqcUWVSX3/jz/ZUu/FBYaiZ9BrMnmnBp
0nv0wpxaED91nIs/iXdFdXyAO41YnugIEx1iibQ6c117ozoaXwHkGztuWN+8B9VDzRMc3/pyRUdw
TGrlnOkio8eTJkttZqhfeCfdYc1pLmsIshKLa5z2vIXoHgU+8/UOWUFHDY58HYUvQ9OYjJwuRqwn
D9rX3qVfJb+x69BzeLYtoBFKLA5OIarPz4SRNhfujAl4bPhO1RUa7Lv64Aeho8zXi/daltWQNBl7
dA24T3zQ+hnkauJHNPWFInWTXnfu/qMiTOD3Mx5C6CiDW6mrpp1XSP9Tb0iAzYJ/GtBvCpabB66X
Ib+pPzo2P0ssy4QO3HpRZR+gQS8qWrRVobmWkmSN02GH8Cx9zcrjFkNdnGGKDvmCrz+352Ym5EuT
gSiFQmiCdTcteP0vZYP6dZFHoEBsIKYxIS8NCkePJbOPYw+za4oo0Y7i8j7F2vMLpGZ/g6jacH4G
BlKM2wDQoJ/HW51XnfQT7yqqWUFRXbhfdyV48O/exHmsOif4j1w1ia8ZfKfhr3fZsAiGcGI1IrxC
wTV4LLVLIYoWdefvVH3ywndWiKVw+znfCXdsFxZ0g5PkaX1ldHFW4CItRLHKSXWu6jbazEBLmZj0
Kn37DeJBncZB/x/e/xQGrlAdWFKH1SkFTxACatpcbvYFp2v87asa+Ikh8FQdVt6sDvlTVRdFgX2u
b3ZkcHhK4yyYVrgPWBmVXd6HNxCvmxb4n4xyexrwHeGLCDVtkBjf2wUSkeDk26KrH8/SvR8es5tK
ZYpl5BNsO/vZLCjpLJJaESAgIetiUJZVe4MoFD2ybKjRNnKvioqepVG4u0Sye37C/tRMLzdxn8yD
OlrtIqhV6b2kPc3CJZc8kSYUPnW/aQ3qcgfV4uY+TmQujbAr6pvzCu/gSJCte0ZTFTzw+ACUShdO
vHEVyeQuqW/TWtStkwKX2caE9tRTcdljMVxV43OZXkzXyf/j7n0GYIupiSz7g3wUYpVo0u61vhA9
ulW5+eQrRf8wEBcC4ExRfUlgI4AkDi5Zlp9kQQYAC9Nl10k8as6C0GCIMMrZ/QjISSVTF5wucUWs
Ej7DC4SwuSoUCQ0RKgJpfQTwOrIykAtGktqRyP9Jfa9prX4qS74fShWBuI0FQxgUeKN1RB14OdVB
I0iFd35y9z59WPbG9XwJtr7I9wRlHpNfHCSG24H1PipQf5DpJg9R9Ge/BvE0d5VcunxSocozYqUt
pzqAWpSApvUIBMG/Vsnhq/jpi/2917UAyu1hsQoWonWYerfeOP1HU2Glwzyl+LQ9rJq5AaNQONuS
qF+e5vvswiayCOLIr0jIkD3VjIEJSheQVkfPny6hOqprE/C01xJ97q42kR4+bwBKFQDnq08dnf+u
/MlF9MLz1/qna/iHLzY2DuZJaFJemxWAA0d2uc+j6dSYLyIhbk8+8bP8XUSGqOGPrJd4CmB+OhAB
rU9x8OK59xPwhA7FNaI3svGAufmGVhUYZ6M3+h8hPjLs8aAV0UlRrEbk1hmVDWD4skHYV8FxYRcK
J60lzjhrIsZ5C28e2pNh8oOf6ZGOlJwlCxHROJIxkSw2gW0J+wKWeml7ZBCo6RY7D+FVvQ0pNgfj
xoxvwcFPGcRQlZNZbxA25x6+WR4uQkve+NQvrFiVsHN3rWXfN3bbLRc5EldnyBoczZoO1/CIdERx
0GbXVCGNU8kaZpxvMrU21/dhA05EO2N2hvDaGckTg7QvQAOL9w4uIUDk95s9Ifn2iHjuJOxpKiOB
usTh2InbmKQpFUo9iyZZ4+v5aWxXwcIBZA51AxPHJTchhkdEm1B3kn4b4HcjBo7LN3UPzM5gB83p
2ERctYeSsG50IpBiOy2QWaU/tyajVRC25LXx1YceEAqzZpRIuqB9PFw2JFlkjISRrSO6JoKJsUAD
6Boigk6/sfXOCJ37SUS70840wssBxJNNRglCUkAYxqRaaHrq7mPoP7kIIN7zLCwJxzfdJa5n5Gom
Oxp8KUtACMA3syl7dpGQOt6oaPCSfHE7jvnXc/SheS8GDHZwlSp5FpeLfvGXitBphkSu4a0cSG/8
jVLf/1sGgMz61BK6TigWn/2trevUFw9xEPrcZUIdjY2rIyNaQuWrtv1z/lkj/JosL78Ghut7fRqJ
STzat9holk1o+JZU7NPMBUohhPhMK4lwYjE80Cko6gFMVvgq51yHkT2bxkiVWJ33rDpkC237+ufR
iZsgBzAwm/QPWH6ldIo7q6WXugZNsmxTC5Ft6/nqAUGE/hkZM7H4Z3tldqUXEMpHItBn4a16XiXC
v5FTH+I9Q9JQD/etEQChgkBUl5UYuvcyBBzBgeKnrGbMRSOyHeSWTXwViNuY7jvTXXgyUEUD3Bpw
5sFc9Umu+vfcaC2XuuzMIF5as7UJWteakmia5Zkn+wh4cSCvT0S/kuaZyzV8ld2129AjjNSjSGJk
VXALjyyL3IM7sBAav/IF5qH/hfwvn4YCCj4MuXxMvDSzu4632GApKX6RtQ5kMkpDgzTSqpnquKZg
1FQEUcXj/czsuMuCjY+mmwAxlm4Iad10udPFpyzQu6BGFXeWkKkYDadw4Wu/v83aYnYLpH21BX3G
qtQiQg+X3FcZU/lu4Kb2B+AeaWZ0wVI5Ul4Iia1CT4DpXcV6RKoxt/yQFk1FwgalqZU6O4Ktjaj8
kp4vT/nHb0JSskI4hlf9lL7BRqHEykCHC5WN5s4H3lthjXCFIa6YWd+7RzJbhu7/JfkI8fZMnSh3
HtKHkI2sFQYO3dBEyanBllW2BtW1ZjlUtWiSf54fqrOY3wBunCHqUbohoJZB1uzc0ww74eWZl+LU
8X4Om0Ansg5SGL5qFWslc2AxPlciMd/Wf6ctVLlfc3sNHncrsxidvoI9Q6122ZLa+Zs+Y7ErWSAS
SDr738VmOH1UhFSz017YPGwTxbGYmPSXTZVPdBf96udFM+QR9bWnKTdogY3B42/QeJbJ9382ZKjq
mHE0/q8Xy/rjc8+q/XKu/RvQji9XLKG9fLbmEFP13M6IYU/v+9vsOBY/ze+UwXESBEeekljJ32K5
iSc4FX2yosfaxO1brzibhIsvmMz625tbdIrArXogrNFCS3gIQ6KpQkErTMY9kE/EnuwxQYjWmb2T
a+zaw+JWxcuG+JafjBofS21pRvkathJNjOdAgYsO+xe7+8L8GQ6lx/5SPX+yjvk/qQ9RrCMg3Ssy
g4dbuzo9HoSec/WYTykC3cqOD7k3aa3dfmIFhEXViOacog9OE7ENcUTxCsOvl21JVRfSZy/qGydx
8pciEHwCZesvMgfQK0ornFQSvsn5BOn90we5/bMU/cTzDZFMYt6Imx0ZoxzJjtmfT09uOw7CUliO
FB1eCbIpQtLzXD8YE0/3CbBixo2utXlMST6FVSogRKp/2oXbEIRsMva1RZ7MRpudEIfagUVxeS3t
I38Nyuz0eImb2AlOVVEeFn9JRQ1gh3nMt2fQtw9q7kIgrh9AXSbsy9+/4vVVWp8n/9tGg9b8l0bQ
5F0Nwye5Mmp6vEOlmdQZRJHXG+w8WsPEEOMmRw7ArcMBn9uEnu68jmirUeghzED0MDEY0/wkiGkm
kTL9wQLw8WbUxNM0R69Gl7afoITuIbAgX9S3IhhZhfBMeVdhE4XA5KxolGuIzGkeSIFz23ViOwpr
AudoSECtLFGUbRM1w8wctgrgtiLe59FfSL8kDKrreGvKNYea463bAA8JmHK9uV9EJ6hjR8orVedy
u8hpjsLEP5gXJFsXDVX3PsgBE3YEJe/M7yF0DUJYkF2zhDLDAMra9+H3PGZn3EYNUNVNhaFlea1p
0ymXIHcIz/I3DmoFb9KZJ8rgwPZne/TeCehZ3hgDJUSYlsosQmkUD1L/HKmozVe8l0KbuZtqFZWe
S47sdUSmDmnNaaOid+i+n9Ez8Su40tMxdRy51VDqNREJQgYNigSZLy2WKiyg3I4Qsmm0wum5KxYf
WzMtIsjtdf3eEEtsGEB85xNMUA+EQP4bjdHz+obSyxQsV1fkrOYySKlSPq34oUaIRDUrfuDDGRKp
c016PgzkpjvdUwT83sOeo/BgQ3IpFsgmyUPKBzhGvVIkSiZJvAR8kFiCA9tG6QMNhuCaXu6/S2zW
vngTHCs3vXVinyvqn19kf7bLhNZsQYP3jMMfJAzOMZkWBnOJTfbn64cWtzLk1a19+CxjVHWx5GW4
dyPFfwSqdmd+mLATDhspDdfyWUBYHvkusVELVvbCMtb/o7VNfP34TPSgWg7nh7XP7MvhuGXxidBt
mauZ/5XzqJuR5Zthvx4gc895Xql5/YMNLWt5TyrelHN9Npu1dsqE/TkQR/VfOu+BKdxL43+uJ1Mg
EMNTOv+fGD7r3yqNjRkEBN+MrEWaSQtPeZrwKjvxgHTpkr2GkC5lkUIfwGal0Kw9girc2jS1eEaM
YZPid3CBg8l78L5lSPbbetq1mxMzHlwXWS4om/6zPWI8c27Fc7P1+YkgoeR9CqQlWewM43HBan4i
GBV+O0BcDuXHBAq0AHunTpo4W/ia2+Z1wPcNkMpZEtguUUoytkAmWbX9xMxns8eaN+EVCXZVfmYH
PpUqOBnMRyD78cO8Cv+SNEkxpBjfODalMtCJEvBUhfCb1r/BlDIyBkX61sgRIcGfoucwjBFcoxTC
UJ/6Bwhyayohx119DalECi1fkPpn+iCRsUt5oGJWGcMIMReCt8tOWM+Dv32fYJrac+v1m217fEM1
ZxT6ARck45aQnLV6oG2khJzIsTejIxfADXrkh80zAQhjBND3h5kO94gFPpYQLzttAfiGUFqEHtX2
nbvIU9CqrAHh+S+F2ztVRn4cqqIseaseAwv4eVL5y9Czz1KD7DjMv0MzGSgjGhI0T/XVE/a02Tyc
DuRSONZkuWQb4LauOr1AXuRN/GPNUz9vz5eRFMzvRhkZ80Rrc+cFWA8tegVhT5/O/Yxy4021mVOI
PsJVzt0yVGaP4J9QAWVBCnB9Iz3NJy646qV7zjh5xF/aNqQQy2L7aw0Qg9sscEHqk+33yBkARD6y
XJ29ZtGm/1LNVZ7keyNXrc6++8xVRkBFi2cnY6+tXS8uUp1N5P6FFIg7/fx3Lf7OAM7gFxBFgC5q
zzX3U97GSOiKi1yqYAqKwx/usf11vvQMQfVrJylH/znSEi+J7UYL03yN7gRBVcQ/MclYe0nDUvWz
/1BH2uzzlH9v9P5SlkwsjxtRrlM5gi/j4iL3xQNn3EuiHPQv7zDB+sro3eRQd+afy1TnwcVg5pY2
o5/S6WRZQl2GCzHzi7w+dkyZPQkDCkdgjIxKyjk5g7Hd7JZU8nJp6ryzuYT7tbcDOSam1dwZVXEX
xXULirDIe+4hgso8CBiVoxlRatjm0xyXp8+ji8Q6kjCVuNBR7FGD/bnbwmE2Efrls4UVFgVr5h8Q
JaYivweCORX5AFEXsBby2o5Eh0vF9WLl4YlyAsC4nlVu/DlXUmzlERCvZwxUVpQxkq0TJSBob36s
lcYhi4dU8ImIw/6ofSkKyEprZhnOH53rS53pgz/JxYoRKg5TVQ9yohfrvuVq2uSE7o3twHVyDStx
PxLy9sLZuWN04HuMLRJAkL3MuitiAOO26CEGbjm1wC4tK2J27Xb9oqfqfpd8+pkoCGAQKlrtaz3y
e950grFmx1kBB39SCDw6XoaRY60c2f9sX5lLfdZWGpjLcexCbYzKBCaH/DGDmYPbwpYzBYe/Y5Rc
Q7fuqOyxVqruMgUabBJycJf3OcU3DhHZHF5y7v4VpE1lHQjQcStNniRPeLQRdRVcbQX+wIzRU3yI
tga5G7JTlobwtvUYE8YrDVPnHLIMuECu/8BRgM+Y3b0PvyoHIaBmCKMMal31TR1J9vB1jh5GQTLo
1qwlzrVlOu4IwZXvh9/SskA9GjcpP5WFVLXGw676Ix6dQaFRBuejCqHuexlDR7q+mcEhEOqJQQUp
LuQglzNLZC/GpW0wXSWDWwl3gcsH7D5eruss1uE84a9E+Lcft1+sKIiYHw5pcnFh0mR32kZhiwGA
U3bKP71NykqK09iwxiVXTOqheWWhiqB/HFFGPmB8ab26IoDFQo7zE5DJ17vQi5uOKw8RckH5j6PH
o1o64hzTXHbfPQTW60QzPYbAL5+c1gy47vDYT1iEpExzWk3B0FYTIn/wPr+AxJJDvMKtDzr0LY8f
MEkKqtJB8vKD8weJRSWcjtVb5QUPtyIqJPOj+CAplgO/vKxfWtjKtlwQuIVj10Q4I8ATElrOdc0L
TD1GoYZuKsuRZt3w3ypRvTNTQJdGv1ttpNRgfsxChx52gSgcs4ZR2thGn0bCI5Lg3AjiLry2Ayzb
OmqKmkZt//meImg+I+lkvXAwNiD/7OlUMRXE8OtCZ/Qzc5zaOL2vcFFK5lvTPpxIeWksOzaEj3uK
14FPMOpAUMcPvD0ZQ2GWE2WMtpgnb8z/987VGFe7wU6a9b1P0vclWPtAB1u2/RdIx9n8hAw0Bshz
0fcj/b7SrcUYcIQL3iKWmhsqH0/YszLRrDqAeu8ksczq3t1uQDUPb/LI3TMWDrOcbDJdbqLDXhqO
8TdO/em7gEtRowfMhgSS8pELTyX1XPKglRGnA0e4jChWYdffmfyRafl5MgvRAewQ+quZZh0U25hD
v8JbwMODoWTWY/M6CsZhIGerCoI+FfVwjlRvYSt6YLV32UTF5yoiZXFujky6bdGMOwYhj92d7Uh2
s9Qj79M3fVlXjTxnW9PSV3SDAkeQNECRBUIjaNaH5FDkzicCaqZLlz9K6QTiWoa8YYwXDYkusnvh
Fap43iBQjNNsayzogn2r7nhQSo/kbKjEK/fLtLOTy6qat0w8kJ2mrrMjVJwY/pc7BIwmmyacKhGM
FeUvRVDUoAinlWDjCjMJte6fI6Q//ouQ/djjN7b6Py4PGKJkHcckh4d6zPK0OK+ZN6qX6xfCvUnG
PK8oj4SkbyqHANh4ZbPuR2nFGDleiZ2oMvGJ6THw1zGM4SSeVie1kP575pqTcKQOfJP3qBWpaQbc
ymjJUkW9VIuK6tH8T0B/9yLLL16Nz/ocrQYx/nWFJLp3w+hMI5Df1PsA6CIKRI3nz7MAPUj4ynYL
XtdxBYePwn0kkIq14kKPEkAFtXijwvAXELWpF0BXaIrNIKK7HV3SqUvoxwfSmWD6aP/Gjs1/iOIU
cv/wUHuuiLJ9nSuIrLF/9khRdkm4E7cZmeh7HIYAwIkXBAgJF+CFhShps9JOrKffSEaSRPcL0FXA
5/E0PVtMNkZrfmEgEUJxu7ELIPXvIR0iHU/DrZhbfO1NECVgKDvL9DNVSZ0B1nhz9uujNKLQTbsV
vSlz8bCFoCfmBAT8R5HipC+WZe9FU0AqflLETrxRYcYThWu11R5KZ+A7vPf0vP4Snq80qq98w9hG
Tjk8APhjRgHC4Ww1Ujm9AuhFGAT248XPKO3PIoUrHsKbTOtxpUG1Dr7ZVjTOzfWtvKGlXCFoi8Q4
SlFm1TwtSor49srLFQlW+wOlggLwMISvdhf6NcW6Buu7pl3+rkYkDeLRte22JcvRKradKfsKkXoF
7o3I+Zuf1Lzie4eqsrysdMtcT81F8wqLb10slnJw2pag9gQzZgQaf46/HcRjAupmJxJ5dZj68BL2
3tAapAYkwQ5B8kVtxXI8SdzEt6FCwsmAMYm9cU7ZM1cIoT45VlulxsUaVlgffp1pZrJkddnfLmU2
bwjf0NytaXkP6o4V+TbSgWNzr/a4hbcwfCjV7fekQoTJHtrnESwrx0fAC+swN3InlxQZz71G79BJ
7MNCHdo1gUEU3Uqgy+N6bY9LC0GvTa83eBuhrG1pqrF54Kwyp8swfRNj4B1Bp7tt+DkJKPQMWOqe
84eKmyKeb1nzelxF+HP+O4QCUg7FpOkS6jsb8+5YTRDwSdfEkmP7hn1qTjZTFapjfApnOpH0T63T
/5veF9i5EGZvD5X7tOnDQCEehqfcfG8UQKMnlU65vG9ZtldOcAfAiaJcDXYTLa3A8yU8+0F20CRh
DGCEnClYMmfFBKd9H5UPJe/xXg79WagkgnXj2t8wqF9/BWgA22ySNOejt20B0ZV6DVHp1ZVG1LQH
mzjWuVsQpdSfHlIifjpOzS324UsyrRlvaUCocD8SVPw53QIhqAjLUytbQ9u4SNpAerHG+RDMqftZ
ma74aIijJXArND4B1wCjqMQKihe0ztNuRA86eFXRtYgNL5hL95anFv04o6eARN03K1iBzZHEmF8x
emzFXRsCgzRl9/Xc+1PmmcYialN4tjPx7LREAoVvq0wqwsQLaEp4XRE2gtIa5Yp8B/xUQVc/vI5b
wqlnB6gQPczEYOPmksLHwWQ9O5g1eNEOEejFUDdZcuEGgIBEHf4x48uTEA7V4m+oCNkj38GmBCOx
dTRgLWzSO0+aZ01sf1oWqg6hmocQmYwrvrvDjo40laXY3lospVLIbxh7uEiyBVXynjEVryZGFdtw
On6jQ9y6iM/57Xtqe4VzZEELj/nvmg6Iff1rQgiM1JlqVZUC9cAbLgwlyXQLockW6W37ZXQhDvil
I0lw0pFl+U/cGJSDM39YTzN68lGCEDgrUx+OIMliyirCycAsYMTxgngbRnG/h3OOhkcUJX5N259M
tdE3bHbpvxrr2B4+5vYWh1jAdTlPFn14b2JnyIMZTHesGIpkHPNnA6s1zE0lgvp+GaiOn/VZ2q8G
0eiKLVzACr9TZv74GMT2+qOylU7/orDrWOVGxxjteIBZN3241c/DceqlxGfNYU8KIvSjmYKcFoLf
gqK9lmNchauxFowMW2O6yte28oQ9sRkhODRsYmbSxSuoZWmqCQs3ADp1GXsQtaOlC2WEjq1c8Z8c
DBM1UMAl67cHl1UnaGAN2LPpRdWZ/oTe5hO5MCUbzWbXsyzv0Ju3uIUSx5NEKIfowridsEOUyc0Z
9c7OGxYyY0QoXZzIBtFUEyMq2VELLwRE10D8r6mlwa0g+pHAdjeoS+ADPW32EVnNG8qEFD+JcZNZ
EzxIh7cPKK43DXidPh+UxFVBiVQ8AoXmX5hWRXcVGAizJDYA2i8RUJqda5sdign4xdC4mTiQiGkF
kv0fc0JKE3TkyVNwagB2ukpBAvNPuGh0jilMovLXktUb0eCUXjV9BVBUJHN3XqaspSHa0ws4Ztv3
tEzDXjLrLN1rQ2Rc859cSLNeiW1Mm0b/h+dBbgp1w+lRVVzOu+KTdD+d77LEQV0co1Ez/z0/nQ2p
EcugK0Jb7ScpSlmRP2ZgSRg7HoDkrh9yayhUvkTdf3siIPSDTyk4f/G/caHvnjp0VYEJgx5YYHlU
vZvEkwMjoLW6lMQPz2QsenLOdNhMedl7u3ffpz36rOza7t9nk3utSXxmTYOwxYEusfbsWaIMjjsb
+TVGqGdHWRtfZXl2BUjSA2jTyAVbOWdUfNVeB1b4LB/bXCEjCM3MwyaSfX2yoWZ9Ba9vgXh1+YZt
zewcEwV8xzjGbnWSOawzk7ccP1XI4aMv+lSMHzC8HVSsBzvYQ+eea0pP3/aw+3gZx0qn5x73lvrI
1TJjDM3xL4i/myBSQAWY/ilMO9sIhmgpYZY0y/aA5vR8jG20Tj8m0jFF/u/67HCkG67hGPCH0/Su
kq5fUe8FRPXdS1tX/KYEb9GnVfpupx1Xtg6yHKd1IMGIYavJ1naerFT/+J8wkwPfxMk4amXFqMwh
uqLyt1gvg/2csS4WG6t0PyiFpw+N2vTmY693MeA/U/8Nmn+/6C5nLFpgoo8fEFKMR/Io/zf2nKEl
6g3srklyn0eKN6o93MiO/BY9YFJ3hma/HGv2Exwdtp/jdmjjpO3vht6DyTvNnX7SeKP5AhAlRD5H
O734j7B7eq4/bqSC6X4zH83v4Yb3GFVNpk/OigzvAY2U7+QkRHF5SFte0bDx7L8VBKfnGpsJG3dh
EpRAZ5+eQ/GxQWjAe0+MO7hIoc52dHTJv86CHQ6rvauamypH7bm2LggDhTKhYPkXeI30hDtcqffy
OkV51ZSto+qI26Qzd2ks0Zg5SbIZMKGnXEEJl27lBCPm85oE1ApdMBSySBKEc44mjMENn6zQ2vyS
o8of292jNWbZ9eOmLVr1P3udaYYlah6dcJNvwe4XZ0pl86RpDjtKxiLgKbwvYkLoAPgeUJEL79j9
4xVHAeX1//OWWOEPGQaX5MY1tQoOE01bKur9N4xMSmEewicrKs5WkpSSa+stinRvjlbRSI1V+Uo7
oYMRI2GFiI0T/Br4+kI+y900Z90CEcpVv3n4ob8NYQH0CEXdrKrSnDt8gNrVkun+tJj3CfYzUr85
o7UB5y+kBveFVh5cRc3N4OH9MQeX6p4/Mvnhg+OQ8ZryNwSVtg9nXY62MpoHRiQSoe8siqiyJA3u
uRvcv/HP8bB1RecWE8uwZ61WWCqOL9/CEEiCecOgVjsM9D9STCgAJ6iWXPcmwRh21Jf7tbsbgUnc
UolNLhyUEGe8MF6/I11tO/gM6RZIGtJphngVt4Hk0ojHJfdA67lEO9MrMFEecRxe7H3iDtuRQozY
mpuXtAPDiLoay8BgZnGTDfvzRI5OGDJQ3cEVhUxUu820vcHsuIdGJK2ZDGNr7QI0+qM3clwiEEZR
eyG4UTjIOlUgZzu58UD/vcI05l8LhwaSk2BBf6Gu5nH+Mh9n8HEnL7CAMkHS7QdLXS6YcVeugdWR
GCMin430jSiNGPUUnVLNFByFOmbavp4VZn3a/iUE6KU5MTiozU4rSZQg+Vo88MHUtLKOIJeLO1V+
hpr8xfRTd69pgTxXxkVzepOopz1Cnf1ja7Xc1XFYKjL4czy7GGLaQrOdDa98tNYMZKCU4/TkM+Qx
RXuJqX/eyu6twdhMPpH8s4xSqunan16yS/ctZ+JC3xIhpLi+6AKv/d9hOKTESFbt58o7108ynm4T
aJGPcR2gVYBV8OLsd83TAt4ACLAkHqRekbmzPYkCudECikariZEmRKIpUHifc2LRp/hOoksx++MB
K+NmeTP183DRRk/yMGwht3lI6wQKKenMXkdAi7Yf7gbWvzDTSPnNRLDcAP3Iaw6fIqfOF7PeUjGL
CPGgbsILTOnuTTMiDNwRTS0dL8WXBD2shsWbyFRxwxwcuhPZCqORsYDTbom/4Cky/1ee2QCBoaKT
6ddsQrIT2Q2MxNfTTEDnvyVBuYTSrI91xtB7LkD7qA/S9pSc13ou0MoWlCvygWNfwdA2sKncMBgC
ytqO7NR97pZHC38E4ZoGIGAva8KqLB1krI+j4oMRHESQZ1eQyeKI9vh9vlp6IvgG/mjpv6kgiAI5
RpdBRwm18mI4V9+8bHuk8WZRZ3x1SHlTLL6GLeve14E7jqTEYsL0BL1gcGl7g75AyBtgG44aLaXr
TH5+aADZMFnQLBTTs8T09DNCdFNS3/mfpcAWxLycxUuU75MFTf7ABvjOAEUmua/bfRmYiu5rWk6l
XzFgiHJXhvVz33aLWOjTZrj04tyxypQigVfemNQuKme4V0Qr5GQxcwaDCd7oxVtH88eOq/+BldP8
fmzAPUUeDTRlFh536osOt/h0k4C8wF8FD82ii+se7ik91TSTnUHfjEZweB23+BQjePok8i6l29SG
lCixonhOY05JM4jyIdYuv73escBZ2FXLPKy0lptQ4gqBNsQWhN9laL/OZmFs2gD9Q+VdjSNiMGcD
iP6GK2nEv9IpqmoAfs20bEP9TA+StQNJ5Zi9A9cYJ3UfLlmZu4wSDmnl+8GdEm63ZvXReTpESdMx
OhNrEuIJszuYz286J3cogzC1DxKwen1A6pKRQig4nr7mTsjr08Xy3mWK0G1dr5ERMO6wYA6MtGq+
QX1jF9zOO5g39DiL0P8ga6jUWGjNd01CdFVyMOlIstu0lNhVkD0oqu9xwP9+efis+cWWF/cGUOw9
im18kGBS2ZpSYGMZcUGXEiB5H8yipFr5hzYn3ktszmdXVjqIb85oUZ06GFHUWfsIp2wvpHnw+rFk
w/DyEiDbaP/SCvN4DUUZzRR5vWU/xSN9kkGi8bBke5oKOyQ/RXormYd1lRbZ/1SHo1882xRH4jsz
4LK6NuDFp4FSj7yqBJWBKEVEpcS3wlGCgW3TqWDMjClX87PnFhDhVaAlj9T4HeErvl8u24XI2WWs
KAc1t6UBRqstoUSt/9lBPyx9a9B9Y+SLwiEn4sQ9wJYpX/mLu2vXRQRgO6F/aLUA2otcz7wuF7hu
NXO5Es/BkTPuPt3T9g1Kuc/Ut47u6tukrd99S1BWivinR1G+FtRQQ5Y/+YOxF/HZMt1IqAP355vr
/9jibM4Z0vq3TMKkJkPVq9ms+cp9icqNl5aNKgj+A2NW8beWYLwvy6bKr9y1OJ34SJhryJsCCN8r
gUWS8Tr62cBg/sNQfNhu0QvNFhBfJHeWdOVyk9fp/IqRQ92ykxN2Fd8OWCOR0DtnMe5C5q6qBPSH
XstCjeDPJNV7c/1zM7zJgh31HsgN0Hv31AhpBr2fGxJlSUuVrMsFdgdmRnTf7DakyzMuM5nnVR0M
LmYvuXTWhtGQVGz6LYislj8ConV+rxLKwc7a7Vt0CORxgcvnrqpWSsr548HJ/bvkWBABRUK5uTCG
+EY6k9RHTa65suCRnv3CT0PQP2gv0z5iTloI1+feeHQcJDPGs36hT84risgwBFi0PjwN/+w4cXKp
4RsSQzBv7UOADBZ9fBtci8dcQMl3wQvutswEA0VlRhMIHs6jqd+SUWPa1gCXTrbCKO6S8PRY8PEP
Ju7oDeaeZm4dryztXzr51PdKiqV/5BK9zMZUIhHPlv6D+ya7Rrk74ogrjs7z5Ib6ZyrIGZ/qsVnu
iAfrx0jvQpYTzOGj4ufWzNYmijEXShWJhRUCZonNKPdhaHfBOz31hgqXMjrjmC6AIlDMoaUDHhOP
UzKR3AvIhmZr1Q+fNDkzOZ2D9u5ONKxxisryHLsObVWrjscXemlTWoY2Q1tGHHYAxrTgBVmuD6Ec
A7eol3mRcniW5vobIje0kv8GKfDwq2souoyiYYeqKyjH8MfZOuXdqADeHn/IblqxWTG+R/Ep2tS0
TvjBPRehY2t9USa4Mn5c77agg1whSMwSlZTn3kTJVvZ8n3Htt4q7xwfqoUc/xNhVYlSoOMpm4S7I
IjXcBqG6LVKTnAtdevbbh5vCRf/oadkr6ZZNyoURnn14oOpC05C0HawjXtibza+swTK9KHPgLFS6
r27EloZFKf/2WcdTLNwE6QWTFZ8lzd1Nzi7/hqn5dyBB3zbPeNzpTwh6Ytvv+50BEKcvCMU2+ORQ
Ilycvj0eDEVYclM4ZBM7dSPKM1tF8dJlsnECTqtPSVcqkQn+1p5u/4VJSkqfEJ7dgbGUAjt/Sdwl
YbrlCPS/2c+8Io4gcLUQEzFGiSuK0OC83E4nhoLHiWHnx9gnxp3aVWc8N0vVmxeqUuqkZypTStir
yiH2Qt9LaKCj0w0GJvjZPC0JVMMEF8+NWRhY9hzHb9igjYvlePLncgSfr6lxHfJmlwFBrOeRwpq9
KElPgGk2w0aXl9HjnLAvDoW3UB3nEwuv1arnyCvQ2CFOAQqBijcZzPXuJmeT9bNJrbCyTaoqGwua
g+2hpCxXFhG5GdvttP/PQwsDWugzg5M+JnPre62tn9fkW+Dbw65ZF6Cy7GB18h4XTUcmIS4UK6KY
8FGo33T0zOoVzYsQMHJK/nMWG4V/UfapspFXbKMg3ycF6mVS+IiTs/vlPYuCZXKHD3lQuzv+4DxH
GbMUj3dBDyXyXKk9F9ucy5IzLzg9FV5nJGsKeN9FAIwEYzRGPCVndsdiZ05JGy72JfJWM7uiggkv
Jbip+UfLibQka4fQ2uCi9lxkECoRFYaEkpD9tUgiir3x9Ck5YlZI77E+11ivs82HpdQrUn3FZVXF
eBI+V8ZxHO+K/UCVIjCVzecDoaR2u1wgC7rf90gJxct83pCAqTHY7iV1gnaYw07ueWegka6tvfnQ
qVtwjgseel1OyrdqKQmK73+ZyrXwCTlW1EC+5M039i2LYBIyjGdN7C3NblvcWQi+SqG7I5QWiDdM
hALihzH9had07JcPIQvLSjsu/3XB/iNo9m9q2tRHyqSjMcsnmciA13jYO6U3se4pnH8d34F3GX9B
4orYAMOJvwX8AuPSxRQRCzqXhM5QUKI3RksYIlyMNOQoloBmm1ZBxvAA2J6ssS80rbUmc4tQ4n49
wonPyTqzdJPsp0Iw2GDkmNAdd0T03hcLy92eLEa+tmT7r1BmDSnrEGhlL/7IBWvZmNW17UrYuy1v
0t6GYz2J4W2KJnVUopHg1g36NJx1qRxN/HMILhP8bvUltGSSoPOs2+EbVSnSguBl/BKMa5ZPW4OV
UHB8OIB1OwGg0xkK8aHkYMpGYTeRDywNcG6oxSIXGkrBgaRsPSG/kQzbpo9vFArzHCL7N8bEupw+
ntinfrDVF5F1JOS01eUzlFUp30Ouly/AslcdXnZnGPP1T6hI/Xwwar+0jJ7PNwhmy0dhBSmJWwra
FMB7+KlWYfuDNmv3TQEPJTSkBz7l2pn/vbwQRRzBXh+jQK1hi6EEGswnIgBBRZLOb/WsU2gPQC+H
fN5IJ3T4RIO//R0Wrjy3p34YuPE1yaog8iZYqFaJouddbKOlmifORPh+J3B23skX+suEO2C+jQPm
CqIhHz8nUx9rX033I0pkcHD6RYJhRrAX8VbU+GK6pYGWBGh0GMjC2RvkuqAYZNrQaETtlM960hyL
lT7nZnRA9A8WQmT19+etcQ+/yA/HYE+g1tJP09N4A8jQPQ5bww2jOAT2P0Hm85+SyRXM6LsZAhbk
9YuLvMrFADOqbCo3GPtOJqcQGxDkpQLW4shVnrN7bJkZQDKlxDNU1uV01xLKdzp2ql1tD8mW1/fr
tooyGOIuvcTBGOx2rKcLmluefdSysHOZVYolmmmc3NMgcvO3qC1Acpi/W9ppZEsoCPhNyltEfW9F
ALQMmHhft4EBz2bHw33UKWpSsQIZ1B4RpZ+7aRRodtinkdXTvkZNK92N0xGWcu7T/ZB0x5dNjsna
TOatc7BjTuYQYpfur7cLkS6NAUANGvTZe52cwaawlfVrQalU/6fK2W7uj97EJMtgJB4jXrckt4QM
kr0dakzVbOBAIdEqhEBA8Z9eVi9TovJ4dhPo2+x7txw8rREaPpd8ldMp7geqK/pL4jUNMY9Rv55M
/IuxAKuBv+qpo1uibVy3TW9Mr24nq4u/SOiMn1Bl+bzVKVIqixFUx8uQm1XEMNyWudBuJzHL6vmJ
ZzEf5DyyHirOQioklJ++cJx3LiOnK53dBEbNFOg5/NbOc5cBKcAUDlZ3sE1xvfEVE5RsHbPCNo07
nJpaOJy7geRNBemEbGkZATjUovOeB4ZcbTdLpt/Ilajy4c2k2zJ6loLHMIHdjC0LnP0uYV5tiCs+
wRKJ/xxnZRdkSKBdv3vxY+UfJx3DmF4UJggHzxUPdsCycV8HupJfMc5uMlHkQ3Fx+NsJojxdnxKI
2KPyaeUTvqACDZ9yVuc/WArxKOo3ys/VVd50JrGOm6hPE+p6Al1fKWxXSGeMe8wC16fQE7PJO5jt
JQkjyJNgdubj1ZTuwBM+tLW9Ne67cxEpHLlE0MSJGD0VekVS/uiGgOMouDVAzrtmpU1c/BZ2FCrH
MLzU6oX6GpQe/9OEaku9LniMSBILx84Ndg1UfDV61nZ/LPt5AXFzDZT/JNESbr+Anc3lOio5/HeI
k9opmQ+WejJA7NIshz4h8d6U0833I9adDcfIUH5GT3CFn2sgmd4kDcE3Wp+eg9UPeGKapSnNzBi4
2yNvOeRalV9dVADvOXsutN8sWPX4I2h7Pz0Xv3bU5X6FXhzplC6MbrFH1Zdjw8KPuDT6t3VMUx7T
+KGovqNveaxoTvHvkP2lpNgU6eBx1CHzrGxnQ+TBKmc7ZHD/JOD3A2sT/PTS8YbLqyCgeQbzx8D3
snFcZQagJedRHrBhDD2VhkLDfaj+JNCF1gz/VGxdzyQVUEIZlJz+Gh2dHdSTlKGJ9sFpjfdzP5jp
wqw+bPaXDdvgyO1e/IV17DX4Y2MRIMr8WQQu2bstjwCMkNNCJ+L3TI0aB/bf3F8lk4Y2qp5qI8cW
rYySA6HUzj9UvKOM+cxKVUWaGZGlHqBQo7s7aP+3/gRV56Ib8qIlBZYOymKwBjg0OrB6deBCFA09
cNGUcQw6U62qcx2fjxwaItWY+TWVBSJThvpYIl8rmbdLQd6ezTx2/CbCMUJZyO/jjcE5VruNk0ow
l2ic+78s5nMPkDn3KfHO1RlzFvsuXQU0OIyNWeNcaEAAWUajhgv52Gudy69hd4nf8j0OQfOco5cI
ejXjX84h8RRfn5qsAF6nY8J1/tbXB5Uc63WTA1zPf7WLOHxWkay+dPFO0c08g7aF4MGhtH57AkCA
ksWK8LGxQ7Je5OX5E0sOBnAM6Da4Kmh4+E9CgQ+GyvjFINTP7YSRNn5gvi2kF5sJ3Bguwda2/nLZ
LcwzYIr9/qKFOZj/GQQeWnzEcb0Im+IRD1K55M1tZ26nh2v3EFftPBLkLkHGY9tGzoO0lNtTPuZ/
+yq1mjichjJUGQDP8du1XFXATVHs/W1fNujzR3pYU0hoxcsXyd2SNdCNkkkxsJq506FGSXXdosNM
coOGR/5Rb6SN+3o6gq4cGsjbSBplm17lg0juaE/qoorqmR+qxqou5L7p0AUUgSF9EJPz4tCJjOX3
b1/RWmGOWnw/V0CkqxbDbSmipchv9iGTTNiXK/+jxQ1RdL+/0WuLuKVFHuErO9maltCzMUef9ARS
1SWXOWWazBBRMo0EA5uZ83QXNFxKR43YtPWeh4CimC39IIKiB5U5fUYkgVfe17Hz/8BFSVz+uuBR
PZK3dOx7s0FIKmunf7iSyjy5EE5tV3MKFF+a8FgD0N3pYxOGL2QrQboWjggiQlBSbOWiFxaW3REa
eDf+B//nlfDDgulnyBinLKoWZkrK9KdSAuuKsaIzo9zJUIlmSndvqtDacGzj8FD8r7eyWEa0KDmt
R2w9OpfMCuq8IPp2ccj24blkQzzAki6NsAvBvGpbnEB0n8+3TNfpPhPwEzf3baUQIxjDi/5Qp5bv
BwN04KYymgWHsOOHZ6DQw91zG0Uex/m38JRW7LQDBvnqBCJZJMmsQxMtYmr9+W1j7Ecew9PzdoMs
DbnryaIhmgTpU8nO8rJiSRSgjntdfOf6yUeuR+B629FVpRbtKtT3OG17cVgjrRcCpY2Vl/6/JJLN
PaQ3VozOIznCw83cYhqKNX3ajwh0BXGlP9n4jdFVDQwpKvJ87EBaewBxE0kjLm1oKIT+ehJIF5SB
8MBWWtwGQ4ycmlGR3WyWb9E0azILxdVzcT3xRM+MB9XvfwCSR3yW9os3oRW+Wroaz8BkaGAK18Rw
+GFnsBvE8Y8eclyPx+LY34gVptGpuyFi71PmmGUNEK/kEU1BiclY9Stk6qWf5km0RgfB+wYwjxAZ
dEF08Q45rsjXYicrEoHCBPwqUbdT9tystNlE9zNBDz2WdRNBugkJMRaZ0UYHLB7h99Yk0KF+0suJ
uojid856JZ6X1gmnlw77pUGk9nv0IIa5Y3VoIhw3j+0IHJgb/5D4oRV54XVayfuwbxcdrmjGhFhH
c18woWg7FY2jfIJzZiduwECK33gB+T8ycg4hF9jWjzmzlPixqGIXK3nyEcJGT8iAVjhMoubYHiit
jqqSOGVawkLlKhVDzAhmMbUvzBOq0x52VAxhg2WC/UAcX0D6+RbEZTi3XvMXh3GfiFwzblkJufZy
ZKtRdmQr5CIjH9bVgEP3bXcwRrx5yY8jcVwPZ0Rz/YgguF7OYaBJu57TjdeH1q5hPWgi/Zrc4TVC
qYmhgKx+q1StZjpLOUz4F5dXTifA2o+lr9cKy4Lvj/866PItrVDvl831UwkHcXE2cBIN0xOnHjBp
nNdZ0ZOQH9j9FBvFvUhEhr0gLR3fIUKlnNsCc9wMAVRDKpkfOAlIZL+l72i6EuKQH9vIjuo+oj9s
eFznFzvQUr1qgZam2iuStkzSZYstRn3leOUVVeiNSCn+VQe3eyB7CR9BsOCmvxLygKsjDAMZhE8+
1eNO/vqr9ZvM0EPVLDTMOKFY3UYK5oVDUFJwOd6XO+/DD8Ajrwuq0TXd9yOsYvc0Osp34GdE/vuY
5OYmWamgBF8hZcdHZ+q6HrZ6qddhR3wOybXwFg29i4V8x9+XOq5EnUSUt0BumA7ri0BXz/dQyZWk
b+cwQEn5F9Z6cR2SFxk8JTxF43tXltjRWEtGHeM2z+FS/xssIjcMs9YL1lOsqZVdXtZ0HwWAmmEH
ecHOuD4Sf2XWVmoQSwybq8JewOIBf9lCmkv6RLAvFqV8CYqQ2JYkiYCDEJ45lAhhT7YcsoxpP+/R
iO45JXt0pm8fWg2Pm51Yk0PMXYwXL5WJOBVrkdmmfFXUsi0pSAha+MGp+mIG+T94rGU//eLP32xM
/cT8Fa9ArbM/Z/CmPwQoSubyIZIjI8iwgCLNJTsXzyk/dXa9o5Fl4lGgIL5nJ+/DvF9tJjDKqpI0
bfW4R+HS9Xcq4ifmMN6FHRk1DOynGtXC8jnF8J2DrEYDencrZ2vQffW5YDq55aI2K6i+19Qnkfh1
08dlSky/bjkXX+WCFHnAeCJBGodnL5oGMGuEdPWGiMrDV0+KVyaiOM0FqhUI+ZBYq0MS0eLcNH7t
yAvfdFxbZSFn8+KbYhr8MN0OgOdMoK6h5fzE7jvHs9vvxMdW9mJ2m2oz4QqJ6XwdcIfWBQ0AyI2l
4YNF0PwlbqDypdTQvepZbo7Dv6VAatOYVLme8bN43udgOg6L0ZsDzmuwxXrHJ/5SjIy07H77m0Gn
kVsQElxINT1UBrzo1DynIDWn5iWfnH7qEMKbsyILowzPe7QEWnkA8HO4+5/7rR5ZXq3tvffDNpbF
V5wo8Wfjcn+Rj6Zek8sJbxieV3UkiB2p6Nbam0w6umh3ocf0nsyrefIeAXZ+71cOzmYK7UuHSiW8
UshW6+D9097ZQoV4x8lNnq0BlPTqUmOhQ+b+tX/FBdU5dMtV7JWY/4zRu0TtdjGyywaGu2jDCxox
Jqy2KsmLhmbrOmrwLGslAX+kK+H/+TDZCckQq/lVn83CSn8PqBjnBBHnYIdmUIrTXWKn+G+HZmtP
of8qzJgxZOzKtzi8jk4gCfdf7E9MSvLggDmZc9GMR/aZdHolZR6lAfH1nAIHOY40eBVVJxXeBYei
Zgl3THCUiHsq5FWdOvVfjxu6jQeAD8PP3ov7vtBGDoum1jrwmsBSL/8ZvypfaRNq2O9lxmPTmofr
dbWHg1HHNy/c2lmlTizTf0wU4aDOL2mQTa0qHW/2H6gcKCg/GLE4sHy/5XSX1l0LkvW9gxgGRsBK
4AhsSdrPjquKR20Qu3TqN70R9yzX4Oot8T5lQYqch+gqojmTtplh2PjynpEenKjc4NsZTft3mfZg
v4iJxwOH8U5RzT1quumohWOq4Of1q9ibu6vrpabJiIxz0EhcFRTlYo+Sfid2WbwHlPOWoLDdw5Wg
24xgID0IE2hRkRb0iUJKJ8tdBAvbSx1GGzW0FiUPwMK5FTSuynQ2vDNyknBPebLpGChWLxC4FIqX
utzUofWEUPdR0Bg6cOF5BOKjNU1YFxp/oWPBkm8LjYOtI92kkPLvZ5N2mjsVqbb0345Bbm0KvQOV
ew3Onebxt7gdb6Z41DwXIg16ll6ZgIz40o8h4j+xXk4VlcBwkZYncTBguEq3yMVdZ5o+Hd+Tk6FI
JFwDhOCsPotlvH7xgcqcDhRf/XxC2kFLStdXORpng3SS9ZK6sU6Cx2/gFxCxb2i5VsnPWDsKfASE
iHn78dHZTajBbjJMK3i+xeAXJkmyTzGLmE+Y+dnCSnR5O5fdgAWCiUWIw2txyL7R0V9eWzwBv2Qc
YxV4ocvmKp9CS2P3FYUyZeHYD3EmK8KdoP37xYGrYnw4bWy/qNcdApcFMXEUGNayMwaogHHsFWKc
Y83chyyay0jzQOQJZk5g9aLxnViSI0pZMig9o0pyZgrRAbHu13Q7b7VrXPIdxsf7QBjM0t4S+9mD
n1DRFtMhZRznouKwDgeJK19i1pAR/f4ZtUszHsDTEt7yK1+N6+0iohQZZdagDCCaaW+xMau+rAjF
hYyetN+7F/tJL6Sopi8nZVTtvqfp5TllhyUyHGVsPLPl4Wplo1K4yAB+w1MRk2qz7XdbiRWjn29x
fyV1rQTNd23c3b+tyvElTWU3v7OKLtoM1WEX6pVn1iKkCdjcw+g5AMeQMMu1wH9qZu5P4/hBdVY7
ZHzcsojH8aAhavQ+dijm+DAoSiBmTxSWJ/OMkooA/VfgXuzPOCauy02aKePr6GXlC+UlJ/4ceaY5
cEy9Di5gWMBJYee2p46o7P7LC1xYHR8xuREp+3Jjf0Wj7A0rnXzThwk0lw11sBfyTz3MDl3fBmGy
rWKUP0Kws2tWQIx36MOmHBjy/5dG3VxsuPghT76T+UwYfyhl9eQd4htit+hev1fM2BEx+RRv/BPc
l3eaxEPbjn/9J3sunKAKzcjBAYmFMugyyHg655PB5R2nQGB4sXABL0CO43DdgUisyE7x6G9go+C4
0KQLYhvA5nofqiBtRXQpV8s1rKmJimh8M5Shatt2opCg42+eDsWbxWCywJNTFCGGvmGamhh+k8/2
qZwAupy9hcMcdshWjVpt/KdZocVVJE9nH0/VkghlsVGloH16hgr5Ct9+N/4q2QbwK78wGhkOqaDs
5ET7CDrSJ72ATCDwvBDia7qKksP3t32+PpCsmL+Ob+rJBoS/VQmmDWlf30a9tFECNTUViQqi1ES4
IcaPXx5mv3a+MwMeOlanng4TawRHCG62gCJpX8/gfU1rp9P2bFuF0avawqseUd7kmgXQ8ThLMoUm
ngFN5kO6MvIMPF3SEi5m1IDMNX+OMYCratRdjvFHdTnd29N1exUNvYfvhC0ymHs0JBIfbwbbm+Wg
S6Jmm38kG0mzvdfyfYRCQYNdetJtpFQeE1ZIepq98MflU4pzHMwygB7Qs5oxUIKC8o88Rhgtdn3W
dBAAOdRj8j8ZgkHQLJXu1leolwsMWKcLO7pdEHcQjqUljntY2utNnvgxmlRC8KebVbB+YxHYwmVx
9JK6VOy+UeB1qr+p6b4doV+2HJhdgRsWuhFrBGqype69opGLpiq3m35Jjl9VYIbR4MnL1EVi7LN/
ch9Wwe6oz6poiLDGdV2JuzcNStqcvDs0u4fQKnTzqrJ3BRAcE5CViTxLUsqG8sMV4t91vTt/sbgT
Cxc8w/2ykBSVdIJPdadlGB0IUEs4qo3yVTaVv4VWbqgxcMIcAF/bX5OICnmHWwrWDo2tn2rNizlp
c2Wg9LRIXEM9hRRpOAnEFFeBFTNramu0OjLVnFcwqjyz8vO2vm5fwd/FiCKzjQPGBCj0eWxI1VCB
VeloZJm04nzQaRsSKdU5xDQ9OVLj+aQg4cFS3nxti3/SmzfdPh5p51DFGuUOysFywmHxjA08xP3v
RyHZF044zkiMissNzKLZ7NKZqf6+yDvmFlbLX8g0jaTSS+509Vszss10YtAzn6/nYnGFgIAye25w
Uzz4tChAG3FLI7nPEjLPjkS3rTyjojz2yYBsW3MmQ8hhK5a0Aw+xeWgw2l5w+ABmSAna9XllO+bA
xZOq/JmE9g4Y0Sj4Z4BSpivm/dnS4keZZW30vtZSfLkRhKv0/SdyLXAqQGMFkrHsNch9s57UsZsM
tn/mt6DpiB5qEaQQxSxlTm31tKB6Toe+ZayyBl4Tz2n6Cs0kQkCZOnNzvhhny/RjH/1h2WN/B83N
HQvW6lJvSjarj9WOf/TuOMdxskzJKgK/rQapkVckaf1IcWZr5D2kzlCee2aCXdVCLVc4J7A6iUEp
omKGgc0M5QWDUrkjLXeIW38QlmyO3daBJbdEssqfuPmBBpQo8H8PiIWuPOenY5BeQBy/g+b1FdRH
DjijnXYVj1sj5yRoT9rdzEUUXiiOyn6h0OkjpXhfsLnD30uE7zOsOrvJ/JxStWE033PW9kko9gt6
CGarY2Oxcjl5a1bbew/Wn3kzsyytmzING6Nn2l58MtjftCdDBa/aYsbzqQYwjPvIhru0Thrk/skI
AhJimT6MRsv5zojhGchrskFVPBPA4Qa20+km/iy37z8OdGbGPYxQa+ZWYpVu6lM3QLDxCpx49i2l
OlmSUlmAY44r4M4BM2aK3u0lgMuo/trra/EAZIuf8lLPVfR+e3ntNDjbykpEqxz7W+9Vkij/9Yjo
ytXlhNordOrBLJpzX5zis9Ei6WWZ/mW+TIxkUwwb+aag8m+ST8IX4wlyg/nDtDlCedBe8Y2Js/O3
sJqZl9yD6RVdGrZAOTxC+b8+nT/k7T+Z+JY+tJqhcwCoaJd1LUNdKd8d42sDovYDpCt8S02RsG5K
i84dHSuEvT55vw2EuLfyaPgSac4CFpbhTm13Qn2pSWyGQL8LG5fe2QiM3eV8eXOrDTYDTicnKsvB
ZOHufqBBxa17PNsaPm9sTEZpqGFGA73OvyQZT8S48dOKtT1CKE1KNJRYg8C6U0uHN752T3KLJfpD
nrfRqCOcEeqdsVYirYtg53f2MuSaoS3xW4A5zRJv0IASANPkVZqgPGAZ/dCpCJGb57VgnXBEyryP
jvXtQjhVKZq2Cfd2MuGWfCOISOtZBHlbPJX0oG+xlBeZm9LovjHOFezTt2Zh0yx/v4kNQ4RDJxr5
tCfrrNHMDxI2cbgjaZjPFeqBscq2grAIKNAFAM3ehQ1hd7D99gnb8daz4qxNU4Qofdp5amkqCGDl
W/XzGyARirvTHU23AEgIuXjpkB3ib/us9gHb3alJeSeGiLv2VnDVAeYiCuHWG/6QdfdillzYeP2i
mhsz3d6xJzVHwZSnAcDP4J73xC290erdIhtXfoY/LDGgLuiYxkb1LdIqChlc107saqJdFTXoB8by
LZ1YBSLMp1K4UlEGtGY2dSu53/zCZvbbGYHiwhEvqEoFbIN06+O3MgRg+bIoXaBOE4YrWRUppX45
ldjXMq4LN++Wto51aoecfDO2LHEiyKyiIf9NXLkPN9kgBNHjYWS0YkcuLSjHWCUqQTsQ3YOlO87W
zRnuP9+kb5f/iO0ftCaul7k/p00RQ3L3+m5zf7YfyP/7VJDqy6DcGrAa736rYjC4CUGPr1YlUNhZ
No9Scb0c2anKLd2JQQ7F/Sdp8Tyt1cg1CNUhkHc6BFqQnzWcFlYH4fOy/hh9DysDJNye1d5zEio3
xudRBb7okrW6hdzMMAmqH0Ql9jUBIzGk5YzmUKLfnpFx7QN8MLpuLaq+07FDamzAtTxBdZuxY02w
syhMmBEUj1zdUBboT2xhFaThmoNuxCDt9dcObOxzliwdT77swX5V3ToxZBlysv6mUAzgLf+H8BXT
awEtXOwfEhs2xtTl3wGQkUjlGGWsEbgLYiAJTnMxm8ZBvq63oPvLcYfiQFPsNBzqkj2Hu6bnTKo3
a4G2Y21rbhQrkkfogIdB6IYIcSb3K4VGB2uzLY3um2Mi1Ur8SPxaXL5T/DrYc5BN5+xWIiKx138f
QNPMWdsD1MFlCnwDZcUNgnm60/960dGibGBsZWdK6kWiU5FIMkfg6ulbfQwXqhXNA8QDjEZFZe6Z
hEoRj+Mmm2dL6uAwozRII2mRy9UzEn3AuYdzeg1gBTE9Q2YTOBWYZS9wLw2dNXRU05QdG0GQDCsb
a7RNezl9MbnZuZuHpaJ0PVNjJs4yrBu5//0mi3UgRxH+UUVvkgYiXjfnUA2f7KzJ4UTXzM8J19AI
v1QtNmAOkDBk6h1pT7/OCwtVOl5Dm6DzAVE1APa2pnXn+CUETtk7uJ7z+FZDPYnT2PC3mNzBAlMx
N90zjD2JTEKco+QZjzOB0Zy4IJbiiUYcDzlhIYP6zXwpbeojkPc4tkMTv7QMLvSUvp76tzgZIhvz
im7auzfPK6WMe586TFBBatV9PeLBTE3AqnIgVjZ/ddpxMLwAlP3ayW2NoBEa8YhkmFsx6k0P2krN
0gIJqe8NO8i2dsz36/uqLfrWySU8HQd9ivYOnKRxPeRBL+4pwXComS2iPganHJtow8eMODrQs081
GxHTGm4SPl7SWzKQnEoNLP1G+cblgB293+yxr0jyjuEUfE2njb8JUjeihyJuDJ+RnQMMchXlSHeH
t9suTQF6xkV5vxdP+4PoXMsR//uNWsz79WtdxairdRohBi0yPiFHuXJ13nKatIuBc7jgnaYs7Xxj
K2TDyZpksEkHO0aKswOxnckUgEEOBNpcm+RFhF9mo3EvoSRHpsr+qRvBclRYcGNq9YGu55OgG5ma
l/R3ckLyfYIBv518J7u8Nyt6Un/w/657Y88/rS0IR1w+vb8u410/X1SlWzZZBEfbt1g35eza8Ax0
7EylD3CpvTmwOBNpjTw4z/9dPstxLsnXO8dJiJ6QEA9c+ntI8/QEXPArEwWPb6D7EZv99m+kvAeN
N05kpgGna+AUrZhD2kdgCZYrcyjbi1KYuAHpxKplsbdGj/tYxPC6fH2uFCfxcFW0UztE8Oif8PqW
22PoGToD2+qg6VF7oaibHYL2ZODYzDfwlKCuKXDW6kaKqxfD39mB/ThhCbImO4XP6IoAUT+vCZki
nikcQGjGEs1GjLRNtGdzF5pjLSSXuYQJpD5TBrSFmw8sp7i39w5ADSeDDsVMeV3otph2T8taonI8
0QwZRXqEKfDCPKv7Fm6zoapfOWpIG/fKXX+e+cwG+Ml/H+y/aiAhgTJV6pOYAGSCkvKwlwRGCrMw
M1lSJ93BSX5DBb+kUth6jpVTD3N7B8CAsM/gslZY5Cdyr5khlroSKyd8UNqL2Ekgg21Z2JlNTXXa
qGPpXcVzD8XYHDb2pYu1LOTJRtd3sz5pRI5K9reJJVL9wOHQqyIiNCW1R54V8Mh8Z3+oTdHHrb5V
UNOh3GyT+3RFwrqXS1erDcpU2MDHcKKOXVb1ikhET2f55O17g/0FzDwHzaXIG7zsdKZeWLcYutG/
cOGxMLRyGBOot3TcWnk6MqLPTNsQJPhNTgrnElKMfANRyonZmf/YMtx377mqKEHuDoZxzN4BDiFi
E0Km3neCUkdKkUbpSFAXNO0B8CulawWdqX1hpDPqd/Ngf4soFjvR7+BHTWQHMZyvT5ZDgF356x8S
qwSutTViFlItACom3VmBbyN1959VWgFdb1JGGfduKHb5vKFzsD0pVqsSaqPLTJZ/wHBnzImYJj0I
b8J1OJucYRqeE/tSZkoD9GFVnMHSf4BHVxtYq7X+KDoHwKj8IfX2TOpt0fUMh6EuqPHwMPMRjH/T
TCoGKpMO82zZmdtURhKEzMqtAdSW8d6/uZGP6T4/YeibYy/p9uNiGwOY+tJpxj4D24YO43d7CHQd
LPHz4PADFbBwXbtuazbFLDH1B4TxI3U8FRgBtycOk9veYKzLdxfL2JXJ3UG84QOg6O5RHopGSVnI
wf11EVYBxkzyX0LLrwDtP/DG//+ki6OR9IpxJEaFiT/l2Nd3qaY0JsaE6aRIH+mJxHYqANlJRt0/
/3jOc2ONeH5ht4HAyp3Vwh79TdBH116zrZoMMIH/w1piArW0ffh45jY14h88joaaAat8IKdxvSta
GYGnASDxl1i5EgeC07nrhhxqgWcpKiO8pT4yr775AUZqp1EBHAoddcRKiSeM1sBINwl5zN+5qTwW
lg4ray0mfMuiXuJDaR+PuYGVCP5+LEgKocz4dnrfHOg+J2i8ZJUWA4tblaisapdKwJPeRcqMroKv
G01Si5g9x4pkQOMxKK2VyCRLDMEgIo0iCUW73nHkZICjc/xaOZYqwoXPV9WbgBWlGTyaStPL4Tbb
xJwv8vu37JWvtfNUCkH2JmFR1AgKF/WgfjApwHvaj4CSKZhqxpzQzu9/hLNMG+AnC2Er2l7G26yB
farBaId2XMmxbOc4XlGoifJTklaOFgATzv6845yyXoD0EF9AXVeJeSKNI4YQ/8UA4UfpcLjaoUlq
IzYvKjLnlR4HnCm0v6qCMf/N6xANUWRBH7hHae+Xt2Isd6QoCNOfLtyK6oDrxTWzdipl83CUF48v
91hyEmiQyJJRjF0TkAMruomd/ARyz78RbksSiDdGtmMLaBZCGI2NIY0pC76x6Nw434UI1FKNJ4q8
JocUCvykVDzuaquGq9N8wF3rZZNBz3ulKUAUZgvvO/QTGsX9a1z51YUb2F5M2OkfzOfNtUugBBOh
v9CBWS62G3HFGhdoUFRW7pLJZbQ9WjojaNIgiuPW2+k3FFRp1oq9pat8KJ9xsBg/XQVR8AUjDYIO
4ZP+12gBj8oFxLyvSGzp8kpky43sPrU7gA+3nen6zVxzUomV/tg1sZwEn8yxd0x7NLdsn/+70N0u
/qEj9VP6KxiaiIbHCJUuASxb5uovW+vOCh/fyys9MX6D/O5yc1ximuRuDlSfm6Bsjc9na+ctB2kf
DrK2/Ni/zMc0YgnbCSCvtu1xntY8f/zT1apZ3+aRCtomxdAQ3XtTCdVgMYiMwSGD/YFsJPQgCb4Y
t0qfcc/nVQeLw9tPIlgG0t9kORWZ2nPkGWwT7MhrGRrz8a3gYZPfB5AfA3BlZQZb9B/izVQ8LR/b
7H9bEDFL+UfTaJEBd5gZ1gQ35Qs9e/jn5nJq9BMzNHeKXUFtiRgZw1A2KMEMwj9giFpB5mMmCO4T
Eadp65j2OlBg7g5MFac0Ic9UhOPZrcjIGYiK2V5ufXmZkK7z15YqzNUZomKdHGdsKM+S4jzL6aSf
+keIj66Vkt2jWqLKDuu47Q4Uchv8RAChWxvCvPQ6R7zFJ0vs72eFnRo2SXoikTY9UbCusaBXeF/n
YfBjfHwArkDMrH8tRuMJUtPFV/3SIiKo0WlDrWKFDh0IXpK126oc0G9+FlWcT8nXx9Wm8bcYB7h+
ohWts2XmEwvA+hMy9/LuoyHM3I9l77VupeUatz2gGxkq5FszWIbkgFEOplW5+EeabgKL3HEjOejl
RFEBb0tqjPeEQsD62KBfn7XaiXpLmiaGzSh4Rb3dE8FiLNNwcHiTCNTSLAhqeS7VvKNsmIKutrTZ
5TaZdtZFAf4h0RrdOMn0JfL0C+PTHshjFMWUHlKfFr5cdUfdR9/WgsFvO2jULpUSIiKN8EYFHixr
/YFNO6ai5f767+nt6l2fnX09/po6o1MAXtBmPPz23rJ5lkSok6Fm3N//U/IV4qxDZPkSiIEZ5nlO
VLtOAg/em7ehOl3DiS93M+DpCifWhgOVNKEM0P0UTiAQoRLvHfXEY0jZEcTnh8s7ok1RQIXMXNCw
Me/w0ji/SmxZLGQlNGIaU/XNNSQSR9BTxaw5yUA+rQjYlekqmLcvJChv3qMiztvDBNlaMb6yQTSl
pwWMJmRSAvolWQk2rrWfvWFqaLGXCsNgUJY3zmRhqClvdd9DNFpUNVXQEF1b1zndRQy14Ot/dnr9
TK+jlYlRd3jKEcl3Jrt6MVxl7ZP0KJ3y2aIZRVmL98/bBWxTDt6RyTsMTeNGq2Ol7hTvVb7lj2xu
0FDlAnJ7VzrjRDy2gHGbTxw2sW6Q/p3OPj0vvo8qqpD+UWbWLI53K8BLNAbgq6wJg28/d16b/xeB
JRzzBTKLfN5Xw1RDqYy7DqUABLtXtDqnSHjOH6/ZD711+PW4Xk+sXnu05qnYUV+cpQ0P8Y5dLFVJ
AYgvRRd0SsfS6RTOXWfzHD5yGQswlTo+g9qpPM9G5SYdlnPb0U0EQyLfQFAUAdyuyHHmjY01yDdD
7NOSxnO73i0vPgYcIpyjM9nJMAelWbLZyb8QRJ3hrNYJnMUAKI1AgzO3moIJT2qp7ZEpgV+itTcw
QYfFjnMSEigjI53cpnIY05x1Or2BrNLGtzJ/mGRgK+u+sLfy1zxSQc1TuDLhmn+huSy7Q3YQZZ9I
eCaf4przOeGaDyh3UZhd58DwUskg++vO6IdhFTIdsKOBt3gm9LbkHdRA3E8Ata73+JjPDMiH6Lc5
3gfsT0gEI8fqyJxD2ad0S/LrIQ4Ixi1J4wLpaZVQ3DZ0CTSWQIyZpxK0TTpE1HHQhx8AOBXmefVV
S1QSpl//cDuRCkLS/bU2qaFg0wfs19fC3/YorsCvjBj0xPdPv4f722YQrRBGAV8Rnx01K2pHxlY7
AN70h/jVB4cnePsNNePWegg9s+fFOLiokWz+KVi1d8156yuR1Nu+23tjz+7o4+QNP53Zk6RrA6og
Oiy2wWqPK3asASV1J6J3sZbYBi0p2ZvRFfn53CtJLPOqYT3Q6Ja9rqMhsef6CAfFMLoLc9P8LZf/
6KaWkRyPi5pJBCnH82MErbf6KWsimNkjxRMNpBNMxrIbAshL/D/k2GNDOmnyslCGurSur0GP8SBp
aUXuABzSuW1bwgzjMaBHXdNjXJ2aXaXrIsulc3ErUsCNyfwL56svFe7pBR73pAIbykhNXydCncoi
etU1D6v1oZG622LG2OhvZuS0xbHBz5KA10B93kmmiwizx7v/uqGiKtKz9fz8aSx1nWy/ebVYKKS8
Y7x7vOurlTv5LPbPvrG4A78nLtWwbycIGl18HMCZC0lcw6TrNOM5LQwL/quQQgbqyJ8Q4n/K7OMY
F1piyTwV5UYQ0Udl9aC/Dhm4u+04A8VDVXu6yl5p4oiLWJAMpBiGgfoknOvTn2iTjVx/G9/NTp3l
Fw3iS9Z5G449FhS76Z//Y2AdIfniv11BhEJDnjVY3VfKTC5pKaTJJyHBcjpqPp/6Qp6DJy2y04XB
l6T+EJpgqrtafSwTKo4B4ZFV3IuNHEvIHflrHr+g/RFl+j/U6ZfCL9DRWJW1dJZbDkP4KxlO8bY5
/mrLtrhxfZkJmeZ+u9fnmKnw1gA5OIOs53JPw1ZLby5oypEyDuw5BFuml/XzOKVu5bC/s/Ov3QTv
TgZjvUvh92qL4QZ1Z/GTkw6LDp48yBE66qO81QJHcgY9sZS1liuLFNX+hOlIx3FBLEBIDVtJam0N
ewrDqM/9yOQFMMvUY0qgLzGHPDTkef7JitNCvx48Md9/w7dqIn1PZ2kdF6uY02QKUh7EzlkubmUk
04dlhQLe+X3rUdynRoyXc6ivqldWfY2YROvB1V3Z1UtHSEW++zJAalDm6Sru1+qRUykJO0hM/d4U
HlhjJjY872IxvXEXtGSo504Hi6Yu9hsqc8/z5mBVOCYq2FnEvWdhizNwyI7QNXlWc6hyB2HpxL8Q
nC/iL4j4SWqsQUL27X09+S4EpoZGh+jFV/F/XWytW7yLY/fLXVJBujbYJO4317laYkYjPln0TCYk
6+UVkOEYGhvFf5rjZCQyVHsXQLsFW22n5MaqF2zCp9Jl6R9gapRkzz3cUe8+zEH12KqlVV2I7pZL
pH1jQYBgDEitw001u6vlOiZ0eD24R8JCigLlQ30m/IBg+qy2mSqtETomO4ywaMYhLuvdg0u9jBcV
+ZABmtzsy7ZHieTm4UDmj3fP5wsOGx554GrHFheED8RudQ+944jAfpyyPmF1WC6PHoAsDS2OgRQp
XKurXG+SPLhdQgKX9a3MiXxvNyq3DYKED//gAjkMYoAPHHv0ppO6gh2gIkF+fZOJPKAIK/vRKKwA
h2z6ZsH0A6AtucsL0fuT3S0s5MHMMisdyONzIfv+VRN1FiMKt/paBMBgpXNCFPmTMb+OEcGLWMKX
V5LRlgp8Q+c8/N2qqLwEl2XWVIdE98KBvR5aiTd6I/OQZjzcx/6j9OLJTaZlD5ZB76lvpGLWroiK
OTGPOEvO2PwgVxwjcSADuHG4F3X/+OJ7g/66BAtnSaEdJeTM2dwLF4/j1dbyMr5SqfZTomAAFQvt
s7fgeLkPSfadtOaX97fxkqNbaTouudcoG/xCFgbV9KaFVYVaptpXwnvsJsTR6UEWQ89u7u8yPH60
jBR81tKh8ivlHorUSPit0d7oJMBPmUampxkbc6uZjKtfjckYfe5TQssw2ZqI/DH9MhgCjScIMO6f
dO+Vzx0TW+zEy+6lQHZ3BjcgCp9/xRGwWiMh46aEB3vWQ7DwxVmCtuaEqbtSgJYrxQfKAIP7v/V/
9hC2L1RUnjZOLZqREvnavuH0FV3mq/wLOpviiTV8Zg/97GD1B75aahW35LpDaUe6AoAHuoN+hou+
C+PvIxjvFabF62d6tU5WziEfQgrYUYia7KSgaMn3ixKkZUQMW1yM/73paKVXNfGoGcEMpk1zvhuN
WvKZfpAOkMt+MqEkm3TnVBByMjQbs2weVe0u3Wzu6lBXR2i3ZMwsue9YIBANTWhfoXiljjXWcCgy
i8rpurrX8ay8E2royFL7VrTb5DiixC0bEoltkbYgS0W/qt1qnciwWTI7AOntW1/hCpwEtvkzChiD
dTUswHWD0DXqPrjViC4TGQ8GsoH60sbQ8rxdNs9qS9xzHOzXXy5k2zyS+npUGWkEoWu7RPUdljAR
d/lgC9u/OeRTm5aA9iOguh9VK59OfWydlOqazNSMQuA8wwfOJaNc389X2DONlmLC/M32So4UQRSo
xObU0erLaKY5jAnpoGpdf6N/Td6lldud8QX1bSECJ6AYA9eXCZCkgtqM2b9yMVfVsuPqtKI8+hbJ
/Loai8MxVmCm9vTUk7mNGi0J22IFv86FV7MNZBGU9jJSDYhwhzUhPvghjfW/f1VfW6ttD8ulO7K5
Opa7VLm4Vm9Asn0Cv+JPWzreJ3e1/NeV5CsclrpOKcCsAE5Gx+lTXGeyGvgEXlDH3J5Cr1PeMRky
JkZhbxn7txTEJ82ltYFBt2/qaitPZiH1PuYxOqOhyxW/FN9E7JDwOZI3hjeX5R7uF4mTaad1CT3Q
+1IVzH1LtXAlrynJYM770yJ1yPhgFAvX9C9r49C8HXUISFcQsVxHTmlb547uRvAGhUGCDO6XtGJc
bY358Ln94y1TCmx0Wn4j4JAmy04leQ4a5X/E6gmteIUgSiKznmU6oZEOugl36lgSLVsDGJr+Tu+R
pV1psQIMiByAzY6a+OBjPtQ3XkDAm5MubdRe+sWUPCKVfrnDyv1FlO61qjqG6DUYnumdEUmAhgMw
tAy4xSrFR/xIYefzI9S+66XxXtWP/QgzIjhy/hK6KY9RGDh8GCDA6GNsxNVYNPBAu8dS6h/J09zZ
uslwlpxYnm3tZpcy9Q1Gn5XFdaT3FIZTx0NqSSTP6URrktUDIRJNef06RAKlRR4mCclmCp0VE9Jq
PlZhLEuyH1Dx7Cg+jtzEMbs+CMRnrPRcNbaEYFTSvEl5ScSR6/B0OnGV47Z+iUW4stFjAwhFJAAL
5nEfOYjxfW0HvnqLPmFJgEx50RjxZnCmnj8cHI39Cmi7SeS1nrg+8FyOmQX5H8/OknURQ1NZITMl
gj/z9htri68vryPOodVcAIi/EnoOSZy5ry8dT2hnZLaoZ0/jHeJ2sBKxdZ2Zf7Lb0Qn7g7pW6Vty
/Gx6YxCDNBMoKsLcAdSLYOqCIWgDEknbgAVlI2RTAmYfcFVKxFbKOn5Eq6RQ+OXAt2oRhLY8a4+0
/qJn0worN78r+4WhEFZgNqEqXNPxp5Gb/uwQw6SgIftYHS3xlL5Y1V84zJCjO312V/qPTw/39hqF
fl9wxsKrhEAfIHi8+rcKQEZUaTrIN956PXFkugngjwANfV/dnCz1vIzcy/BJlh9Ff7Swc0zgi5Cz
14ghD8XDzDEKXKBMmAptHuT3vhaiHzUx6DdLcGMHMvHr7tgZ7ho6hW97/3kys2q4MGa6UAtV+bnO
gfymz9HUgCcXEHXPGNZg5wl7P8DBYMTIf9RJJWxVHiyqlz9DBks2mYWeg1a2bck1xZ0P4QoHRNBf
jRb0FKxd1aJ2OS260112cWLQSUcFOpD2zYtCj/O4H1xE1qVc4m05bvy3sy5UHz08HaTdyEh07AJg
Y5cdM+xEhoVBctLfdqXuaroI4zpGj+XwHI2ALLGf73jV8sYVyLd++k+uWfUupEM73/jYymUn2t3N
kaaZzS7wr5iKtlwNj9Ptk1MuW3wlNw6UGK9QY7de5MjLHsoPZydw0mZLNLCsXq80nCIOEq7rKCos
SUqh9Yb1PtharVu20BDyC+40gFNo6DWj6ayHilCWtbKOkPpVduQ4KLb4CZNDy3GV0Ahbpo9ZmHgt
c+776SJq0ofpABaOmpDu4b7m0gc9QWfTjgCe/8VYXbKrnKaH97FpMXee8kobX+hrc6hy2AjoG0Tc
tBok7r0Y2FqysRHDRdyc/2yNPVlMgSOXax469MzkMzAc+VV77tx8C8JhskaaVEG3wDvivqSKvXfE
pF22cuzBgERb4eF7iJvcU/+vZnbylOVd+B3NHOYs/1Z2Mzyf8+fVc3h691F8vqt/Vul8NnTVgOwb
uTx9v1DfPwkSdB8ICqY76/Wed7nUI8+1W5ihDpbHXg1N9XF8ZpIA3xZWCxgNy7YF7l6dLKe2mbGH
f5+jCZaiUI4ypCxE8vgrM4wrK0i6EgQ4u2NCqhoh9+jIauXovs04iRjWdbUczWtV6Flq0QXckCnR
P+qRU/ki5RHBxYZ4qXnJiAaPdQzO+t7boaRLVV+T3lTJ0fgrPNq4/vSKdYMpVEopQ2DLHbehtbxP
+1zkpvEtyXwDDkOCnMAcRGhLEWhMXGoYpENTa40qC4hR9VNUh0lc9PDrhPwu/rQp/aj/LbleT53R
yBFr56Qu6aS+g/+391vSyrfCvqUCgJyay89RMWKokDRDhr67I/pKDoDQAheGzVFYtH4uqVwQxuoJ
vdOdV0NbSyN0hlJWfgZzEeinXsGdZJIAoyviaqr3TtHS0Cvw9uyHPXJHTo7j7N2DhkcXp9zDno1Y
/9knxB0SeppN8U9dZfxLKy3oIEAkH7VCl9OKiAwk0+9+GSj9MqNOFsum2pkeHDMGvGZ+gewwAw+9
9ZP8+G1+/x7pmsRi0XlhQhDmazrrYM2NlLyUiZLFP0p6eIUMDaU3P1F1Myq480Sk9WE5ks+6jmwK
JxSyirKgEy7pqFRkBzV5MgppaYyIFTUZskbcPGjAj0YuJ9drxrNoNLZvA1wzraVesteXMhIvhTdl
oGeHg2cfjsVBYVGSX/JEH8mFhrV3jMK2gfLGmn7l2EiyKbW0ZSZzaiLCwkAaYtY5nrQolDLO7Tvx
rQgYiP4NA93qXQKLrFqLOy+C0fRzrxH72zd839o4AEZe+9l/PJs6wUxJ0tufIF3BWzJxR65x2Atg
66RA7IFOBmPMs0+RqhZxPWBAEmno4fDjTJbfbYPKyq+yQY2CoyOZroNa9Ppi+Gm5weedyaFt8CQZ
TmAvI2wjQFHalsmHpsr9g89r+mlLS36oyHTbwPUXwd1WzcC4BCtfkJt/ddadgObkHO8iQNMdXdNt
8q5BwuxE3+QpgZY6yDDRiyKyC6WmnN7efUa4mukJsEoDt6uGw/b24hsAUiiMuWiiXtw2KJfhbN9d
SQJ+JV3tZ97A3A6pzxJWtyLTq3pIEfB9zXbIKQAhd9DfIsDi1X4b0v/IJ0hsEfgyLlx6xeyg8Tow
fOu2UE5q/UUPTduK2iAilEoIl9S5ZfbIMJb3UU4shJgoK4URn4bbyl83dF38sVFYOnaFM7kCpMn/
ejfqCxBKjhniBK7VbvUvrHZEHC0QsBazOZyBTSx6hTOmxxw6s6RKtI2UnU44OUwqcnvMYgcTVde1
qCKrZ4JzkTnLOaLD5uIzFCK/NiR0tXJcXDiQ5A2MbWt+jkyghEZvahSOjQvW4lTtMHfOogdwVntg
LAUBZl2cz/b9E2Joskh1W6xPz04KMOEqn8PFaKSezGZ9wQwYdl2bL8WcfvL2HrLed2tgaTm7DodJ
1OooghVs2Ia3bCq6dELPPwxrQBXbUCQ9qgRXP/6ZPMi5NxJimcT1di8GIcRytomvMUCt1P1GJAbF
bS3VcDtTOhMgYrC3VyogBz2dJ3d6OumOFKchNrRjUr3CczsBrllUwsK/UE471zr4HGY5FCwK/8MT
PpmJ5shqkqruNL4gAl2ohJa+Yp7K+c1u8hcbXr2QSB0gGxW7bDNEohksZttD2CgRvWp21df7aQVI
TufvATEMDK5l1+cAf1quOD3cL2zUj39M1b/hEf5E4IUkOy8wta61fqnDVEO8cHhTaH1Hcp0jARbk
YNoYa3PKwJfXdrkMWZvavtpASswaFDpaj9Mbm1gCV2qdAA6MsudRrdVJdyil+eQMxDsI207f7Bog
+ETq20YcYohmFLko45xQXE9ikY7Zv9ATz7ZtX1sfmpT4uK98L5whOweu8KwbgHzmFIgvztLay2xr
maxeHPusnfEmovMB3TefJcye9RqwjEFScyEqzjd4gOSkJyRvWeN/x/cSrgN5TY7ZQVSgqK1qMyla
+V4kd3L8+FnqZaSolhMTev+jPFavFB7mUS+gZZu1noYDCm68LIDUXDb9BLper5SzLC7rCrYNvTYV
jUjzyvsY/pVkraNMybekFuMD3AIo5UX3uKDUalhKOSqldO8uBe7xX/QK/8qS6u5Sij1D86DOqvyX
bsTblun1V1PBjJo/Ha+0/2dgM9FI7XCuscYPmeKHoG6oZ7g9cZvGUOlStQAQvMxtfib20cdLmAfF
QELkSSLOq6updTqrLDkfgjHlD8aX62nGHlWlBz7Sxof99w1Std81Wpbiq546jALT7AOwbM/9MEV+
fjSzpLWafSChan0iA/hvBPXlXuc99+XyHXcGoPFIzyvsKM6hTZkr4QuqHGMwK8AUvlRbPFQpAeAR
ZbUUzub01PsOi4SXVZsZXCltxXLBGtStA1jDGo7zCLQ7LAuPQGESFr0hzCbu/asjuvGMFzUIYUMj
2iN5CrxDDjPI8nvYIQKRB1UjEMIN+yCeROcYu/vnlkRDsHqc8583K2bu31lGo+ofOOw7w4g79zYd
nGJLFw+0qrT9YbTRfIgRmhtIY7hnjasiPnI03TOtBwN1ish/KFQHYxksj6hxuOHzhN/1G2WxSLMs
S0bKJf5yGjIJKcblucbx8qktdfS/mbWqGZIjsYipih0cTO0ZprG/SCyBhmN5wZSUOfHYrtnTPZrz
hajQZlqq6u8sVS5ercDO/m+nlOanpGq5innejtH/0iv/w6DAaxBNjNpTuoFk5hUnLWPycuH/dBpg
BOe+jYAB9mHCtTPLXWUYGNGcR7W7MW+LxIe89vmclucJxj1xtlaAxoXADHYWfVZ8I5XuUs9ogu4m
F5XKAChGuEBXPRd+urE6XtK6ni8hvBoIYT/i00guEGqFHhbLylCkRLfmvO177DS4er0WglaXr8eI
Gs/58gjZ7gT1ZcUdZ7RElpMhcIuARLrNnVRS6qUvzYeRb3agQRQWHAKq9+so/SPLZNxNocTB2IXr
2otdWE2TtNQvezxndnJS3Cm50nk7SVtbVfUT1Zb/W73RrD8Opgl9VpKreM6SnV2CQlPZoBLmhUXk
P5QiXp7NAqZQt2Rnmkeempp588C6qpss0cUFQ45fATZHzuy5nFd1iQVChRE+od/2ytVzDEPtA+zE
Dgguh1GFFMVHz/gIZF37ZA4b6E0N+2kgvR+qc/GXXU04t/7wA8PyL7AJaEBt/bLHByN+S5ongtle
MMHrwpokp9AQozLkRy+y9wc4BrD+XngRYiPAhAAHigjdkCc9fmcUz1/qnHjI8R/+iw+H1cd7BM/p
JkmpQJwUZuhn63VHBRhD++W9uewsUBPHUzl4q6zOqBBeobFk7Cn29BFLPvja663wh0evzdA3h+MB
VV9XwvNowJ3lnF0yLjtkXY94tlmO63ts3NijpoboByQAQhtYc3DScf74d7qMyJEJWfZH316uivuG
qXwxIh/8H/eedA2Jv7m98c7BanIk36IoANTeYEA7JDnnyiTp6PcHkiC1eDhocEDmnEKwT2oZkqvp
za7siLyJB4e4BHVHCi5CEmPeFhEe7D/CXoDCfTD8NK2M+rt53bkRgDnnka+m1y6vwb4AAIfGA2Dj
wdCQgfiFpAyk9V/nmXaVCjuszYyANO9e0UhMOBO+A5sq6EpxKFvIr0XRSo9X6WFRTtLpBK6ouUht
d9lv7ONfjtVymaoqSdww3Fqh0nm1zwlwD052bacek/aIkrZtPl83tVo0oHTeX9Zo+IhdrtGQxKIO
TXhnfRJHV+yz4O8V9wNKxIlWTPykhCBCpFck+bpn238Gj1SL6x+GMkN5X89uvYSWWpAuETogMSHw
HcW1F89auOZDiTgdB7S8CqvSg76HxbvBUE4M+aYQuWfUg0sMTKvR5SNhkHJ5Y2ZSu3f9hMwH+Omd
lN8KKsVDk4xGq0ehE+g0StwkCVXUea1QAhp1h0etALOCet0E7ervqj3oThxcic3LK+GucvGFsTRt
twT7dEXKUTPg8aUwD3cDXNXy/duaYc5P08Uq/c3ZCTR+/Acj250uMfJMQ7svic9qqD0x8vX790WR
JBg1QMdI8EtPSJUVqjJQtoBmX6HbS/bJLFoIRkXcKngc/DyNDpWQGcoXEJV/lTEPTZ0eKHaCtmHQ
HRSs6808uXs+bDU5jw2u/S5vvb5IJXJqx2LpBVTidKVz8+lRHdoA3z0Ai/FEifE93zOjUVpwYxTe
J2Sf2RHMiMbehhNC/e+ekmkS/YDlAcAx/jfGq+y5T/H22Z+MxOdfOiyPkmbKTFie1VqDLpYQKWsF
5GyPoNSwn/72JlOrTXZEQeYS+1mh82Qx4dmgjx8F0FlWT4wdRqsb7VWUWgY0t6GQ5zt2i8jHeWf7
o06DnWHrYSUBbyj8rCuVauwe01Lj7AcTGa77ZkPY2fUmBWTnEQQIvBpm1kb0tc1WaFLv64QIYwEh
UepmGuBj57CKsLT4JQQPyTxwBE0f7uKiNdI4k2ZhBjKAbk8namjjBLMVNIMsHTke/MpJj1UuGFcD
qZ1Xy/acxN5ESGrpZAQj/sFRvigT9/Vh2f58WzfKpAf2GX2PZYdjjEMwf4bIlz5DAfuqmGnMnzTs
lG0//3VHpRMQ7w7C44h5KyJUzFFLSiSr1QlojV6HOhELznL+x4FeVJIlF9qzAHBWzdSXwbX73IQs
5JX6KkBoVwhRfP0HG3ODCbdQdDQgsun3SeyF78okR8mrpyRRzJmkIKDu6KymwFNSfFPuDLzxS/He
+AYwj6H1QwRugtFlmm/h0jAazwqYachwqGsFgbDxc90Ssjh57i9GZfdWUDX9qjtVTdUF/0nIrZPD
rkNWfvAdWW22TeNJXGNADqdbA6b10li6ltu37BMNeaItTEf/XQUxstLDAJhu1mXEwawaRTNqYpKH
fNlrQM28lDvL9x4OsNXeipvgsImlLLbc6TXpWdhL0EZYia8JQE8tqTnewy2bsG3KBeDh/HXXv9lu
lADYz/re/E9fL58dSxEAjlmFNi1aPtbWjcOpUTOSvyage84t7OerfDPz3p9luppBVXFg60tO0yYL
HOeeubFV5gPUFnjT0x6HvXhsfPsRTGf5hjB5Ey36MOm5KGaUiX/XdQ7lGfT1BhqShhwY+TdDmIJ5
pwjc+D1b3dH59mLYDK3d7X/hWXRmJhCKLLbzO584gVZFgLXCd1s1iir1rF1kOZZmf3dx6hFqm9Ti
TSqBENN3nOc9rX+77AFlJZYHM2ielPaYPGTneplRoozZIq69Eq9GuXlh1oz+EBgATa0fQLADrB+l
jlfxiWG03FQ2gghoupFVEX5P50cJtqCPw2t+tSF5r9ISJd4QnqeJyob8aMyidw/EZCpPSZi9UyQx
TihK9hbmHsx2okjX30AD7EAYwXtuNoFP1EBn9gLF5+mBhCw1j6FzJYQaGY+JFoomYOWXDi4q+38j
CgPuFEVRB7IqHHUgslo0csk0y22RvR1zy0cWLIrbbOrxJMIHBtlTNVIOD9wxW/KV4ilKqKyM5xdb
UYyJv2R57Cj1gbPgswIBZ/jxklViSTBLXxkvOcJIpl6pGb+P9fJ47he4lWwoUDyWaeEA5CMptjpL
YNgbrCFpa7zYU7EBh5WGSVhWbdFCSeuSDEYG376mJ5iJgov4cC++suWNrOC0SQXPPlQcsSLxsE2k
Orkv6Gx3ILqmlPiYfg5dcY5N8TT6GkSLocNiIPnml35dfOHyfOzKL+EKXP6XsYCVUd2TRa2+3VX5
SdKgmI2DFxyoLfI1BXceUMP/58UJJFAemmTZh5zYJIb8gK1gABdOd8Q/9X4XTnSUdb9LKl/YbOF7
ReX6i5Q/Ds57rplOmMrAMwlRGSjTP9GCd5RoKHcKit0WjVMb3aefBTaOL/dGx+PF7gLylOF8kBQp
8mEET4nkj9O/LQtNXJO5HcKl608eOLMta5Uc+BIQihuL23QJgzZ1aT3nqz3StlueeZ8Ny5A1koaU
H6NhaPk2r0LhqwPK9ZkWyjCrVdA62W2C44Za/TVBuWBr35rfWd7CKcqsmqWv18qeXtT9UXJ1CE9V
Lc4HlVxeWQQI8a1qeEiu7n55GGP/O3GcmJPWg9toyZiMOzXltqwYvNG57cl7K/UC4bA+e2i0fvgn
majH04xDRN5eTJhGZH6/Lr5vDPOpNzrUJWkYpwTqJxCHstmf+mgYUIApn7SZy0LWarwOROZUfJ5t
uc+gtZJAGtKGv0LySVLCqUP8efqy4sGpG82Rr3szgVolZWSLENOv4hr+jBk/xEwb6hxWkq5WU93L
mVcfR4MzJ8FU6Lor84byMI4k51QLSo8I5vT6Iw9G61fR4VzW9/ja3oprm2rdAuEwU3W//h4mIIef
r7uHakeCeX/14fF+ZjDit3rYegoHOfUo+l1mIO9+Zpkdi+ZzNf8vaZ5KrQpR3ug5TBdTmYsAKOmS
hDMmmAPGnvlHlFE8dUsAtixBQMl8cTKyaNkn8XVKRDVDc+RDtI5yju0h3Z5QteXerw7s/O3Q1xpa
aSUjGf3xsJCXJiz6VewZXq5wc6TLiVohrbC7QWiTRsuFucXoqhmrhNr+1nY+ucN/WuGsy2wHQ4ij
BvfkBJoCdBg73V8gTw1Z5BGx8AvoZ4rw1sCsIXG2D2Ag/FPm42978UZ+qf423vBHqitb0yhKowzV
TsLlne5qMP82eecPj9j5U+rQh6I6r498pF0JfMwFwJlJLCK0/BG+zum8/uVDvgA+1v49F+eqsgRN
PwZLW9kgHJ0i7ba0gDCJJGI7TWqr6R/NDv93vrWLFsjQb72KAA0uOTKWAxbnCoYl6Hmd0MZqW+LV
X5W4wbUyr5hVV6JNhk24/RvrLfNsbYor06irDMQmg5R4h/4AeFPkNsBRm75HeOu9LuJvuXZ7XnFi
VVWYSJ/eWLKNLFimyY/DJ/dE0AmiHP3Sk8RlP9hCEPHBIp8Dw0vfNtc8mrmmVhg0K0wl7RFvi4C0
B5BAadhox1kKPeWOhcRbKLRBFXaYOjqvPSDqTWN3KhzhS4EELlEbixa9qWx5FYjExcQmgTJYC2LJ
xqRmZ+Ult9XdQ6udYoFa/9DZjzjOu1NkVR8DH2YXzU+OZMksXyr7zDTpbOO0qKQ2TxjpYvgquxbE
cAOv7So/3DFQ1M8A7Na52KgmNJNcwZujJMG9BXT6iaaxy5ye8PYQL8nR204uLFXcgudHorPc5qXF
GNYPmJTmnBnBoIShOnqiDYSUKsP+Ae78RSyDhTHaYiZ31HjIfa+jPCONVJtzOE6hszjfktQj1D5K
9vaD8SrLnEorITdIrz1e4/Q/gDD7NPtsaMGMTZ8wbgBxUc58OfVeTOFmuySKMVXYaHxo9LVC8s+1
9Ac359VBu6Fu+nIrSVGGU8rlHnBfyboiahcJgEgDso/sbvWov5xq1f7nD2ZDwcwiJK/FRbHg8GvM
QZZJrolo6YpT3hNxJoPrTVuNYt/hfNF321KkA2AghFhYVfy6Q06L3WibKbXhXl+Dh1fsikcr0Tw1
S2JRl0egYmzfM03TdPQGcQNcNB5nTvvO40Ab4Y4q+u7wccGOjWpF7U+J9bK8e613DbiX6TMAxpLH
fk4qye+Z35M4wHOva85o/BPs80HwvFqyFDd+5X+JSdsmU99I7EZsczNyb4BQdi4HE7tZ3V+dBfBM
7T/NAgb1pxHN3UwsuXPk/Fx9rsw6TpenYI3ix/mGTG5zyNacxRlDD3LfJ/EGsPP7hntVUYImr6W7
oT7jWmvmE0AJ2c9c390GltQc39ZqEp9xfbaZ9ntV/UaMAEZniPEKA5YC9eQV18FOthfhQn/Nkpz0
k2NEa1CQTtIo0186+y6TwEZ2Py9AZjP1zNq3DbPrxH9krpp31br+A7e/05l6NkDThlNUkMKulvTx
zXsTKADb21rUT4Ro9yB2uS4UJJ2aAs9JLd0jypdG1qFBNlf6IEg3O2r9SzeH0AArCa6T/YSZh9Uj
3MgOxZ6sMLINbotBzvD52DDYaVWFXtRFBDpdEw3e8Nr4ofTG+sWNHm/4ZUIY4PPu3gXtleLTdpI4
BhZUAFZPixp92pd5fu9zaEykLUPMFX69A3kMZhKXIk8OVHGY1MV9I+NzsRN3s+iULawk5dBRxhBi
CXRiojJVkGmkgMrv7IdZ/qegFFmJ5wJjkrBr1co9s6tweZ5JR0AP5iHr4v2PETum+5e78OJ3CRAi
46nd/cv5mWyF2cqTAewLK7fu7SyoHUQquRZN0TthxS5MV8bdk6NuccU/2u/shZgUOG85b6hxaNKT
HTy4gz5rtKIP7Y6S/tnNfcH2M2m3J0S9r6nbW963qYyaxnsDQ63nvRDopEiWafEbKXE6h0L0GTVl
TlFbITVmNr8MtY+BgG5gJazSUQ7jZVxCLjS5LdAs4BSYh3HM3dcn+/qsEp9c9RWlFjMRo+8FPyIR
I1LySRrJFUaY525V5u5Ki0vMcvvUNooAz0S2GIP04YqrSgaskdyB9RExmVPz21R/1mt+RhHnxol4
fiwqu0C9F/4jljszEGvGYsUCQlM6s2y4cpLOmBMHBFO9kD3pDmg/QO8Q7lTX5EBHA6ltzwDIlmCI
V+9pYljeqKVWkRgJkL0c1sNbL7mPJIfd8kacS04OsKyKwRQYvl7khsueNd5iZnB0a4Y3q2ghD8qL
8boZ9cxkw37Jwrl6gXKcliJcMb3MPqh2jT4w+DmZHqGoB0OLxOvs8g/ybcGvybPjFZhCc+PkXwNq
RZ4VODnefHHACnwHjYx8xnxb3EmsVkDOJoMDmkDYcVL9FQXElLMJq9RaIbFJ7GizN1mpUG0t7QkK
sXRh73LochJWTNdZG6DTxnTNtyYLopCnIrpEUdId8183QEzW0MfB0n9oLmzi28SgYQNKTNQMbmsZ
qz6y2PdLdFKHYmw+aP5vqT5oLTVb8utkhZzQs85b5span6w6FV4ou4I88D/bs5XUUYEc328t1Em1
EGDHlJ7BHTFNDvYwEgZ1n/+iv7h+wxkr0+zdykp3GKHKADD/iIghbt5whfsDphHZEEhG6daZQ75Z
fL0BGFh6KwT14g1SdA9B58Ft0Jv6NSMt2Yy18jETb1zrwXSs/3y1cHqNl4uUmsF5/Z6Ww1hX4MQr
5QHpc9kkNsV89Xtyxv68QRboB6kwiXB9IsK1TcFbxJ8NTUbOfwf9t4eR8epKA3Oi+ATeY+rGOXLb
ETK5w40sVNgP/ISmtn0kdpdkjOBF2C7gmjWQq7mxJcpxLFVUQSzN0qKWI/xHVHoqObXwTvzuMmOH
ZTIsJ5kWuSjDqjR8YaLaFp9zjb3azFEVBAD+eNb5fThs1cCkXEAXU1/yBqSYPkzX5xhkNFeyCIjf
EiTOBo/IRCTeb1w5q/ts2LUpdJzpnOht2rQAEbD6WqPvOEhjE1PdDnyxdil7fWntULF3JlGl/yuO
tIXb2iu1z8x4kK7Ic57jDINYAhC73ZNNV+NNgiHeM4jDe836HU04gy+UY6MTocIBWSo6uPOabrkD
myVqqkHsDDyL/+EkJuBRiKCTlSJuikyYv3SIZ0jt3ymzWzKHVfDXvRSgu433tmyOdJRb48Jm/Udi
s+yBzGYoUEbUuIXrtNOm26XRl4DLpeD4jJZZUCl+TDesWirCgkiiKYszpsx2OY6R7kypDsMQqZaJ
Zpfzr+GFnzcZWPNpy0aWz1RQXdFOW0btb41MSK0yu8lA5P1tdphgBpy3Uyh3Mi7mfeEPxIzJJSCz
Mst64KeZd6RvQP/j2+XXPiIZdkAOT3l9Wk7AIQuaRpZJegQO/eNFXVrA8snJvzfH0cILEn+g8HAj
sdmWIkgaT8HWVg2G0fQsmBJT9tmSJ3iJidfhlbDbbzAC3QghpyqgCncQt6RNQaDE2bJID5dfSANc
kkuTTIYBivy6jlLsoyuG7ShwzSJ/QNrJXhHjZbjD7rtTMvJCH/cyf+a5sShcmMuk/DYEaznZUp8r
AGCFDGP3WKO1XZJ8i8xk2eayHy34EUArKfG6mBrhkIPzQ4FmOMc9+80FySeV7vq1UsAD3hvIW3nC
D1TotOkS5QYSoLQE75vLSyIP8E7VR1eyiZRtQ1hcH98C3hgoySd0glzGxV4gRbChH7YvW1NqNEQA
jWyVxGr0QyDZYOhXTnIcsducAd+pHPEWa+pBaWLOqEwC/1Fh7C4Vo9fJsoJ7GC+Cg5GTkmnnYNv1
Sm3SwNvIG0cRgqMNDtJc/kPo/OUftIJycBTlgUZU7Im+VAZnjokQcOset3RJGyXqLsrzKAtn4CY4
VCOadpMe/GY35/mz6IkonJ6AnVHN3raTznqwxGQViE4GVRBz+ziLjRPZ589H/tiPW+vc6xRmAkQA
DMy+yagoN4Zrh2FRs2MEH0RzBC10Z8MfltBbxNJ6q2eATH1G9XuMAXq6Pxfoy4BhWV6jEgaMbNYG
J5SW3Y0bwCFvzJoadYt/cFu3Qr4ROSWUMtk0Fb5GeskN+U4pXkx5LnwqkiC8SMbm5ZRtgKzkaPst
wF42atk61KZMzOH9FFq+8E+rqmwowtQN+cCrSPjK3at4yEOyTCeXsAgM6eBve1QCknuoUN3jEWMM
bNHrAg6L/IaV3nBncfc794KAJnjfYmwzcPx2FDSuirNWZEHMIVogqDieMC6CnO3gMw2yCej5nlBQ
Tjo8w9m11Kb6B6+h5V5Y0KJxgdd0HWwznSErAmGZ7L2NHE5ekdVXdEhLuLpvt7U9gN4Z9ev3tqwo
mtGatBojUHSbzJDxK072ybT2J7DlBXPTa/jsH2/AORMlSL1vksvJo7Q2fGUiKiXD0anDVLxg09hG
kkSgYsVUtnxMUAD5ghgEhQrE7CiN52gRbwIks6jGy1UiVjc6NkZ2m7FtFUBT1msbwlFVNa4uHkYU
bFjhn/+0cb2EyGAkn4RsXBpEQ4lqYpscOyq56fgznL/1CtPd4I/vyd0pkpREkERS1QATSCy//EG6
VrpeZc8JMn8hy3ebMUzuYgh+wXEMY8hbitB0DmXYBaZkqu0YqBzCE3D8riiEqxJgE7v7xD1pAtK3
0lQbI6mqSwv1SAqKqbky02OMFiprt9VhnnpVL4RljnhRna4zn08EpI4xJMIrcAFh5519k8hUdT/g
gOMpwwLQNGgiAdzQ7ouR5VU8R0n2sPssnHr3X8mA2uOHh/DG7Blgtwv/HhwBPed/k00kYRzdBlfq
Af4YrA1uNt+JOuAVkD/5vl+kjNJRVeGN1OR1Z+iwh+N45Lhnv+e7zfq3guobSaYxliIZE01NqIsk
MjevoFvmGi66hCzqxnGRReXLNNnKYx17QgvqO/fMOdhpNiyM7sKEZ433yJKpEKciUgKBh6mLs+Hq
1UnDrQF88SsSNO1l775T8Syc8Ooz6IE6deHFyvcFpZ0zyAubfmzlP78IdhYS/GSd67NEmgQ7sStZ
YD/I//vAN/kfsu0+UxW494XqcZZi0TQUIAsplVEFUIIqBl7jscnAm+T1x0c0eWO/5FF2KL300RaB
j/aTx8MCbyj5P9hXQrEoB3DQ2cb+st0abF5MqKTMjKxCP6U4xe8tpIUXKyKvgPuup8skkgJi1oAq
BOMRtBke9rmEJ+7PsV9g7eNyjH0X6InqQltHjjzHLzFn6hqieHpaw1NXMj/tO4viPEb/30HD4KwW
L9E9AOv0d8xOqGR3HDrGPeB2C4Wgh0NVDRE/xjEldqr08ZEkm7ZPmiwTatE4TgE0SA6hUboF7jUi
aqg2W+hz6P86meQyIdxpF8KPavY+iwng3doem5Z9A/PU9uelJO5puRnGH5cjPqBwUgC4Dts3Jpo5
xNhMMHmueflZ0RGMWimnvnLvXtIkDlFPq2+CSbDwb9+JOO+aDEEg2C7pe1V5Twzxt+Ffz6DJ3NZ2
B9xBHq4F+4ZodKg+meHh4wTIhhO5NTwelhm3oUUHqb/yWfogmZCTSAPbTP6QUHdvm7LQ5zPld4jo
uEU/OoXXJ7wLtSIQeE5CSCNl9pw6pk7hG18LGoOQYXDm8yz1PiBxnV2NoPz4E2qOiCr1qil0ywHn
6L0hwAJB6Iz/jGWJ0umnzLMi+bhMbr7Im3k5SxBshfir2wOeT21Cpc9uZTB81Rxaju2aUbWOk50E
qKaC7rHsfuiR9RNfAVTcpiWOYxUrnXbS7hETKIqhw8utYVtKS8+jBT8c5OmgkBR/52V3aj/aKlqs
WePaP5Tw8QXP10D7mTZjdNmBhR5LudpTJzHTLfPCe8Aw+YICZpbi/cYoIwBOHk9PCDECuLW0Gm2M
Bm1kEr93+AKDTnBckYfjFPnd6UIERZZ7LLpIDJCAQ8pivswnHLiA6dTzeBi4mGDIXasaUDZbtucD
bPdOsYOXbEwgyJrZKJPN3V96JWLbmf4qqB/o//hvaRT3l7zq6L/cYB2PafCREo9mDzbP4xfjP/Jd
o2hQL36B8x22+zUCoUmNCmp3PVNDT2WTG3w8v/t+uoW3Ec+40AK7yMTfLgsHFhDbjVHvBoizueCC
57tp3UquVK4peT1YuUcTmIeL8qzVDYjA7SviroF+SuEOn8EhaYKF6bo5Mdzbf9u8QIVO2GwLTZ60
wcP9apLAJQA89YlhtGlsHTzaI6Sy7YJ0qupqos164BHfP6E6SsM8O2XmqcisCUChiRe43Mpbkqip
O7mwA7UI241sGp+kJ9Wv17T0Mgx3ivjYrqhkwkywIYyUvOq13C+kMYLQttlz8ReSOowXsLShd+aQ
Re6FFFrdcpl36pcpaE1cnOl06d0wABFPU73Z+XscjEs7ErTHECn07e0zZaPhmWaViQcB9YZjRdkz
IRIcQYorzLgZ5ZUNemYumOcYUvcaBdY3MwutE/OlzflPBMhTaQWOZtR4u6vhIhlUQbaNhhELy+jg
3DI04MXWnGelRb7ZJpx6XMTLA1qpVEbp48m4DgenN1+MS9Xob6Ftnx2C9X97YEt+lgA9Gy0l1Yws
cOJxkc+SrUGsjoAjmJB8oUEon1YSoZQnvg6ZJzjkQ8lNBHp1pEhoSy0ODjYKZMJr8IEqW+MzkS1H
3S2EqqNJFXzxx7OkKyNf20NtjdtefYR5wA8f4GcgIYJiFudME1QW+wDLznQmOCajGv0qbfm34fhx
1pSsukc8kDTd27X3/hk99wJ2uaJyvrLOXKXiAzmkL+aEhVW203evzK8TGTJ3epWMDg3ZYWa8piTQ
2oFCrsumr0MqcZxwZ5EPH4k/7oyys0YxlDx60W86yDVN/ltlWPvALDiPNH8k6vRqK1w6C3d53rvu
1QVAV/LqiEPNGRle89pQTv9Ls5FxrcQzyI8ku4t3W1OphrUf1fx0GxAR5N41OZxtzhUfRp7FUmKc
HN6gWYIzEU5OUe8bBTTKnOHp8rZ28VdDPrl8+n6Nvpictb/Pk7YQg+6nBofza/oTJlXKOmsu5YXD
CHQkDZOfBctC6WXPN4ft89Eld1s52x1Jdg9E28/X8VucmSoEUqHr2/uy5nCGu3K+1uGSNNa3JaQn
9RfbmsPPZSLBGjWs/U69KS71fbWG0SdDuumYJEcjVtm/vpN9TV3lZ82GLNw/DU1S98p5RUbPtvOW
gtwMeDmSaeXiKK4C5FAHpC5oVteGZ1o433bvIYUpWuhqbOCWt+KuA9dy27ge9X6wUSgp+CzVsFIP
pMifNH7ddLYZVXJpo6HrFxfDl14Pw8wLjIpZxoQAsWq09ZuTa7Sd06G0y6CJtoAqs7aCCSJW85YQ
Shk9tiE3qTosf/SR2BolHmGVUOYrJVRPA+RClM0uVaneLSLwp5JzhAVfWw80BHnnpe4jal5swQFp
EM9/cJqwKZ13RtRB1ERAEatC6HOhzjLMAZBHa5YOJj2RNE2Z3k8F6ZsrWcy55n+rFDy+04OSQ1nT
9yaEKN/+EC+J1/bTyjgxuDR771wNaJh7mAtDUMc2dWVRdTjtnEanucaf5Ue+7A1KZ33x6mJ2bp8e
8xNF69aBC7P/5hMbJsKdD7RUDV1i+DC3FooyvMw40WqQRkD1uIpx1uumoOodar8wS6Z6kPJTwwv1
OQ3p1huk1fwcJnF9CM/hx6Lwglb0S93h9ERQfHGMtGQwAmKKpwvF12HQZcVmfsn9bI4LwCASBqg3
RM/1cgHrJ5fbdwnQgX2IRzHMCBg1nRNOLK5S72oWM+G2O3RWEShl8IFji/0EdbrAtYTMGhk0RtIN
BfVHP2+lO9aBgfX80zKU6CYIcArQ3Ttx3REUVlQiKWnHnDdxN6T1uGnTMD01hDsU/3S+pnXHYY9A
nO5cRpGGWF46ttPSt1eM/J40y3MdnlWDuGApY5ecSeT/8pYh8XPOBQNNfZFFaod46YcA8jc7sC1u
r0xExLQOfCPfqOKX+T+3U9OGm+0NdqJn9ksDeUOs1AyTJ6yBXP1aYv8rW67xw/Er4+9xzVKVasFH
Ey0LVIBmJkDS6lR5PWPUb5UyTmDIEJ7KGLjbqcriH/rfDHOjRvrae4JW4T9s19/3AiqI2E140GbQ
0LgxTngMS1EGhp21/McXwMgzNFQ82sFvb2Js2LL+xgl4BgheMVWujYirQW+a/OX5qmeh+eDCPA9s
4pxCULLiueQw7havYJBRkFl0YlX9HwOg2RFMFPgqxYevNSr2PBYZBqNkF2brwXgA6ZcTQAp9CqhX
fm9Zd+dAj0ZjAGU2ysb8YBE6vYZ0YwZctbSG5WmBoYNn+Orp7tn+ij4JIAnLv+4bXcekAKwFZNwR
eFsFQF2ny7LRtbB4CD4sKl7GQPjVJ0G/F35pvopC+665v5JRx4MSfrwDf326MQ6tj1vtSTiYEoT/
Xn7zF8JPF3DdMA3NOoS2b5DZVu74MvnqXqe8pNyc7ZdCznkcukIuLb1EDqL7GKi/pySHZySqZYM0
OnrmbJfPiG5z2vA4Np1nMiyDJzS7YfjYiqiWregasqKXjUF7KHZTykuC5QikxQ5d8m3QWfMcCzhh
98D9dn8x0qjWg4fqSMYDz7uDSjVp5j/Fx46PQAyFhJcehbrMRw4SRBuaftTjSjl3/E91eo8Xx7K9
mgyRQ2B+Rx3ae0aZtqI8nH+qDjIoFg6U0tnLFJwmOP9+f6e+e6IUYqhMUbTHUuwU48KprCjqODCV
5fY0SavkGrkbdlMXVIoF/CCFIfd04nn0a/XK9uZ3U5LYKdTiG79CCDvk8cNHrL4MjLPXNUJUqazh
ybI13asi0oMG8TAONHX1QI0CIyjuuxbpdAdirK2t4k5NWH/fW8AmzYDg6dBYUPrBV6Z7DOnD0RO9
seyFHykYuhMKdfBHyC/Hswqup+N8XfQfvyX8yIhv2VXQldD1zozlTdrpIEolJ3a2l9AKMWgKOIwv
mO1zasgV1kj6vF7sEYP0qsyBBUiSGsEkc3LaMInohtVatiGh7MmmP6faVVM/zMNgmhsDqPrd0xq3
FGskXunaUhBBviZKr07Shuw+VZS47FYRJhTTP5x/K6MZBKYLlGu1Y3npjzpiEOOE+77Gy3tufUcu
0cidDDqV9Oe/4dJiBHw2ZlUryv1rMwbyPTEo/vJ+lE0TN5rPaX3Bhj4fxs4dmwNgsPmyKdnbQ19R
pad3Ar72QBHwYBfBj1blqcDSjHkSmQmn9gHoY/8f2lJabqyZwQB9rhdpnib2qA3qVsFEK40QuWpU
Lgo4ScRx+ipmMSUHkuKWpRuFj4CgNjHrzcxtWRLdZ21b1MM1itACpT9/MDzuuaju68CzxyBau/tq
d+fMHh8804VtceUG78SuNTdH1EJvGuRKiLhnF5CL+UBaTdIjjC0g/xMaAXwvtjbouSM0GHN0tRlz
xWiciShAsYpZq1Dfq+BG/Nu6jBgD6B/qMy6POpFZus8vnt8uL/seVCYo6yNXeAJ8xOMGMAZtsdxV
6DRHONJxWME295bMALo5cZK1UQLZ3YvSBpuEw2VXit7/BNb6sj7Kw8Okv0Gie+/+GVX8qgFVlYQW
6xDXjiMrEyv6I8PVyUAHvRdhIvfCuk5sf9tPzwmUpS9rGxow0Yg78vEKfA5RX4du2+4mf7AHJOSf
kjB5Z3Dm6JcbGRMX+T8IcKwGc8V+iRzlA4/LMnB54Wekp5Qps3C4IVQtpCOdkOQMhUjjtdYEuMe1
7L/630+XuDXM0g/DyRTDWnnN4rYXLHf66v2Gzn+dSHQhIchlOArC1PBGlfGgXnSHvyVOVDCaHEue
WM1kjWcc7ncCXIKeB1xiTQDMpRuu6+lLmjDnXgbBOwgiNFOdjrsEEwqLd5ZQnFE7qJniR8c/24PB
I9FPReH/pcuAqY9KTO//ikq85REVXPN2NyAvIYdmqbdIALHNbi6JoTGP70inwtYxTUmFlHBfN++z
lD5u+q/xleGGehEhFOoMicuaVvqvfAiLpkMFGRYggKCuCajP7IFj9ZgCodk7orjVybXRDDxJoZh1
82SkMSucR43k+zg06PxotV3mSx4dGsTJ5KlkA6xVNZwKb6rE/NfHu09rwgB9NAAHhcdJjYvsjnpv
bs2h+mmcswJxSiySqMWST2wAdCqOSio+eiHZ6YWVoH/SThsy4KYZhqvqyTmJM214/6jwgtXyl2a+
s6VM0DYlB/Q88tn6IGnSll45ee0sN9FZPH8yod1gxOadwfV2EA3B+usz8pOrXQJuSybkb+GCgs5C
wwZhuE+Bw+a9wziyiN9KE5p9O6Ka794F6uhZ/4IiHz+Rf60Un45fgd2rCp3o18cUQZzJD+ZZWwG9
GajFbd1HvQ9VerNEmRZpjN0cBj2GN4+BS2Afl45A5loAnx1+RKuISBk+nJisNPKFoFu0bfFzeawj
nki9yOij6SSxBLCo39xFA9Ko2jDGkvn3myiqjGeeilGrmsAOXBK43kyHZBcBViDhq9LLmZ/Fe2Co
Pt6ZakYeKk4MoCfrgsnlXC895AHlDtvleZ0feo+tzBG+i9KjfZoNnLyA7WoVguDo8hqhItm+chMt
IX3aUF/BDp+e/sDR4g1x3F0NeYUtMWBKqkpUCbzBPYzYgvW5V6n8O00wa/yXUHz2lfwmRIgSjxDR
CWuhukBlVS28I8ftn5niAwX9XHxTB1R5ktIqIlHbQI5W6xzOppXLa48FwUK5I4iKNUR+5Niy7W/5
+g+ZSjRQR0WzbdcCFmZ+3swdXADoS3UoNTz0V1Dogc3l4n0ADyYQuDuqtuwQ34cXwNE4Y5Gmr8Je
c5hWJ6BjGph1i331cUeZpCPTd4Qm4PAIzOfs5ryfGr9zo5rITnoQ9s4fr5j3I8SY/94MuJLqXVPU
egIVoS+byPMr5Utd9rlylE+nj42pH8xDftm6otqce9EdUEWa+2jYj7sQkn8VxUN5voqmLyuTfVRj
pusbLaHnm8Z+Y3w6YUYtsBEthFZI8y4RDQ5447DYICmcTMdiANVii0Y2Rrt9hs1h6n1MfpkbnPMK
WcnlL3OhyCDj1CxjXl5Dlf+oSpl4q8fiT1xrbGh6ZEHELXS4GNbtwb2rSOdI8LnO2DsD2IGi+0PH
rQ8L+NmkS3u8kkUPYXcsC4zOxqBxE2dW6vtdY2KV/uY5dK372LFWJzBqj8WoXMH6hZh04f5Q1UAv
+euXIiWIRGDSGc4ttMqTDyNi7xqoFTu3a96f9Zy0IS2pbaC0oKgBZdf/VcZ/48cZ7ksq9ZTBBKAC
JBEp3RgRDOzW0WZ83IdI2pANTeaY8xhG2o3CRTgQtKrUaQ1yDY8lqBXnVcTLja1sMktcu4yldaaz
ZwVnNCmvVufS21iRpOCg4rDdsbqDqx+rO2Ns5J5OHEyOlfp1fdlZTVhqX1d2uz7FTlHaHXOIFtfZ
1H49+drMi9xoZUD3oNzeIoC5dFwdAoG5fYUxTqahmLAQS0Oek+QVFTw2IzI5+v0JFvAfImI07nVq
uyg2OdYKxd1V8aZQZ4Mi5PxwgrjmEXUYAXNTHQa2CLlUlwDPiO3uqEGOXEiUuWRCFnq7RF7o9eAH
DT9uZFSyyBgS+AuK2uRZbk205dgAIzB8BW+0Zq/rtdiIvcQCkknqsC0eGePERG87dNROuMmdMJCr
UNFbIgVqKjOlC1M3Fh8PLX1FdXUuhVbPqgJg25/k/1b3jVpSvndrJcFsFNZVEdbq3m0uCd6k6akS
6/szgSAlsTUAG/YwsXYRe3gUJlwB0Ck18MuHnlb3HhiUFQW90o2J3RLi777ajcmfdJFVEQU27HG0
j1iaZTY001fuDMFAQwMomiCTkPShknCeFOrc0udlMpGqkqQXyYndOvVXtWWfHaWz3+tkHOfhKM5/
LeSorbQ+xYqYQMn+Eep8w/Ka6PGMx+STsZ7D195SyRf88c2kM7AJWRARtKfkRnZApHW8SFNiIHGm
7lHO70KfDdZcYfrjplSTb2ys5wYhVYvomvXur7MPPBnsZwJomGtAfCzX5k+428kI/FCBcHKLKy0c
qmf7jdSIN5rd1y2S2/DsvmUE0g+umSYO3i7QL6F3JsVGh1mgx4PQJziObfRImYWa/CiAcxj58pIw
XyooXoWamEa8HPBtJh01mvHSh5tjVBmS5uLXjWdzFvJJ1wwRMOAzQnbKrok6GJGtDl4pnm17R72E
L6Db8OLhjib8XKKVlCbNDPTv7PTK7kDlz1P5MwLhJ0o3wAAQg5O36/J9/pnlZ3Hfwy424JVewHdf
Qrw/9vh28l0DJKahABgQczDZvThAXzk0N8dgTYdN6IHnm0p2j8nc6rYhmwJSq6UcMkO16iNGfn5z
koG7O9bsRfcZA/caJqRp5hm1ozsIZvYiXWR/jtxkW2s3Z9EUDCp1dZeVpTNyqX60dEwmXNiJBXI2
3JS/rmEV68bHmGEsEO1Mk4YHp20iswp7quXxJ7YgJFf1Uuzyxv8c3tPD6JuTDZbGixDzjugIabhI
kOWVEIz0K3sRRU/A5y5OBQJtikKAE2M/CsC8zbV3F7Z8cX1q7nUQwr5cwbj6pA8qEY1z6aEKc50c
AfIN0ezfVjrmcZreHA4U4LdQ0zf6u80aeNNwwe9qp9OBdx/27oEBU0n8bZNCZo5msTVSs/QqXfmy
D4Nbtj9b76r3ACmjW9P2GNg1Tnmk6+8L87t/PTlTV1VKBOvQVxJMCBqZ9jXZ0gSr5TR3aEDNhVYj
+8qb6Rcf6djxYqL3lH8sdHUlc4a9ijYqMoY2fgiCN9VPMok6m3LrM4j8kWnik0oIX2uxNc6en9O3
I7uY9N8tfLvN5YMHkUjxq9pfaGC78jSghpymPBEPCUPHnlYIndbXmjCp9Yyeb8AQxje/3mv8UywB
/Ee/7tR4CcHcQNP0viBOTmI8Yigc7hiqBIzNtULvZa0zzDg2d60Abkjo9Leg2H+rsU9dpLucU9P5
oc0g9gxjY2FgoF5BZEbKuIOBkQ1fSazvyGAsSSHmVSFrXO+nsZF+iLZoS3rfK415weQ6G26jz7g9
SU2bncwInCNK9ujhksgfHjWfqA6uMR2cKA06wn7g5z3G5FCVo8PNj6FoLed6kKw/+VPYVH7UpXWO
RPkTVzLyWAgEHPjCYfU7yRJbNibbfalCtoeZctQUj5HbuSetWa9yZNIznXx+eEOvCL9NID380lFu
NHM1H8+fb19lONTRWyfAOTcj8ud4cneeD1PCClgg7V0zNt3EOizLq6IiWTj/SG2sAXsG6tbBW7Xw
XmHlGfh3Lm8/VSv7qxJz+nOqfPpKhNjiKvlVNJcXha4NZNjvhRjj9pRF3qb41OXO2sGSjX+hDKe6
oHHvUKMYN20vpsK2k7xW+p3Honmx82quC+zGkZJRBwj0gus+rc0aqZ7WFaoeSWhmA8LKwYMycB9O
Gpjes1TXbLyVyxUgq2LDLde7AqC+G0/aodmuKoAMEqswHwMqmih78UiNYhfQFMwzjAyMPgZm6XwZ
JgpHeVb0iYou+tkWdvY9a2J+mj5y88zKRswb/F+uCLfyTOTHLfFiOvUvZzdny2l+3X7/tpVPyFyC
hAdPVE+1kwae9pgbnSS8hBVmaD3pw1R70NIXGI7chwrbljTeFVQOzlcaPrF88VswH45LQi/ve4tY
ZC2lE+67Aup1L6c5c2c2mfvDHqGpAgRCYnrsS+HP7ST0EBKwGEctThUS8Zt13UUx5ccXyeFO9OcS
zOtNwjQ1FhayA8O+1mgXKVk2If5TbjTv9gpca3UwmqiDjij/r3thaDtabUFSHSt3Dnp8iYshE414
w0OtaQexiqmJtn+tqCwWzELEoDit41QvBrMwCPxVK4sr3WoaemtLD5eEpASVqCeD8sZznJgGDWw6
4esZ7fLwwi+PsFsl9rxPsfdNtpXDYjUP8wqf3GUmFJDweT/BmULYl50eEV0wHCWHCvahbaam/nZj
YO1gBxEB4KpILljhXFM6pMGjCJFiq7tIjacNDBkJcRRc2xi9/9R6Pb9OU9HWj91hY7kKPVb/tY1h
f2iFoJ9r4RjNXdkntTKwJHmDQsSfgqwNB0je0epIVGHG75JI59aT1xxolKzMflxIrMg3DnQax/oL
yMy1+0/WRqvjq73e3KJhHK9lrloG6HV0ZzNF0ycn5kD37JV9p1fCoehW3kGsMgJGHscmf/ME3ISP
sGB5fEA5C+QQ2fx0pubL7gdA1mgG8MY5DspgPwxPtp8o/0OZCsHGSKw0WpSy4MloywQZwoMmOI9A
h5U4Dve+tINN8JIp/nkydIOJ0QYNCL/84PbBLyBYEndSlb0/c+RN7GxAcOHu+IzzPJzbaJhRqWj9
BpBkRGAWhF1OkwLqc5zayQVECwakIA+XByXWZWWNQNIckvqaVNvD0neSncHP/iCAbaXNFICw8SX0
jW+0RKuIQY2VsB1ZwtuksQPU9tYDDvDX45j2VUxx748OzR4woXo/cWOrn9tzdvwx/gJZQoItL+ka
QtMEgOcYwiI7TPhnCayWvsP219o7G9WbTqOqZaqQA3AW1TdAOIk8hTmuNu9KV70DWPwVxXYacKKP
kgPBJpPFQeBCx+xUEdQW8pmjI2F56tAwHpwdx0OHNGvpyy3EKJMnEOOOoJRh0VR8YyZi8Fpeuec9
0uxEXqjTwAhGdsl3Arx3rL/lM/Mzw9XZUPC3C61n60eOHum2TzQyWYvH94TvCH4X9QpM62wakvR7
EV/+Iao7bePDmva7H8F0mgXwgTAumlEjbbu2cjNd5KmK7HllO2iAZthSTMhAqjcDq16F5GnKFFFg
AD35JXvVD/q0BOIg9g3EjROEXLRLi5BPGy1TB/WGmiHDUxTreGRRmBk3b6Z8Stq2t0OeSvWjQNhD
u8WKx5sFod2l8iI6k5xTFdAo1/O2qORDcxy5nGV2ujCwnhpyKAivpwpsf3NGIJ1WKuDaywTv/j0G
zAyCU7I49+Jilm0tW/9uLJRGOQYmsK9i4VEa16bG/mKjyN0yCtYCpLDhN+I90CNuKxkJYOHeVFTY
Rl6h5kPwas39GM6dMD12oG2aa8urNDK8MJm/SmGG4t7I7P2YMvd6eHEk+jI2d7j3MpgBzoWFZonV
N8xdtd4ZI4e+GJ7SiqdbzbCml4Zd/cZRbJRn3LGL/Yc7lyXFHoS7PJJ7zM+y1VmVGdvF1yQ99NYq
5E/DmU0tVPZkLxLZs0KenE8oE8dpN3a7LRl4JSHPVDlHIASaic91NsqMb5ORGiq3oywB6H3X3aoF
aNvczQD+0ZIDyE2vCE7++H8Jp41IO4MZC/Ry46J7t6HPUmqzqRpRLoOX/6KoSKMsO1s4dSBuGDDO
rb/l5K7IoNFgmt5ZPEaXV0I8mu+tbGyfH1eYt6IKbYTPX0Rfmyifkk+39IISw4csc48pbt2v3td6
TgXlpn4DhZTGCjSuHRCuRvJrp1P0p4m0FNwNT0glfLLvGNICO5yvigeYQFSHtZJ2OK3ajfnPlIUE
elAaIpbq82LiDG4ACGdup5ERrBlQyI4JZ2ZLGulIB837Xcwrt5ms/0HV9RQB9kMEP2vKXpxt9a0h
ab2FK7jg5NPZ0TB0Rh4QjmyqzAoQb7bD8tcCEbbyXd1vqHOF7ITbcm0UNv/RCiyqLHoEWWPXnST5
UMsaS4BOCDk8Ye9sjrl0/aqFr1dyqY9W5kCfuArC6sG1AXV+9fnolo/wfbgJkx8YLjYAegaU3gQ7
dCLG/fV0wNa89fP73RVKTxpZ+e1gyAZUCbuhJXtysfdu45+NILuAkXA7p8VT8hkJBjQrYEzbWE4Y
ocPX1tDacvLaEyMlSZh/zsRRJo88Km5bg9PcjnXx2yl+pdRCCNXOYRUens67cKU2I/DbwOA/pPgI
cZGD7AW34rCWFJesoSaGaJ6QtvhKNqG9UOTtJbbGOigTmEJIhao2ui1/7kCYBDXZPTF/Sb84HXxW
NlTDAScx9vmolcojoglvSgnLPHp/LGKHMc9AHizyHMY6d6yaQ+sHT3EY940rS84B3oJwa+GcM24r
wvAwT9Yxj0IiQ7JyUCr4Q7sqQE2DFCZFJah5fooU9DtsgC7XgkeJ6CsxZvC9TEjA5HWHtuDZRrJV
nEx+n37NCyYV6/yek+ZedrGx7x/IAUh6pR2y7ab/88uaAJ7mv3e/7Bp2bKjmmNAwo2J7nsXstzSj
eyaMcbCkkoFLBewK4Zy3OoVjoiR0qd1M+kmxrprDmPJg2dIdZikqPcHSbJDhSC/OJT2nqk5dvoOs
myBussg4zeJyyioEmofWWpnTY3xquyABLKvGT8RNsa8bcYaHq9gqeAFVeJU/HKHqJyG3W6RD6onp
liBNjAU9K/gYGboEDSKk38vJv0OIeKTiVyNRscAw3qDdPqzNll+luwvNQU952ypojhXbVrd6T3xX
bthB5T3OHyAGul7JsQYOqAHP/MdvZfgIBKa98KB9zjSIV7OL5Zx7DMvntaCSec0bjwCWo8pgFdie
34oANv2QiigV5wBNcMEDNCpR6mm7DWTR9JNnjMKl+vXI05axqhW0OYKSGXS8lCGr/GJtejMA4PoN
M6CYLaaqhgvXM+UiExqCJ3pDKbqAPTT90Sje2btxKCZokiu0UxAeN3u21A41nO+T08hrQ/Guzuip
as0pG/0YBCG580jiqFha2K15ETYZr7AwJtFNhvv90BqF089tq9gmvRuNQHrQOdJi+FWJNSumjLRg
RMhgP4ynHKH1qtUSnxBDD0GWe+GOq0l6o8bC92ThofxvYoIlln5yhjl375/DCiRLkm9bxkV6r2OP
luuYXNDVyJEVFhiGg/aib2v+5aCYA6nicQXOa+zR2tMsvrGEwROeucB0wdS4U8lgX0kxdgvP13Qt
aEO7Ec8aoWjPClaNqfF3r/J4QMRKirWNrOa9hIW9S/Hwh4hTU9wseE30f6ChkKrHji4cnyiIYxa2
MHyqyfVJrFgTUJEuViCb9rONlRnxfU0hqHorGwTsd53BU9YIj0ck11z95QiRX9KCrlgYOkKNnxV+
WNTNab0KJTpsfc4RctEbJ1ZMIK9vNuvXzrm47GOUwU9xlHnl5lNl38Thd7dbbm0X8wcHv/ZK2j3R
hq9tk7xaQxsdTNSM2OkfFwwuPuFjDRVOuwwHijlJnRl7tM/MU7VcgHmfrTIUrNhdgLzOPfPztlHX
HrhI2/wdpaZyPbRTrKr7Z1fR0iPZO+6Kc2Ys5Gzk8Vcrs/UXh7coei2fpnC8gvW92JR9sZBfuhG5
Lmgv2v8vFC8k9Ru7SahdlSdcI0SJddP6SYhsP563MEDW8w6yyBIj2W0ON49PDHl8Ry72oaQw+5TN
xxH+Fa/+eBfCKDjJG8GpnIiA84kUA2oIRUURTnM/DaK0m026vXg9n3B9rTwQXQK9wKo3qFZQ0Ll5
c3JJnmKw/3wiQlhcBwTdjK2FbAlHafV4qXrDJ1rBJ0Ps3qzGxddTSSGmRwgmPo61Gzd0JBg6bQ2K
mGz9k4B1EA1FvdgbjPSUqK/mw3/3+VbMv+huKOdQbKT26jeRX8QEW/q/VT/PQz8wKxqWWuGMRA4G
S9qgmhx2OPabapqK8oO6kwTzAAhkO5mSFj/oBYE/ruer0ABI1pP+fhwqz0hlrUGMPuaIWEhlQN6x
KzY66J2YAtXjXEaFueb9//k3+xf4G+6nUN04vuR9pdaA3GKHaopLfFs2ndOB5HtVqxz0d953RGVM
jPXvkxmETtmMV6dyOszZLFBEUC5i643nO1qURoLRmOwr6eElryhcHFAR8kALT5efvzjNPgC90qgH
TteCqOZF2/rySwg3duF3+VRzGVDFGcYWR2b2zw3qXbaCdRyAfiyJTDm4s7sJ7SXVx0eq54pqHn1+
V4ks1/0Pk136VvNBz74IqNwfCi6s0IuSNYvo69pmRQEusdrQQE5+0Jmny/jxcgmFNrMye/HH3Xob
Y8oscIZL4YVw2r4Are7OXWe/G0rKfg/8NvbrYD7kFQO9bAcigGAU7SKTW53L1merIoNjKb3yj+lT
teBH9JA6BfOu8o9A02gWGmTmXieHUEbMQ8G2BLHbLbG7zatTC1MPt7GJZZuyMxsjYS4VU6O1o8MD
3nduD4WRUrqOGrsmxIbagtfgOpe1QTGHX8kOPQd5HC2FKVejURrO2eyC8cZWDrKwGREptzN8TQGa
D1NmjC516hUhPMFfZi9G859sg26fxmBj/go6ZmJ8VavzC+98fR2nBubuFxbJlPSPju1NA8k6yvE4
S/Z0q2wpFv7GakYgMzzZ+q5Vzv3Ij54YUbCml1yebo2cEoaxbyuZHEx7f+xK8UZ5ge0+dWc40G4L
oMSFPODodiHfPUrlLkivKoH9BPihd2CaN32WqDHARA7238BeSgghRFVvY0Mu4k7PR/oQ4L7B38JL
mtrfuOwlI334VZEuzsGkqaq2yMvGOyxRTibPwcBYcH9v8tW0pmi//D+pLyT/SDxXSq+TqF6xhgQW
Zuj0ekdn9ma2MOZNg7WHav/sJNfcCNl5F3xUHqBORnfWNiEVq/NXu9fMMijPJD7hfW6eGSHgByKb
DJZu44CahNjqk4HYOT7KQsym2AC+jwU+3FV035xl3vH0wm9lL7XaJ3yjTprhjKryvQ/kFlHu/ks4
jTuuvVyjIH7/Id39k4G+FlIqTGod6E+crqgPqUTFF0Aqnh/QifdmWxQK2A5jgjaJ1q2v1eADP+Iw
Z70qzT71/Oy3N/wENfEWJ2N0U6Raf3oySVEDfVUv8C5r8FqnriEvYLR8E/0eDTYQ96KR0fNWt/0U
GE0BiYl2gyWkAbICp3nUe1Wctueq+px13a2VoOgXqRIZNx5cj6bT51Z07na2aaJXrses1PrXzHIA
Tq4xu81M68il+j8ILZj7BX9juKilExaq4Jhcqa3XuXCZxo+mdRPcji+fMdFdis5Bs2sIJFXZJcYJ
FSiBNe2ZxoYyg0SCkk4gdBOr7RyTXa1GTLh3hf+0qDVBGJtJHX658Z5utdWJON0Mt7ME+8SR8myY
qk4X15dYafDo6LLTalGpCV3BlHQ1TAFkHUUWaTSY4gRGA9ED718ICIXI0FjsQOXFeHCieGxgbZtH
vB9SKAKplxwR/BmvLb9iSwVxXUJ50cMtciH3FqzzqwtTTM42C/LCbXY/8DhXikvv45nG/4/GhC5R
FYOwArGxEqrj8wv0Oc4HkWjFiyims+EyXngPFyawyTUnFRIYNUNOWX5cxRjAgUI9XyhVwC10Twpy
uiwP34qLKEI5/a4lNJdHRKW9HuS98sj+oeKi597iiKhiH8QjWpKVDauNW93fI6wV9MYNR8dOwjgr
6BfR4cu27rsjnJOr09y6rfQDiirKVhKOgdaC9/+JfJkVatA0LBLDg9JuRZcp38eyhjBSh7VF8nl+
af/I96LPhMbf4A8eEK9sJElIG0WP4a1xRkVuax6BaKF3l8qmflCvMZo3Mz0uahjQPE4Z+w4iiiKI
wYn54k3BYSkKA4iu0xq0jvWtuICI5r6oHuSGSB9YKKhEbOBJ+KwWE6CBPBfdE1VTgPrN9fWseKKH
Dv22cUAF0xm9XgkvPOPXh2CcMHAioW/QPrs7LsGaC7s3g679H9Iigqu5j+4Pw5Ub4FzKpJ/s7z5q
FOGVbqFs5unXTNLAR0ND09GHoXLvadCbY9sKpK7RQoAsnBj/INcVvNMzWv+87LblDMSCwzwc++jM
xZjQ1scVy+7ocmZBH5J8zDbZ6eAPppxLIBSykU7cMAZbFgYiCm61RcIqjOYjaDFAUuhG/yrpNk+3
g67Orgj4F77WVPgMpluCSMhP51UOGvjFBifzA8KUDcNDhIN5RsS5vkyD4v6VzhpvxYErKrj5PqnD
WAtgsj4cQfgqbKNyeKARbu0B99i5ydbEMHhWKT1c3eZF20m6kbBOKUaBjEvl7o3iIxq4NrQ/soK4
wdUyHZLUuGg6rGSS2luvvuSFqrvIGBOXI4uT5t89835r8nAxtav2X/97K826NigAKX3ZuT/kQStU
5OyW5Y2ojtDHZAAdY4DN9G7hhu0Q6ceKPvm1FM4CtkTyB+dxGp/QSVQxGy9tt6Qp+cQFIIFtwCd8
eOtdwB0qb5XYadGAu5fN00bxYXk2LcQfz5QXq+MUPciIb96wIJP/MEpgYAtcC2rmEeJd3qTbzDMo
gSyaZrjPUHHMFxXHdexaYn6EdOmnMw3g7cofs+ihw3RH9Cd3mxDbUoerNxr/2aCt8w2Du/XMwP/B
pzNnDlMTjopqtrLgdOnRhtewOvVHWFNrH1EVfEukFAnZ7c34bSwL3rwCfDbD4nPDPEdTKgd+VNYk
VZRecvVycj9BG0ouRhI/IUvJN/qQtL0NqyOHuLC+qAf3lMQ5wjDeC+sIYw9IRlKPpxrUsFIInRUc
JXRUEXf8zUWMD1xB63a0MPD0WmZzifZf9LYnbZAW9LE4GuUj1HsoZB8bXP/stWLmEDGOEKiASv7u
nkyxe24uRS25FMwFnho5p3c/Mhb27TbgSbLmihPcZ6i6UbKHGTke4FbyjT8noEVt6UcJmRtD1z8s
YyN2LfXFQriB+BHw1Kc/k8ZOcKjjWCfEgA5+D+RTaMjjenOZGnEeGeq/a1rppQicp4ULrAIr5i+H
c99g0a69YHMNZnFnQHsNzTNaeUOA+R2lFjY2JiFj43k4EUFNF+THnifjDiGNfvbp9cKMezH/ZVPT
cE1a7LJgwhLZFYOzvuut6Wwd77V+gp9+7WOSVzDU8tzFPnA2ESvun+yrhydrLwt7MAHRzK+FqBFl
+ZjsvzV/5bswwyjUaXEJFiSrk9XOyKh1x0FkFEHqMBui6UIqJOUgt7EqDGM3FjSMgSgNx+Wqu9s9
Ue1qbMQXCnk9V86TCY3CxiS4eC6EY/4ia3lj3rW7fBu3+JrhOoXjeAcVggJoa754SDQvpIw5HmUT
sdJm5QPUCnuWjuA6Q7xChdB9YBwZ4EClTxRiAWw7ZJpgE001m7wKnGH0juQJUdgNIgLDRd3BBsD0
KrqnQ2Y3b0i5cXjqbYtiHvi6AGT4x5FsHdZO5xgFxbJGuyXSaetaWfq/H/c/z9Cc7Za7CMvUkx/c
8mT9E+teu7ROERi00iUbKUVlZT/Nlkqz+rzvVdxjcY3Ng1pSp4gWBFMUYghW8miaQpY8IVUQLTqM
D4K91ZIGs6bOFERY2P2HXZCtoGC/mIqFr7aXXchav2rFzmaYvHRopVFymJyg3qiCXU+WTiEPOOZ0
Laa4ZG5Gl1ZT1YithcaYLu1UlkeECn4eJR7wTpRCZsL3MJM1obri49F1cUhq7a3IVoAOTc7wFlHr
ZQ4XMPilpX6cUA9mgvjhJ5Q/mWTooFZmjsDE2Y1NjBfuFtdi9aPNNLVlHnYSnfEnN2UN9vQVV4Zw
/aZkciUkWGZH06O4RrSHtSwWEuyXJ9nMPbTiC+F9Qxud2UnoE1xj4WphrEv7Y64kJlPHpTrtO2pD
kqU39uOqGGX6rE6XhYTZOEQQpJdAAQE8aB2O1XTi31qoymYmjTa/OeD2FOxzR5ZOBlRYnLaQ0PRo
vW/VHAsJyzpySfOZo1yHh38RbJaeWLo3YnEk577GCsWB8e3ADDLk6iqbKIbRLZxuwUv/JBmlvHa/
5cb7dZO/OdStuKntQqOCw/iJsxbSvoNdDVIghnDuWfVJdnkXfZSFkwwVqwg6wOjd7rMeax84XF5R
KNhQ+NF/Z4rNfmNdlLiPSfAU6uvjFh1zSBBCgzaCk12x/+AQVaQlgtFSR9gFAgbaxUA6e8QIIVPk
UWvPhUWBLxUHJhE1whX9jvcA/h1nWJoevrBoL5MUo6He3Gw6ucGkTBzBYkrurAroRRZtfM3LtcpM
wTFPN7K7K7skqLCIv0BPLtwI3DNsDNAgkTDn1j1iZTZY48gP3cUfsof9nBl50KGBo85JKzb6ZOfa
9YRFomoY3ac/OJE0Zmlgo6lYJtiVQnLUzEyYBiRq2Nu5lArOQeWxQIK/iV8yFaIGmLhqZsWU2VSG
GuFtonFcWyz/t/SdF/TSQ7YB+/aUWVUD5CESLFRVNJeSlUGuPZfabaL9u+cTU6Cc5GxOvSjX4bQs
EL6Mawmgd8lxjBY7EGYmpxQRB062ApRlMDzbKCqaNh6rTJEyiupknf+ZxItsJomqke1pWzqLSZg3
WgQT9B83ayKYtikUGekgAJSQ6X+8Gzg8dxUm29Ml+RBsdQUefqQzhI79N1eBq6ESX8hbS5EWShLj
rbJo/QCEVIH2C/JtQQuFhQZnrHYKSv4I3uAxxzqYIPBAAm2qIvJ4sejHohyOxuIF2bT2Rkqch7zj
EERekdaJcZd4F04ArOzACcsTH/hfrs1LWo4uwNnQ4q6/DQd6f/ysbz/6AUPyqvNgRVTJDjVqeVm9
H4kogjJJCZSGwRv6b4ktk2L9o0PkPT3sw9q8LZ3UGtPrFGFgkYKoHzJ4AYCXawaWZG51T+9s+BBW
v0md6B4Aj4E8ydOwWybZSIPXDkRGZ5onIzhrV3NB6Drv5EbcR6WpGCtmkj5LONERlYgtRGIRtbIB
KlNamoomX9ELB/7yfkkTqaxww/hSoXLJAQ98ZvXyHUjy+cETZzdEdVfpKr6iUkTqhlFen490OUre
r+IP59dwUhVCb8oomiFBBwmUI+qqAQjLcDRolB8Kb8rPbylQMM/SrsyGIKTmrTQFx/O1a/xetAHz
eh+EAcHMflGvMgj1hruO+vyb2ELCYi1cqMCaBsfNAeCurXlMm7IqGIRJ9R3IAZnL8M9W1bp59jhO
DhITAKCwUPoMhkVqYKEXy92IDMFWCHn/Dd0FT+1MtXCeqShY1PVzDzZvcDtL3l4DIFyWFgacFSIr
xinwFEbdQzzfGWJTL9iySvcKxR9ez3/nvt42NcG9HVlI8w3WmE48AGs8gOjNdg1R1Q/2RCmoH0YN
PVe5sBa8N7K9U036KZFeXho1P03BW0SnMFK+FGyvel5d1n3u63z2QuM8p0tWCWRMee/6HWQ8DJPL
F2snbU/eQ+9JJXP9QU1yJKT14iW1tQDRHvBQOS06ed5v8tNLPVyTKVXslP7eLG3CaLwLmmy7iK7e
RdvrZp5cfGyKGAMX476/rFVJ3rO2UmKRIvj5npHDsAboZgKfbGp6BnHGHPAdbBFn7mpfZkvFq+/M
NE6T+wS953BI6zek+JzNHMyxjZHAsrGJI7SZbKeuwSQPrSdYuHRtIlR3KnrX6wBk+B/NYfMxUWKS
x+gDL8cBuo4LP+M6fsKH7/1Cdgo/M6gVkeyEBgxfvuZzInqC1EKpZmyKvm+L6a2U2EdzLoaHuBu/
ENNlF5tPfZ35HYhCXPkX8VWGdJcoyqc2I7DXpG4kTYmHO9dCOH3YP4q0xPecXPWAqeubnA9DipY+
HwGIKbo2edW4ini315ZIAZ6kFZJu55S+LvJqsU+SPtJGrtwaXzhBglA2GiWUa9DXq0Gc86gUDpLN
3eTTFVdaEoEABPk2wGrWmiqw5aql7CLqNvCammi3kw8+tnKAWC0LxsCe46Sn2B5ZtGJOvB+oH5EO
Nk7GOLCH+TPgPW/mnuFu4PUZKJ600soJMihnQmrW/EJWtaMaW/3M1q79+81fit5hCR8Yp24FG7E2
cvXsPUuBgxh60u2UzcvJ47D/7dU8+6wbks5LGINgGnVX5cOCRRRPUERefwQOs4CC1FKH9H/6VTfZ
IkiUOsp2B9UZDLdltiDFSawkvpXAPcul7/kh76x0nx6e2ImBvYLop64vIXOY/8B7wvN4tpGzHaen
DHTQ9KzAcdu0E9pB06idgLNMnJpLZx9tIU7ncKG1fDfJa1FilYyvv/Glvsl43yN/A9XfLTJoUlBq
2g+VPNtLFUsSDMmIegoTlYjd72rufhAD6Sr47uXPgR2qU/ppJlbMQex+2it8ZyY6VTBUolo6UcZY
dMsqUtwN08V62h7yJlx52YxZsWOI7p+6/VoVgJZjKWAaBKW1jP/bm/kV3Ma+j7zG4UCBbRlOzSOq
mHfWAEVmbc8EFTo9J2MxOpK0RcZ0r6SSJlWe7hBYXVDFjDZsYvsr7QOCAeCi+lg6BdgZlNKHkV9S
EBQEhz6f3IoAWJFSPBHv3PlrK9nbeJ/HVRBc7qlLRp/TOmdso0Nv+KKCiSR2DYhG5GgP6S6y/489
+6PZe8tcmBtKJ6cg+eGJMQMYFks4mN83MaLwDCyKcOV1ZELjCVXrTWa+GsmRqDGKeH8zrja5U1lc
puWc5NXLoKso/rvzVqcOPZ54thTILfUhLT11ZpiQAFh9o3mmN/Uzsu7F3AsiBjJVEyg48Vlcg1+2
jHDKvxeq0PgcHjhmlAYaA+wIe5Rq7Dc1sKWphwQfzwkJy4PxaCy8u6AvsRoECAFb+Ko9qHXVkAry
NOj/LaEjfvbDHW7zaByWHiOZ5OTvxuWkaHZXD3g9fbVSWamQBN40vb1291Fc0AP/YFOiPVBSbgs0
+c1BGT7Qu3NrJu2F8kvX0blZyze47FP0c0LsJuN+kyHWKZfHFg02YM76E4xe56eLKCsgALaJjAS/
GGneDVtpk1VlP9cz/ZLqtu7Ke6Ud+/9WyR2/Aqa10R1dU/jM5aNnVUWaIwuuQ/HueFfMUVat4dTX
7e99peH3BAyOKFMPVwOuHGQVS5VBNTCpCcZTmpZ53YLDNvKON00e8KJmn3YcLQgYcf39BBbJpQ4P
jyVUBHPRZjdICG1d6vHcZJd9XUnScIhVe6hCEd3NRQzdnL0ImmNfk6+XQsBmbsuMZB60cAJB1U87
p7w2s4hksPDjzHIH7MBuxHS+iEYad1HICWDZFA+Fbe09CqnJcDXjUy5ioPXMmWPBnyXlaZyDxwax
FtHTbekIPIkQuGFC/2Sg0XroaR1UvtctB92rDrm427igB6QyUacnbUY/3OkpAgaKC8WF1MFVkSxS
6B1XsUmPLuhl16ZUo1HZtqyyiInkjVesqtn2B4ffnjHfKOVf1REB+XHUnkCfwd0bYfij2iZSvgZo
lrmItmYwaIIS7QETUUWSor7eQ2C4e59JiITZ5us9JlQ6M37MEcXmufaDMFnALluygVKGSKqBEUtl
oG2fJdiMXkI6phoykfXxtbZRP+zUwqdSe7qi6/gPPb8GkMItSNKUQMOCartguL7ve5c0BhiENLB2
KNCzD/4zTjVltZKmnXLv1iCMqBW/PJeM84gpSBpw56UZ5QXrUHW6L67oTgeT073R11vjV4xsIYX2
RaenCVHsodxYps4nBQ4YuU4IhBRhqvUneRLL6sS51iNN9t89EG2g/l1+/W3/3UST9fCbpYl7QfJA
6Z3KHOx9MgmlzgoAY8n14H34d+UlVthphLw+xZf2FBRDoJEUdXgrO+Ct9QT0kJyMlMwzxXmKxQK2
uCbvuZPgB+VHyxmOFF33c0hOwmoX3gnz9FuJ1zEXsvvt3qn6W9PGF2TblgSc5FDB9Xk0U5pLu99W
tkv99zQOwjza2p7o/3RC6VEntjjJS42+BMocfoMJTv3ITSOQ3e4YYNIR9bRvakbeBRY+ntUWhO5y
GNPP6UXQtVRj+GuZYc6KfC4o5cM6p5slC/exvjQxxcSkC6NWa6SqLoivie6oIOwxmIzwzYyV0j5f
1zXhloEUD/82L4TmgBrxHQ3KI7NnMcR9O9MyGB3jKhYJXaTp2Bb+osPtC8n9aAdVw4I+fNbKYwcz
SigGG2Q4V49uLZ7z3yu60HgQTJa82F/BkU9n6HXrYld5ewythP5Xu2t4ROxty19cHVEjXuvhMrgZ
0ZHkEmK+7rjmShPw672+rfkjuuWe4QzSnPAJ8nUabTd0BVTCeYXFcEyS6QavLon3UraGNnDNFxlW
E59MwFFwgauJcIiJXWAQsbyEvaxHNSkTJ6obDuZ5aeGAlPf9BzL3VeIoqorLNh2NLOo9QWW0v3RA
Wura2ooNUhz9ebpkkN+1AqnszL+bpEkBV7Kr1kFB2OIonn1dyP+y9JRzOl1fKRoGTpe9tlyoXpHv
LRskJWGSKgunehtpGSweTaV6foVjrv4WDHo9h0282Tx46uKl3yOpavIVVxJybkl4BNyemGPKrZWC
f9+SYxWCGjYpeFBvcXASH7JiWjz+E13Ys2tapTii3kfIaPBms4UmBi82oIeJZ5RB19n+0+0elLIl
p6VTuylbu6C7HNzh5vZD01EY1qKJrqc7v65M0OIzKB+Cg6cUHXckCFf4np7EAed6c1kB5FFAV5iK
6kHkKzI65wf8JadEjvt6CtDlAQauyfT8G69hTT4I8l0OgSH3m92jpuex02JSuoMqTkN9ZCnWROU+
RMh4HX01b6i5fWdfK/w/HlURkXAJXuU+CRDrdMZMP29dYNflyn8NFYGWTHqmWUXX47HLxnofHxns
ctZeuzRkPZ1Ywt95qwzC9iW25AgwNXzZJmwrJ8kCN2agRy+GZx2df9hGRKmRN0uPy7dWvehBTFZA
idDmzUeM1wyfwvFM8HKWVvh4doXr8mlNUE8255wT3fI49Q15hcU3SldrapnITaTmJGT4dcPG7GPD
1NlAVAeZE7wjIxrKpE6h/OjROJHT4Y9wqkIi68k+mGNevVUzH+de3u+6PmbzB0U0kIvp8RsOWwzc
PWPHbbR1K0TDtkeeGqClkEfHBzIqtSxIOvuB53QAul0EIUrUM//WfAGVNneAoR4bIPsEAIur9O7h
xETe4UngsUSyrmY0p82XjdCXrlvU8MXt5YxhW8uEx5fjodmOOzmBo7qTwoMP2yqmLrBHISqfoyhB
4Hu0a6bS2dlpqgpLO6GkT7HKZUeFF6O+jUGXm/N0GLojiBoew5sIQFYvMc2LibAcui8T9OOIfiPV
ZyhhiV0BpYt0eg6cAY4uJV0nb6M2G8hN8e427ktyqlbERIWDo1xP0f4fyigGXsFhvXmgdfGHMJG9
WM2hPc+EWXQdVT7tIiBevDS8IOVzcuSwXZrBz8G/TYkFaSNt0ouBcgtudfqnwcS6fNI/AMxU3i3R
epHJR1bXk4+eLHk46xqgfRstahQzGPzgWI8YxSO9T7Z5J4UGo0LM+5NtgC2mVyyOuCzADnTb9m0i
Puwv8dZTiw3TdVom99FH3YChqs4QZif2AVnlBJzpcVg29Kms0InxjI/PvSTxiSk1qOXbPG813eE6
RUMqHFGDo9XYHb9yagj6aq424+WsUR3A2qOYJnoIPzsoAY/Pq6RgqDT81178R4AKRjvcga22eDHP
E0V9ne4h7tFcYfW3OVcuFjmizBojD/BTD1xuGBCvnNJgkgbtnUKErlsgeukGFdeo2liu0b4ceiPW
E+2BBvAmCvsoFRrzhtGt5Woe96fUDs63t+UkHbCLOBDn1aABz0WDqzypqoBFCOxQ8mxC4OrbPRRz
ktWAOxEkxfnINn1AZGm4ry5NNHZUVRu3OE29DRcB1xe08XX+C+2KCSS+ZS1aKSf0F2fS/p1NzwPM
aPTjRBGBKv8Pe5/51OS84xN+8aksQ4bpbnkovC6z/hO42wIn81z8f2NsNuzWsHcHbpkIkzuBbH0t
2m8InwNzFgBQi0Hq8IFODRtm2oxMWy3dpP95FJiidBkaHCkHSe5wCqjf/mrhbMD0FlN7mTRuwBKq
i6JBVN52Zy/6FBpmig5EFkzSrxD9qQ9FHb6Ay0EXujZEzA7VOQqqSEjyaYXkJBRYydQyxjWduXBa
KkKp1QXXrwnMQHHMKdxbUqXnNmFJNiuw7Zju0p8IFRytoa2PYD9YsvOEl4h8S832DTRm0Qg/Lrhd
Ssb6FJdvotR0NROM3nYaF88eZSE9e8Yf6b7YQG7EP35w/Upntwe4GnMIvCa+UwmQBRVcVEvUxexp
9jfR0B93pdhyfPsIpoPHSjyp59X2AwyvShqs4gFirRZRWTDONuILPoXZSTZ9p431X7MGXKiaBqXl
J5AZXs3FQtlDB6ZMIh0jaZYhaJf5hRs8UXyS6tne5aU5cxxqh6AemwyLBvlELP9gS8UlJfGVaPiP
M9xbNgSYx3ulGTR4wkOUj2GnCRBva8zn0lqFeYsyoq8mTpg/PFVsEJdFEB2dM3iguZFh7EoKxfer
zg211TPtzcYXA8s1MxTk95EGhumGudlZxpfMia6o5fwNvdtzIOdAQVZqDKfbomQlBAdG3esrJwET
lwIRgx0nsm+k2aYNC+7d3kW8GfF4SyiErSfKPVEkhpJ37DkQzB8BvtBJPZNklMMjg1pQ6uPum2OZ
b+zDC9/YM+vY4Fblu8chGJicaQTCOvHAl8FAbnft33lTe50+UsS712DYO10XoWMocXWCIPxz66o1
26Gf9e/8wX0raTy6terir9zVmuSTJ4teJqSGeammDyv3ibnHlOyNypGnFHNjN/i7o7uJ9VY8rCpK
ucGV29Jewdn533vBqzajKU2381HmbAbBhVIx0JkxbEmae52jbVuNCWpP+CV08zFT86OtXv1j+oFl
fIsdR8ud1fvpZF6zzZwcCs4Uf18eAn+xlMS2WQPQh+aVOYfzyVK6IonRdpEoRAuviO74Lxe9hq1I
3ymiLpvKYq8jYOGsG2dH8u2Q7IV7CZG80HBZCgDKCUJdf49h8Ng+pTOoI7fchhLiUu+OWTk02h/V
OD62nas/llvwbIkcuhRjukyYqHbARMSbLGtzBQ1k1uYZrwkBXC1qFVO4TeDEX2DkmP2EeNjLNv14
1KDLc3+c1fcwdJ3zBt2l5jvNiOUzeCzVzipnIEc6C4ojaMJe7hA6CItYkoK13gFgCbeuMmrSWO/8
u9MwBxysqWMFNbVjqeV/kw7bqYFthuDQdg6NkbsGZ2h5o3scosztLf8wLz7gHYeV2seJ5stWY/8r
nFcXBRm5M7K/EvmRVeoc5CAhg1cCamFI5KScq4XRZEGGDjip0Bq5GJ62natwif/JcQxLlYrzXLA7
FOQ5fh6kILHQKwCncxugXqdm4lKbyLYkIqlyHlk2T2Srcb+Dbfk1pTqCPtbaTmsF55a/ruNZktfj
I6EfJD9PsP+Ggn0Rbj9OwGkKoFXTOhuhTcg5Y1IbhiRMWpCqikxZs45foo5t7ft0IiEcQZoB3wj2
rhQHdPqUjdI+fXyatYpVZQk52J94rEX8U9ua6mvRBxQfaunn3FywIAvLPrMWlW0Wla0LnVzgsXBr
j2F4WBIRW1m8PqLq8iresMmD3C5MdKve8I7tqKSjUqNLWPStXRJZ0bSYflkmCQpa2IpZi46GEHys
YV9O67d4nl4GxsxPMeZfjf2X73bKDqV804aJdydQoLn7EYjCJ6VdIAwQ7EmURsMh31TquB2lNwDj
facU4VAkMjUqMsSFjuNOAH7yxD63WpEQdPd19HNZdBko/e58XFc52CoAycSKaiHlwFma7LnBVRtM
7U2NQ2USWJayPivSI4meyZuPlQbMYtHUdeiJ47nbXhd7CDjmaTfS/kkLnupZIMHRj/xTIhTvHMLZ
5ZTdrc69u/1Pft5/vTdzD/R4bThYbq6SoroBeZHc96JYMJjaEIhZF1XunUnrwGOhhRGfvmMzxvxl
r6D4llWxWlTOasUCM6HHx6hm/+EOgGJOg17zzRwMuXHXzgqhxp7sc2J4HtPTHyqgCYYuWI8TbcpV
zj9D9ueevX+ziUBY9hYqdqxtpzJPB+yF6aKlnNdwP1bgv8ZL5Cbc0/rcD614DAU3GbVbahNVja/e
edzeNOV56M/ukdejdM5ITDCyCQlp7d7MJ3Yepr0boZkY3Y/9kyKFe6QWj164wWmh6n3sVEzXKHw2
HBUVPV2iQCQIGnGkcsYrugTGYTc4ELXy63fL2np4DlILQS2KBYd2cRhWjx0XGu2PxCoibw85pxy3
P8eCL/U43JQFl5N0xw13PZYNvJCgiWIiVFKjOKTKLC7HX0rI0MQtSdVN7oLkQ8r25ho5Gum+1uGP
Av4jcHHbfPeCstv/c/twliiKhbvd2rzU9cYqnOe910WBFS9V+2f4iw8OfnyjWrihoa4SjPYJK+z4
V0nbA4LWODiOXTZTRGryfkzbkA44sWKgq3npluqkKfgYIwVg4WGkjK62uyZmSNAuLcSxvJGyRH2P
zhDOEKEjG+Keh1pfe7FJBZr3a/E8U5VqQfEtYnTltTAKk+dtY9jH1sLiPkdN0/Qa73p70uq0YSJ1
gfv2twlUsOvy7P+kahJp9/lXE3oKazyOrtp2+2pGOBX4MwNXO/gmnco6hLd5B1p7/UzUSVZfuDMp
dqBvD/R37xzkOytkCMyLC96ufRpb+McX9BrCS4+Fe6WVkwKGqcZeFUp2U54st8xmG3WEE1xbkp74
492VqCeueWNnYWkFRhN2tcjZ2mnjUzArM+DvVf5sdp4jRoPxi22idJ57r0c2M/OsWnszHFGTzpv+
ndAc4mq4LuPmVA4oPEsbamOXZpFO3enanWg+Pd7Pur63NMiYz64tFb75R1V1VTbzE5CVpGvb4R+q
i5C31Z2IYMO8wLga5QAe+JlLqFCWa0hIC3ZpKY23YvmcEJp0PqT2UYwV2yIi42RjaHd0x9x4T0W1
BHok1Acm4clUGciEicTyWuMhVnV0lHSEkQTa1NXGaP3WTBPHe+nC6YQZYLAHJEuvrPmtYxjbUJP6
CuvTh7T8kc8nr7FQtwLogLk+AIOMaHHDrp6HICvOAooDX88jAjrOululD1ToqMFMK4gOm0VUJ+vm
PDCXJRSuMHkDK+iodjdpbFX9HFfN06LgLV7G72ffuqxm+JnQG1uehK3+6MC71hQM50M5mnatwugM
gjKGCWyp8DjalKbiXhkNavylPRMEBmTHBL3QKH4jX3HfPgS0rB1sxZjQsEVPtVeEHdAXg62U1GTo
SLeZlVdu6VJgoueuaJvzikl0zDV2P78RLLqjN9J4MtcnOhRFWZ10i4HcuRgl+iN0TKAwv7wMpr+K
PWcI+D91W+A90onrvVFV6dhksqudO4/Xv3DfcrKK6+KJ09OolQs83XvR6A7oOiP4RsahOzfV2QHJ
+9A/gOvVmhSfA0SMiwY697mTa7kt2ztDyOloyfu063bNCn+Upzc3oR7jB7ebi5lLiriG3R+IoM5x
43Ia1U0V/zG4K4HthUEZDOa9sTpvqvFcZ/Z3E6hKI0lLTT2Y6uTV19LeZ5OBKs+y1UkULDMqfssk
h7492vQcvq1n3j+oiwNQhGlduCK31afF4EOuHUbTfLD9H7Z3AR1Sq8xkAPC/VoN6jHkaxbqQsfir
4p1NCeA4a9bmgIsjs+nY0ARroPd6DbU066qsupSX58ybWm4QoRpYQgXs+60k4SImprRW4/8kZJhY
jV6B0pQtBMwEtOE8PTfnkhVg9y0esbNGbPGWg7Vrypx4NyjBUb2b7jKOVcwHGTQqfpsec5cMap6y
FUSvwTnrxccSAFFiR+lDgaDuEmvGcUKRn2ehQpzXSxQDBTruD6YCE8OH4lwjwayYdcKOZl/QJ6mE
dd5G2HXyApkmfgNRmg8Qav2bilSx32K5HKNZ2B+kB/YyNlK8yDMHuqnkpE8oHisNto2s0E3GuKt9
vJSThH7AOZAeLIFYi6mWJH2EJXWZtsBIZ6kATEl83YCg2zulZUP4Dm8ejlwss/lAqMCsUZo5zZuV
l3wQ/SEINdYIU8q82b+ydzyvoCF+tBAYLxfJEn64cWPY6MUw3f3S5N3yd9i123fVBPpUTxTSTjBm
szUnkTnUpOCaFzL4Ou554qN2H8rHVPGsxg7yii4bJvSabM86KoppD8U6O+joMMupzDoeAYypdoce
ocn+oD9fo5H3JNmxLbCVv4/Nnzg447R+VUQ0G5Xcboz3hDHD94uA7PYkwYE/Y9h7tamqZavjiITT
5qYGcnFK47Ln0+jARkys6CjmfWj0qHRUmB404Teo2g/uN3sBpahE4zqQYmJWWVDd+OnQBN39lXEi
AUuroa3WEtGdEjjst+rU4o11W0yR/XAop+AXmkWJV+AVjRlc8Om1A0Izo3jR99b1s2Xqa+xzD2RW
tB6a1s99ZWLbHjBhbGFLm37TVFJLSYtGF0IviKXt4ASEHMfqtqfLrb0kBTXwV0ewedJ2Y5KUEIxA
j3of4HuUO1/2Lg5JJ9/Og+OdyyALhGzF+Kz9YzkhsG92aGtcHMdZ+DS327LpPkVm5ClRU5V07wTT
6ctyzukyPp5eYfTbv/iiun55hkvM8KdVbcAfMt2h7ipNpkKTMgvv/tXqjOAjmj4RFCBNl9B49gt+
ZInp/YpdXLYDwQVVqn5sK6UJZ4Gzmqya7gInExyEBR0Nga9s8CMYpDh7AZNHlXujWQCXuopu9yFG
7ubo6K9jd9gK9b5BggfKYyj4ts25wOjM/21PBDzGi29el+E01o97Hhh2XAcs0Clj3cLheKbH3d0G
bbDBl4PLWX5ziCmKXei2RmFIt+X+SAQiVffuj/D+yVzb9r04uAMleHzrrzza//e3VuiQAtxWTnJd
V11oMaygkCQ2QVvM6aceOjuIBe+ChJp4OWdsQ38jdLnh2OOTq8wtOC2YL8RYRNN9W1qf3eNqhPy7
DLmQYDRqKR8dqZ3pOFSB4Qq90OuW6DzaD83bWo7t2VYE7ILIAaPIIgIXHO0V9DQnim9L51+f+c81
ddWAMzwih0Wv/OcozTd5Z3Tf6DaW2Ai4wKYocICO5y7xMG/iKWNXw1/KWfWAQ9Af90QlRz2FXVe+
gPrPHQLFV7MdFgZafQYgeAt445KYJTRn0oL9JHhqFExnnSveiUoUUjGt4fNeoHcvpoht9qRuoz95
C6LUEwuDmaEY5nctW7pJVHtnLPKGj9286sU7vr7XGgmhNNPId7EDn0YnkQWU8bZE6YUKnkw3DGvh
1KYmHcCn+DrXQyTnfDmCcL7eTCI38bJmP1Ix70A3R63mUrX7lnvH2PvMhhBI/0Vsio5dfKQTDxws
yoN9pTR927C6VCXf7YhO/BeuTbNUHNH/5/kX9H9ozg9y4d86r4M4uaRvZoOSCpSEJwPP1QTVQntQ
+NupqCW/Tc4RR8a1HHFws9+oxjakwtvamf1sNkIvw6PL+WqjJAi8AM79kgGzQ9LPEuE5+xvrhTwo
fuj7BC+a64726Y1+uHP59iEt2NKih5bt/32REHgYne73SoO1C6FUOeGwx9FMejZAMWN6vBiigCNl
WotD79stvglAubUmduTYoT9bgKudDmiUPVed2WTTM1hm5dKA8tE2SQ4nNlKE9FaWnDoLFpYCrOYz
QyDExUmRTkOBEx2MFSsuWc2K7RDvQkC2Vi9Uk1feDoP0sLYFyB0X8amcAJsgJ9zxsg6ZlkAzhEBI
V3nV6PwkuZqHxmlt0Q/Nk5lCO1d/FWwj1a+zQmGhKOXAGm92xhvDWQviLtK+l6pDymixOuBCTw0Q
V8kHmS8Q/KkwBvcOGmfSyZdKlWxV07synCOUoQBUuyHxkS10VM6phbubAe9Mw3hJ0zPTXvpQSP18
rT+zmdSeFcmjF39tXqO0FsF0nBtqSQQX55NVhdlO4arZvX/YBudIR4pIZPDEeLtQaQAvml7Si1zi
TIeaKnNZaudHgUX4StaK8kiV0mDyYXkVvjMtLDkiDpaDplRRl+5uU1wAizfuGFPXwGCSr0EJ9YyT
xx3U4bBjoTVMjheUvgyJllulaSdWND/YqqRxq/18vUV3l4+bSu9LgClgnYiQPIt59XkJnJsJ6vV0
TB1XzJHrKPE4CXrBltOS1W/S84P06CBfFMeElEBzuE32HnB3QJOFKTe91s5GiOTYjAcaVuqtDXkG
ZOQYmugVxYxwY4VzCvGvlEWVEZKl+oMjCX/HThTn8epjbUAnh7JjmSz+CVZ1QmkPwwkZwZa+96RN
I7XdOctZYsfeClkWYsqcVUJ2EbhYdTDFZn+oItu4CVqBDuVJd12tfJwAb6RjqOVAdlEzPC3apRGV
bLz2PbWzKMKlEfWFPhzQHHZ/XYA93HyD41uQ5z01BPLDu7cQyo1pFt8EAsomrNI1+q6DJ8lmNkRQ
Pl+WYynwrdMKzlzvJHl49Bhna6BYQ9PVt/wlXRxgvpo0GoCDdxliyF95ve2ExptbqqR4NN/4IGN8
O+m/qHbiIzsamg5a4WY7z0RnNKDnj+OwrPP2Julo7SZg83jHfJq794lVd40jt+CUPgqN5Fm1ThNX
nSaDALqXa6o1eNmLRe2icwyeony7LssmvXqyvM6rWbgcYyK38Cpx7tRJmI5NUEMIRYZIIjEbDCwi
aD6sR8WJWQ8NFRRBxA2+332H5gisjGrO4/R1OVzuUN+Ia+szOrh3PZz7OYGtl+BEE22CZlPrxmfw
qUn9YYpo1/N0w0F9ag1/AGyojeLUB9BigoBANNCH4jIVZB/0RXULlPYBxySK9vjaTQU30s9OqTIU
R5BEmFOZtOU85Zt7iSujS29gU+C38+rGjVJ76f+BMITrDz6TQgfVskLKH++CUFgJEaAxu78mqydM
7A9B8xfORl90t6N2SXZ6sf+RPsl6c43RvoFqFQ9EV0QQibc6UqNpeDQec1rrVazipJJhu3IVMFWI
2NYq9GQ9dMe1G5bz7G16F68pdQn8Bnf8WG4wvnF8B5D9UWeVssYF5c+0ey7lwh+GpjSItyL14eOu
93VHagNOHAZ1oWIm4UACjiTbyYDmo0Aa7wvjub0sUwxBU0739hNbJzKJi/5yZzvz4ZmxQ1lL+VfJ
dX4eAizd/81WkyEFkscvYj/prlgPptqXoWHZaMDmaIUKkfNwY6BYtAEm/ybnxHYX8XGPiJ7z+G54
nOUFOTbZYSTFttfKB1mGBqQh+zsTUuL82jUEokuuhfpOgIS2RsIWwoXF6KohQkzV7pKkTvwjm7Yd
QY83kAA/BvfbGzLY0xcN3RftzqRhOyyUtOI8RW7oPpeAz3oao2hoDw4//KgJw/3pBn6dDKXXMGu9
wZRuESUcehRmhFHOEg8UqwNUkg6o3OLn0yuyZg0iC4HyUhDzZah3JVwdNhh7a1h+5JTo7j+1e6y9
9Vyv+MhEARWJqZuihdG7tEl/dF/BqxCuXQtPEO4Q//JYrlIt8rjZmjoIwZiSgU1XvBPz8cphuS4w
KiZ76lbYu/eNjxMzQ3wYlO/mABkfdW6vpp+7mhKN1aufEC5KaGND0NX1K/MCXVg7cpOOjxli9GmW
CUzy2gmSKOEorkI5/cgDGvDZH1gBqCgIn+w3zgQcxtfAG9b1vX9tYiHXhBblBVSXDSi1G+UFLsBU
KS8EbVNQnBbKuQ9bdZYZdrbmYHvBJG60hkVtIsI3iZtd6+aDA6kk87dcjXjUj+2J+c3kg/PlWGDM
0sw0ohQZllKwNBBtwdD4ov9H55W2AHCydYDNPZfTBRNNa5e87bzcxfF6yQC3iTaE3eEbsAr2jI4R
0c9EzbbhEzQOCguhTZf4K57Vdn9KOJya+UzvZkFswwGu1+QxtfGCFn1fXGNhpzAObXdGwfHXnTL5
RYVK+ONDKa60vnrhkyCPUg25MZqOi4Y/GbyxDhnxrLNyFt2YdvP8rJR7qwS7guMHBNWrCRsPR874
GFDITaorw3krUcCSGMYmBL0j4vbSFbAAiLufKPrjUc3b2UEhaeGo0OAhulj1Oll3K3pdZ0o7kGW8
PX37wnebPdGryGFW6dUTuC9FHZhA/ol3s0+nIgVb8w3AP+78qeuNv7eGci1uCUREv1qAgHIJ1MR6
JZ29eLLlv7+C4FM4qIq01Y1BZVgViEZaAC38wUE8FnR1mKLztqine72CqWC7iMkv8jNYTiCWsVic
fosEfxF8ZT8D03Fsg+xq3NwyXTo5QVB89tIoYpuGghTjm6sZmhRN1ZPAAMxdXkSAGLGdA2s3/e0i
Aoc1uiZSk9zdYH0A5pORN3TDYK6a7p38pjG9tVyyKHEDBkxqJQuE7gWxqNdhokE975rYgudoGSRw
kFoPbUhXcBLa+iwQQ3eVzLJMcw7JNXd5ZEBYVK6D1lchPCn+wokWlSFHEZQgiQMqxrFnDPnadzOw
sr66sUMAg9MaQioCfdZ0UmHcgQNke9KjnpOgj0/8mlwSxeZQcQ8UsNMzPsyjE/7iUTW/SwLj4Zic
hfAk1cN7L63ILxUALIJwvEN9ozOABsxaxsNiZi8nnHb/GGXMRHGBaBWbArEF2L70l9GHOV4h3nBO
fkUQ2dysKzKziMjI8fg1EmPwBZ4PdHJdi2AvNZ3bKT7peAmuztefIcQmmgVuRBh/AA609Pkw7EqY
Cx6NCYog32NiCp3Sp/ovJJslhEBfjM7QILeqV9lZ3Al9ONh/nGoPWR5RnwCOWsnWN2VCRPyRVRl1
Z97hkdx+UIdUS2PpzVFOg5aAQSpadN7jX02Mslf1Zu/+E/fjfegunzimdM/g+2oTKDncBKWrcnxE
0TRXSFPyMaXH05ogOLkHV1gqM2r9XvQ0H4m4NBT/zluYSA8bXhNSjTiSJZo4bw7n3xAxxBLmeU/M
DV6E1MK01B71K7BvpnYvO40l9Q5iAII8aPeciO1Hu1rO97gwX+EJJJacnkz0LzduVHHNHS8A+Fzk
TRYZmGMbaPDmZq9vtnJ+LLMUk0mZ2zrboaTcAuZftAa6pXilF3R3knGNPIr8ssgyaGzarKvcHnGC
Z5+9OE+VsN0Jluv13MsiSpCE2gtYpHRDsP0N4Mt8nSwfGLuMgCfwy2mHE1g6yPXf3QZslU4KXzd2
xL7ljk2W0KlKNww7d58lxRIrdIYTBxdpWj7CZJTVxGbRJYcGy5X+0FFI3H/nliXHH/NwSS5SsaBB
Tv1+sAxjpgW3Es1t2JzY3oHlxnj71IWPxxbWpfousUHYo5YxOhQvS8UnlNfUsJi1b+KgFNo0Lp2P
cjRLJPSMiiGFsnDyRdVE+qwGsChbzT+xk2orc0TnvIUpepsNoqb7UBv0MCLnZdqCdRpRVidlWvSA
kWQ0eVxV+FIl7hNHtaZVHubUkCU5Yjc7bCqKGbhLUz4NKxqheBc7bfcCxhSQFUbo1pcUdW2CJfso
O4F4OpB0dDQwHCMcFBviNFr+QBfbKMKfCg+eMx3zNdEhnHs9cjlQwX1I9Zqe6R/jKL8LOA1UZTAc
Ec/UA7nozQUR1LTNZZbGpNV8UpwmRpKh3bhSfTNBf6618yZI2Yk6TCR9Se/8uKOj8B/0fbmwVQu+
1wq4hSTfI74tCbyMjy/BX0byXame8wYjQ4Rc4e2WG75ezWjbsRErB/1vXUPzf2V6WH9bGJq797mo
sDlIxVFeUbS6pf9K8X030AC2teWUMlEJhMVClH9dDpv5pO6dhK76y5YuiDmz61bl1rvPn0Wo5JN9
z8eQ94KNyIM5svhnCtd//V7Z9AzjS27SuRWW893MuRF+FRL+scoqjwSOV2Lj5klBDnsPrR7J57GA
whqWhYJBL/q6Ngy1SeVj0HOg7IqisO3j2i2Ga3Y5EmSOFBx8zHiovqsv+fpIv+Xrsqiy1fI1WedK
36JcXQWE9O6hinE/Vvhn5I5pRSonuss2MzBTqSR6fFf4x6cSFys3O9dYdW7rA/bbRs8rIffrFxkT
s+K7JE49779uWnWJ1Q5bu75ZnDyH896btWItJKMtJIYNzu2bXU74en1z7Okl4pQiB5ctMW7lha18
29KxjIbnTRpaCiBVHm7m0BqeBWmYrI5Q5y0xWiUC2SaInjEnUDPc17XTXG8MxU3zVfmFOIAtcNH5
/nbpbfA/FG5CYzZh3sgRdflct3evaxTTt6EuknY9tXJyZ4p1SN3WefJE9Rjb64MeGDMIM8F3cRhZ
TevDqSlcHFh/YqGPbSA26M1uv38NvN+KGHmb3mTdGRqQRbsjUgm+684fMgJR/CrUqQwR0Z+YASI2
/v257f7Qfx/tTnPJv0pT6Od7ihpQmi20lB0/SnT6VMpuFLhm3UnDwM5IcF+UfZuFg/iUAAdz+b6S
piiQvSJkgYHXgtDnUI0nKY1qPElrXxPxWfvMFMi0RJGyJtbPTQdUJA9CWSsfhU9pnuNoImvuRuZr
NK64IQDLpkQwcbGLdj9OFUh2E8DdfJtOqMTZ5PJSWmbNhcLRgsMxpsOUT8AZpBVs3+hVR+IeJqBv
XLam7aob4eVoKCfPkFT9S40fqyMBswqb7xNMYR+jOBstuJDwZf0sGgBGlTk8Qi7mgLiUpK+7Xqlj
uG8EAZqEJE/7bVRBETHD5D61A/Ez0tUNywupXkSuyANeBQHhPThDnh6VBb2OxiaU4kL8Sm8EQDEU
mYAM0P8EA2x90pA2zmOeVuQjISGaLnfCi/8R1+6nGaBwMRppS4e+HiBmtE8b9c4Mbr7BCe6kdcLa
PRuZDRRaqSneeY26GfLPXIvfTVSo8tlLMghzDrm4lNMqXiXbiD7ajrkVm+zrSoXYzCCJVcnInxO1
13KzyevD9cwsRxGuDL6gY3rbkl3ebn1dchOCxBGROjHyBCIszA8c9icF5KrQkJoAl+tou62PX8+c
XKZcxhnwPSqts1nKQvIkuymVRYuPQu3u8rZMPr7iY3WAUIC+8HQ5T8NdK7XbBAq2VRAJq2KQyG/I
kITqddbEek8lvbpnjgu1nBPT/i7OnaSh0Wxvm2gD2e/mG8qxGC+S/OYdQFQim5lum7PEjTmZgKdu
i4cfg7foQqjFQgx+X8jbXqWq546HKdohgRCuBsiV7n9OxEaUwAPkyu9kBIQcDpy+kiQKxobwn9/G
nmUHP0JNBT6XL6+l/FLesyZIaAuMuGqg1RvzJv3RyQ3TL3HtR1Ao9vnzCrMZQWDnUApNtaZaVs9K
D8tf/jJfBG9b3jvb2Sl3Z1jMVAOQUxA2DW4q99aTcYqRkQ9TpAYrb8siSODCHMCKAw2qpxL57xCx
y95Jw99oBvEXY5B5npimzWMGEjJfMFbMUpKK4ry4p+ZtwhFD3V5Ry7cUXTytvuruxmjShVJcMcy2
ANaj72KfcLCUByeKhw3Y+AHXaLV7ETPCGyaZ82DvlSL6hE8W987C0iWEWYCspTXptFyoHWCVVrfW
+ebM+8Y1rm3fAnmejZtlCJn2r2FmAz7QnpEEicEAYfzWQ3ziUDqG972iFR+O0x5jzTaluLuZVrIc
rZeTVaLh7QShMIpJzfnwOBZS5Y0VEmGldz+/GHXpZXqTVMNn+a+u1PGZOKYpXdoyFFLsIr/lW3ja
2lw72OBqwuSaGs5+bus6IADNxF06XqIg+U4qyCa/K2dDodG+3nTIRmPgnW/gg+HB3517lfyraaD2
azHfYNvIiqn1+qNwxttaRguqTH4/EouUzyz34Q8pglOE+8c+JrCYXkeFY4GiNaZD00/v2LlYagU1
hR3THlEBNIWnw7cBpnk2Pk34wkFjmjra/o/rOt6hITtSjIdgOjyIxu5Q2w+Np8HsU0k4Rp7mVt/B
O14XNIRPh9juPsFo7MJ6AHF4UGzrXvgntRPWCHv2bwCvYs359qEQHMNvonBp+Yys52gE2ATE7hvF
3vMa1rEqOgmpEd7QKDbsf2NAkGz+B2CIOaduGBqXevIudl9uF8DgRSYt0KcoEhFJ4JeoikrTUyIW
3EdFU9h4IgboCXB+SXuxK8Dntw37QOsw7Ohuq3I+qiZim4da5filcDk63GW0t3vcpw2eJiEX2zai
0vA/tyuRb4yKGtNQP8MzGpRWNlS2BNrnQ9zfsNo1pXrxHcwafOrNdDhDu3VEBLtxkj5OEgs0z6/+
+syebOg2gbjUaS8s4qH9Rbk4Ke2MfJq/jbmnSMB0xSryy1a7OECi3zTcYg1MkHEY9El1oO89V2FS
JQyz5QIbns+LBPx9gqqgmPsl1xPa0VdunRxuUo1d0j7841ksc8bNj93vy6mCWbh7UZGGWgpApkgR
ZMFdZ3xgE44kp3KcTPj4Zs4jBsrwWgsonRsZN8Ks8859lnVmX3aNAcOhJ0j1sWInEY4w6ovMAeWb
JDmPIq/Jnn9MJ7JhCyX6zMVijKrUbQKAJG0Oo6HREULd28L7rL6RzlAlXc8n78eLnvxCtL17vadT
IKiNsuIH9gRBaC0D+i8/qHH2PS0SAj6O5yGMtO3iB3YEud58Pn0NjHk4f6Iljr+bN1kdWzYflFPQ
s2M4ymrJlPksaghpCdgJCMh2hiJANeiVA4sL82pWrh/ZufOF7zmPjyH9L5UfVORkmZ2zqKxRbFPh
IQgwUZb/0ImGAwtnTz3Ut0r3VQipe3VI+Ctr0/Uwj2/Xswjnbaq/kiUu5wb3/VDZPXHEnZX2lsyW
cjXaSqaBhmqm+c6RGruoOCHc9mws+268EUy8bvEpytQmMXTxvu+TlsRHTEjsRm1po+tqQXI7xX+r
QXKPiXwGufeoG7d5ZnwjEJr9ue4ejvMSJnKj/SX3thxU1hWGwiyxyHUvoWmddoLVuqmYLmthkQIU
PqXBVHt1pfEuZBt9yoaZzUnxpUM4dx6Guavw8HJfHTyS/4wtKKjFIki1xcum9AEKZivRD1URCoo8
Zd+JzrxRqWzzsAKEPSboQGNlFjmRy2H02+yVATDFqWQMi+SHzLm7qfwiwSzqi2b6O8UW/e36ecAg
QyT2yuysa1oiv6CexrFcicMNHXaUpMLSCQvHE7+ljhm5XoxPx4x/Q0qzIZnWkDGdGawyzTIZefk4
2OQ9WDYNAktpJhZrqqZ++Q+ZnJD43Z0iDXTRzXaUaGk4tRyXI7Ob1bsl8D29p3PTw623zK/pNGwB
EmwhiLdYMznZqKCEBCyB2pO1A5BiQVVfk/dQxI967AGYMeMyiO6TaPuGZYF+/ea0ZPtY/3y02Z+K
F4CtZG31+qPtQcG1aXX3p8yKB/9T4Abjoy7uBJdmqS/mYFhzt9dPMsdjsx0a01XKul+/V3g3T6+q
69kZfAqyfPc/00bMDyX2qvZFfL0gWD5cy4rRXHpfobuxowwdOc0txCZ3eXFJ06yFfCRPrjv7OPOQ
DMKs60+70srp14iChf0vWFVxNWedu4/v1qDF7oUMKb3A8aVr7Uk+Xn/2s6PhWktjzHcD1w4S0Ioc
jn43r5xccKYe8GWbANLtJLMruzasnOc/qx9Aig1fzgWULme2eReL9bq8Q0EZcnlrFO546AT3GIA+
7/D1BSY9LyNJAtLvx9avrsyhp7Eo2SSP9sTtvGVqdnw4vxp4URGuVL7sk7Ma45M5J5/F+RqoBqH/
PjWF8Orwm69ddRxTqq8xg5RL4ZH8AEZudqJlBHJLkPcbTnKEmz/ueX65EfwwAsj/WiQnfByQdN9m
8+DYaPhA6EyNgcvPZIb0AedvutoQvG6vND8AzhcYo6M1rZ0Kvz1lNeyzzlU6WNXdvvASJOsOHPT1
j3z9yvE9Cn9ZAKBXl9o4aqLtWbydHMW0bSpj9FICMDc0hSAoETVyvHGdTDbq7THrwzQmhK1x14ex
BDaFnfNbcjxzBQJuWPXntH9OeinR4PyNR/lB8LQ5VSpvxD3LfTo2YQXo+FtqP68f8ZZW81rwN1hm
v75huP9JOwbsRsjtkSQIwAt5crI+tL9ATq3YCv+njXvN/Ace9uuScD0HZXbPfDoMP9tRk68FgQ+V
YcBWxEeq1McYkcgVIzo1fSBAlNwa4Cc8DD+qjVMXwZ7AZXsKnWVxlpxbr0Nvf1NzL4tEfdxfXv/4
zTUmyRfzj2mhWsQAu+0u4QboGkTyWs64vOvHpqaAaBBgGn6RHSuzyxvj5QnkQ2eZ1moVeuGcw+XX
5R5i4/zh++sCMbhVSPJMh3LSSfUdyUwQP6SJuUkCnlfupBynq76W0n+e3Gk/0c0+36EFqJIypFwL
1GPRY0qYM+2ctGgSiBOzM3Qo/hZ9X8tZ5qRslWy0MPHwMuUX12Ozow53ScH8eU26x/GckKybJFEI
8TNByAZ2GotJDhIVnebnpQsUSAOoHbDHXATfogAzYtR7MsuW/omfx5XBSQAvpUJQqik8UFpyWXJh
k+BtxyRDEL0yHdsq8Su2Cis/kX/7785o19Ug9H1mAPcSME+PlQi1Hloq/MiiKwSX3MODYS+7rm0K
7vjgAzuPf/gyaPxVEjAl+pJYWgf9GrSwoUUNLQTMBg7ad7m+QIgRCZZN6yYMZ//JI7Un6NEKThKI
O1NJZJQhwR1X69CHXMDubqyVjVi5zMSIJbzv8/ypqNuOVtKXnSNz4JpVvCsQzIcnPg7oCExe3QMG
coihCWMiiAQUqfRpPb/POcYMxSGWXoqkh5SpVHip61NEHag9Xpe66AdotuMEivi8tvnM/Cn5xMXG
sUUvTIdexCN7NgtiYGb6Fy49jWEOKA7IpXUxaNs7m+7FMDHugbKcyiB/XtmyZivxPVb2haawTg+n
jPjh36EVAcA6464GSm/PdNJjUn81Z8nuYx2YiuYn+avtNGuZoYs1UHdKKmmzX51uVS7lkXICcS4D
3N/fJMFs56kSORyPrdyU5twKPscIIFRfwvT8t3LhmjAutoSRUNvJBV1O1HgrR2fbu4iezvlZ636R
3wGRajX0e6dCCTLeEdHJbAowC5XNeod4SmrnTJnScjwPMwhVFvBka1punzj7pAXI0yJ20HHhFY+q
iu8qnpeiwyVuRn2fSAoKJQIggGqm9nJ4sJzZ3FKuUu5Lu4Xpg0fb4vnm+yeKmgLgsGqz3o7lCw2a
tOBSCpzIz0aR+D91lrdatQU0+L6FidBGZTCUpO43lqW4HIz37ZQ7JSCDKri2iJyQykNiXGMrP6YU
Y2UujKPJo9Hg+ZOED8L88RoOh5H8L8E9C6B7H2Mkj7rjWWbZ9K31WxhjzaTsHaI90K0DBzHqwhDL
cGQXkpDm3cB5YWyBtFPKZ8cofusxsrmDjLzol27rBYVFP610skwEDr0AdP9OoI6DK69wGV8CEXBw
847bXlDo+tuOEDQdVk+OsPS8Qc3bh+Ra6Ihfi1NF/9rxyDR1N0kbw4OxZwTlyPfCI7WY2Fcygj1P
VKzvVBFCaM0z5Fp0IN9lnEMIlcvUq+cRxoorfGRwoxkw8sN/nd9vYbrGTbBj2r41fla1eEYZY/Cv
YXVIoWCiXYhNAIpJUaOEruZiEDFhFaMxi+gxuc517FfUbqVPLXfajkjQFfcQ/Z0wHj/hO5r3zjrb
dYcGRvlr4OrKvFa2goqWBwxMxtUJTuKUbOiCP7MduoD9/T3JWzyFbsmz8j0x2lOyB8Ui2VU2BDyf
9W3y0BD8tQ9jWznZc8q3J6LsSGIxa85Thg/sBZJYVN45fRduckTGmFmL5FgCvriZyvkdiOrR2bpN
DEkZRtO8/8/V5auMtc0sw5PnPh/2SQKSqrBMBijE2aTYb8h6GMiCY7VruT87SlUvaf0lvCtYuvAc
6rcOYG29eNkB9WgrZCpayHsSFzm/t9Xz0zWBsDJ5Q8DglfVfSmxpJmQ3sFCNjTvMJFMmsrCfdoQn
3Dj03dhcZwJpqJbYn4Fkt4OJxE9uisQQWakR+yDboRzf/wt97K23vz2xc/R5YEwcjXIWc2uHWfNq
saQCZs17CRSfvSMA2eosoI2N88dm2/5nvX3s0LLRRM0vImqLan7ZyIGnLXbjI/rd50jbat+McwHD
Cwk2Wmwy+YLoktqI1SUxaz5eDBkHh5ZxOJ8Fudk8OT2/sNM7ndhK9xHcSbrg0sPMDWPphPLca9rn
UlX+hhJPirVKfAk0EgBMqQyECBNjj+Hkc8wEqJPAQhpAVIDKq5OoEptaNSJNoxLAMHL/y/kkvYSf
L6p9N6yquSU3nDEXZoH11cTzQFapIyoVvlGyPRw5Cup3/qY6HQkrHn2EBYwXVqECbu3O6lL+5T7f
DKYdiyMendvz9UoyOgRRfq+PIhAtW3Da0EsvRIYhZlfY60gTXXTFUb4wcH8b0OKEa7YpJnFTXIjG
RjzQ4Ex+83FYUGTWz6Let8LUiD+afpdl6RK4rDn9/QgmVwbdejQGf3d5yCRiUU369jAs6H+Gyf2S
g1wHbkPHXudHx32N4WMuA3YKMPN5LuRbZlQ2MyzfX+/dh8+3P35zxITGs1dTc5XEkKdwyu42/0Qc
Dr5R+kblHQbyfguF+IIzPqvRmdTLvHLOEr98a9wOyDM1XGqITdjfhAB8JNwpRnV7Omzro4JzRtXK
Bspoka4WBuWm/NGv0E4vfM402FTNIhIgA2ARJi1TD1MzG/vgNHM2FPJxcxkfzhQ5LOUHkwo39Ygc
Rgwd0AdUrtis3UJWDdpE7wONG8wTt6+YntQCAxLo9AlV/+le+AIL2HRljsOMKLeTeJhfNg7ETHPm
Lyw4cjZpPSRJlV3wK53VOqcYf++BeEHR0Gt9FbDiZQRqMef4zxxpF1ZNiszKltVKn0/96bFrf3nJ
RxS0IVzs2lDfr/Y8WTiS6/9q1n/qp5Hs5AECj30n6gRjs9/fbE3ZSSck/74JUN+5V1PTNQtgjs/e
xSRiVU6sgE/WzxwL6FVxcvu9YRfXSBmB8BVjTXOHWn+/rSPduN7aIiZgE8bPLnN268EpJY9Vcv0T
cDmfvLX8pEmoqkLAA8nCaqIbHTBxtZO/H0apltBvIPzyiJQDHaWfJnrCYUJxip51DEQLi5SEooz+
2MYMczNquPWy6M21ONu13xX2twZzwxSeyKQ1Qybzs062jkSVZq0omv844+kR2Ltiy/EkgL9AOWi1
0YaSBz98J6tOr4z95ECArGapsHYvQRT8R3/i7IYA6SiaVq1vZ51a1S2PL0K75+/GSCBWyf8qQjbM
ThYfmL0dBuUWHOrVqESKs/rf2jDjh3vuU8OeMi2VRxWP7ijxkOkAxdJAlrfFt2Vbw1AbHbwaynNp
sEE4AyIisiXok6E4WreaAOpNPZOAQ1CUi+vymujdx+shVdbS/PMEEtS19szvf5tw4hZBZYGWqUK8
QdcL1gyzcXn/vPi8AUm3ar9lcZfJjO/8+NSBOTi4PT+Fr0bj4LqXUqlUgciXQQRIZeyK/aGnWkGR
gyRGvMN0IHDS2JlJo3aS+RRVjhIYF+g0rEvZCF9PTO7NGM/hNXHZb6+ucGbr6kjxFAqXejg3d4B7
k+n6WAADOJfPrc3p9Jin5o7A4ws0P+vgXXH39u2cUinoq4F0LV2cf1R9s9jxWQ4ZzNjACEBbSEV9
R1WGpkJ7aXvqYQlnQgyhLZlWlIyw5XAWjIm7JMgljN7l+UodInJwDjRXCuJpWHFdZ56FSx29VjT1
TwI+050jp15EJ7pkUFLH55haRVZOVdSx4v1+YufT92APdsupN0QDh9iwnRWP3TCY6OsBWriJTHK4
Py6NmfGXw5/loGJpTQ5XSX9QkRBtcTFcJMI5v7Dll2FeJDs4JRN5yKOr0IEHzxA8Zn1LDokDz9z8
hvQmUe18D5QsdWwZUT0QzlJbHIddzvxblM2DlSH0hRpDbUa4d4BToyA6XzIqxZw+lfudwx5BHIaL
8+saropTmPyxRDtOxhwPq6lk4ILi7i3NAK5Bqd9Q173DqYnp/tpfJl6VJiaj8ogRKyO0ycESONNl
KL9wPhTzuXebeSCHRqEKofxvrcfZmSc8smmuwp+6x5ORSnQ6zzAbcnQ+uVWwVgiW0s6FCLX/Dl5g
znBSE7jVtG3aaCvQlIBVFzNhwWStEhIMkz5cwzWubkVW/G5gB5w7WpatSy4kc/+8PHzJwi3Ni2kQ
JxoBjWdiq+8iF8FqsckazFGsajgYrEq2PQ+1KNSJxTfAu1c6j+3lDlkXWJqwM+6WI8qcrQYLCcP0
oKGdpaxIIGT2TAJ5IYnMXd+Y329gm+r6cqb1PgatqR3xah3RgqW3ChUJpwJZWr4IzVZpJeE3I70N
wVqQHiCRi8zbQiVd/Ug+P1Xv1Y8aFxl6iQWIfVoM1DbFP8OSZxA1G0tFkIm/mmjN4wwk4Pdo0/cR
tmakxAmg4j7B2kNxV3BWOa67S++P4UpKmTW1luhywI2YOWy9A3qbENvPE+OMcnYvOJiCdZQ+u/fn
0Y7CdBqGm6LIlufV/AchyTlXQy9lP3R8oHRN9dbUj2E+dppB5dfhPAI8Uo6gt+lckHuOjGGMJKiZ
iYADJ0NzfBQSgEIQKj0+kZtqha7frkpIO6GancDk7K/snTfR+WZOBoEOpEYRyDafQUZgRbKSDeiH
5oc+eLnnQy9dUOwhYCloPqQuN1RXlVEndD7djvySOj0RTGElfBk8JiKaym3CATFsy6fxP91a8udW
c8cZXSZ/fboVj33Lidaxtnz7jlwRJOjun/hJrEE4FomNVa3Dj7XPWH3OeWzQghH7L64OPcAVfBJl
GwoVKVJmQtaPhsWeHBUqlEbT243idn18r7oHZEsYGs9yamnzSR3g3JCd243Wfz5fNv5eVt9J9XCZ
1xoCCczkSSHcnSHWRQH5V1RpxHJVD0irJRUfscURn0UUrTuz4HSvVwP5EnJz1CSCb+Kpn4y6jyaz
TIdMaFeuB+siXyP4pTAqeMgfY3zHcvDJ/lAMkbZ6TY2Et0P/sg/cAMrccyBvuPJ36FeAYtlh+mp5
7kZnLR/4HxjXNAG6MUEwklCMUpLGa/eVqSzRm/26AS3nwpoAwQoyXfq5MlHma+/4/0FYnI4om4Wg
6ML8F3ArKP6IUHkf7fNMFnWBUu0RL5LNtWKfLcBjQkioPaulKfoFkFqG9vu9QgHen0mEf4YbGQQx
S+D4xTBfJ8UuksqPuxAHbUsBFnJKg6Oea4gmvwSMWoOFQDytyGVeoORJOsO9fkuW9iWjMF9d75Xg
OlTbZkbMgqq//C1Wky4KztMOT2ifsW651I1OhUCMskFfaY+jyn1gJ9yMPXG/zSYTgNz8FaawjZPY
kcKhXxgCjFVX1QVAJcBsF4rW9xcNLnOHpxT1/2jz0X6lHOS9MpkMkx9UunuDXDfINEjL7/4wRItY
tORm2h0zSwCM7SfNK9cqq0M97vNvBzgFU3inYcesegPp948htvr+2ib4d8H0tvz5pwagXLYbRfzY
V3VlO9YlmLlZVTNm03mcVqorcUHZLpz1GtpRsNrqg0bNn3pjFyXis41/pgzFG3rQ5Ew18bma/ewo
OsmQH7xeucEPylDr3uMecu/P7rgYu+9jijF+sd7cQ2eiopnXsnGk6Vj2aHB/hzQXHKz7GgRNF8an
BRhCvlxbhF2lkHDmTc3doy51yti+SyDXkKuXw97q132iCqIHdUKs2z+yfkzzT1HrIKUI0DY4AFWa
byDEu8UkyafIA4cuEBVl4qlSGmB/u9BfXmFaYFl2modnn8TZRj5NkgTDNUrV7iXbT3b3DCVyZ9I/
xheDG/yqC6mXFN5Y7/086tlp1cK4byaP6eTt/FwAqwhTicpUaBUUdc5We8Mks5y4bilcXastXcjV
D3Ibx11hOciWYKPHXIAyAdSk464FxKCW7gOXvb2LnMf8BDb7Zb5obcBSbfhphgFMDkXD1LgelkU0
GDiss+D27k24dCUl8yzWpnC9CbK+O1olBUBXK4D+FDxR5eopkd9Ko8t15r7OSCBRFqmEXhAxkj8z
sf/5Wi2dge7P+Nvf6kGrvRF+J8WpcFU7yFMSzHDjwHG8xt2cHwZnpgwuHg2Vjr3Y3QTKb0RlRMMj
Egoniwxgf5weHkM5nwlqc11RAJdduoupjO8rYYjMRd4l1nrvadu//R/JFUxu/+cnOdnroIE4ZeOy
TNPqneVi7WTFPAh+Xns+6AmMUWr15h2FDm8CAsq2dRS6QykBtGrk3tVhsx+K6/OP8Q2wgyNyszH3
9oPoUb4RXK5tcTEefDsHEze/U0O1I/otAZ+f3bw1vbuYOpG5KcluO4dPJO4r7Nk5Jj2RVh3nDuxM
g6NvzkDfllKobVEabQtvfDwUnwBwUoveTdmn4od/UDy5FbXP6uOx3g1KzV3D+rWQlGgw6znq6luw
WO2OuclAUR/zKJXwEfs7qsOSTrbkx9l5o/8IZxtVh7jW4OyWX3yYl0H3xSFS6k67cx5iK4O3gFbI
Cg0Kd5FCjEO9Ty5IUECHhb0Jyq+ZU7BaghwJn8MO5jjkFhir3wrr3yNle/4gHUjl6EplTsy9FnI2
LEmRsEiSL002F/rzWJ2GretJqirKu4/epf55qm6QexhnqmAd2PJduGaUfl+KRPN09jPS1I6fya2x
otMANSePnROB/SIyJkm5q5GksiJQgffeQAxwdc+7s7L59qBj/YQIEKZCWrh4QsemwjbDV9ffL+JA
AO8ACTMVwPBxikQTJonMlF37Nt7Js6tYdPgTapDwxeR7upJ8Ir2392DF0q5NhJAWcQi9pX1cRBz+
Yi3c/SHWg4XK3GOp+ywuIGxvgCV5+FX1c+yLVrgRkJR9bNF6zXwibYDuoxVdR4IMYdzvX1yEidic
3JpFLnJhL9sa0+kssGoKei3XjJRTku1mfgPJa34UDXfQ6q7jJ6rYnqMGLFPMzGuzFu9CEPZXm8PZ
jni2oqYw/bf7n+4+yuh5NBNOH6HuMTw9QBX6GrPv01oe+tAzDYlarmGP9Nv1s+KCIrE/2lLlCUZg
BUPeAhoRrwJPeKCSpZHCKTr4T0+efqtzI9K6fjrZFIl/LpHB9KxQzuhNxLZA66hLl76nkNiITzsK
B7D/0TGsJhCF1dQS5Cc/HAfkBwVMKkoX+iPmyXKVaveiKK0YU8yL0KrX8x8ebHgV4TCkoyV0+l9d
B5x5zDj0UgkUYmF9whUTZLUYPtGXmEUqov/Du0i0ZvF1nn5gNcS2hWFbxEJWN80/xoEZBsd79B+Y
muG2Ss23iGPXieoAa3iYOtGKYDWJfT/TrMWTVIrJ1uv/8Q+LiU9ZJwrTuGTxmn6Oe9FTwEBdraYr
u8nxTcDJ3F5peedGgHk67JCEwP9P3Ut2znksYx9jScmNA9uFUsOHgQTnsfTQSkvQC+81+MdIYA9a
DKiNoU5mYNxD3bF9+OfI4AxE8xfLCHxgToeD6snfYmlleA77cO0MLGc53+6ZjvNECZ4sqkoN6JC9
j2n1T+z3kM4QEpYlR4RQbm2AALc2pwEcSEfvr6QouXUNF8EEiOQtPyzrk/Yk/+FQrli6+82prLMi
BWg4zn+Ev7MX6fnbkxmMgUlDE5y9mXoT9qTtrksafW78MC5tcWj3D7U0xUpWqcEYTJZfX2X5Nll5
NkRDeft9RkUmVzK0Ggso2BWiw6pLPVB2J5xD1GqvlJzkXic0flhUJ7kcjM+GtL9rLhkZtAvFZjLf
jvHCp5sE/+eXx+WrgrwX63A4T+URtJPaPnufRrYsTYAiweGaYxlQS50vASPoPoZ37J8GynivS3oO
Hwj26WefmTZUl5YnXX0xppEKLiJ0H431f2IVTseLdgUbnNOyTVnz/7aNcDMAUoUfFijh+Ov6NfD+
2mNbUvOYosoG7KJ9fpZfhcnlaC3d8zGlyodrOqfekYReJ5oA0tUNKfz9TcdeTh4zTMmSf4LHxcjS
Gvq0tq4jjvF9hdHXcpKTNJ3qcRsxL8vTIE2v+vwIFRAnuyMI9LqIj6XniQLc4SHZ18NiR0WItu3T
Erg8k9Pix6OCL6hUFSV5TfAA/gQFnzAONI5vxDg3cG7veOKQ3HNxHyxgbHJsRQ5CNGZsnKDjTpPP
Gf7mNloxL8lBua3cIoCIDRpy3eYFxGARkWEx3F1r4C9LIoVB+zk/hwqjYFsTgjYXwcOnVeeOrcoe
ARVV2AMhqn5R2Qlzq2KAC4Q4C4dqU7pKwr0De0tkeNNetQOWyYfbnvvafxWiucN006wOq1xUzf8O
7vS5+Ky/c0TxVqzyCbdBTaT6CTjCdzjOKAjB82f+JfVB9Z0kTWcsFAP2VOCmUWZlt4+raSg9Z0R2
CpKDkCu3uTNWWecnzH2LhKC+2tmEfaQLCctH/ad34dBWjbqDMbSAUWfCgTCgtBInmYCRrVo1UYpH
qWPMZgVjImcQI11RudgxeakJy3lH4aqKKj2NSmsFtrhQAp6krJuS8Q1QBgDb1UxFvlkRmchnHul+
jji7krN7nw4epU+y0ZQSpBxWWVX9soWSwujqUkfatIvY1RU919D6XbXL9gnbzu9QCXl8hRgO+Iyb
QfehsVm0TgODggAsQsVZ61he8ZdTVMhmFtfnrQdxpGju5f1KwPx4PDS7BS4j2KAd0z7wwXb2DhDb
4mZVeRJfVmTlWj7nZ05lp6Lb8PfuyK+ZnE6wlP+uogLDSrQ4FmTuZwTXXcXqU5J4JmASuKJzyJ27
ueURKSKvviHxnYOtgbzgSLv3fXrGRMkcGbzaNDo45TasmJtElS6nHBMVxSQjF8MW9HgGcXNNzREe
QbpAogv4hVj/WO93QyJ8PXfDIEV2OwqB0ZYo+McmbunTICotWtKzf5vkehVNJmlmhLN2Jh6wIorn
DVGa3VcLsP5aIhVDml/ZetxXCRU9NUxIU1sxjLbdaIr6cF7FQnAKams71QyfHAD34S8MaCfDsoYv
/WJBI3HXrWPzeFe0/krQLSGHpdwKSaabgBH69/63reiwZ3f3nRGg4LjyxbzEIjGHxwqlM2iz4k+s
ThzyHg+4NN4EuYNCm5+97CvG6hP2CBkAsJS7AmT/uXT2HN88uWPTcv+6/Q0wPO0yzjLo9TTYIj1b
N4mSC0K4LRYDldDaF6jG1p1HSjlsOLK/UqyhlcACIZHsOkT5b6QV4YLuN3VqAYGKAUcg/OeP9RRf
g86zwz+FgkO3MYky4mMXIkf5cWie19th3JrrHgt+ebSrzBS4szHVmP22ImJW/AVGRhPi0t3y9eCK
1zrJTO9zWGw9yTyjzODsqer8mgCi8hM6TNsd8IABMwzbARBsLRdwq/s+1IQ9qF27gy3z0+UUq3nQ
m5okLMpmXN1bXQiSBC9Bd2v0C8XOJxvK5sX7DLcWE6d4PwWcVwQ2LBBwWuw9zNUS0fRYTZeRz0dh
MYAV9hHLtjZbUzy907OWox4T0uSN9Vea680xG5B8mP+cAMVkZkb2wgjJzyNZ0wW3WjZrMZOMbQpY
sCQKWRhbGl+HIagyc9GTpGI7TGbFBLadeXNqReKNQ+ZDL+icIwQwjSAWnhwiCLQjBDqYcjDFkbbb
8KA39pMFk+o2cPe5aY2saZOI4PgSdHlY6/Xce1W58E2+Q5Ps7D0GCyqxWicsiEXVRksoQjD7qOY8
4BG5Ca9s6FpQqKJIA6dK1xLp3SGCwwqfx+TXCTwxK/zAC8Ce2i5R0ljf6KhZuPckFEBm8fuUkPJG
gDqNZshRYELr3xAavRfMiioCLfWRueq1IdFJd0A+O2eeELKWeMcb80F15n6iaDGFHCY1yXIS71ka
OuIWvchBppYSvJNZBOsDpeVem6I2qLoXyDTFWoSyYrQk4Mgn2VObAFys227pyEUHMOVCwGHTZKoF
nHBvF3x+L5oLBtTr1KSuIUEwVYucDTbVlYjaZHKbemXCfn6ZUYUzm/V1/elS7XbXSGLBvod+jmf1
RAGL3+KuEA4F26fhDNgmqwaePKX0UI1eNvyqhGBIZtykZb9dxgTKFqdg+LF7DnP7v9+yvBX/6j+H
DFFB3Zk6NpcRau1agkco4DUMh3nKk7TbImATgN+FdsOBqnG1Nw+DXxbAusvNH8A+oftM8xtibSwa
4BdePdrmy5yZD4PWsZuICx1M1r+hqT9MEScGtxj1XQ+DjZQBqxTY1JVpfiWufF9nUUh0AaNeDEtD
2FS2R0DVK1MqDbc0OlLnKDUdGtPlzzC8KYxa4uRv1b5uZBqzavFlwo/Dg8KQ9O+XCbJzwsT5HTE6
jSiWVEyNTIxr9K0+xazLqiKWQLvxcsM8yu0gkHDtPM84TQ41RlqI1LymQno8IhutrsiZFDO7ykIG
zZpxAoe4eiUiQrscHvZMF4Y778lwZwJTKkOXedh679IjT+2M70XcuMdzpvjN+0+JVcHE7Vq0Be+l
zMJDfZtJiDA05N/PotwEp1fOJ2p3MK3/n7pIe0loYQnXtiG9Uai5sl+OOD4tkcbIFoXxYBRz+dgJ
GLdS52/OCWOguUu8fJ8C09RL0f9pl4DxDTy3YXAmNaKNzWNgTB+B0jmb+F5q+VgC5gVwIk63dC4G
+EH9UsEfHGsaUXHfFRsrSP1vJhKwV9bZ6uUCpHdEGFF0GwWam1Mvkq3FwchQKPtM9WBDupQiNR1o
m7MAzZr08kZ+w661wZvaE5e8FFlcyePeXunZyAOt1niadPZPflhLzM6Y6vhXqQi3zK3Z8tHiy6dX
FzxMIVatat2Ws8BXP0TvRq4dyj7aUzC7H8pelRWcRFtFjfHSv006zeYqO7JBM9DlW654JSrLG7ha
WcLRcmC18+BmAobDbydYhKJtQbh6+++zx8KgZbkWXbaaukP5l1SkYj19F4nB4BK424wiunGD77+N
1MlO4B+S0GDwSlS9wQ/yzk04roNe8GEjKastwO8QE9Llr8wlZVfHksEB/CKQqa14MqLCWbkXvZVd
Uh9gsabC5x9GzIL+JZ48tdcRqEw8YGaXQ6AJH7Wyt6GzATj9X11gLwBOyhdj5Kd6uXB8eHxaIyfm
GaypsO1iZEjxTPMHxiI3n8AcyRIMB/ldZT1fwkx0xtFAvDC52drxKMJQ+bsWNb7vtblaNE1wZdwv
xW3Xrd2hpGgIOlfYNgUL9xbFcJwrllsOuA66anWZw1zc3cGhulITE5178QGQQFsGpJd86JSCfAam
/sVrccBG6UFzOWCjwwlTQHKNiwHDiLJTWJuaSPK6/wN+r5/cwV3iQaFcdNjwwAFci0L01fj08kJl
NX9QiG5SqsDuAEUneiCDgSXIWcRv/4I4rsgvVnJQ2o6fthja7akAStRWV6KAygpS/ITEpfwdzOWf
G73OXaOhRc8xQwEdZ+E1A2sz0zhlrs34QD4US+xUTZNJSM1ntv783TnlO3fyLeajaTF71s7enynh
le5NHISAwm6yyZuaq8jjYvCUNZHSzLbk0HFUyfiVvpBa+LhXsxeo+X4xjzqFowYJQaUqMMex1Uwd
E60uKEpfkpV8UVolXAKKd/pTgdTULU6LfPrEAe45bxZYttrXbOHrVGZP1mKmIHIuoCErvX+tpm3/
pjUNjTQYc/nlDDlmGCuC1VRjny5BuhWuED7rX3uxQYcRcgm6Ml6xNVPV4cZx0wiO5FBxxhJdYmni
DITUj+L9fWo6/m/ZONmCfV/1gSdHI9E/8eSUi/YIY7zrazPJmhq+mPxPPRE9TG3383AeyMWiXmoF
Js9S0axF6tZ2bejAHWwfEfdOKFFZjdIdzVN0pO+bs3dLiltE4N1oEBLJtvOjBfGKNBySCg2CXROg
93yBLPP7lcsTFTmqRJ7lfOSQGREBYnWj5hC2dX2jp+jTJ9auCQru9EUWKp1FjcyOhxELRW5Kakcj
eEsHT/ZkXORvA1MftJCWz+8lIWnE9NXAHgcy1b7PHgTNV+cbiNfLZy1xbeKy4r7zQp2Jn5bQI3sc
HOZ55piLvmEBMJhlalUmCIjKvC0izJqKxxud3biFR/1EZUbjXdzQ0/fZ/hp8uIfMEJhACOSdv2+C
4ijOaNfZtSIbgoCPulYNUOeeVYTM8Ej1MT996vnUh4MKd9CJ3cfB/Aznnc5/1tCqBTlm/FPNn64f
uGuswnlMRc6wk1VI76E1tt7LsWV7cbZyRy0yi6TJnFItNhgrk6TGnr+w29QYMXe2ROZrWBD390eX
jn/tNC56CGd8wwbIYGfuSZEbb5NctiUYtNQMinIusS0yX/0AQv58tR5TVde5JRZKRVKE+pYoYLtP
psuHz0VLtny+rtO1h4/Ku/ecBaPIDrRcWInoLP/opS2brPAocmB5bUxvSR0LIVMiv7PSuwzjUL3E
8K2accKdqfXbOcipTzpSIFILVqGm/flmALQ0n0oLnBn2R4k7/l1r/1aXR5XqNs+9ZctbBG17MeBN
QtcNewntoWI/DfYh9QXBXSt0yBUasERx+uSKxbJTpd/lGidI3KSkBI3Zs5aC3e+rbbNx28ORpLe6
eHOlWMvnICJ1GQ48a6k6EeuoPp2Ip5sTkl4u8U8t8wvpTGmviz5pekt+Q0THgODSMdvCcwcEeQsg
0nvEHc6B9fMv7HBQj3vbaZSo80nOymo8EofSDrT3JBiTgdMiHba6mToS2t/9hO2fPuoe2fML2SY/
fqVBnWSclrLDrGTGpU3X8ONoUZS/h9WGxfHE5DeTAkwcvhSHidsC+ov0QA8SCFOYhLfX0flwt8QV
D2f7ow2K9aQUwkD+VchXMP4On6ny1bO95/kF7l6pC/xNX116oyDV+uPoSUGE5++gtPFhdmEm3Zov
12+0QiSPkVn1ssL53ddJ0dn47Dh2XhOMJKuXtKWbF7HIplE9AWw2+G0+73Uc/Mw1wTQKvfOnKjId
AlOa/JN+XWmtYM+KkL5zvynFDIO38jcTYwuYS/E7vQRrrDnJvW5qyrZ+q6s60TNJVDISYGhG+Y1H
5ut6U+UrMIJ/RYWpOOqwykdlyOwrkaQuPUZw8Jw+thVQLmxnz4yrOVwVqQo+Qsy1LIP8rLUVFZVe
IshQ4T451jxgDe1GJhVA4d0sW6Xhfh4hd+a/MUXN2NU50PYIFPj2BO+Zb8um+8nH6zAVloaZtMU0
6leKn4/hHeG/MeXuLsTfzBxQIWxNU4ZLkcZn65uhqrKZeyE1O7tF0nD6hQRbhu593r/Y6dUxpAi3
/XT8lzqJ/fah2mJxVs70L0/M8ROffuW0oaaxJujVAXo5I+e3Xqmm01i7i4yqicEhK4GcSW4G8Ljr
hldSE2XdReB1d/+qiXHn/j0/VLtAGyzidqPnLHLwAESuWom+9E9HcakmLTthUDmoQvz1F5mBK5jq
NqDp/3V/D88Dxi3wFvbffSoAC/oxdwIlyFbXp20oDn4jiVQhgMwmXqhNBvG+3VsJMGivhwiQCzAC
katX6lYOGgid0O59j5faF3SFLO1MZ8QbI/o/PZucqtvCg+/u0nzzovjfgSz6F8YeGAwjA9WfI+qm
H24Okt1Y7yeUKhdobJeUwgBmOFU+CrkjI4WThbpc+hZBhBNO9UKWq2L6jaNVnya64qhhyF4fzwLD
/SrGZUzQGIp7kfAemaeQ/lvoGGrzsUgsa9c5owHvfq8rws8VnzlwclbUO9lzAThW74WsCSCFeoyc
sLJ51uAPcM4yT623n4C5eEM9nqLi2qIpFnVKXiL1qcwyOV1erdicFAx4qvOqcQsb1CYjZi29mffC
y1i5vYJKm16FRH2KGLk6Oev1iE3iZ8SZNjf6v8uF6XeZSH3eOIXcReVlruA5BR2qysv2ePLybZP4
ZvEJ/S6wRWlDMTof0EWlV8HvLXRrYX+BahOR7KcyNOxeSRHxyZnqngJSffAMAnAileZRYdvrY8ZM
hEaahK4WJ3CtVvk3P2D9/c2WFHw85xA3mJ5ySYRv12y5FFWDamsIzpqkBSKCss9M8QnZ/YPTlQSE
+GHKAhgqUTrAlaYBNsH+YdXlL/1USv/jSSaxqDIjoPMr+j0ni3NEADIrAVcIiLbg+hK9WExPyPUH
fqPcEs+O9tf2np+y93E8t9IpHHqkbfVamGdMjFhwdIJ+s9FCMaXt7BkShGZNm7HjvXFD5dqyyjIw
FQMvP9u3IDY9roI21dK+B3i0JdCMjX468jljLP9VFJ42in0FM6a+OSfZjiACx4IfrYAiMZF5sLCq
MJj48b85Z7SSC5GKfE6qCdqHQYUj/qt8Jy37cJxJWspXAe/DBH5fnrsWWsuprkZfcfJsb+tvQwbQ
9j2dixwT2VIwqVh9wiDAQTn2J3Kf+UCSlvvy+bBe2+ht1zPbWmorffYYgEb/dLI6W//qSg9aAbxT
rFjzmU4agTk0UMbSOn0eMPAWibJOq9i8oM/oySPdlToMnSjEIgdKkEpm9fc+I2MsF9cZUjUIbvMd
pQgv4qsIEUivZNayixDaSao2n3dyeqEJfKnYvEtlC9eo5nyb+5lvgDIvDUxbV94Z4jtSIA+/LHO0
vjqv2h99UC8s+bhsEuji9BmHi4EgTqEdzVuiDem3HC2qcMorWAf7CLHr3Jrm7jiBHDKYHZoIr8aj
rDW3rTywpsFbpv9lilLIUlfRQGwu4H1XnavvsBy9X3NhtmO79wzeeVyCsF2+UyUlInvWK4YMvjy4
JGlhTruYsmT1kg6H/r9ug/GWDQrZBzb/rMcIXI7HvryFf4dkX2qSKPwyEWBs1H7y8BuJmV+iZ/3r
KYSx/edxJ65GDFmUgj1fPQw6PPnH1SudoPMz9MLdglfTggykuAgJiAOv/cnCMcUtVwNy/oLfYqUd
4vJw2uI6Zy62w0j5d4nQca+Gg5pLVqUs05aEuJd6JamRDR97txWTK7tiaSHXNa93Sdld/0uAOm9H
3QvkgV02jjA7F5mp+GpLuVb2exeWoKB/GyW5tGTSErSFbMxRDgZbgCj+Cps6+9DNmSEy/k4zsyJX
lwMOvJyKa8cbAcCY+USgIxYpHo0VUob2iAjDxa+Y6KTFPl2xbn3S0vf+2WAorncJBPJ0LguVSCXm
fkJCDjMcPUXt+CL+jiqSfcHjNEcSIkiBF8vAqsDYL+1jIz+2+jqW+1s3BvNRZgL0tejw/sIQILbO
pFm43Qvt2RgM9c+0EslZ/l2fGrzfEqVVJt6W2PA2BH/sJo4mooBydLIW/fndVC3AAynQdelvzW0Q
ug8ZnkaGsF/j+u0Ws6yT7t7S3qcfGyobHU8BFEHd+0AwHazQNi6sOAZYvqLp2mKSK/nTX3oiYZfF
X+RaiM4K9X4SS+MDK+bDwXnPItjapBXVZk3YNd9OSdHL08f2d8PjpSLQvdC9iJID1rEZi+cMVgYY
maerku0TEroQdEe4YqBRfPpHRJtdR/M8GbiW07e28KTTlyy+nDRRdzAhPgXaz7Ch0G1fejs7jyZk
JI+1UVGmqI4eR9JQ6YSfAKSVulfDbZCIanoCXxQjjnUmrcAI+5VncVZF+ockUszAKeI1fSmZq4qC
fyOwD+NSNQLqCa/4tzGC21OUrrlrndKjHoXgjBStZ3/Dg7/OUsg258lkQVZA5cLbgOLSG1LBV5RI
tnPK8cblKmDNcXpprXlwo7JfAd6Q9sMRFH+VVEqCEm44d25e92v/kZ08v0exf1qvxx2FhlclCrst
U3LTP5kyPOBPZMLjFpzttUHjRmow5S3pZNQh8xl/YZ2bgthMkcNfKsw4W8qEnozQStDqbN74Ariy
ZwMTColSIExetP83W3HFGgvYsuk2Ylfw+RZZSKO3RsmBBIR2HyIrlt3QyqCXv0WTmaEc0eKRyjdN
bJntsY+vT9RIBCMgAsEkt0mzQ3NG+5QHPMmQpLWskKg417nHrnN0z0QywQBJCmh9FLzfKFXNXlMd
frA0cdkGFHN7+7fQUbcJL7Id5zgk7Ww/MArkxIjbnddq5pH/uKr7R3GojPjaKyvFi5W0gVAsY418
39TqHydnBmoVfGyf8byjl+LA6b7D0OtGog0T7t9EmJFAPe48bQR2MBJ1/N/u8qKlFWITIQ/gqyMw
oz2dhe/5G2cw99LXNTynkfV0Ir/U3EC85SHEL5YifbBoMKvA7rbCiDKw5C2xEfeEM25H1sOUr85r
DdM91SwUNtnOXxLCjFbfdhZam9UsJdggioOzGl5U3RsUQkwchibaKUNxFsflGBdYDeICry+0G9/J
xSI+dGPjvzp8CIxSao9w9H9rSaC0gzVTt4GzHIMpu4fRR9yInLOx551Ulpklem3fNVmtuMn8mApj
q4XwR1zBUjzhpqQaVWMvXsWwSZWdeTeoQMSWCzhDx3b1ee6UFxdWGXl6yWRczpuXelpXGQibSC6y
Zd50SzuI458h4Jd/VZayPYC1pCh2f4HTLub98q0+D7Hl13+BwUdd9ACQc/fQaU7dmMeeQonrkUwV
5X9E5gVsbVdMyTeGDz+YnfoiyqdQW1evpU+Twx6ZzlQuVzIAqizXPIptJywbB0Zmle03NirskGzd
Nl82/sCruK9roPg5E2rs/1/YTFrNrwhZqNiS8xJcZ9mHyKsI2uIoKOzrUiM46UGLwbJg6wzETBYW
CkMlGRxCqwx3pFOY5fO5hkOdyS3f1sm43DumaQixpm6nHXNE5amW1WN5B6j4hKa2ct4alRwrrYbU
fTg+oJ8AFKktObraBlhBl124VAAWWmXgE0juDYjRc6rq7IvR/DhUdv8JBajOsFIduRYIwhYQk8kF
CFevYg8qZIsjFGpzYYhd7ResYHW/NdKIbwMes3JyPR1b5T+YtKYQLngtZ6+bvwUkCSvFBMD1YIMx
23+FIZkXGI/v4Am7Rr0HKmxpQ3lKM856rVGq85iAAzgl4kWM+Nx0YXW6KhdRE6fmd7JQtn/2lopF
bo48hcdJjWL3rtTa/kUoTckz8KdSP8RlexVwuDdXS3ZveXf8sVM5hW/lKo08hmtGlXQJVHJG6QiL
ZXzwBArvwKEQIbMcZgRa1v6PfeI6clR8B5IsyO0w1Wb3Y9c4J+C4Rq/UKIJSWjh4K/iJPdizD/tL
uXZnNalZAj8iRpDGzve7zcXaCAR8Aizg+7T5KANrb5kz1vGU3EN5dFo1T5izjEt3EXTe65Z5k/Nr
bjPhfvHYdzm9LJj5mGiWPzcTZaLT2qFfqNA1/zY64aMdisA9D1fDAsFMmNNKzRo6IeCdweS9NaC4
FNJXHnYrCIqtTx829F05+PynRSpHJCm5X+a5HYfa5G+vwmV+2ToPFuZZ8HCQuSfjA1snafIGChbZ
wmPCxyvUlqxfcLTfZ0vVyHFD1ZkU2FQKlyNW6IjCQR4TuOC0UAzOzfv1gsGJeIc3FXlWUDJN45/j
6JUb1sUqySIyLfMcKbGxP+8FUWs832E2NVA3GC/ULhE8hHzp+1Z3DYHqPCYXfoMK8tBqEqDThU8q
Tox90S1gBNCDbD5276Or2Ov8/xxdOfWM+LcxiaXT0zi/RXB7PID2rFMi0KKt0oGZ+/R57TFTAqge
FZ2UAspDRYevn+AENx0UGO+aMPkigYStaLaXnYpe9qmIn66MSELf0NJSQzK2gi/dV9L8aBVHMqAT
IRpQTpBc54ZnkbjE0vPqEcCTSovGlqDEcnIqD16xcyCl9jwMsk5zvIJ+d2tJdgJEy/3FedvHvjbR
wsDLpnwsj30GgkIdZHrW60W3OERIHUsGrlFriSVyK93RM0t6285HMr6nYMVZtZdNx3P9sZNsN9i7
pKjQJWvmCXlLVvVwQTkwScllWYoqVmd1srRDEIgFAO9kR0SDSEiHW9cO8a9y3CU4Tv2HkRPlL5o1
lU/1usdz4LyWdjNy6lK1s9jtMpFQ1HKuLoDMva/oQUAqEjYda6pnteAhmejj0lUg5wGaKGwtzJiw
B0zbhU00/jWl+VXVdoRuCdi9E9x26RPCiPPmmDWnWUTH2lZKtscB0ho/7pvpvz8tY/ty/3b0c7lz
DPsUVeMugvAlY8PICoJ86lI8ECUs1Xvjccn83qGgdMo/I72raqCoUmN+RAstTpoZjjXK4R+OCGlr
/wGlNn5Ndi3iaUM/0IxLDMNJC8XKhnfZxsbxaKIc8HN4OpUwKSwOOWa6ZIiGXmEP4Xjdz/i0LtQl
ddB4lTgSTJQmuFNKkanI7myONw1xoh1S8U1vsm0yRdOOj4OpbIFPpZX42h4cjF98joIAxEpWDuCY
8YaGxKUnN2nsFJCK3ZmWT1pYmeIKiRX9cx0NMuQEqvnLLSwN878cVeGedFZoknAgnKjIkBARozzx
ar9EIwHhlft3GEp34Gr8V++Oa9+B0UpYEve4nxqFbVEmIOHeOX04pSpeoMJmR3hbKkTD6VDmU0Rr
KRDH8SgJXLWQr07qdat1XZiouL+tWnM7GGEWZeBZeYdSibI9LEBbLRLFfxZeuMm8bSFj6b+V4B3t
pDDqgU5UEbmod+Irp6046JB0BD7LnWKgXpRZwkD+91wpQexJDVOx7o+gRPsFmIJsaT1Ig0wb1SM4
n9Y+9OOHbqqpMgHydIck3uPgEe2FUKHwpD5T2WRb/KeIpHZEbxJYa/htqZV8SyXRZivkRpPHV9pg
s97qgJPrLG61LEMsKLKCopE0X+0wgXObGo2ej+a1gJmqj3bQhcLTKVG4a4eCVKtlYzD4JYelIhN1
294uVrUK9Adxz1+oV1hKv66AXhmJzM/plaL0LFkxWIhCChufD9jxKF6V61LrfgQNeAWXoa6udIFk
bPs7lFojX/znFYiDNdntJm6h2QUNehYkCYJGvUFDZatyDPAIErT9VW8DWeZpdiL7N7kl3A1WYYMw
LSG4O/J+j+RJsCZb5GkGsiIfHIOoZRAevWAjsV7kRvfZ/IHaNRFFBEXcqt4f7k38LIqfOD2beerI
OSE+FGBxrX1oouMNwItOrbUM8PD/hYN0lVO9zrv4IdqLlt/MPTIS335xUjJ3KmHzu4kaJb2cnhTR
zPLDI7NwK34ZVjtVJn7I+jR4/ZDpnJk0ss+MSZeRccIkj70cOnNcJ46D2FGpNQxnRuB2ycTVDfm1
ekUPOH6+Gve3pEOWAmXhQpreWQ7j+SAimMX/xNCeUT4N7z1Whw89MkT38cBs3wVzAf7Ll/nzC6ih
KWwWctRq/J/IOAnH/ra1PS/EET13NLBv5LtjW7/VppIQObRjBDBRsBZiui/ckYmsU7PL/e/RMODv
JCjpsYjM3KYX1kNnH5WfeIgcylEaviJGTI5VxVOgx7IJv2eZ1Au4iu82zFcrM/9HHBqRFfMshZ3o
SDi/kxvlNVzdIBnmE6LUOjWNCXyhH9/AAUXupfuPPKx7os/AQTE30RsXo57HtGa9GOBdoYH6Ik99
JzyASdOrSqghJWkS9DOTNTPxbJpTpaKrxnT9zV/M7f9hiljPdZPf+udydRmUEukhK1Kb5Bh0yQrW
BuHrW8eF1Jl6vl54vu5Jawj1qp3U287jdIj41mjamFGlbopfcT6yDBw9ig2mm52I/mwue3hpPYvF
4kGkcquE/X8Ho1Jdl8tMrotSSGHu7/ZykLkpEDo61KFMIaoLx7zb6cCENeWooS1EYrBh/vwmxVE7
CiygFKZqP+tHw00h8XVcitKplHhsNoHsc5zqWKaBtr8NPAa7Zbw3ddYllPeeVswUou5mlP8wTl85
btcJNuqZ5FAA+Zo7KK7y6vy0JaQTij66q1YnFslgjdxpyQljviPQZp/y7uMriuKOwKbakFyoVL/Z
vHZM3D8JstjBqKUudPXA3fARCINT04UlzYk0DtWyJWEgIH/K43seeIW4VSi05BtGmY0d6+/knldI
JgbyBAmOFm1NOr3NMM6h3K6/qfFS4KMWlSQ1nnYGytsdxkC0lVB2VGDy6vYLFQrsiks+/Mb1wQ5+
Plpsk8XsT5pQywAFdj9x+b+GoXfxJdx7aSBtw3jJwPCobR4vl79nrgDh01xOdy6zvPuNJw6HTXhK
k0gq9Ij1ZqXeB4JoCoxrgRCD3C2QiRGBVdtzaAX94WiX2uSb0D8e8U1ZvU92XT1WXBEH2bfCp4Y+
PQWmGauPT21i/TlSu4oQ2DcJPl7Rxn+6694n42FekT3mIBCH3gtDmu6y0Y0QLJZIanxJI1yMCa49
zP/Mx6Rqy39EPJ2HTAuMxS7HKFsucYzYuxfaWxYdktwP44RIyRto4L5Dpk86IO0xJVKDASmAvzHf
xnuEfKRNmvgFDzyXRBuDaoeKkN2jZA7a3qHlcQ95zQXYO1JdrrHb2KzNkpQ68M5Uv0h/vk3xG54g
NThaPX5Ult2cLRKh/49ZQ7c97eozhOe86QxwcQLsZscBKyHyo0Fqn4Mk5vDXoydOTSD0n+6IAAZ9
QBU4RwQ+7cCRYKhGNUo+JHtSLjEgFndAB4LKF9uavgSJNpdwffQoi+HZion9D7TD3HonD9OzZU5T
Lc6rh85ih1BI01Pep852QM/MsaoMvkMS8gFsJDgYob4+jk9zSiHsx2/WeipDOe9kX1RyiCqe7YHu
4RqH52AedhwGyNWx5UKNY4RJ4ega1pLegl14crLvuOQJliPJZSt0pR2qWh1ME3c5EuJbGwEfNOrn
xOHc3fUWl5cf4anEmJpDZ/cw3kCHrofqtkbmaVzizvipa2L59qNIvBdZv4LwVWr+5eZvP2QHH5ak
ryX+e59pQI25Ku1R9lZ65orChBS/C16nE9y5vOkZ6wGzCeT8cU6Cgt0rR9mCuCibblJEJbKKSxWQ
uiTXpKzJchL3GLdn7/fBC1GFdR/Te5IDkpDNQO9UB6cN6S8ufOVKTgbsCgnPMJCGKvENbde0ssjx
Ov2v60QQO0bm/QNzxHb+Hwu/xQbXXS04ebFB54tpVKmFsymLuGGnbm+W2LS31pxdEIpovzbpeSjs
cUM8uQWLGLwqATNF8u2DknBrSRtIHw90YSK0losVJudT2Wmi03qoI8rPxfAFolzTirmeJRCYnLp4
NzaUlhXyVHrIxlexLeKyBtlWxiwY0wsObTXYXHoAYQ82cFLZ8UNi0oe+gxYWElYLbFqEzqY+iRBo
yYlRCPbH5XNObC7ujCbPfM5ImzjeI1XdWJiDv7vJEo+4G9IOCbdhblvxckiYW3+k00YSV6z7lZc+
ogXYkjuV+CfRpKezK4vuuoLexRHMV/FfgSyj/17KWcZDIwHM/nEix7UUKD4i3tBbFSlqWiqtFTLP
GhhZ+s3V5/joYM4ni5eGdY/cb4M4emQnyPVwf3GHSZ568IhvK29nuoLscSlo2kd3Wuvdb+RNZ+se
KOW8mPKER1z3h39m09Pg/DVuJm41xKnYj0Vr6Hwsxy1UGl3J6UOmXHFwl9JLYOYoChihcQT+AiE2
iakrYPEAlfuPtCuCyUvPqlPOS8cOONJAMlg9xYi9GKapjLZV/uVwZWVu0y9IiXK/Fb0TzvGEEWuc
K3riGsClOjgLu65fWi9YAqUXoPf1OAogz0Ni8MDPPqQzVe7rRQxtAw4XV8KUTTWInO8uFlfRGEsY
v1kWxVfi1pn1x5xcCBCJaaFmE9xmjVl85Kg5DJWe0VmJcxhJ5nr+OyjBg0IvDBaGGWB+62FnWEnW
+uVOIp7wcC9JTv8MpH6TAAvCuSgn3floo1EruwNl/ZNtTRzh/Rgvg/S8slUbi2vg56AuEux9UuT2
uSYS6niCNBnqNruE118CH5i6Nz7Yf5ZMDr8hzYoGV1sxtoWnF1/6EsLoCikeQGNd5NFZZJBIMCcZ
uhq41pQ1KpdT6cutglw0igBkJzQGXx0+lK+QYUckMXq5R02WJfPVNBXrWQGwwtJmh/8jscFnewW9
Yp9VOwyd9gkkymtcJAksAw05/0qYFlgKyKRpMiupNSMhZ3uAG68uQjsHL396eJATc+qdr+N76926
9UFIEVgTRSEKyyYZ8pGXEi4Fgli5MaXJkgxhpPECtkxH2QmZQDHmRilTrHWvtM29297RLWp7qrKr
WhOQWtDK47Vg9EjleCQfGwIKnJFpUmUZandA3LEauthcm/VMs9zJGX+aSYC/jMJK0CMkz5wBHk5a
xe9rTz/+S4mbOS0kyTnwSBFxcIjeFQPb5tduLGk0vkZ3jym1MTHJWNNGI4HUe1MiLN/fSPLajooo
NbltOYcuVwcHPpid9lr0sYofNZqa7crpwtUnBO3jsf/L8OR94LuyK4E2lE1/VXDtlzTW9iK0FVVZ
5m/YLfQWiuEmezKd13WuYMpoeFLXvj33olGqesMiUiyNhxI23t8XeTHj0khDSTGSP/Me0ObfC6RI
tyDVBdori7e5UTGnEU9ObuOfqK4nisHadgaKCUfAygb46XxAlEeghb4UH1ux8Np4IC5scyhS3t1u
AZJ1eEEawT3gRTO0f0PEC7MPpq3tC7k7nVsd/0OoZEfQz6GXClQlGlSGkEF3TxSAms0sokmy4xjX
BX7bdTNyMVD/ewLhrMazmEPO3Y2h3ZirqUsZrLVSr/dH0z+SJI8uB44s5AfjuV22bYY3dXKel/kr
MjqfaerKhcqnEZmJFhzpld2lwx4ka5xw21aqgItBJOl3pc891AM1LuMpmlpg3NDGaQJLl6hoS4H7
LWNcWAqVmCs9ohAcyFXqHxdnCPqPtM8vwREtrxj3CVQIC1u90kcD2yCrtzY2Ks1YL0IXRtfQjrWT
4Pep3Uq9ZYB80IMkeQAhSSFXjUxIRiu72934FGXnGsy5+JL5+TS4nJCOn1kqlhPUa5abZLHOc1Dd
olkuyLgwubRHTPqDmhOKDFPRIG6x6yhM3SWhoHVOs1xhgzITO2w9Qj8d5eybLr7URd3NRjT0tiLb
yV9PXtExHAlMVtS4kUyTOZHN07qCouXR4NBPKhgdxQFCbwY3Isf9FQXPX24pP3ZokrIqmPQeJ7ME
/uEL3AWXEuq/dBmP89/oR1IxP9T4F0kchFJ+Ocq8uK1McKPjMmVq19HxTn4F7Q75gZ4XwLAcX6qF
ojrPr5hCh4SYDpj53dOvgHXyHMWoQYcKTjzV426e+LCb7DF62GSXX2BFCjauJ+kDd1Sd/dRdOGvI
ur29pQvkvQtxC+TyGY1P6IBU984ieIiVKu/oFs4sGGk821+TW0CxoT1+cXRruzyI8pJhkmkQ+ARP
CAV5FuhiiON9IaYP88lAvUEHoMih9UJ+lwePSZGNSGs4lS5c+lx5fH6B2jijgTAUHy1NbztSH+o1
2kUEW9KVf3lYCYdJyDQZUa5gG/A8CoS3nHfj07IbNxRRIeD2XsJZv8nyYgKIePIDqBvavxYGcaoQ
ZzNwxDMB8FkHKtPbnE3tDKVHnXKOCBquX3sDasFd47KDVvrybn5iCIFlhtyHdR1xjwN6VN/HYisb
PblJAZ7lAv6kzhlGMHfoSWwxhdhUOuQLWr5dF7rpda2ZYH10S8W4OonS8lN3ZSt96FWvY9FknUdy
qJXcrxbxkQr+IB02WNCVVe+ZyGP3A4PXI1h7TbqVhrVV93fv8RlrokXupfSkbBsXIw6MnhEcBdfb
xTsvb1KgAy8iE31+vVrq5w/rsZwhK/0+EvysjBUakMra7CrkiHFz/Axj2oB8EnmUj5WXWT6Yjx0Q
OXqINT/6efdAIg2V+LFBzBqthPuPlvwP9Hl4ikP4uBAITG4WNAp5qiARU7wvCjyoJLUuFNn1LQix
Ga7vNIN4Cefq8FoQwz1aizeuWVG0OgPHoDUNctF3pU2gT0/aABiRIE2i1teqqywQt3gEDlMr7kwe
o1zC1w3dXk7QAy0ZKyYdh0SUf7x6iC+/fJbBW13ytxo1+zmCF05Q32+gLsihr3++XqZGbij23+9E
KVqvE7ePkFbSzQF9rHuRdm6aLXCtRNE7o5m6xCXRfGCZQW0uePzQazGJhPgiWNzMmMzK3b3HKrA5
ktCH8ifhWg9m2R9jIsA8ENFjIVyrB6C/3F7vZ3UQJK1wTDIC+uo+84B1jbhxdtraOOLCG4d2NOaz
W138Y06TTRq3/9VnUtJ1ogfm7qBzetzFrjYf7g1rDDXOALnjQDtNUvr48vZUl8AV8DUiqHAoEdmO
SXkMUVwu4VDc+m1u6zrPsA9WeD6A7umz5jIc/AF/8Hjk3xIftRJ5BWzCaPRYs4CLhaR2SYAy1G0z
P4rM1hdXYVmWbyCSQtNJ+FzqvITAx9EXf0oejfCSvqQilAdQAMc98NGGTIjWvFWOkRHuplv0FwT4
Sima0LN2IlBV2SJLSSJ4LEpf+VqHbDaDVck/BWvYCBOH27+WCryj+QxRpooyzHO+K2cFBYmxPW42
rGmEUoyeJ3RAtjJPvqDOw9iwp1Gax4uip3vN/bLr1EpHSic00+tZSF/cN5SCkgV4hg9h+0gVxcgF
a7ACo3aHR+1p+mkiJQkaAx67DOJBUKFq5VV3akRCxZOApzbZbZhnkYKJKUOARPLo7XTB8KHf8/Kl
V3MSzTWJyiiia4urhbOeNRLtjFtkwl85BRDpEwnPIBkZQv1/AcS2MLdkxiFeY4hB/puuq1Zg86uJ
epBuh/F1iaXRcFP9fyKZKd7LWdx72FMX7EORqtVRLWEGeAlAIwyntTGCejQtpp2xADX6bcUh40tV
ftBv0tJhQCkwg2iJwEHffX5wVk5rZ3oxszcXtWTb+OivtFiR/usBatN620oUf2nGMWtucJB39S/F
k8FWMPfNGpggn1N5Mnic+MyIJsgtvZloaW8wk+c7q1en5Zoi4/CmabHZhtuNRCS8Yp5TKuxKblqs
FxNBy1yITuaD9ZnBhbkr08F/fsL01u1I8x/bMY8UAJ2FCgd3FytpYdAz5LqXSExJCefAN8tRlmfG
6YRB8VGv2XEJ/LIb+5+sV6A5MgnF5lXJIb+/JECg7FheL3iWIai/O/bPb2iU0WRM/5sjflEy+1WW
YMoNvlZbyoKG0PJMmoxCJEDc1MFl/SD9eY48NJ5uGYf1raRxz+nXFHNE5NxJA/Hh07y0Avg25Xcy
DdljN/hIi/V75X2UDBngpeG4GzcSonJKaRBVbd0vvOQfutJeh7vMMEuxYN2y/GFjp+ptoRu0eu0Y
P4IcAJg72bY1heGiE8daSyllUb597uU97OF+RLRzsATaUsR/uUwz+PMZsG95/lORid5uh0IVqrKq
QZcxw9TjLo2y3NkAPO4sPIfeho7hy9expJ9mAabEO38yuqX+c1KD7T4IPZla8aicNhfH7SBKbrms
uiBqO9CGHqF9rsELw/UBAVBH9kfCJFtMfs77RMrHZFxn+h1U837FafEln/GyczHk8foW51Ks70lM
ugbn4kDGn9Y43al4Np5ubOae3l4ApQof16jzS+ENdigW23QQ5tq/x3mNnBcmOo3rsEavdtX1K4Hl
1wWRxkWDLii8mA+Z+MBCTYkJ3pda1FAzvi9y0KAxs50YbKzqCq/XBeVEOLfFzWsHQ8BU9yorjY9w
td7cL7gl26McJDZEWS+SOQ7czEE9MtCr56J89CMOENEyMoWt9xFmVowCYygzSDZSOgCh3eRIJvcd
L4hqQvi7drkTWBX73fqkqqb66zSOywlNBwPyorUKCjA6GZhtys2oZfsrdLQ/NCyrkSgEet7L6a2M
WurfgUpNXk2awH9D4R/YRZNjxUnUvKcaNGEF+ciWyKJJ/EKXddJMF8gE4obZOtvcOCrlRju0dj7h
4pn1zCHqb5g9Nc1ICCV04Gl1du/O8p8bZHn1NE719U9j7UDxjUy4Q8llCHl0CnjnjbOVHGxUlCHj
LKqJsx4SRiwL/dcw5VkBdf1owZdLHjcinTmWuHlldRJ+WqBBlwYGNWKzPfc6Y45T6/lwpguVLnlw
nIbcDE6XMfrLYLOUrJmjQ6sSfmbnA6l2rY268gF9HrvofB4fIExRRsBYclOT2qtZo2mzQ+tanYoM
gE2Q556OhotHqnlh3GGSYKtjGG/x14n88B7Kwk4FA3a+mykNM/nEB5m8QbKAUm/04m7iqO5X3nBP
dHRDM7hrbWzlgn6NRuPRqxc7VZ0AL4UrUuv1zGlxMVJNoCKcT+1EWWdismcbkZTscFS7Rzijsf32
kZb1+OUciNard1+wSmczCP/0gqenZfa/TgwQdDIWuG8xepvz0yqOPvuIycaLqXYXy9pi3bzABgAb
e8JBNCNV4saSyRD9xLzGssc+1n16xqjLIqRsdAt5iPBjd2njcAS/TL2ZcQFzygVIpCzrMBElfpiC
dq1+3uho+uItKzXquOY8YFnp3UsGgsAreB1D1+BMv3T3t5gs1sVcVQvUqGMGqRYOhDoDwdrqWVWD
P0g/roVCpZ+5ALByFaACWrJO/XfbQXp7lHIugQXxaeDFfCe5WAwpE7oMj9tgxGk4aueZfAmaabQQ
XlmCB0P8OqSYdSN377+whIr627gAhfEpwsyq4mERO6rCUX8YEDcLHfHEfKddW94a8N+gYdR8Yl/X
FItwr/fgaC75Slf+N4CccZ3lP0tYaaTb6/Nz0//lPyIJCtALOgRIG57EkXMn3zTPcBIYEDpfL3ty
efIYi8Jp7Gs7x4dCB5ZML/kteojh/fBoYObDXc7KgNK4SWIv1eWA0NSwHVpPhag2GYkGEnCPvrpo
Fs5GxL1vnt2au1kPAfFUxmjRYvNQfXMK7b/6JZkQLj09fSrwy3bky/uU85baZuLFFl9jkfAAXetK
BH+m1dsRzO35Z7xjUkfvts4L1bY9iG7wiaJg4qCvf/20/gAoQYhDLFmp4POB39vb7C5CvLIXC9zs
4Bz56ujy9wq4rqXCz0F0TLJBVWDC1VY9pKPUhfACt8wQzgdpSIcs/Gwpjs79Bd5+cSPaGldXWzEa
P8GgLrMbPYT7KA76MOvjIVqEpt2TBy0bE+UWTxGl+023uA9Y0yg0dod+42z0pJynAXwwDM4O55av
PZoj12Gx4nOnsMwq87qvzkeU+OQWkUXI6khbM0TlXiwOF1PYC282XhfQE+gmLjUtLM7RVE5/o4hq
1HBrk/cidMZI6GiGyX6g4dNE3Te4D4E2RC2IBZow2Bf4njb5lgB6DqorWSufxLNohdI/MP5yXFyT
Y8+OJEBXQzLd/wCexvcPa5Np/iFQfF5GwxI4hfDu175PhdutaRhPxzjZavPUJww02jpotlytfymD
40gzvwnBso5+bBnrIoHA2DIA5z93xwYaaqUFCkYTYJcYu4KY/WlhiOaJNuEmVHsLOcsl2KLCHymJ
iON2dcpIUI08qIVRVeurrlpW4slWyJdTDffsU/op+LWutUGfescs68VAkrDu2KfI82ga1m/chTm+
nXkE+R5DhZCCkftgdBDstHXVZuP2Mlgybo+FKIkscFl4QQ6MoRqPEdlAlhMFM/NSrHQf7vwk90G0
LBdgjfrXN8q/9vbVYnsLQ9Mm5TfSQCbrheXnRGRg/XnCBupqlxXvp8pgp1z8p8PTpOkvyM5CQU94
Di49bNRcEf38n2Qrkd38C7QifWlunRUnZIJrmhE9TxObTCHcanRNgwBSoyjaJjejuT4hluL9BXUe
qSgqy+REyzZTe19N7zSBnp38PpXW//6Rz7ZL/+qMNCXd80GPnVyrwszd4cNSd+mKd6L2Nu5zVBcu
usynaUXPy7ibF5c/bwVdZQGbSWQ5GKvi4R41RO4AfvbRpHTptEYsTOTBUGo9lk32tC98NsmsF6pU
VV5iKtfmEKZMFuGBoZoHPyuTsOk9aoxvvzR7Ndt39BXjjcapwpK987VLpVKtuSe7P0wkVNSEGwVy
X60dZA89g2lmjH5LXyz8cgZNIyL9TUyQ9eO6xnilabXokJ1VOdw3KsarqsNdGl1Fsqv7qoOf5dTs
imj5vLYKPL+rtdjIFl7Fd9elDASc8UnOTcYvu/YJ5I/s4jTXcz6Qea/Q7Jhx+xUNLTQ1tLxpCD1+
t1muNj0acLiknbIN+iikahNCJhVm8N+VOPgWc+mmql+99eREVdL3siH3OluUZLJmX2DGNlrgBwvi
/cBe5Gv3hW3BlL4u386g8ib+WjbR9uQNhOiK7XIwryOUNBNMkKHRSugCn8FpVaTR1xUhmcpnLz2L
m7AwCAxrOt4w3OAeCJD8jU2uleUZ9KkIiLIqxoWtDk+Gko1HBT7+zTr1tfCcUt2saqeWrcr0Mmud
C878JW4Q2HojkG4fUcV6FlqJ781A7cl+EcREipmG6F2n3ylmHIF/+tAZNi4m6gUbuYmwaXPt1ic0
UDul3TdgnvjmU7+miACaKyd/tm7EdRPG2nQmDwtZvqUBTcf75+FjaSrXtPGh7A3+G3P3SU3djPbO
oWz3MmABRKNbyuB7tUoYQ5V4RIxXRdRfeOBGIKlUZM2ZNWC9MaP+RbZNb+KeCDZyttKZCBkPqAgw
1XaKpYxe7xY9TwDBqcy3oB90oEwHHElkZSejkhnrkjCSXu5SzSY4nSyh6dFhY95PzAaJKyFbsdOU
/zW5f+P+i7FrqEnHrkYUzJeWbssVksgW/3FRJ8zWhEM2CcqulcXPeq63/Qa2GStUiczhEHq/AsBV
fz3NVup+0Phkb9lwZHVy7t0VLERtBooNQOiEgDoUNdyXllU9d0O8VpFrJ+iCT9TgVZyeT1NJcvJv
2alQByo8W2CUgftoInHeEv/kGaIegdaPhz+JKj+uXXNmD4o4DXebmYqM9GbV+TV8oCzQG5U/xYbY
rTNcxHmd5hytrDlJ1QlyyY5X7BvSmXpyT9FDlbyTY6VfIn7JJ9QZn8IG875cgh8zgkEm2sLkZqg9
rh8y4PfOD/gdOl7IOgLeohCe1fJvIIqRXzyXYeg37r0I4Xuhn/4k+nxs/UEYlSJZtoHZ/DiJIZFE
LTBZInpLXg4FX0N0iW3Shx2OPyG7Zv7vqM6WA1T7vlCrYuAaNlLdY+BrSDa2F5JBSp6UITBiE6i/
4R36iQnfg40XeAwOWR0JJX9AEZzc4pexiWIrMGk2JHk1P5BJMFVQHmzTX0FflIGsAwRjvV7DU9bh
dlk3e44zNhePlaGXsFkt4viW5rWOzhPnaWvNyJKrQtMY2unrnS91tO+mPNCszZuD+x21xi/lHj76
aKtsIBxO5RP9WGMMwF7XZzLDRYXkKEJgCplMDO0xsD2LyQxBYfiGT7+IAMlHsDitgPM+mQK+qlly
surgS/GETrR5VmlN5EMwNoYQqa9daeGGmiE5TN3hlBdIghD6gCdxA98qVFrZf64wREqVTnlQweql
oBgirEpkp5nmhkUPGbh+RRu0nD1eJ0Kp2qE3cw+8caXojSrJ+lKvI55/VEl+zAD0p0wThzLSnfIt
ASMuJES8GJEmMKSFizGzT/EVu63nmYcLMEJw5jDK3+Eiku9wL7O6rirFk/pdvb9ei/6FhmI2h/qP
SMY0Xs8PM6fKAnzmmxw42SpwKpo8Hz7UumiFUlqrtWJyMiovn/qUGhrnwLi4//GiA8kGl/jXBIzx
GoE0pDBkWRvqFE2M5N2xgjQ2MvtVa0f+a2Jxf5IOoWsf5GnFIOvYd9O5gmzk56Z5q4xSedygN3dU
p1IHSet6ouE3FJCLAEvpIhbrlMM4HeHv0L3h/DjjChTmJDXyB1CA2SSVhEDRq9I5mAr7XJcer0z+
u+0AhjG6D3ALhyMjulU5oA0PUld0JvxUuPqv2ZCphaeT+Y9PhgDLKomMkl3RYzcvlEclEDONqbZC
jDffTgR4tVmYXnCaZiMHSVxYPX4KIca9fx1gHkuVm4WEf2wNAVlRfQrsHNo9bYCiKKRMSpT/E6XQ
telPw/DGtjZkW1BGOrbGAqpC3jN0YbOXHMjBLm8g84t1KyE3iqTjWYtP82dH3ZLQTU8H4UjeWGgm
gEWgJTdzMSjP5WmPEwPp1h/2lnpyDYHMrDcJ4XDa2ttxgsgNWOJ75AJPRigC7K6yFbGOYLTTook4
AG1KTCEkrsX1mP+uj0Q2Ei4Df3gH9AVupj6QzFVOKA+zjWvG+g9vVG73ZMqqLHuzC8IaG2mFkz0U
7/tIkX8/21lV1lljLCf3C5/bNZ2St+gsFjgepBWHx2Yf9KgxOoErDeoEvtz34QJ5ySUohmYVcBn3
VMWEUm0pZe4Fy2oBZzAndKZ+aydk7VpWzRZnET45t2WnOr0nLmt5jCQxY/Au0JqP/Ax3azZ0xRYV
vx8NxvXLsDfns5VP1NUxk30N/Emr0uyZKJxEOOr4BAucuc8euCfNVfK3KQnK7KC1ZK3lZzfO0WeI
oIrZW3zxaT9lM0fupAZe/RNYf/9LMP0xi+IYHkgSJBE7UEGEOwrMlYwaGPMnRk/i2cgHRb4PISQY
VdDepbh1Fzt7cG/awjf3dNgoJraae1BAXejSdIIkgDhcWWRmwBgpxaimxhTrSObDsm0B5e3HM7v6
vnGksNL7LElD3HJmdpRAFJ0fPNCMp75QqHKtbVhKHtxzq7usc4rGRlM7TOfAzc+R862rc/oTiK1v
f1x/jKOq3zOfWAkOkjHGg1Kj96sIfV/hwQPuHQV5SXKmS/+4Rb6Q+01jdJvZ3KJyxiQzPSbhlogw
ETEWtnQP2GcmypTzoXALwdugjOk9TmMqVpeT6I+aSTHBMoOa7JMswZi9ZWuVo9qVr14I8cLyV28f
URxa1G1sKocLbdyVbdRhvqLNzNHCVkK+UpJZBJIHkl8IPPQVYDVC6ti9GwinrkHdGHDSX26EqWBB
lXa5TmowwAxWIW61kLN/tFQZ+VNaFosCEIRpHpz4dU6tvxYcrCdKn1eA30LxG9OQ3Tk0HSBaHGY4
v6Gu1rjruZ7Vo7G1QzLlFwlAXjpKXp4Nimj6RWxKKgTEgOVId5FdEFLqarR0nNmkgiQBO0psFvOl
EILMKr8sMaptN8gFN+twi/QDBMoQyH9IL271y0X8sLg4hYQvVZUXyi0XNCjISwMIV6RDN/L5Tj8l
BpatT994BqW1gXrWmPwu9g6QR+thGP2jwJ20JrREQplz+xQFeRrrTorKiFQBMguTqu5cyMb3vDOQ
mvM4Stkx4DtgrUkPAtUnBk2AzQrGMMzUQ4RStsFKyQ0PNNXZ2tX3lyrV6D+wlu3sNLIPRuQmAtl4
kI6qAwvV6IlelcXbBAEA8MVEy6R5fW+C7426MNH68ropKBMGZI5pLGelxURf83IOdhLkgrRgah1T
e1n9xHO/hUdTMzMgWqP87tooIO0g36xP7bflu6g6QNI8bz7YA6qu3VrRr4LydC18hhJtXyTiWeNX
etHGqJQd6ksON8Fcjk+TuBdSSsQyB+q7joV1eDn6cnl5IIcedrI1TXkwKFcwn9ePqWJoIJXfF8Y/
w2Szs02Egv6wJwKAo29RyrgCQ3Vj1Qo2Vybq12a0DXmgsVE4re0gKNjfAr13JgxHtTXEFVOHkE9p
IDDkwvGGNL4ZFDtdELIJu/WehBWIGNkOEhnLAaG3muBJpeWBuMQMKIAjjqUl1tXaroCIENgrHzU/
JWqP57YyYmg9YSzosAKEfIGxpbC3EqM/3bLZRKkDVVZ1imY7neZjd207mNrzHIifjvBNyzk9mQRI
xkT28FERZX8Bc1KV0hKk8BB5vT04N97C9Wov2z+jkHZMiv8MyY44SOJvEb6e9vtlgQUTqf6Km594
COGc/qRPcaqBOrQOeVqidIcgCnMKlp9mznXYTyrpwqq27sHreUfdXL3LgC5h73bRc8GkgYGx8mTD
TB0xEiubOTk73RlTuN8WS+7OjWKGrjho9/85AzZh+7wOCMVhbpgc8XoCnwy2ikmPeoujczQm7VFx
CXBkrYcMRgF0alWu8kqWDjBNM+edd4xOBWM5PJsaBCqv3BCOxB+GRDbkFafd/Gl+fhXJncxC080c
m9XzVA192LHRVx1tsmOVREzXj85brtvfeg3hIK+fZrTiz6ueGAo6P+cjSPGF463Ik/zdJlFR4hnK
8JGtfRyrWPxLCYvQCi7aEOXMiBrsPXagllHa9Ke3S9o4Pi6QfKtA/paVaXtsnuNPb0Mcvuguo7f9
5oN6oVRans6V5eiGqA4iwPi5boQ53RhK9YWwyw0nQeSLewI/gcQvvn5xy99vCnJyQDdyL1XUrMoQ
jJ0gVvMMuo0nuNfiKVJoFPb6ic+UarwzeV/kTnVrrEJiKeHYkIJRlpxX6tsxcu01FZtawpTtkHnt
5Rvnh4/sTtLhXiGlZmsuREc0Y7Ujy/0N0kwM0xKMOXRoMsGNmhIEBUWtfGNvxXTYM7OjLmfs3HSD
GJV/FaeWYvflroBu6hb7snlSgPrjDNT9V81nmWe9idNy6wWpQHJSspn0XXAH51U2lQlRtlFqBf+s
dNSlzdbKGZ7xSbCanWJvcLPQoBxw7eBluXfqE9hQGPyImPhPyo/y9g1eghXx8NUwluBBk/WyIALE
lHBZj9XtR7+D74izVjtPqzV7gM1Gcm3SijCWUwpr1EHNFxaXTV5GnSgWiKJsLwouUPG5QNCWecQF
EzmE0GhTXailUqPBaXT63ln5BQfrGC16TGRN0cj7DnqUAvpdfUdWwfHcWjsvbqzg1mogjGFYiQhG
jBAgr3rnGsYcD71xHWqKcnkTUSWIRjFl9JmAqmwMDX7SPj9AB9r4T63zXe5NMTr9iDyxLS5KYbfq
xqWVcJ/u+5VkpvnZHpPgPm0Av5uSU111gzXB173rjU9dHcqg354YFOUYmG/z99OSdsoYqhG4oueT
AD3hRKuWIXl80Uih5AkS+dAXzPaSSHtfHQ+Ytecqeo5kL4mojVGGomZkG6HPfQIhI1aXs4smFQkH
XTh/LCXoWEFAR8zL1SZt6nw8jRqIQCjM5VKpVEiRb5wiCOjqh4xOzVYJ1um5VY8S8csASv6+eNSG
Q+yuGjMvYadZHs61emIZOsZngFIAZdNgbp+ezstN0h0Kx7Itx/VZcJqH20jXsLLyEgKXgeYM+wdj
HFm+I6cYN2mqb8X4bTPjQ9i457aePMq40Pxn8bJbe4bT5uIm/MnoGIgloKjTFh6ELSU2nJMLNgiv
KJqvr/0pda5GQ50UZrRlgU+XVtF9KorXEMDHz7JnJW3PFDAY9/219DyB9QyASrNV28Yq5cUSquFq
VMGe/x5SP3acsuF5eU/oELufbaeLbdBTVfxUpTdouZUX82Yty2LdX9IRPZXlwPvjtl/fUeAw6YJ3
NLq36dSBM/s7lZoSG7ifPIoJa7jpjiFteFe5FaEFkuUvX9IpRcMW7I0GWJ0t6Ikg9ceL++F3nkHp
auvQ31gLVMiH2qELehIHmReyVJb8qK9kbCqJySWTaKQ8vKfStJur7J/ngvMSt/OkM2tZHVZmYpA0
aZjI0ICPzDNhlp94/6xe5wzpypr50WtSft1XppD7LpzTYp6hloW1xVusOOi4Io17EhXcXITVFZsU
b282JO/u2P2q5a/zo4p/TEI5RCzG3o6kZy+J+24G1CDj5do0lTbV10FOiS1YEcFeYOHc3wssVJzg
8NBjUR4vnemzK6nMoYCGwQ90tcnKQQWz1wbv5MYzmxvxnlvBnjSU8i2nA/CfzjreOEMuzmyYdAlJ
qXUGoCYQRwS9VSoKORsZSBJ5jrnTQsn6eD61LMcEQQWkuamSTisudabepzXR2KfLSQrF4560fXgK
wiwVaYnaJldcF8P39L2vUP0bR5bgz8AT1djNlxq28UE4s32GbokVxSJ+aUY4XxlNZQdW5geoNnEf
nET5H1RGF9pdb1TqasOW9/DVJ8VLHCHbo4HBM0gO8lVr/ka/lcsD6aJhONMTJULi/LiGIbteEOUO
ore3uEFtngMIzVm3L20Am4gaAovNqSK31dGEA7hY8FzqFSsSmyTpdINrhkN5O9CTdi9tbpJ8sFcq
x2Ub1xznlMy6qNgW1ghitagdKzMAJGqV+VFYHXq11AigUU3orwl9bEwLn8wlEGz3W0QKF6qH23s1
X3ubHG0I8S9nv7S3vULEE/9XA9ZL4RTJvhCU9Ar/nprj639I7hLDCJ7r85oyaXTTzqNg9eNHT+xI
M4X6yNoEROvprWQkBi4FKCPirkJa1c9C27Mk+SgZBF7iQhmVlnv12Z4JZokHUnN0I3vXzpBHsqFv
an0FpVkjZHxkMwCwFkE0jGoKeZZwfdpdYsv3hkD4gyknbYl4C417ClHN5mJVfJJ6oEAyNpMRU4Fd
TRVMj8dtQ8lLwaw9o51cvdJ11eS3HXVa+YQhmh2afHHbV9qvSZQzE9kgTQn824tlmKeCcjm4yWFn
7q865q7qzfJsES/pKePL/Fkj/2PbfOotMSS4RbtYfq0QRUAsQcHyDCX0swP6t9drYwMd0pO3a+Sr
6Ygs2MXsGM1CtRXjLmwA68Wfzqhd3VmE0aGJdDgr1ttJtv2wJy8cgQgxdq09t+n2vv9LWOs2a2HE
sKM771TPDXLlCOGR/Xynz5jpZmIe/FKoc1s8GQpz9zVVsIW7T5CI2ZzT+Jloa6SWSiI1vqIjqOQE
9RyHxgYC7eJQmzRwgHxYu/1eR/+f6Gg6/Upofm3Fcj2svvKY+udJq6Cup9QuZUF7mcO/27kZjpyw
T1HHn88hnQ+fp8igBJQ2B/dsuuctHHzWr4p1pcPAdWmDWoSWcrUcPkMxHpO3/VZcCN/zqMLfR3re
KF59K9NkJUyX26cCSZly00NwDrctxjUfZgjjFIlmcbKp/TZLdDKnggL3Ba+3G06XwzCV72rkdiS6
0wYIiwaah2Xbu+uHoD+CdMui9bNegsaua+u6iRscbkTh+RRVTCqabWeHjh9ouQWmhD/rJ1LVC5lK
yhTERLG3Eh04who9/4+WNCfvzBKSb/jMtzFnzR7veSN3Atbw8iCASsEy83+Q8pF2QpOIhcP5d2jK
dEfYOMEWfh06iQj7S8Z25drFmcSXgCg9gxOQ6zet5v7OwoLAYtCLMsX6e4IXkS1hPB2frOQmUsyn
JEtWEgu7N46aGOjjvhM0YpYnbGSnLIUOsNU7dQk85E+LJdO5r2DbrEwg6y8JcAZppBN1ANC8ZqV1
ZcMa7aBFkLgYev23BhLdLRA/WU7fiejz/WM/XWn3hYDUK7lpAdRqHFOJCiHymy7QduXCtvymNbVw
rPU8HRpxW1XUpWV48VkRQL1bmh23J0KVv3ejFMJ7M2Y8J1ziq5fVnMFimEZZLaFGSmm9JZnBvf7m
w35Df8EvZ3sysbzGl+LRhrO1saqCKqMe7XzU4lMnH6lIV/AamIzXB+P5OfUPM8B8eeBBg1byhfin
7xBAfywXJnPNeIjFGWfz4Elzuw6Lp20fCFKHAXEqGbE+KH9NBbR3k9Ctc3ENE511/y3L4gEeb1Ks
h64vQfhfsf2lQ5K2s2evL4ZBem8ohubPso3Vm1NaUt1BSwK5+GQoOz8VvSYgI3sZNY1Q5uoreUzd
bc1/fWjymI6yl+CM6HcvVt4xFMhbfPMuvTDXuDTZp5iHsyei/cQbyEfCGYxqmwFPXE/heYPZkWxy
in+KOCFaSWE0dCE1xGcQ+7SMlS24+BFwbnh//B9Yd7PUMy/r0jEG5NS9cXLohlZWLD1p7yJxwGzU
aWjO5dAZgvxyRXpMFLCvxHi8ePbEp44Np5p3wecSykFM16foqbqnsNblV3TcRd2tC6qZfnsWixsY
N+kJCmFNTD3K9Ih7MnoUq56fLIxodGcmkmYRjBVZ5sU8acS74bgrQB2CkmKIjzB37FV54YZ6/MOl
Jh6kSZBUcGx05cy62BWySSP7VF8vRKqpWAyx5cMPMVAC+8UnTBlcZhoT+6UM1Xmou2OkmLHpBW8h
DIz2Di0U10KWP8ht5w/9ycrN0spCLFb3n14uvZn3RHrrgPBu7zsH2j/1K40exGq0PdLMV6xNa4tN
ddoLl4DM2wW3+vSaRAumDIl1LHTr/gbwVtNlSnzvTB29lESTNEYN+h5WG5s+G4S6TGeP0xf1IKQY
FzG1fhJ1Q8N39U/Oaa+Bu4HdeBIgyBAB+w6mP5HGIgE0kXgXWm2TqAkD4mj9IPpbkavWO6zXpekB
M3Koa5oYknP9Jcxrqg8CQ1TMWO26LhQqM2Ji1whWtcEQXbnSjLOs7PC7HOceuEHfS57lmz46YH8n
wC87GjdYI3+lUr+oYuMi5Gf77ae5+imNgZUZlNoZ9891U/GjXcAynX0PSV/sMmu6xdesGzYMGW3W
5MAhuW4HXue1nc8fijSitIF9Y/7aXv+MdDeK72H7m0YSSMt9rSJk972UsRSDOVW+kn5FEa+KIQwg
XyXLpjE0YBC/uiYI5spRTSKNdT90FUqJkgHQ9yLOVKFxB62nendjCdP0hktAIOj9p9MUq2z0N7N1
r19jDvysF/Icn8i7ndWTrX6IWSWy8an4EAIBgztaYlOd/ObRpuUpZ400nqNYcDyzS1O+CGj6ZOus
o2ZdZieu/pcxf71MOFWz6S4sGSczql3RRVWt2/6i8DeG3tXx74mTYE0K4JkoWn1Q3SAhQgHtV/0T
6td73AWeL4fygRteGgD43Rb6dctcyUe4v5NBBoLxSqbP4ebfT2kIXWLq5wEbyKCZWezeyizHPqcj
Z5+0N8TglEx2Rvm8uPy99GXo3aEfOu/D4mMpalF8bQWWN22sehod1rfZvUB+dEDPSk2SqQSS8Nvb
HEGBxSdArCLsz3/S08pD23m/BTz12JYCaykFJ3OUIV3YpTnnH3elqTn1Zx7jHt/mjCNHY7A1rFXd
ZnI1YUrFkauXaidHcK4VjTYjsr9XRkDge/LU7RtOjfuFBsaMrnyMykT1ml5IdtcnxwJNGASy3Ccz
GEy374P1L4jsJHueemdaym3mMJDKmZJotieVmJpA1aaAK84ymSO4wS3VVIpq/XcqtZB1Qbru7cYq
ozIssFBjnUSFhcs6fruuFVqUcrgJwdyOIBH3pAnXoO2hO5XuXaRW3n6pQRPiIwc+5stI/0f8tijR
6oLScXO5HGQkCkl7LcQid3CqKu2EuX6Y4qP8RQ3N5O3rbKRYXPGXl5RY045zkHxZCxAFjOUwWWZu
4NQ4RT4ASGHMDIOrVDfK03RQklwdmYw7+0YNg25Y7AuHkbwm2zLLQkrQ5HVsTivGAbvOOvqzF/9A
QjiDQRvA7gcVeYHuLE5Cl79pQEDc4Rfcjtl+1IL+pLraTGNoZzeBfGjz+fFREat7GI+6SfnY3END
bdjr4SMe2pX63cWb8gsLHdCDqBYz+wHmrlUIqJLicacBAsyRZKIgrotpGyJsaK/SZCSwLNWBtSMh
/FRe011Mn2akclIGLzBWSBouFzMjk8ZgDin/u01CJMasTyTOt9l+PABKR/OqJDliTpbmvRnBsCev
bskebb+vUEr4n7XLC65i0xDVzG4ifieX1pUlo8Qp2IJAkiLWBVm0mnbKeitHt22UOFAuTBMd5RKo
PHP14zMqrpxbUa5b0hUX7Wrtz3eWN5ytk6B5NwPGrCbb/KW8UMiD3IPPlgvnk3u39P8TWWSB8JX+
J3+hjZ/vsXyEUtCBrCsuclf2gRvXGj/pOoexs11ZPO+IzshgKhi0wzoQ+Q/j+JMSHeLqSSIM8mdx
MCr/Z2YBT7LSDMzvdTTQVqpvHpc8Cv8vX/2lLZRoFyU4t99dLj4qYVuT1YiOJYycsJ5RG2y46LeF
ugHmj6Xvc9Nhg44KLRBob3FwqieBwzFXQMcW/Krww5iiVqJOUUxmddEHW/OuCUAqGB9Z9PnzY4bo
QesRuj3PgUqmeitbmyieEbGGXtqABisawjuGMAb+1DtQQ9U9lyIFB2Q6FeRrw9/PyD8BhFNBqvF4
nsCPhVmu27LmSeKCf6rf2AAPgHLi7J9Ig8UHXRP2VXzqeqPscCGVemKDkDp+cKnoNU4tXvvKA3T8
C+AGqWBbqIF7fEslfcFJuse0Zq12pZcyy+n+4bXaYxmjG9rhDGwcjliTuYponQN5TucnLV93P4p8
hCUEVIGtnIZ2Xei+wzjIir5ugHGXMBJhNFBUSBFPb452OzcjxgDYFWV1AmG2eNR35sILBo8d1aA9
OR8teVTTRW/39KeZhRsM7fcoXhZArrqU8Wig7wJn3AKI2Ca8gzPrfamiwGGIxC3NZYQhdaMxfJrQ
qIuqbOQ0jSRnaAb4JpZ8isyyvg6enWyY6Uv9LWQpVI1SNfJuswaCvHX6WH1L2RuoaXoJ9mN2V4aS
IcmgCFSVdGtisZx77qS8+/3ttncnOt0Fuhw36nqVVXxAciUBMNJTjhXKPxHj6SkAI0DA1TDMsTrf
1AmX8UF2tteKwDLWVnZ007eYCqkPQpFA6ZACfjeyGkQXXGuIIAjhCYpReCNN850CbMG3grwaaqM9
fXm1dfHAnUZVs8ll2OmPwgfoagjcij88Hekvn5muggp+K4IK4NuLd9u+0xaiuf38jJjWC4ygZiDR
ISmfhzVMXWPgPEwbGKrB93yYRjSNQRX7yXin0t/bUqbrC0fb4f2rjuGVCwrq57XH2x2Pit1elcms
B/zW9+S80d+joqrxXmt7XVKNPqPbgBzdX0RhbwBv0q/29sEyagIU0774MLTzuSW/R9h7wjVB+WCe
H4LM6bfUb3ftEph4W/i9CZ3wh2lbPkOgY5W/wXuNPz2Dlc2uw0mzn3LleSgEjNnE9rItsZDrguX/
WX4VxBecY9oCRjesMdDdp9Aw1ryh1dTpWL9/OovR1Eb28PxFDk7793h51poySBrsLae6iUyGr6s8
i0jecrA+Sn2BXQl0MgPkfdCFCp5YMEnn+W63ZXlJEXWqh0IshN7ZWjQYPXQaLgYnP2Bd9eDZr21X
zFVaWSHKb18rzGzI+mxXVwi6itPilRgQvMoTxTBMGkfwySBM5OfSAgnK/AfHoNJEcG0loUJaUJBw
ZuQ+6eYhXJ1gngbkF0CavD6st1+36NqIHYZAlK9eQeMuDPVgbPi2uo2fTR+6lYqtnU7kRq9UOoo8
Q1CpHZ4kN5CtqayzmK7jntrGsbZqUN4U6gTsgjb45fRK42OYvrzguHnHwjjksaLMEabm9bGgeXSh
f5mBDvsPaxS17kP2GLoxVMJS58VEyM+huy9Og+69meqOL6M1auDGanqD+fZqQx4leHPAjUdlHEeg
2wK38bLuaX31Mlr+HuNATAx6ZrpJlQFN1akwWuSlPw7YVwhA6C9FJjjoqI2JuDIbhw9kXa2Gie/f
tJOkuOgkBDItLv2LyPx2orrCqXf+GWG5br3O2/kEt5rBolpEUjsLtl74LOw3njGF9KxMOocaFAAV
LkOCrQlFOg030gDL+0VcHESSogVOJxKnuAu9+3W6yyAacbfug0iNS7l46BU61tA3IxuAWKcvXmni
XJE0HYpfZlEhGmUV8F5vbG959LDutpqyXJ5iYIawxY0bMdqXg3otTd6YTgTgE+0eCpxJlbzqhZ/w
5IvR7vIJ6YsjO7GlKnp/MDC5EYXUKmdZCQuGDhbQ28ScvNe4smjVrR6OF4GKGekWYApvA7KtMuBV
aavBqhCAgvf/yh1hF2oOwBM6GtRrt8XyPam6U4nwJUtDbGH4YoymLJgoI+RDjz+FC/LjGVhYWI61
IsfnFHpDSJkU6z7sam8bPQ4ODh+rVtcmNVfoQdJshgfVfasQpNiWZgKtVVEwxYGvYIGaxs3hYykr
64Cz9CeCjDSlwwZT2paEha/+jFXWnzSgGtu+oN9fdhTGfXSj4o+LC7nMsDowtmBPcOJWJwEDnJ2I
WJHi3m5ikbhDIjfiS4WGsKWBuPdT7nb4QoqOxSpe61x5HiPxhlJBnrp4Eo3Nrts/drskegMFGPko
NOrVMgsXyZ9VLtw4j65RG6JV6D4ZCUnhE9xnrVAQ9kTnyDy5+KDvWj2nxYMz/08LfdJ6R3lHiNe2
FQjWxffTQeZcBR/qAwPlklMEmLnsIfaew/44n6kljB6W3cFPD0Jdj1+Ue9/E+kGnjBWh0WPYQy7A
NmFE24P6u1s+ufU+uaMLaFze5AD/rGvJJ2vA5GhaUgHE7TIx04o6smTkOGGAgbE2Kaf9uGGSbbsw
XypdD760KmKomxKwf4E97FBrqbtfm4fwR8nvr60Rec5Bu0LAuZbUQ9M4BeCrq8cbC9ipbr08Fs3T
QURc/1nSob5pbr89pridOrRX1LhrIhOdU6mFVNabFUkhlHioUkN3cjnuykmrf5EvK8z8leOGf0Ah
kjcVluzY1zcaL9H9ImIK5XocVHNIg1HUZawhBuWpAKzrx2Njk6vUy1eTpVkNEFICHUBaCOk36x85
9XJCxfEpeAWBFK3w+MQdxWOxJUEFNQ72DOVK2sfL4IaszMDZzUBFnZ1dvEbMBPG6nO8JySN+QdV5
zcRj2nn+Mi1lngEAzs9LvkKOpF2pY2fIg+yr1RbBkG8eFqlpAJyHtwoQhmdKe7YklrIJDltWGznT
ZUBm6WJLtxOb14eyPRRoI5RQzJOGNStVdnlukC1F1E9aJCDu1H+2ID8d/g7biLDW6A+LF6DRQwUJ
i53kIsW4ez8bVILeMY+iUbIVyhFX2UI/5Jh8rEbNJyFEj5U/wQg85DO0WCuIm3+85PzgiwzoCetz
BvKUrMpJ8F1D+2wI+1ZSTmS2LitttOaRDwx6Lfax1/MpNMAugnYawYf7Hhbfrd8XgFYXJuDifoap
yTWMKY1aREhL1BpTmrtfN/hHfA4/Oo/Djgl669R17piXFC4hc1F2Z1WFoWEMsITm6ilGrVqzQs+f
IpMS56K6CJ8Ix6hRE61BObk6mWrOV+2Yt06wfw7bDYvb7ETcOJsIezl0mHI4AJgHpuZeVXbWBC2a
m4IsItexmVJGnrBi+iGE8lnMEBU07pMncOgJ03/86LH63uPlOfRvDkpKmjik7AepkhYbIdWj89VR
7fx6Jra5G/8i0tYE9MUW7neGDlgT9NCV9YN9J5u2QLpn49y3NNHTfq/z05n3gas3rNiTcselBCNT
B2tDznKXKvnosN3EyxAywa//lmwUMYRaQcnm26o0nMF9diFEiIonaZlxTfclRJBPK+wYKWh848lq
L+wN0WvnkRsg3TqiHIkdtSXNUlKsRl7q8iy+N4pcso1ev+7OkPKCy4GYkm62kg2HHMBPqQYqj5Ee
YfUBIh9wuhxQ73TmWMmnz6wEEQaPpHNo3eaZ0lNdgTmWDdy8/oSnHn4cHPRYMckFUsvayXstlut8
YhCmOVbjZQ28vRhmf8xz8964sSs5c1TUBXoX4X1LgXp78ihmfew+1HevPoevpZ0R0D9OfqvR8Qaz
zSVinMnb0eanc2Q/A02bW80wo1xYXYgrd3MuFyTEdNtPRty4r4Q8BXTBzUTMUgjL2G8dJfYi7XjO
NQmtHlrWxl/OYJ7LFXrdSRxh9nnttoBkW8uiTAZOTc+EeukSB+uezg+p6zL/GKiFuNSGiXhERIhE
fpSHdZoLUmZnWGoinfOLreC/NtzLQov4Rc8wUsjVa+ZQpAp+0wKgdhh3dylGsQubVmFexwz0ut/4
KJRbMcRGQYttekyw7KPjZOz1nMVYt7MidrbhpL9nDE7YmyN6au8yeAbzeJ2y/fAVZnFd8TFIrgw+
A/xQTuJWo8lWY0oYY9WTtazzVGUWqhg49wpthGImNC8n8Q6inctCIYl2yv2HTQ0fT5/x6ziAGGxt
nvx5tE+fvkIsFSa4xB3WwyNlE0tAx2ytZ5jTR1GRqNNEiBOVV2Rcv/WPPIe/jjqBF51wRZtY1ZTO
js9yUqPCFMp8DuUDYbTc9auCF6tOS3PJ4X3WeWQIvsr9nx79C1uoF7LnlQ3iBlnQBDutP8RLET1A
PIwEOIMEyyzOtxTxHNo8Htb5fKCH+kSEWEm0xg4qFjirDsLvN1MpbqfGsixMx9LMAfLDpRvGPKWp
IMYzkpkI0nzWgVhExyevMsfaA3SsuwFcVCwRF6vf9ZQah+AaB4fZ08Zxtxd4xdSPM4pP2SXEt3np
pfxAFwx+feO3Nd+mPUARseR+jVEIlRMbMYWmX/W85o/W7KI0j+f5IN6Oe4V1PVjcITJrWi0gOLEf
aRtuV0ZnQNJnVuyZdiPuKwHwbiJW9s28zGjkdRd3CokamCOOENhTXAxhpXFBvk8s6ovRgdymXjIL
WTBvcK7J3NpuYYtpEQa/cPHBiqWd62ktrxE2gS8ocqVCJolZMHhozSl6OI+ag4HaSdYvxh5naan3
Pms5I0L+TiGj5/oEXkBhMUj1h1dHoU9clMoaHoqvLasF7YzCwO6rB2WoiFvToYIGTYZpjalRND1h
sWORaAKvsAwCwd6E/IZVGSWZe6ruF/204RiP6ZF3wJpyHViPlJh+6A8wfUYCJA1l0Q9WaVTIb+CK
ho+XDmWlf5j/Hvm/V2LdAKXdYITZ+JYLuxAstoc1xeRXekVyQ/ZtrbLqc5xIuDblMnDAO/XU2xh2
c/cUOzSfrVzJiQ+z4xM8FjCPi5wuxx5ULwXYCTJ+BYIvDMBpcnRS2JUI9wXhV1cF0l9QM8jWuy/A
mdxaapE9pvxy/YTd48ByRBQx2qLzPl4/ZoQ6ZXlk6q8l85YIMShV4utofumNbGXnTd8h+pW93IfV
URV9rVn+t5RbMB684M9V/UvCu7Nr9WOzmjqkYPD9VVvD1fO8LWZ/kS3yjUkDl9PZ/KbTzcK/jFcJ
UhB26VNEdQqqK5L8CFqvkyP0UbjRWlIhc05soHMtjuutUYWLZs00rO3RyJM5tWAe3TIQ/Hp8Fdrs
DVxXb2fo2O4XVtOvlFZVW/PuPL/S+jLXa0JcTxv4ZgP87cRWt7dTq8LlQqF4x1HYSbD0rP9WNzyK
u24yuSY+OGFj7qdajue4g5po/9yIpA6ttbbwy8rnGGOWexaJlPLsAA53RYpLw7gMV+TxS1RbZUNY
sNUMHOS3zpQrXuYXlBmHuk8Ji8vSwHq+y45Noqs4v8T1KBCLWFhHjOGU9E8s9PeQFuWVHIDSLXVb
rbCSKHepEPvcPzrNii1ARpiTqMTDHo/H1FeB003/TrXsk+zEUgPe9J8L0HzMu3FtbuZYa1/t4Y1A
pfsJDeAgJntBBMUuvCo/Y1nYiWpDeCBgJlK/Oy/RgsX3r9vg1bWCfCXYJEQ/pEzWYvSEMtDW2fOP
H4ctuvK+DwOAnC2B2U390N1IIAJeu+OI/JBth4bkY2DxO40cqiJ9PwVzpoLmO0Mpf/iH7weXMRt7
CeoRRFahCPNi5MJDXaXpXCwB5DflTVhKGVMt2/i4Aonv6Ygz2GMZxAh1cUhog6DpdU9pK1Fyg2Py
uo1cs4jwHY+sFDTpcIlW7syjK+ioD04BlI1YZ89xJlXB3fQ5wPQi+sGixiGOPHV+kqAIp0nj5UO4
C5xTfpqZYoh8+e0Q5Db1m7kl0rAmX3dlNshPhZHuAcG8Gp2Bjvt2wZbivyyP50qLffJNhzK4BZGP
aOobCjGRwfq9CZpGRw7Y7GjRY0tLiVRteL5NYVr11tWbwUBBRSXsFELlgJz50KmYKaY7TQ/r97xv
U2Qf1e1vO4tCKV//zvOoB2A9Gyhk2wTl00+qm+6jPgAov6TOLAbfWRVkv2EddepQ8bJB/9tr5gvp
pJWK0LNJfgAzMzDTAdd/wbvjveLK7Wu8dhbNQADSIqafAEiNRnNprLgmy0Ou/8DOMq2NGa6cL/Du
89mzLs89Tfn8Zg4sKlpuBSy2VKFVrPP6AaS+eMqLMehHpudJvO2FYQ+nwEQRFNKlHZ0JAGDRLWQ2
7HvU7ztAW1WMbWox0jJuQ16wIHfifJ7YkN0Bt2AM0sMMESeVI23y4s9IIO4L9j9JKz9YWDTulhqC
VsWM9TvVEnlAHLnJYf+iqr2+9q3+lxmib2EetQx/LdJdC7ZmFgzXpwsV1QBGr1V6mykCchz3SYCC
g9bjN+9nbYSr6dU24ul+erROiLyjduRGUvUvx+LUJ3Eg1mOVz61dV1emUBai0mu/TLMebsv0V7Yl
/OhBTnC7sR4HYLeeqZv5kCs3RXla5FnlW8aQ9HHFtbfHMjr0ObJNzdFoWELB4AuMAvvgr3WEcT5n
SAYzYWWs0s1iDspk3feJNHh4+nNkoIoHYoV/ltgzWmTpUyon9ZhcHZuB1ceLNTIZMnS2yUEV/+AJ
9wa6zUWXULx7c1pZSkDC2jRBiQXc/n1sNxS8tO9GKv3RCq8jrBltRLP4fxapt+/zjXlFutKX229D
2xDC4ZClTL9C4m0I5LXzgr9/dn3KYiZ2m5KZd+qxie9+XK9i7bTKjGvtlP4RFFfDnmB2PBKLWT88
jo/tGL9xnbQcG3UjCs/2HkUiNQN9PZ20lMreG1zjW2rP4D1Z0Q5aZFdSzxf4KI4NqEvxxbLCMJbp
fSuJFjw3rwp3/tMzhb/OllqWvMMr/1Uqt/MCLnsT82BNkjtViBTCNHzxKzqL5xyMy1QhebYyrizB
to0uY92Nu0JzUGFdzNIfYxZwySELwzE1fKHwTnV/pk4Bni9hmMXk5/QaEiQnLAcPM3Sgtz2JxE8c
fFLV9qQSXQaJDmD8XtkLTSKNFLkx3ehqQ4w035RKTumO43IhYpGnQkO4pQAZGn3HiiqZxXmjr6Px
HXjzc1EMwjj7qx3d2CcqvsXnJ9RyTbOIFAGN+8TzWTHBhWTwCsvfxn9N5BPgATTMOgqmnwC/QlEI
gv8dSnJEbLamnzSN3K7tpAjgAXsZW0phgqXrzc02BGN4PcZcUM1faNy+PLRZAjWSZftMEgIK9ofh
4DIAYnAEjQUs5dCIIBNEjVlO4RZzXmQrW/vsvCMBeQf9tY1Z8ZCH9ofxn5sLRDS+TMVyugqampHQ
A6ENrAuKSQ3Zu4plHUvO4kC38BTwboVzMCe7eACzEYtMemiGRhth8JqwrQrRjkhRu2/VwDtevrY/
OIWxgXglECzN1LDmqvIsvjM4u+RTadFnFqaAnKrrCbpfFmDjkhfkPSKPIgl81aKUM42V82MtntcO
t6w1t4xSN/fsnzGJ0N101bRpwA+mvPP/2mxio9jo+uScNJvcc+tIYnVl6IDiQ8W1taPyEf6qYfsl
k+2dB0EaWalaTnNiUZceaZa3m+uzkQF3VuQ8aA6kN/d37RnicK4wVCCZomdwv7ktgI6+UtBhQV1b
I4veoC3Mg7iYMlnX1WGmJN0sfON/REjKECWzVrCagxusMk/l2oA1b3s878fH66QmOnsUAHCm0Sy1
g5e3t6833yVZ4X5mX8gf7tV1JE5dksCaKvwq+aTulkz6qRT06IQEnSDcBs6dssLqpNsFBRuTiEoD
xNooGXOzEYtQyZVbtf4dbCPFHSRNvt0QM7qe6UXqF3WVboo9WjXmvrbir7MoUjWRp5MolTwzox4j
gspuyxrW6OYRgW685LUNDFjUmZF1rHTgNK6I4GhOr0A5jhACcXOtcGbClIfp+UfGmKTuvN1s5TqZ
HSSMiK4FpgfpWauwK+u6JVSSEHsnxw18bcakbWYPKP3OsXrTyg6Ev+BsfHe19Y0i/sFrcyZbhng3
YouLYcMQg/54uCL5zgR0NSw3xPQ41XnziwYPuRUAoTYAhc+yM4s43xwQGAKfm0RgiDP442/WOO7B
i8nF4bEI+KOk+j6PKeeccjIQLv8FiugBQGJEQaNDt/cIyuOr9YTrfOfoli2lOsm1N3lJDfs77bN9
O0E55hKuDqMybrxwvcJnhXn4D3hFwKPbV23PR0AGa+4TPpBkkFGXe7uhVxZ9503bic4TJVW12SUK
uU250LxLXBtTpnHnk/MVzg6n3ZB/HYiGjgSsE7VD8DrAyQmV1/dBKQfQ6zvXTUDdhgNE6vhrROq5
aIufy774iJrbJL4IBEwMtdWfzAoPfSjQDLGLHMRTvvyYPd8KMJDNR7rGF4/B39VZ3ddz8Id0cjPe
ERRX5j/cXXjcedvz8XvKx+nVNCF3yUoARBtfsZjKwb/VsO7SDG8399Ll5aeTJ2XZPRvU+Lg83vEq
i4cT2EseE5CfZasQr37neQdluM0N7yviPAFOGw8MXV1W5BEEjYc05LAb0NFpewF7HNRuk50zHxWK
BktcVDhRE82GzdFD5Sz+Wmq3ip4wbB5nUNLiBS/fsY9bp75V4BFB9YaVkmPRdyrwL8CeeZf0wuTS
WXUPPG6yrK1hXPrZx/BMLjh7zcN6pO2MkdYrC30cOrlwcHR0nWjoovqlMhZcDTv+ihat+9+DqDE4
A9A9Gi3+UxGfn0YAG0+MEAeffd5KscZub99/owIcKeW7uGUL0ZVildUAWA6IRkLQxD6kLos9/5vg
rEd0yM5h2BsvJLp2zWpz0QtZN7dAL9fg3TZqCff3CCbTxft9m8S88LOTiMwDguOH3JbaGDsyk6kh
jTZnngnB/tyMoCyEDf6zREfe5z1fG4xdDlFh+2G7kHOGEwEzSmIsRcVC/p0pczVp8TbmnFTJAavr
Yd7LFU7pcqLxVLuJIzqVLJbOZabClQ02HA2zTNTVlbDzboI67+yMUX5I8ePfPAFhpf+x6yIfujMf
mEhzfXyssvs13jrW6sRdwIdWE71QPnherHamZqmOUhUiEGeuqNnpvHAcCcphOeFybGdB02InhXf2
HRbLm07y12GDcqwrtrXuDFKyyRYe/P3sUCB2ggyYrC25EG/Sf/ui2I0pLFmLBOdL2eO/KGkHeq9C
KPZsm7GUicKykfTw8Is77zUJh0g5TZ+WdpCP95/tfny70tLOnEFv0SnLh9BgmJ1sgl+HogVF3tVW
gj6o2C5m/FAAy/2O33qnPBEh7hcVCJ2KMWUXf+r//+Le/TSMVnOyLtHrFuT8OK2eg4F63rU8ohXn
FgBeyBiTTdk4pkUgMsH7gtJLsbUqHHYn17z6ac1uc8s08PQ6QlrNNXJALHXtZ613YYcPywU6O/ns
My0SD3byeBNjoIJ+yuESVg+vC2iHFP2DHB7BHIvcejlNUesoY1QhPs2Q1ckEQMDfcRDwoRVz1yib
mOyLYFVeqj/bASYwXBbNNODuR4g8bebBVq97LWuwEnXrBfw5G78V2X6aYsIVnRMoK/0yFUm2SS1w
FHF4wdToDGmGMEV07Vt0nf9UwbzcTI3+5BclzKIujVL2Mk4+vz65jiszrCBhMfOGpu8vFX5VaoXK
m6RKf2fKFFt8Pimjez2v1s8gH6f2ACmAmNut2ZdzfLvTo54d5Y8cHpc77GHSIzNSxQB7zpLDomVQ
8cUyjUwiuK2HNpTlelt81RyY8l9P2lh2chx5oT5MN3Nnxo7uyIT+PVKVSgi8AGOSfeu7K9dHhYKd
RUT8DtqzS5v665j6F5uOHxHYKj1U8IGcCWZtVg0W0ELUrEU1i6KGuwm988SseimwcZY63EYltFZQ
xTjeBIfWT5WU9j1UwqnE7BjBdlFQEX96s0+xY40k+uiVzS4gYsYSWntbH4TazwLqI7PvH7sz+ICb
Eu0HAiHfRj37wV7Y+teFLATC5xREi/DhYR1OIYEpHLsm9Zpq3HRt32Lx4odXD/LsHNfIV1ksoWGI
Lz+wHUYl4i29oMAEs22qoMDgGXdvSNFOWvpH89egfg9/wl681UZy6CzFSbus/pfNwwN9DeFOJZB7
vjU4NxmkTIwpCVW6QTUTMXQR2DjbXllWc87Xv+pXNjGWxR32WVE/+8EnIoPKWn9J+5bp8mX10VfT
LeWgIOgQbQTb3ghavuhBeKEryzDhk19VMmiWryX4ER7rCR8kYuLTtziNkhkKhO1vq9XAq0d4tMSk
YJInl69U/u38b7bCMD3rGOF4AbMuz0r9hCUvgBTvGdctzXYuXokhKSfFF0x8++frbTOCFk7wQwqy
9T9oyXJrA46Q8/hQPNfCB4OfGSAQWpNvoavkTeAyLdJRoIluEhgnsx/7tn4afoA1IvuEF19ge1Z9
VX+Xnpwk1pJPFgnRAu99X5Q0rNKdVq3LTmGQd0hLrGQ3QhsjNkXWgrzulMBeSQ5+xMjJBjHvBP+A
QW9qGdk0G/3G1n+uyiCUik5x2dH0iALwbo6ivhGANZoU2c8aqwzP7MlZgXMM8Dyz8v19f2XESKDS
mE+71OwHmVvGRUD4ZEgFQcHR1MkUKYkoc5CDByowE7fGF2dCBqCnnKlnvYLVZDa5E+89NdiPYIla
yEdP6t4sbPdOT0yJjeVT7pCQKc3+9hcm9OBFI2sH9MZVcER7+98IQ6LuEftgO3e447/2f/E/4D3f
D9nF/QHzuuCZSFZUUbX0dqK9kc+nwfl785tCiwqMPgFgLwitUG7UFygsoetLsa9F+31sstBptvUq
LHdYoW58K8m/lNO2IgveliUtbZMLR/LMtZvoROwLIDCQrwE7Dz/AXnz25BdOSNm5FZip67li+5j0
T3oyH5hfDd1gn3wMokHdEdyG3kV2gyDsxuPW5AaoHx/9ot038o9m2BXjy5XRkqtdNGsgDgk+mWPW
J2wWjXDxWIVHGbwuzv9hW9CuVvu1kUifT3y3eY4tyP3oriPpk0rbgD/KVfN4yN+iYw0yxDpgn9tO
fB1vxtRwF76+6KpGHcUX0hsrc47tWWBxvRhsfuaozCwoCCYN62F0B1+pYPQQMwRbvWKuOuZ0pczu
7RqdGM9ys+Vlau1JlFapqpFY1HhD2OtwpxAZamDQoN7fHg+C45XO6njEkckM6J9IvEPa4ZZqEIDz
Le8qsbebofGO+rpNbhjrY4mBTR7c9M+rq2gfmo2g8WRChSXaU7H7/2ZX8wC2SKkRWsv+0WBXhPkf
i0OhO1SiS7z3itV2Z7+KuP8s3drZlId6LY4WDKo2TjPCO0hajCvhatjCvlD5uulBYsvKcFsTw9Cu
6qp3unPfwYuQE7UNcBxXMq5ZjEzH841UclGb25/8hvcy/HVEcDXjQDiCdFpzTs4laZcbcS5cingm
/nWGed7CUStr3wlgtuN00upd+VndpyI/QRDuFYkmq+4MuDJdoT1BL0ep1Et8XTJTAjm2A+SViGgg
9XbUJbPj52hReJ0ciETcWSQoWTNQC6V58fxbIuBaMnHBYTwrX6IWojsducbolRg49qDzGJazS240
eoV/ilRsMpFyku/xYTU7ZksJzmq1PaIfbz8GzWePcD12jECccuVKvz6/BYgvHt25rLRC5X9PC8Mu
Uu5/9qQZZ0TKWijWSg1WH8j1bd/O1ND8hJGppmaJAsZPcMRqpdZIzZJQe1PY967yEOfEcTJvFE1q
wvGG7dDbv9/0rXIU5yVJjM/dIeGu+YqvFbvbQpDkXtZaDb6I4XE8lvmB9uT6Zujj9AHirgDg6JKJ
pawk/tH9e7XbgTL3mEYgKMWVBYCarMcLiissEffOijuSwI8kAy78/FVjdJVYHtzDti8XPKH9XqfN
O9UqgwUtKbHiPfeE664IhwchSpkCi3cQoEfbHqRPrFq0yK6DbJFHsJhk/1PML0n0CHmfFvrGuP76
gTsYmyKXtbGg9KBXby09xZdPagd5SuKvfKOjT/f9TZI3e7fs1o4sb1TUAb708q+QYtE89Oe7Gln/
hjnMQlmexkxBDblFJyXMyAILJdilZvdwkl/dlom/JprCaCy+8sZGL1AdaT/JKZAjpHftN/mW3udQ
Bp1tXpN70oQfYnUjnUK/yV5T3xcnD3g5qm9BoqcC9Pclb2svRWWOU5cnQgzR6ub4zzOD75Mu5zT3
Xnu/go3kpW6DOT2A3+BUQTzchTKd5IhiKoxFSJJs3VUAOv5xgJKRe48xTV+YuaolMkLv3Au4Ul63
RJDOWkxOZqrcAK1ADnumRg3IdN4zY4eGGLAInEupFq/m/jy+BBlNa5tt+3VwSuHSf+xXGwSUTcHK
xOtLNNXaA3u2JlWxR/oiDosEkpSQ4e+zmdtR1hnDrm7StPtggZtv21OIhqpaSHOQYBzisMsC16cr
G0syusrTZrqkhvfKhQJ56cGUuUxTFWRhuR2caNDJ/jUEAYNzVCbVMfe2O8h8TqpIErWr/y3X7rw/
4gDGKzh35gMenMSueFpORD9oWVlP9bWelP8U3ymXbPjPB4QWorz+uk3p90epUy0758No4KIewzpe
hRDIO5O7z0JTX395indaGBfPQzw/e4WRtDJJP+8/h4lZVfN7vna9wEPsGHYvH/G9h7Ira6lzaD1U
YNXqh5aLZgTbIXguSXMYF/Eml2kCQIIUTE7AtGDMWWACpmVg7Mxp7++7YYVCWKlOfikYNSrf9Mbz
ZUhANSvlNaCpZQrndxlw6Gc4MJ0pEinlGoBnxNM1wck4kr5lD4zJhREF7BuzaCc0/wX2SeWo7vGO
I6XHHl9nWjMOC6/p3ekLn1Y9iRKIlOrGth449xtL5tdOSkoyXSNAQ+NQKC5Wf1asWJvPX56gftlg
uVa4vIdyEzHDF2THj5HCHwnI4gIUiz2Kfu8fvRjOIUDi9GQk0PnseHG5OcRiJZ1azKxB6q+caN4b
mkNz6xdQTc4ZNLnuXDgfv/ZUMfz2E9IX9XKDooutFKtAea4mIpt8vPZtzB0K2/Lk3HI5ct1AuSKX
3JGIOdgsyQZLUZs2WM6qU3Ee0DDY1G0gz1i3+cNUMXxhVO7GvcE/mTQEOg8GrwQN0pYcA6TvWYEV
3MpO/BS2IGLV4ZrSoans3fSOwVhz4ald3HLBTDjhij6hjilz/FMTh1DrPXM+nAjUl+JV4DiSWP4S
cCrzN8Tkpr1SsxICVsdC70P76XnatuKh0MVdkmRFP481YmCSHyLIkXGwp8xpfsxi/Yt6YGcCh3jL
NuqasRFgEYwDODfbQ+w4jTN7sl3SayW4mn5GZViVIA8veoMXWsKAR/Q/ZrMl+q3v1AwhDIDmbvc5
MnAAEr0jzoRkU6Gza1gpfHbJxL6z8/RiUfCuk9+PQwEjHdzlVY3f/+gIiv/eZaB9Q+l7hl/BJuRg
cj32JYJMH+9ktnRzC6RUsgjupulJuLBWd4Y2cmYxrjY/OXzP52zIxxl6vPHecQvOw9ZNlBg58LY5
jfENpBUvLlLx6wB9sn20PINCJ/mwsJAVMYeNdw7qiKPiV12QFhKuG82d+QzIIKNhTEwhW6rhBuPR
LLUXRYYHCY9wVxKX3hsxHspwoUuw0+rHC8AdHdw/0XPfNPLAY27yEyxXAocNNC39uEv9yUTZFM73
Z7IyDs612HtkpBhD2dgiZhiKZXo2M74FNwWJviQdAEfrQRRIcUjnkkpK5eR9LZFLm4tNo4EqGfwh
LuTm/OhijLe5BYauwrBfPzCSQ0ISO66ym33+Umtkj1r8uyVIaFuY5O/r/xpK1hy4m7rKg6fnU40W
V/YN81WCTLYVPgzIlZtmu6ypwsC08B8PzEepwaOiC19PtLe1yQcpMrGC9fKvFNTH2L1IKYj4FNDB
sHMlx6JlEpacPz2xiAxIE1h6yRHjzFT9v29jA4gEBSIU2/I3gqxLRF6FSRxcyz6ApH9rPAAsGcCY
UK1rzK+CVyn3qjSfnbQk1LaRbw+IbsmEXVnP1x6xkqWL0ozaTfKTiqJaid51bysXHz8ESn7KIEPG
dGalK41lnWjDnAj11o+Is8TwcxqvRi7hyGkt8qKL5eLkHCD4vNRIM0C9XOnX6m2hMSVdtyZl4wzS
PS9h40+akTJhL8oLTwggzpqf120Lr6Ex/XlCOMkyBz7sftPdexIRbh5TyVeIqT5bWs4oLYok1uCJ
mHeE/ik44pMShCJAC0y95/irsPyqXYQs74jcMTCyvHYyG0sH+BjP2+rYEwGiXUkesKAnKYGXYhSL
4zQWbdEa2E8j+OdLjAKCLDW33NOru6V/bjBItgxcrSf4Gqa8TExdQFxgY1Wn+Dv6JzMAQYy5sx+n
dlvVxqDXZSqxCeyk/KqmBo+PsYC6w51fUqtVcqItS6mUoByGdokx0cRJu3fHhAMJ9SIFDzczHVUs
7fKTTYjlEDF+GmuqxdKsaxIHMR4kOOiFhAhbAYBuwNSbGYLWOms6nO/Q6yunsFhQ8Y5HnxQpcKJx
BfdKxnvv1OVOpAVVncll8DyFHtPIVnGPp0xOdQFu/VWh2fZJYnIsp1z0LC0Kbu0pF1VV+B7Z7FRl
fPNPD6eNCon5XpEGdl47pTGF6YoXP6qAMOSo2FEi3Ma74km514f9Su40/yCdtE/In1JeuUhrgo/7
LRPzmJAP9ARJa32wzKVl9NsGJue6g3iWoApwyHbL4d/B2Twy4tGECh6Ly7erLJ2rrWs62Ej/r9gv
4q5Hqlbql6H3C/npnQYqdK23eIadLQk8HbWB09s9yESGYEW6NXTmyaj3tNGKw0ekNUvNZ7+Ot5Sh
hz4vUkld3PkcGe1YmdQuq+2Nlv0ZGGeEcUdwF+OsZA3vkDWV8w5KmBZNzCTFpN8Sh395b30yXaxE
bacb12G2+fCdf8KuVrByPQgEI74fOBxMSzyk+OJ5ToMylbuB3EqtLrol0mWrqWrfDLEihs2GZHYv
gYv7dzZReZ2/wo33vcAfieoYL61dnL5O4eRQWqaVMtGo6Hm4Ue+oCVgv8jjvBGGA8RdSdK685LWQ
RB4ss5JpK2gpBA4fVtZ83vXvXOns0VKJBw+fNsO4JbpyC78+wG2knjSZ7eSoJXLNXmTahGQzXj5r
XmQ2ZHh4uiNs44sa4xLh744GL3eSIlDHSdloWydilf2pvO4jmf5rrxnS/lMRjUMBPbBgTVwb52bs
foc6yma0znE4KAI1cf+4I45jL4l8QXZz0dMO5m62AlHUIxhpQEBn0lMn7CPq1v+keOJ2Soj5Ohhr
/3wc/1XI+1chQmengNHyE8fc54IdXsVCgth8CGx1eecT41J4gFTlxGxMYcsYftZhyq3yANhn/4zV
YCfCddO573CBtFp89vHzwvtTXcXTt4cCL1FG28p2dZPTNJVWLlT5DWQA1LgMfmGEmauiCuLRsuJe
KUeOqIVyBQI5lT0Nm6o08jq5/jrXZjU9pGzRAQX3+ZVPujPyfIExG0vqGRogx0cJR9Dlnm4XAWES
7fMib3BUqMxHPp2nw4XD0h2uVF7BBPhgKbGcyHokzG35voBrYUuLoxp3IK1ihTlLulti5JXsjs3n
Bd/Z/NoNU70zD16jXJaadjEhSlCYAiKL/PzeqjtaoDaSY4V/wjpj0xxNLqnKVns+So6tjhP1Xyk7
FNtHHNlndW1OR7XNwTBf99zfL3CkfVjgLRVFJxLSt23OLu80pQp/RrRI1EiZzsw3cE63FhvXFxzO
qCLsbXmcFmZyKKtxgLTbavnbT4lVhea6kPx2hojmqP0Fnw15eAzh2AmQo5aG4ne+rEt31+qUjgQy
09FH+j2/fu9LADoxsNxb0piTsTYUdt6JQbPJpwDxW/NnvvRQtI57vWOlZEA1bntPD9xqXlbdbtcL
y3ewE+e3BOw6oOejbxzB1eOv4nYmhGIOlK9q2xe+/iphUWrVKOuOECiHOry831IOkcIBzeifKu4E
PRcjsHSpxmV0uVnHDUtWxD43s6pQwpXnadjc19sq4ZRoDn2+e99CN3urjH9TiEgMZ3T0OC/aM9hh
cFtEQypr7Tu+2q+7aD18pJ3bf7DfAH3XKjxKo+iAr40yGJab2aPyyp9daxOzgNs8TatpiUbsOWD1
2GkRrH4HlCpiRqvPgiUM93XV5Yjk+IwT87NBoSxO6I8jpCFnU0uL4XvQaHfUGGddsGacYUzMEgRw
FB9qwTDmJs7hlbtsfSEKl2RHL1Svi2dyBPEnF3tVnqtcRz9oUIrcaV5xFxQC2Z6/7M9ir6bLA9ja
kHw/Vx9xEyPXDBNTntnK6pp6aiACtKOAxKCiGT7AGu9vP5zdTNaDzGXy6lSImSxj5MtJlXMGQ5gb
06CLKEyUaSFplJdTdlrhM2VL9xVVyGnFdnRgTaXVeT0d66t5/u9iV/4ns34pgr1OH4aUamADG4ol
+vxrRxj+rid5wIsTtHHAgvYg5ieffTb16CRgvSdsffK3UGfnDgDL5ScYQ7RSI4PZCSqR5Z0xMy5e
NMa18XryDu0FgXC4twwe9ruegDRX0jB5Ao5IRpdto2sIxnHj4Os4+SZzFtHtJM/2slFdXllONk1Q
TBVnPE/opNeJ8BvPRaKNZ2LCbKghlHhPxrBOZkFiLNDqWNCtTNMf6djrQivpQ+FDzvIxk4okZzVW
jpUysmqQo2E6yBmMRJXceQj8Exf6QhOfRrhZ0KzM+CyAP323rg2FMIdSEwhJlyJ9jcVKVtdF5jHk
QZ3JmO6lbEohYsntAssqKY8rcQMsH3HFpXBD7KEG/8EROoTxSIMeEeVhdkgHw3Zu27Q/rCFleAWG
och2oSqj2hdVTLcCiTBJyMukmGH4BXl5PALV7Etoll14Un0Y34FoyuKRfw2yPxsDUY55uEUcrIxX
ATxb3yrWBtt7eBnWSTW4AM5z3HezwTPAbehgMTMBy3KEBjNotjtKCrrRoBMgQByXpeBBr5evZ57b
C/Tos1t4rPDOmpzfQZ8RnZJQMpgx/JHem8yBCppF3r2kUM3NmT1UO96JDp5ouuP6tygMeWlhyU38
07KIrkVcVD9kmKnqm8dfxR08cfowQf/peuQPTd2ZxCZSIOPvAbnQZoJn9+VNscHnUH9Eqvlvt/Bq
0RmircjsvcRCkwY1cWnbuQWSkqJ1MF3jqKLJDMkFxTiqpJ+7yzDNOo5+kfoIjzVX11oncCd5DZja
efpMyE7Ws2/n1ZNMD8L+7rhu1proAbVkAgIcvxAd05ocqIRPbOA76As4IG2761JS5cBBHnTavJMs
XfJJNE3HnnK5bUtUtLgjeA68WdY7xA0CYHgxQ+CDgEcHuJ21FGvEcEgw2LoPZJmBKRtM17gDpzwW
HyAWv3GKDOBg3NUD/nfX0/fOjZT94zjMl5g0l+cD0Xhch69EIX/6oyeU5jQFO6gJNpNGfbpr+Lu9
QjXX18FK8KnczkkrxggIe5epGFyidh7fMnzDe80KrR4CJzapFEI4ve09WzXLtcwvwlTCLGIjHjgE
ECSlZ8Zr4KN+wLeG7JjxSVhuii5SD0n7ypRRnsfYijpl8l8VQDu6mcqvIAtkSU/ILvy/or/d9T9p
Lr2M3cGyRwpjXeyo8f2KnB77kC2Hzrejb7IDb3oVd2vIWoDydBahQIrYhSfGluChfHg+rA55ddtO
CYCSg5mE57O0RIDwgvKdBc/YWwN0oCO+tQ6Jl6fxMfP4le0HtUOZR4isBjng3KiQ5NUtZ3XI9hot
2xQO6cthwZFom8J4TfwloINl+NPdK/2Ec24vJAPUkptklvlncU/AVF9P3pczh8Y9P+pSicwMJskz
n0kgZMnKamCGv3EHrDoRvzXfzT54m6F1G+A1c9EHUg6Z7gEKKzPP83JcydSHTnISfa60+PdbCRgK
f9klNi/0MKohHtFgXOJItfE+wSBav1drRbDzmw/12dx0fpnBoC5RPE1TrzpAm+PnbIxqOGzmYrnR
PkMHI4Cfg0+CoxaULOfz1JCF4hxkcHd9kyXiFLAZ/15UnaTdeya7g/ZUckBhGm6vs/odvdOIgQKZ
Z6bQYywFF/CkJgtF7zGHI1gYI3qzADDsGyZ7JbxH5K8dNJmxbKmFpbXpi8wuyyDlZELb2/tkuxLR
Qsb7kEcQrWc+nJijWbn2hNJh4Jw8CQ9jz2loaJ45zxahw9J2OPqaHNnEvHrdw914FP4utr5G1CQG
vgnmH67o+bfinpu5lgp5xFSdb+RaUb7CTRWMVnXuexY/GibmtUDrzSODhyrJ/vXKBSxEFXCf0EdC
4wMS0+ba/kBSQjpLNpXk9Dqu1sFuY+IIwzXEzoX1kosnnq2s+sUQvOzDWyLgcZOyxKdoJy7CEu1U
PP00icqdQA+lAdP7V8V7HUobjbKJmHfit/WrS+Kik1XAjeKAHpPoEeGFqKMPMQmYEgGlkIlxCTeu
PhhhxcEkzkGPLwwoqbz44fZucdkGXqVasHkRII1jrAlDrAd1KKBX1HUYrkDEV4H5auHLhYdRJRnS
mWT4iisVmlhUIQEWpTl/zlGhaz4wW+4aOY5rQXV6LRSNqZcmV2Owx4wUyQS/lsnv9mUtwnQygnZs
gVYPT2+wXWAwFwbRnf4B088CrwGwZhRq7zCWdNdsR75oHg0SSuUaR+G1zr5J58lC7Au6ROpX40NV
CnZQsikdM09Os/JKnZvWOqO/3loNdQv2n7UzgwhcCpvB+yCJ6PhWqdvvoVgIXfRK+fKaZfuOt/O2
++fZMdJufypge+69r1mvEIOjyI47mIER+wJYasXi8M2NwtmmGLFGAxDqiqCyFPSnkr856BlLvwsy
21Nu4TQOjGThaSwcujOHKfBHeFroiLHl9KV4cRHn+E+1u0e6is/ITvjCPwA/ONykxgV23zDnLpPA
z9lXx+c0hQ6/HUQMiGl9TsJQzNKEJ9OZyyUyHorIvVgHBM1lGFaST0IimDoox7xgp6GwOzD7+V4O
scgKyvuulnMr/qKikWN3m8xE+rxVQ/LjUiJL4bJ/ZIcj4iycJKg7mRorBVpV4f405NetwTVC+tSl
UJUd1I+GZ8QjpSTLY2csqPUnZc2DaJeYQKONUzhs+x+arrN3IAxO3Yo8EgQKyCPAHqGV93KUa6T5
BmljTFoy0s0aiXnDe8g0cJ80LPy5hteptKOfk0sbh36SPg4IHR4WWh0WdLeeRweeTuVLhnA0hZB4
6snyyq7QwbjeIi4WiqS4OnGkj4d2YE5z2M2JwAG3RsBPUHuNX7lAdpW9gqr6+v021S8jmBkdWj3N
fP859coVRDTQfWSMEgbQq/psnM8A5BafbCEXCDPttCfPRTUzluZe6Fd2z4iP5vJWl5TwejR5AiBL
MDkBNYwI5NO7pcNnZn2ransVpV5P8TKvtxoTwd9ZoGGHDsX1pCEBOrHKldPkx24IdfkZqIvaG41J
KNgx/q+QJw/JHUfMVMo/PSQuoqlcEQJZ2RACJrzsP73wMKU7uBgW7ysGaz+R3FZiXm5aYvioFSo7
epIfCgd+8Xf+19aysyTEA8LEM7TrcDhJ6JBjHUnmkh6x7cxDJD8ky74cTn0A6QclsXalKVAr16k6
3JWUxn1UHyaL3CR4ygySvJiAdaaqWMNuX+cvG51M019YnqfLaW6YriJ6IWLvM72o95C3dte8i58Z
i0hRunPLiYJwmKeQBg+kAT7yXs8AbeX9K1ckf7oOwDeRc1i4XQC6zMeXUarJ/XbVOzt1zKj1gnQn
s9sVuMBcjY5TSku0eDLfvpYMfmpBaveH0D6TnEzSiYj/dT22JYIZCG9fRCb0GD54756YFyJOf2B0
i53f8BCyLY4Bb0L4B6QSwoLLDP1cQwsYgadG6rT9ytRK+u7YONm0/XU37LbVPAQg3nCp0/yAun/t
Rsrj+SxQtngAvpvUNxgxlZcjUR8jk8YZD1TK5BHQtm1Yn+F5+Jb7SPSTU6PgH0o49ItcHIPWGnyf
fR9REvP99Ihm18mJYyqL4vsnMO9gqMvCBDy2znsVIVNl4oD5yaiP1LGvOJQ55H1NWa9maRLFKJWD
Mdc4n5X4whip5g919MD0DsfeCLDopOfS3aPXEuXUYQ3wXuKKMFHhbE+NtL5xeRO8yGsJp53LzGcU
sJC/fYCI5vF3yWUML+5bDqc84YuP3lLQtiLKanIN0Zp0emKKutYgSrmk4mubMSNEgoRW9/ZDvv+A
cyPu2f5vCXf5hizwltaVSfwaKac2SnVxTEldo5YMF621ZDwrLAzA/Un+NkF7mgW3hr2K7k8UIaT2
yznZBjz6blUiUHWb2nv1ysP6tzIdJVo6alzQ994J7XLI2550mXEQ8rc8ZFL2yzLGy4kKxgg9NomN
J3/ekJEoxEI2h0ylkI3AynebGukiO/0HqcC2fEXA58dRQg8L3r0dCd/btd1weQpZiIQGTA1a5K2K
AKgeKVYalNEJHlT+eyHjeeQqC9ay/dvopnRNN3EKk1hLEBuag+Hr/9wRwU5k3ZgrsMjOVy0rIKdf
Uh4Tjp1GnapX9feLXKcnZFNGIiTBHbR75iNVikENW00c4q0rBtK10Vjl1A1y9d30kjHWDjm/8vQY
7mM+JnewwvilZ6Xiz3aOoxnCqRbO+aaIj1IC/naVFZc4aS7deK1YrE+I0lBM+FeFYfNRQiN+Up7o
lWZVXsjCup96Bm7J1yDAofhshb0n+cLCwZlJLNHXq6prkAYzYFayCcARjyyhWOXhEqtT3krJ1pe7
qzvLjg3h3pdlUPifsMEJzreUrsCpta5s8f0ONuUUYtBLo8KgYZu7zkgoatazZtqe4E5iguLFWEAa
ureBFTxUCTyTkVABAf5H/HQKbxkSKsggUhG8ijmd2hcO4w9J/7UOANGbd0tRQz2prLfqjwZhq0B5
zKnj0NsqW/Vknctj/abpyXHtgzde8xL71tWDw7TliIuv8jTC/xF/toBJxTXWzqdHajgW+DoQ4K69
HJqG4uBmHLWNqGjpb81dyMY7sBju7EJEHW/2SlgEGAgH4v9D3L/xgYhSH7RH+mVPzMjK1S169F1W
sgOcfiGbMvEYSgSa/rNCKkBoGvDy7H50ymFEnFSBeNm07eG2Uznqp7GteqDfrlz/X9wccJBJ2mGH
S4IX6/XKbtTVfQkiTaCpNNIxAeX031lm7Jza5jP9Q/GlyHrWmXohyHsaOgwJjTh7Oe7TOEjwInBR
w/5N2ZPNd7mHLPCYoVwBvzMP9AHnAcTcvNoFQRdm81DulBb50XDrZOVCFCd2viM+tbg4eEmcJUs2
KhGdr2+p//GAvLDaDurzzkqNNPG7NTb8JPiYMCMw+Jfj8fBBAlkkRz7thHvP5kzvre93oKkonowH
fZwajTJl6Yre0iQmuA73BDmPHqNh4pBTQTvGexMdfzlFhbBi+MiUUNKovFNMT5TjhvNXOUQ3eTED
/BR9M7l53yVtc8Fhh8DrW2okXo23m0QFOo+ivvyllOErgQwtRwGCXVW/38MmP9dO5wO0uLJpLq1J
Uj0HPWeHgAPzT0BK9MHcoa3wZIcxwBSttc5EK9JS4QejbRDRut8ugUtaXYLCjRwN+xG2AVK+3ZiO
Iyp2lKvw0i0Tij4APf4ITQtam239AGZnPlDoTf+rDG8Bf7UabsReA25CM5a8NxmODpepu71YZpQo
cHwS3WIxW6izt3OcDoZke00B45komMgntMbdsHyZ7KOqCwk4ox+4aMU8z507I9BaNC8xLsiMKR2N
WOcR17qAuHwqWoTrDPs9LpEJYzFbevSFNFUgZ1CZsZhqZ4jo1BL2PueJPpW+DBDuBcgHgguxFjmc
zGaFJ8UZdoC1xMfvj7+eObvC2gWveeNvHFTgEKjZ651VlkLVq39iDLnfwvpUPmUQrR798bAgR6GE
+9SSSWyLoc8HNaLWSU4UvBd1c9XzYQKPi3p5C5aL3sWilz6hd2yF9E/Wshe+XkqOFUi/YidXTGaG
iiviexRL5yGFmL9GdM+cbXA19bwW+zPXH18U0Xg09taMTU7myZZpxc88Aap9Yi47lVEf1IweqpdF
p09zCtj5AOpfam4uVRREvAFSDQ31YH3K2GSSzoGE5LwG27VWzH+aQv32HiNG/U9mouZXiR8ifB4Z
BiTOFU0aXakam73jTorquPv4E5Oe8BZfiBj70RgIQvnztaPx21YAOu97UTT/1UPhPXc5Uw0PjIcD
7woZ7OybZ+/FEGq+lKmF3wnU24MGYryZyrpSMJNsTDY8obnv5PadY7U67MH6m9tf2AOy083bC9Q+
TX61QTxUhz3d5QH9dKQ6QgOe/IVLUBA39ECpn+0FhMhCrFjPvx+El3XI0JIbRSQ/o69QUr61rEU0
6k7b/bhPpQgGLyjugc/s0Slu6J3pAw1Bg0w640WZ17CNoUGpd2wZpDetcAXWdXE1QLwAtYyzUsqh
In6Lc8OnfwTHsOWZD3RBkX4HlADNgjL2IHo1bbMNAZubm2XEMwjR2HlrdsnnFn9OV2/3VH2j/H2s
yNlfos+VHYv4T52qxdbLdjNRMwfZcYWv8yoEaXtAB1E/R1r9X5uKipVpffj+P++IjWy3yyK3gm5Z
lt0wP495q/zDZVWerkI6QElyu6iHtdk2TiMdsZY6fMmTdxYoDFxV+IjTpRPyMXsAYLeTdh/WRu1e
EAy9L85X5PdybAlnyoh/HuMkFGRfFsbZUTlPX/C3oxrConlwGFLbiogZPuU1Dpz2/4mSo6OquGKc
T/uWl5qwDpBzRjbGuGvySb0jYOKbKzuWB1tsSrBIGqykYFIZ8UmzavuKEDR9Jf1M5brHsf6zc3qt
LCD/44Qh1+juc4RrqP5NMDS5vM/n4Gzh2pSajYsN4OydwIVBNebQDymchgiC7NLXDoQvrcAlegTo
fky6unaSdBZVSjOYd/hQ1D+AhoNUEcwj+kzRrwCd5XlICM9wgbN4Tx6p49Il82J233ODI7eJRrJV
hL504DoLEnGlYdtGMWBoLhcUwyYPsLaejK7f0J0+kSMk0mqgPhbPhRo/5zfrsGGIowmwCYpbPy5F
PmhBTqasKoKU2+ctt968CFyFUjslLx6w0l8PNjeCj4rTnUtSq5N6/8jPQsCcp0LTS8/CDt/5bG/9
pu/6dw59FHqqELCHDlzeSVaV9lgMCkWswqfREK+7ZL9wY3yrU1cTnT8ypKd691Jue0BgjFqpScf8
0SofkMqYxQs0EaVnF/y9Ohw+x+4PQmnbOXF11timSCZwNil4bFFVMhdpSzrmiEVb28cL0Ul0dy1p
T3y+dCO+/ZD/liZ9hVIWRz9RmkiO/XKdY8VNsFn5EMonE7cObjdbZehEFBT4P9kyCOfovxZ0AvIr
VV9PA7q25squcQgcGHqwBOcNAAC5EV/Lh8v0/ROWbXWiHTLWpOBAfn/aB9hodQsR2sfQb37bA5Zr
tlAQA6LVAbCZ2tJRZRp577GKQbBg4GlNZ1jnKkr73Z5wkiJh/hiH2IWXMgUGkIPFijWJjrvGlUxK
XfdKtf+NrUkXFpUFg5//PUQpgvMkG9XQQwNmOMbU89TDyH2BIlm46OrJfMl65N3j9WqxegtV8Qx4
nTZ+eHeXhTPfOUal4bBbTXTMSqLHrYpIWlJgko0VXAv/vf64XMdvj/61B5VNSOfR72jOq2wGIbFb
daNRUp3ZIm5keDzUcW7jDr+b3ZuGWOfVUKpRmDN+KkodpqVmIaIDFJIYaKlyDIUw2jjkJgC/j1Gu
temM+5zgngn11KP52k/nNnxhO28kz9uOxb9vr5WvsqLrrAM8cjbvK2OfKcw+cIrOKedsQ8jZw+XW
/z6CJYFZFmCu6rxsoOcWPugVxsD+nwfNqwVvPbfEs5hD8agqeOrGjbtrgTMSqS4gx33mIRI7RYfO
6gDXY6JaQN02HEg4GDT8lgcsv4FqASj0yxzMT5jkZEjJXcxY2XjL75b+X4k7PoQl5UKs/hTCDilq
niyvr7NFYBFYmaIDHAOAPRPMGQ617qNOlJhzr5vnYCgpXYQNMtbWFXuSvwm8tIQSCW3QT7hOPma0
mw2WXKkP7QlU3rs1eBwS7gX75kn2QKOLkNXgWqjFTHzl2NHBBU+IJBKScq318G8bpepaysIsAqCX
PGkcCDrsptWU45rY+2ULQhICHOjL3nlmy8lX34SdY0inf/rkOpuxDPNLic0D35gV9UVb82P4hdhM
w0Pxq4TkEN/aOmU9NwnjQFzBW0YaCkUCHCIpJaLGbKoog9+CHPcnPRRwouXr5/3MiPhtOtuw4VaX
+N+6F2WIOBFIUP9NT9K89tWalAxJIS12vp7xhVR5N+SKjc2W+PNkgw7k9LusG9GYgZ36xDV/3WfK
xoEGJ6kzT3cVQf7bCkbb6BStc0UA7o2r1a0IDUSl9igVt2smS6e8izNBVS8bCLLk3pCJ43jZ1IiA
QWMI3nvD91yOcaPCuD8/2m0XmPiqfO70jbQhkGLvlP01MrqQQBN3H7EFvcQLqqfji3scGzPt9tcn
glRTNC89qGoScgoOqbJm+rHeIqgF43ksQnYmFa23VsM1HiHQRqanoHzPki7KCTptA6emwE/dobvl
iV79tYsVZjMxT/a+dAyQxMHPWKg4iRb+5AVSeeeTmnf9wwouECd6asVUMXa3xb4IcI1KCvfzDYs7
kF386Xc2zNwNML4o3TXvNQiQ7fEmBNnF97puNVtVGKeIKT+jRJl9q0+q1f50FQmZEDUtAC7LxCK3
qS+ksv3GxQvDd2fapuYt+qyndyfNd+YfV01f00ruSgfPc38dvRTy769XgLSrR25vx9B9rVhcGKjS
z6ScW+03JhCBr4QsjaGd+OZFjHIGv3kH2hgvcfAa7i9VSr/YIe3rqcoG7iUiZdAO1bW294SSBzCN
4c2V85IvmstOm+l9FMPfZ3nl6QO9e2s0m+F7lUp6cE4WBEWJUytFJiOUUsDOhLSBG/Aov1IV6n1j
lY5furXXJax2OIon8imDuP12317RqbhjokNdcmyibIaOnyEDriPFzdTPYlFV/IrYhAt2+jNT3T7s
C66X9ttgPfE1ZYmQqDSraZzvpFUv1BlgfZcfAWqY7VPcZItwIGaFBPzX8Lcxy82i9xhdlL6VIWXZ
Daic65NVDapZ+KuZNgR7/k9+tUu81VPwHjMNbk9lYEYNjzNlXSVAH4sUoJowuTEcOMSON8XMcTcu
CnD65F1UxcI+VwulSo/T9sQovzT9bucQLlbM64ARm9S0UTadKA31raMtr1w70c7zWvX4BJNLc3cX
e0OOxvFfUrz02WjKHxseUXMnp2wPSYvagBCcTbsJ3gz75TdRAltCIMA/0kA634HyNvxrvp/axmZK
+UWjxr6N8UvA7lornBja+Fcf/nQ2icWi+b9OWSfNGJ7QhQoHdm+AqU6lNKCaI9yarZtffkw+/15S
S/5oggKp6Ltso01G9cAvnQEv5VeWZYsfLAtO8+8OVDK3Rfq+Us8VPTjngAi12ZUtBNtVzl3vz4SI
6cgP6TlzEUsk4B1NFPp524TndKQw83F0ReHF6VRFRjqk7QK/BUWdzqZmN+BjKbqtDU3B0BtDGeHf
90ZjavkBhsY6+AXmh0Kur0F5TKYNNGKEvNYxQrdeHmCeHYZxnxzlRJ1KObw80+prejBBxnm5+1T0
YWNXLriYgz8jkmAILcO0HBHH2yRsET0sx2RmB0695exzV9bu66NmE4W7QadACQdqvc2vh4UUqaC+
h/NN7pILLDAfio2YDrRIrDrFa9H8SanXtkZ0pXdTWvYYGKc4OTnsYn+W2tV/GOzxQE+THYD1EJld
BrZ5nD6Pb1jTFlLHyCYnYcDcPWV2engYvRuMI43I2JEEgQbHrRFBjgBdnySquPyE7kP+NKXMBIAP
8zw4MZMcbVpezOyDauhESn1p9ao/ScsrGv3Lgct+x3qlspO0QfXeYbRAO0LZeGqw5ythUr7OGSMY
54lUm8tNuar5qjkgVlfItI6WZsgq90c4D6NXT8cFvLF+/WWU0JjDNWYMHIBwEt8ySp2ovfGef4KP
Cl0+ZzqS2QxjVm+LI1bcKm+hNv872pMFmwJrUY0h6oo6zJLx7HlvmMLd8ssvQvM9++FxI6VFJwqG
zqfF6TYEFqsg8oUBFCjp1wn8sMR5fOve0521iD/mbyiFEMzbDKfcXfd1v6+G/hWxqv8bpdy7s72x
BMClzavhanREoGwFVWvh0htsbVZVilLxyZoOEMv+H2sfc6nJF7Wp0MFla7Qm0njuVYKT1qCk5O5P
wrsRVwc5bhzPxb0852zHIkKlorwGN8TbBlY4MnLG4A04tI13gJ2ZlU8D+grlilCH+oTp7pGxUqFj
lbcHHwDOJ68hvMYDhADfA/VLfokVMKZKb20d80VJBncYoYi/VTTiYW6ACVbwlY7ByiPfn4K2xDqP
zjXdH17m73cqR0scXWTCNDyn8UgMJSiGlhZ7Ubj04+BU+OOKmdyzaR+wKgKsY4XvXG/LceDPNwLp
SQuWj7/lhXmJLRJOZs5WEXQfzU8cWXpwa2qHLRr87xUPQYqPRRdsPm21NMUUOlW0M23F5eNz0zXm
eXO6o0lMZ1gkmPnPsApTqqBEzTC+UAYV5+ruBxWIkCEkQ7tbmzUvo9WKZCgOrQROHLHX7kIQzt9U
BVwzzxQQCUwRpIxVq8o/TAW447vTpbu3Txfzokvg8PParY1wlbNVondyBCMjjNgEGzjjeGZPMwyd
SJI7wsV9vZLj1NzKMfbItTzIg9b6g5bMvKMNdOYVWeS7PZ7Wgzhp6NOFP6B1oaHThwAYMiC/wSne
lDUjtP83FErtXLCY6Ya8aagxhZ2nG2RMBjMHPKXjMfMO4ct/IdbXW+ZyQ8OXtPeb3PeN5nor+dEL
Zwey5BKy9sOQAvyKsJKsOBYrI5H6p9MFJRIzchSBzVHV0eC/5fPhy3mg6YIZ5RiepsVpM+M8ZpHG
3xyiomGGPKBNC7QYGS91tlqe/N4xFnn4voi9znH2TaUaVAumxlDCXaHwCZrE3HgPDJuWLfa2bt8I
fiO44Nn1x3te1uKi81tUmYnsLJWoTQYwEZZWAXEX66nt2u3E9wtBH+D/bTTYYcXRhZD0PGJLgFHN
MmEeyfIUg12piftopz4pNfwnz6zwIZMVsn6CQzNT870Pi7DRfdoGqGCc9J8YYsSZdWrecaA25jIz
r8fcT87gHSNUeWdiKWZQISwQFSSl4CuNNivF7oV/UEkj1qRZw1mVG79QGvKqH2U8iCDtnzRUEcb1
YeKHYnte2F7CSZzV0l08CnDhmjFy6tk8/tBPaUrdFeOk1tZPMibi7I5/FOC6ojqJhyk/dJ7gw9EE
+WLqj4c5iaYj7+9zGfxsg35snwrRg3OuGJQrAXwq28iEjyX+ym9UzRu9EeGxeLo7/lSKjpo/o/Tg
E1m7MNWlA7qNFoHal6fpfjLOgQKxMMEvNoUUJBsZi41oz8alYFyuPjKKWSH+e2B4P1tDLHCN5PiC
K4bV+Cs8TxeYDPcVFhipAhbhdI+0laRhimLNrg1K70TDhqloVh0HUqcH8UlDfdBRvdoE3dEo2pNd
EDnv6/+lB6Jib7aNOa+57SSDOSdnyxn7xhh4JuK1EsBmdUtt+dGnolSSQ+R7G6hYAtaO32xbjKA2
yGE6gmsDFif7+QwNoHagwcSx3FEhx4oOKrnFG7XpkgWd07syoziH79MRytyYYnf0BbYdKMYU8r1D
Hedj587WgqCzYvif+gfSUyLHmtSH9ANby5KEstXATEa9ivPjxH4vP9O8cm+jNAYUZPlHfAaIP9Jx
RkQRfoQ3SepGyjl/NXUE9ebvvSuO0oeeYsJYAQ5J5nfoDdMkPgP2/wkkjE1U4G8JoSmDuJrAKJ6L
71DNtMk/NS8sDaW0m+1WfFMaUnFwiP1NzDpMk6iPzmLaHmFqCoOn6cx9hRM5XGZK3jVaxTAPinSr
pFNx89fqeeY/AhXpzXMxalgIN3DDW4kdObP1SPFryC4qYJl5UPHQx0WjFhtxY1pzTF7LunDDrSCJ
8bY7a0gswFuuSgHzZ+9WcLZ767UWb2UpdeDjhRiNsD50+ziycRe7RuWKV4A8EYeNGtqJcUaUbh0J
T8eK/Sof5pPBOfXfZV3S/CMQFsdVIpg1kZaSPeCbDlgImh2MGJOa4PDQNmfedh2n+RQruLnLgRou
wxIL9aDf56SS8EB7tuGSvgMBr7qJ6tqEZFcXDJ3hMlGsMtcck1Je86mEMjNIHAeD7aMt9sRbdfvg
ql/tyB5nEqQ6JyDRLTTBfvLJ5KmoIzVvHOgr+h8GcbEqdIuZzR+5eO+YAnwOWXBgjVYDg7T2MCLi
mc/YCjocEsMkgEwyB2zbt2OoYYBD0uVnOcK9acx9LCg/u1gQwTr2fWeEKRWEDaPb2BbRq3akb5Bv
hEadC8inGk5+7pfVWScRmgvyauEBe5Iabf4kPYBU7ddESzq+7OE3p/ZjrCBWcUpzHqDr5t9us1tS
9p8dLyCoJzWa0iVQ8cKIiuc+O7Ksv1U4l0SfkauJGusYvzrRFc1n+kD50G2nugbLXoBEeAN+SFr/
4gNiP3MFsVdvqQuY+NTfgM+DoOR/74lS1Rm0RjCuiX0Fnepg89oSkAgFFFoqiTg+cvFLT81uAqpt
g5lIWRQ5PjSvNoo1P34/aXO883OtfTjRAOBUYbphB1l0gEQ0yvVaYi2587euGVU7F4gYayKIR+Oc
qTJxmE481ljtSi+MH7l79CSu6gcxyrLOY0dKQqYRVsiSdEtB/P/SfqVPAOpJWwGIyKiJ/k/QcuJl
GC+ywIDixpqYr9hl6fZzJ5JySlOw2NO5HtWr3geN9H78begZG2z8lJ3SjXlDP3IZdiVxWff4gBTx
0j1sy9tk0E2/aZiin5L1i+6nrjMuW07AAi0+XR5UaZTIiA54wNZSp5Y8tRqVMLKdrvOApYBChv2K
dkgdWxgJTFMvzi6AaBerRwJI3IIrdj/zFllC40h444PIRGxezTxaUsi2F719Ao/EKzcdhjOzADcZ
OzDDg0S+2y94SywqcSjSYBsY6SU4zMVZR5X9MF9+NaIlV8c4FmQh9V/nEJPBET68/F+AHO8pRuqc
Cew4q6/rIjd34F63nJn1X12pMkHxjBPC6CR6rl/kZmQgCDvXWJD8oFA4sTtc4xdo1uPGj57u+CP5
tkjjse5BHbsW93coz+3/Ahk4gGUG5p7ETfXqvsdHxIeF/RrzkjkmM/M2V9s7punv4tIMDXHxeS3i
XD6ggFd7XfNtAhWMbld18rj16ndG8l/fZrFVni0e+tIuOH+gATKkeJ8FmNG/Irftb8Qyn6wslPlG
OkEjaIuiGv9HM8TcukdB4XwefSMcchIFLxf/7g1aJ972yvH5leNM3K0y+I2JIMABARfk3quPOeEt
lp0A5SayGqR+k1MCgExvgplbmUYbRYXCIRg6HoXIlb7o0oCTyBzLTiMb3MWLySZHUvpfAfIqR+x2
IQjunVMm9Pbf4novlZkaaAveiDt0N3RwepO4uCnYYoUCqov6Z0kKyDx/hPV+gAwiT12OPc9lV538
m13jD3eL7M/mr/6qCACQLilAT8kt/QTceXAGHmTTKHGfUc890inRusZMYRJpHsuJ0cCkKoviNYT9
yDXgxxKIU0SELjP7U6jUh+3tk+BPyxUdGhgYrD3J4kTzFt9sEKZbgLC021wG6S0EZJmcVVX5Zutq
mQrPiqhlui87djwSrCOUMRNkbuWgTN+jAUMTmAV9ZwX16kYiuAAXnN2oU3r5dFaQlMtUUf2zVFzi
wYs2/t21Be4A2t2klWJZSDjui4nS2TOIDPrHH2Jo6loNS14G/flW6A+5wPPCD/e7PgUH0LUR5L2l
TPCS0nFPsTycm4eVqK9xWgSEyXHI/mGK/pNj94+TWumtl3HfP4tlALwAHAwsZEwoTUaDLc0U6v0q
3y4iJj+TRkukMmZxq7HiHFdkF05CNbXC9I0A5XkbFeCkyV2hoKqwVBmHzq09ZSo4kxgF7OnsyaUf
OlEGxd9VbQqkrY8SBxWR9Y8sQ2DmXuOAy3dO3EM2zscfdxM8O8E1C7V8tTixgNlRzs1FdclpWQNR
Lo9Z7Biwm4+T7LGwBijJpTWuJll3jLGk38iaWiu22SAwUCCpwduYlwIkQzySauHaxQS9EtY2jVgw
8osUHwCtKV1ukmxcp9+7zbLuCdfCP12jGI/hASJzg87Rl2rPvMYeBzHa6N5cKP9fLRtde+ss5bQU
WDEe/EcfdZ4XvxeyLQUW2M9WbEOhRvjl+5XXlUYI7Djg+6STTPrEt2AF26t4KBg3zqc8Zjkktvxb
3DqVUhtGTa5G/QoiclVqSagydGTr8yfRzunpCHCNczEw0kP6aUC85uprx8bQl9HNzPf1mw0wy5nX
wy2PEqcOSVZPZs981XVFQr4oGh3kW+a3H4pabRzAssng3VZdu34TRjbFRRMGu2UPpqb/JIyW3yjG
3Q6+WTFpExlQuAAUGpAE1oXKXIi4nYmyJr7weoZI8tpzM2DXvsb/0Ac4SPkFtutQ6vm9GI94opyI
hg+GI0qqI0n/9D0UHP4uzRhFO2V1zWzFQXg0bDKO9fnzl+8WQALG6O72wrIcHDceBJ2ExGKw0tqY
NxELDFCkhVH7TJQk8+j5lucoZDcAaFrzGfs2uhpHRMK9H2wGFbQDGV2Fjh/F7+EgJKGMyuHv+Env
ezmCu4eZaRj5h/ok19de8JTo/UXeLsjIx6X9B1wBZeDlv62ZwXY6nWdDt9NALAop4Vogf5Ze0ZJ+
CPiSX2WWb27fdA1fOr7Dy+tQNEPnbSjb04uU5o8jMhbwWmXB/Pb85i+/AaorJLjyqrBAIb7sdPhQ
ETqBgH9hZBuf0r1sodeT0B0sE6DV3Yu/B3dGS/quJq07RqUGb2rGJX6NAWlNW5Qg3Nu6du/le0FJ
DhlUEFMV0J4eoZWwEercMfwjByLehN2zwREJziLqSsLAY2QyhyM+1v1HBapFCNEN0j51MR8Ogn9O
A9ugPaQsEfBI6mX6pLUzCI1sq8YCgNVYw73MMu9uMH8t2SSqCC3CKfrLlLdv45vREU5y9tlf7kmE
1HELyJoC5WhlCKTByPejw4JrEO38RDdN2cPZGIZkx41iqGCwY9tI37UWAlm3EjlgBDf5sj4P75Dh
OmYgadox+P2Kvj9FDqrP9HEayoozcuz3FV6p0zJfeLC+YA6Sh0JPLc1qyMrYDl4Mzwpw2bduEzpS
psb8wi2aIlkkQllPhCXP/wEYJ6oJ5ggA3keJBCLn3qHYGPv6vMfKqXwc11OUu0OmLE7ynBoO+Uad
UvlVUornmCStRDxyvtkgQkAUQrJcsu/D/V76KtWC4D7I8J3obAj8zBXicKxk3Fmme0lnrohut91W
o6RGID6UyuMeQ2gH2HgIuY6RGEZXa2mcXK7ssZJX5n6MKme1zXakaUFI9CcJVg0Fm8YMsEgDrtkt
q7K8W1hMIMMsP8ajUwamo9EJ8hJMNekmXvg8RXHIGvQ9RC0kqjTk83kgfEFAofZGkRKs4acz1DSF
WA/kZscMl2nuisoSKcg2+N5BF1AV9G7FrRG0RU9LQyksRc6rnG/5iJCenRMoiPVtyMfzJvoacNXz
bcw+OMt8altpHXAqskuJMpdsObTT790kAQk0/jbF8DDxtElqZapX6HmYyMjKpXnf6Uwr5hz1jXBm
STDP339krkWj86lMPToYs6y/5aiRtq0rjLk914KGlPkMrF58lwSwFvL8CLV9XMU2BPkIomt8D673
G9OQqwNvCarGWEplJN2Q/qUrB7lEQ1tqSM7elucrT3aFkDLjd0NiZs6tR6vnKrF0VKxJzbouopuv
K5pSNcct6V6mDQt3XT6BjmeYQRF75ughQoOY6rTRDFiKQbpHWKTRpXaLphxjAMQWc06s37waOAvA
DRTjqOPsJ4ySK1/6xYiMc+QF9uyYlA5zox/2IRqvMFMzYi9ldSTHNdn52MgDr6/c80o9wybQurPU
ipODtLHp7HKr3suacFJI1EVvoq7Xp0o9qF/npzc3PxykR32dH4SGhoHpLU4+sELzHIwBVg5ESZTD
kxm3E7FEioRhI3yFqwyCFy3S6S0zpfhs1vlR4v6Dewjize7M9aFUl6XGx0aR4wZYtox4Vrh0blEg
yM4LbHpVnfAMFS7aXKO1Y9SHVbCk3+Ds/fE2Jdydih8pLCvAbzpA1HuA/TqVRnV2A2XaCFYQ0zsQ
Y/Q3qi9le5ifQTBqb3EyFI8k60IDnaSyfEKecbjlDgujb6HMtC35Y3Teq9yzK5GbJEfdojC6zv/H
AO+oA7npN0oTOcD12uyQqYHK5ujPtOGwD6e7zWi1vPgggxz0CUhTzODI4K258qGVrlCX+xpbwGTh
QSiFXJSA2vyH8tdipEeh2JeewHFQgbnmQPwxJc9wJjBdZWRfCuRdzKlQo9q2a/cchlHXdkK1lXgs
zEnnZ1ydwtOE9BIly4O8FA4ebmX/Urk1jBFMk1I/WRZxY7sGcPazpDiCeGRB7RTRccmGQ3L8Cz4g
5RP/UfxA8BnLf47hyXOb0bVkPinB+2P9vTJo8GowFm/vNE+H6vvTT1ROyt8Z5UDPYe7wpj+hzXlF
T0qfJNlSSwdl8NfeEFoKfJNYJU5tdcvRi15Lg8X7Xr6EdEEi6158PP5ycgmbm738Tt8RNDJZJu2r
zjlt2yGhYYOl0bIz62JztLNQbiy+2T48GS6pBLfQ/q8Rk3v1LSKrp36fbLQ95szIupkeskL8hfNv
28akhfZn8+qwuG8v/C6GmLePhBEDsAWhYEKCJpNnOozngLoUY8CelkHE+3etMuRIODncQEPBV7OI
NJpasjfAeJ22UHuwuP93xdDy9HciOeGNkr92JzgOcIR3RZHSxGCyKt1w93DngFQ1+ZgjZvOD5tHj
hFbStXVAoXnTztFmTSy74wCRLMurrVzDy/0N+HDD8UabsYlsA4deBwC63WFbs3Jusf1FMpcgVrS/
Vye8pr3IvvHq+3tP2ieuboT9GCfr64TreMzOaLAISRAc6HE/ErXLjND/3K8BwM8SA1mTquzzXdFU
Gsqjs0SbJr4FikdyJ1cVGNpz4vgIEoBkTs1Zh62VXe4Bnd4BefFddyU9ox795Q640TAL0XLgtOIe
rF2m7Q8rwwoHgULiuBV7QG/J4wPxQO/H+s6CD369SGvvcV5nxCjMMpOtwyabKrUbAmButEpeP/0f
Wk2I5YLoydy+AGHjUfaswum5psFxsdPYdCbrLEd1NXkOpSIlt07A71t5df7mP3dIT0G5Ygn0uw3O
Pfm1pxeDnpYIsp0od3Iu49hcH4F+E7HSbaopbxxPd0MOMBUrmKiKZYI67k9yAnbg2Rr4DvDHSx0j
EJeammcZY6uZG2GOzC8YpxhWKZSOUJvJ71UHdntKdfFqX+tcooOW7mjRjqAr4neWFIVqMDNrPGV/
++x1JklOXtjWEtoOa2NjgNtmnnivahB+csJt8fSStD5jbYkLVYdOOQa7P1Y/kZo8ii/Xf0nOfuOt
KP1Lb5afrRaDl5aZKy7KDNt0k1FArch3GNqDVotVraAV1m8KseJm3R+TR+winU9kMAfJQVYh8TbX
D+csNns4jtzBN9kE4zo/4aJGXhAbE0ac/Lk7NBHpEAH5DB8e2g2iAvpcf6Jy7bJbfnpkHyHHfkZz
oZL+XUGRpWGlu8t2h88YH2ecxtgdLb7T5XezOuv+3skWks+lXX/gdriWpkez+2chWmLNH2iRsDKu
1f+6LMLJuKJEIq2tCSd9SBGmpabX+OFjoy+djVtTM702aim5Ml1RJdl0GQP3aUupN/ky573zR8At
Sbl7GTSb4hzkDXxKehQ9cKIGoeXdS/yi5YPEMjKEb6P+wTR6JW5L6MsJuk7BzjJH381buKXAmhmF
vtvjsyiSr2sMghIpG4vJOyZdftmPhAxPIMAbeOrIjRnV5biCJio0Iaq5tuSCh+GB4FKwtg0N05xD
joma7554WgvxyJTcPzlAqqqeRS47TBuerqTznisj+sGxgzyIxZkQEWA1brY24guvxuAStrngPm8k
f2DcZmpE+hNqIXKnXk7bMAf3PJJ4/5ySXwT4vkVbeYwpdyYYY7OU8+lJ3iPb+GWgZAT1aQTYmTpo
afDy76E9hMjN2F6ro5AjyRnTdnEzgAehx+kKWFgvY/iaFwHAs8Emu9TkcagRxQTBpTh4NZuD/NLE
OwU+padcORGJ+99znA9udDB+IDjXGA6EOMzRrOoP6HiyQPhJSoMyNKm1IHB7oofjVhVXDrMozKEB
Zlzh6GwY6xpHxjk5DC0C56DAE9Nhs0mIns4DC7EFz7ptu/7SqCx744KwYjCf7J2F8A2gAWGg+RAL
ADIaoiIVq51hhFWYd8NnH9nlXBOkRbabyrgpYte0LeMbPIqntVutbuN3YFOzeYPxsr2McSqIqpLJ
Jathx+1xmT+60osFL9d7S0gef5XVSJtkiC8hBLZOWUfIUYwyKupyvIDt3Yrc/gRIkyeq0AkrHk6q
RDgYx4o/EiZzi+zn6m/pVo1e+o1eAkUxZTquf3j8yVJdbEzE/HVXpe4vGhct+nGBi30+i3CrwhVe
fDoWPwmkZza+DggrZ7oMMF2QzS+VKEWnoVeLjIFY2FaxJeHRpTw0gh1L68hzsV+ic01UsemdnFmo
Hr/pWM4KP69xy122i/g6JFpKWmSZInuLmwoVJbG43OyvsG6akcKIw96NpWjxk0agfVwIad7PP91j
99mB0MVZQZHJStTBP7h0eW0uapFTcVVcv5NcAgNLEiAaPJWfc9/m0J/uV+PBZLXsjJNfHm7ab1BS
BX0cXaiPZ85shbz/xBGG7TkNsOf18X6L0seUYZFwIK/oicI3B/RXdSUErJNEP6Ddp8s8Ca8yYGcz
3mJ+nclwb4B3b35st5HUkfwkWWyxHfzWLAI7siUgx1e4x1LnWj2PIpTf9EVQiAmXAXY4aP7HDiKB
LC/0cXV55TcmIuiwU/TiPdPMIO9MY0r5S3xiW1tN4ma/9bgFuOvUKHp4bdnmpgRIoIWUnVNKY+cF
rmTK4DKOIa8h4A4teW2RWf+5hHXmraL5nOCSkocxPCCU+H3ImAiAgn1e9C9+77m8tjBlOZZ6lFfn
2Lng61QApkDlVMiXTH9D+y1zMKB4mvIEceeVVQ1rQc4IKhwraWgrEbplGrUgj6yhmYOX8oXVS1Yw
WznHKwPrCOI3ZAlqyRRyEVSV5P2OIFuulHOP2FhwHxpV1cPfgFoCeTgtfIzU1CtWdMeqKMfLXHqj
ytoWid21LcwsRwiy00utTab/0BSn/mNk4iQ13AJsX9SyOvs2YB8HAvjZFk0ZOOf3Hu6v+hR8n+D+
dw6zJCPqEXIeraqUsH3AzW/QCjLXJBL3zqswRXPvNRau2O33vGXakmp3XlD5G3A4Cw3+w0YYe2K7
7aSp348wT0bGm6H1qsaBvN+hmqWccie2Bwu1dtvKS606+aOFCCiGVpnCRmGHQKt8ju4zY/9J50kT
+kJxk4PeDncTAb39USCOjgIl6IfdDm0OlP993a40C0udPQVd5MrloBM4WYWpKNdO7egqVPIqZ3Q1
mjeu+zlRTkEJWX40Xvk+s1RYXMm7EQd+aOETfV2vKohvmH1NVDPB4/Jq+eRAModstwtRlEzhYF23
1f/mIt8z/tVhgqEna1A5QL1E1gZI84a0gVahrAF+6EpIxLK4gXtqmaz7+BmXpoSE0+rSZ/zbxNJD
+VnV/gdNYmVSZcgEkt67qV46LaqpugGS2bA51oki4BpZ18huRffu5QdttYcvug2SmkLMk6ppJXZj
azDbN07tNgxeJMXr6dCohbK/w+w8Nt6r0KRLMH+x6bKhxNAzk421FExOX5RnGzWdhq1tJV91D6wW
mqEs5JolgHBayP+CavVXWrYCwRTqN3vvKgc4seirySdhfB0W4NgSD5AvgexrjUq9qpDw0k1MHfZz
5sGNT2jcSLJE1+ciMRrG0xXCENMbRTaZamzj7A3sg+Mi3Qxi9vUFo7fSllYg4inQE3BQ6NgbJXb/
2FNlbz7B9LmKEf4mQ6+ptfkpkJ+4F0w/M9zbUzJxkklmE8RBDgtkFI4k3GvnxvXtydr+4rRkj9b8
Z43yFcZE0nsQA20j/GNOQ2oeOOUoGudK/OjinQLfBmhHUfTbQwW4VQQHfwEvyKjCHmBw/5AgF4UG
9C0A9bmmZfPMYK0/L2A+df+uJyIISe0ZpWSc2geTqY2Yevf7M+Rv5/dUTt17Kt6l8v7kx5qeVAVL
mslHJNbo+4rPIAGnR3DMVWt+cOiqfnfzJU4u3Cgvuz1agyBK3CuA4pLVAEEaurGv8wRPNlJJ3np5
UsfbJ+KZFdf+Y8hX2MC1MjfmIIxnu/mWnw6l448m3Qe/BP8wZPg5Qoy/JMzq3zI86isb4iyIom83
BP0jaxZiBUy1b+guoxEIvpZWkzqDxHZt2Nm7tSydrFpPSOC05TazQE1oUagAJBcsajSmY8PwropT
dAWmjLV2EN8Y9T4ll8uQBb4Kwi+q7s1eWG5CfdJae1GewLJ2WPgXVLeQ/RB5GPEOGBpkt9om0E1E
4tQQ8rsHCua9ebfkNOS65rUQAjQWekfxKsLJ7k76QTLx3VqjrDzH4Q3NSDrcRzv8tUCWXTAoDe2K
pC2qpDeF1p2NhyPXZfbZAuVNoTpYCNCqqZXmqnd1rwVFRQbCLB0dbbr/xA1tpg5/hGUEeuEpiRi2
Psip6p82gPThMGDEYULh7RRqwv10ZfrBUf0NgY5RB6fa4FYLLWKSSr3Vvyfcwrz3PxVNTMbtzBo2
HkeL13PX7ZynivVUhhxjG1iZpSSKBE7jIHGsext6kBpJsr0NqgtiMKBOf4yhnF21u4XQQNBnRSvH
vU035EiCeWTAnL4i35QAbyqDDWdZe8NimKEpozk+4Gg11axQEs+Kk1FJjLVlJWn3/NM6aUZHHOPw
60GsLBjxo9b8mlD+E7d4dVF8LS6H3XZ/lLDV56jgyI0lkruVU1tYoPEoMjRA2ngmtcwrInUrTWOc
AXSLwJGMD5blTbXotkyzUr0TBNpNmwR972vu2/SZsKkHZPrxgseCqrJLA3noczoufp5t2vMNNXKZ
xebS8T3gZHpN2Yyqh93SJqtXOqMsejoG8EjczkVpPHtQ8DQreiypoRSEZqPcQYBJYlo1eFyny5/b
vKn2WcNjtRvlETSkEnd5Z++cph9JXz38o8ruQm68492psEzEOsJLNAPzz085EH6o+0T+qi+CQWDf
qbrOPOWjzFECG0KYvjGzGXYemXgZnL6ZaGqI8wzXNP2JnP70Y8qK2HG/+cOxIPNdL6QBtHNBf/Lb
9FYVVmNZKVoTcoXmw4A6W4X01sR5oqxuupDK0T579pXJwGEpe0Jgen1EsIe0WpIKndsyNCVaU1rL
dOthmntoWwIUQ6Yf0O/CGyGebyO/SzqtI1d37cybPE8hNyLWOoKFtzkLWRx/qpEcUaih1jujCV0s
PfPlN0PLzS9kuiOD9459xcqUZkzGlGOwt53yUTJzInAGmdfdTvTisxiFh6kZ9AjNPJuAqzokiZaw
nwd0rrd+cHvgUY/o+rSUfau+6vJ479trXa/XvA+wAvV/XNebMjzCP8+LnsnRuq6f1WGUgV7W51oD
NyikuEZd55YSGOWHBGMq6UNnoRGdYMEtKw2ko0Xnj7S7BgkZoBkfkBpdTZcYSknSYcWV7egcyMeN
39xHHqiIGiSFJXtemVl7NNmYilXsBr9XxJO+UpnsrGcIeYxh2n/dFy+FmwQ0h4y/R78JSVh10MYa
15Y0pcdVFetcTKR7MF5RYShdKMbWb15bxCIsiEkkRW7YDrCPSgBQoeLnCWB0m85F83m6kJtow2nq
LeZZ8ydvt8djThSUU+MVALZXSfy178tDirP/2IXFj6GoUFRulAdBeZHmM/X4E+YKpPquun5o7Wt8
ye3bePHWQc/TK9PtJErQ6jvHRL7sDOCXz9J+T8i8UzfOwIzusWfYF1/WkNU4f80AZyqgzRFlwmjQ
TiG4MHtJ8753p+E21t6yEnUE2HjtlphKTfOQac92f9F2OiYlUb+aPovm2DQUHxMREEWMVcM4cY+G
+RkcS0b7NOB58ltA4ZxtXwH8ouVzzXNbhbcBUa+rylNDk29GE8LwmPiGpqUtY7Qt3ft11eSvKkBG
nGgho+LeWHaxx6YfPUwXHTPDma8lmLv+TEro2f6R0SPSd/wHcZqLd5ZY9agzZMGJlpJ5by7Yjp60
dZJVQqQsndVrvxx+ZnyMB3I9FxSr1RBr/0eSZlB9Qzm5qsNhIwrejlo9Sz+GA9cfL46+smoGb15Z
UnwceSNv4FGh90H2Ovpt9KyEBT6zlA7dexdn01Xb1X8hR6opIpa1NCrbyoyp9T+AtJtQHZU2ju6V
W/tEt8nYINqusREayLZa5rcUl+JGXFpIkfF6FbuJwEpVSeQjRbqFdFzmu0vT3kTMzPTEVho4AMvs
iwKzDWC6m4q5aKj6JQzcBydSFZzrFR+NM0lU9iIqDv1R/1s+dXF/yDzdVKNcXlkoybMT/gZdv4cG
isT9VteT5jzGqzqTvTNQDlwCR4ph0Rfc/fj5WawImDvO6yvo843/pib6KZDDhvxEq1vL70ZtDI7l
EE0KSbv83OtD7DtGXIJy8D6gLYz7ln51mrGK+T5ocFq6audLPQ/NVTFJNzFavFp2I5mJiYa9W7Au
wWL5oLj0IsJxdCgRKJXRDmfjNnfIfD+fqx3hJ0r0xo2ol6JT7GDcxP6kHGmDJVxOVRVWIedy6G/y
Xv2SaJf4yaRcmFT9amk+29MvDdgo0zPB1lrlNK94RLkTXf6SXbIsFBmMC6M+11AG3y0mCLYi/cts
Mk3qOtMsg4wBS+CSN1KCHHW4ihkDgxYjfBqtTHhNFaQlXYbKFcYbt3XmIkUa53F2dnpLaL2Tr1ZJ
X5IfC//O2eZsZ6uW9HLnjxIGwJUMoUauRP+JaknznbCBnN/44hSas+OeGPo81DzBENE2adMGjA17
rRrP0VUisXsC8WEqbDLamIfexNYjXiZIoVkgTmWbBSsXO3ImyUTaJituHd7OLd4FnLaW+DWU1KDu
77QXUel1Yspc6r73HyRKreYweLjsqSv11TC7iLrpm9A+XquSV2Cc/0ORH6gf+BdV6zZLiXvWcz+y
iAVtYdswD8zF7thzT7IzeO2YRPLpdWr0k9Mg5c0gXnRY25FbODUzlek9rcgeXiatPtw/8yQIqYWG
USi5HwFzDvxOqhdkCuZ7AdqJGoz+kHRiZZTvsteyA/Ldm3K8ppjD5NtPpW6hYoBjr/PPu0LUn/qY
wcr53fwJTbuIbYLPYsB9yu4nb0BKpnsm9/t9rfsQML6kwob/kc9xzz9KtgTcZHolOn/EBlJh25Y4
ufNFbPxhKtX3ValHkBV0KRPXOcRgmgoULPYTB9jDjpgV5LphcVlu0LBzhBnCcuFm9gNGiZybdL0D
Ogi2DuaFmdnsQZDPqlKKIbDxb1jtXsqKc7HbLaT4/twSVQAm/kQYR1Pj+GUcbovGmMzspdSkVw6X
LcIuT649PeOog86m1UqDX+/Zp3/bqe5yTMFWn25H4aHjRoDAYGsVHQBr39WiBGciqLnlVJdSN5Yd
kxlUVF1cmQUKIvWm0YHYU6X3WZDH1xrOGsvpKYDg63j+EAEIO2TT6cJSS14Ltyb0NHpTp4VxBAOT
JZBKynDt6XrDF3znDH06WQsXZQGA+A0i6xdj7yllEZJ1r73gRRC5KDMizX7SHazBE6ryf3fp8H79
GkJaa88mdpZrnQ3cYMjpCwEgG2PkfYTfSExeM/TeRCDJEMOy40jJDesEhVbJo4/4N7FNM9Pi6CEq
TSJdAj8vlapoLMIPBF/iXxtf4XNyK1YljHMndASAVPpHIPm4B2QSbhXMqsm8HKiFQCLk5Pv3Nuot
+ZM15StoE2Yl/5570Sq9Mm6OemzjiR0HOVKYJm0zD45jITIT0I47F4P66FE6OfO4G0aaYRl69nGb
WW4jWkgyXOvayZMvtFNkH6SB6zFoVFBuNPjs4FBK3gPPAp6V6M3mB1jKVV9SlanAGe2LnvnEa4sG
v3D5oQGoML3YXTNFYmBh/+/ctyeJg8p11WZZrfaCehLLZBsooRdOPinqX8UT0cVmB6RbMmsBnf7a
G3xtLmef6t+lzGpIgZz2+BBC/SWNALF2XcIfT69VMAMVU5ktLaHGTg0HTYEUjfzVo/LXhj/UhYeQ
Tt1loJGzOIAWOpkrzqpSZyNMouLS2E6+KUW/ceyNk5OElulEOrXg4Z0vBMjxO2e8cWUaZ03DOpvP
u1CvzJvtbeUBm8pRkXbXPR46zl/O8kUI+JRgpfBiO+FgbJx5uhrrQlhrDBNGgz0nJleImfg5JroG
ZU8N1/flaNMxmflJzQCPn9Jti9QrG0F9d3mcSLIKH9hALWllqTKNFonm8LS9c2O2sc9n2WY6dU9q
XYr/6PHJA3fsf9vwjv3V0OLsqfq1HpYcw5mnqt7cOXG5JAyzLH57Ucx8V2L0m6dpG+Wf02iZsOPp
BZfmWpbH5++cR0TzZvGZzJq0n7Bnd81Yt/WGnW1gbq5ZMKc5Ssj0vrEo2uoolPo+8b+cg1Hi2zGD
l0iOwB8YIoHiiQsXlLNXHqAdo6BLn15QLCSu0i65K9qo2h+irrFpfRvLNFdsJdpTv/YKGgvZCquL
gSdttGu8Bq93RZdLzBSnQfQnUdSkz24PM6IFp6bGiPTFgCoBN/Vq+e9ZBb1OL/ZKkFRs/olbaGh8
oK3gSNzuMFIjLQgDkjWwiiHacKw7Ccy0/b+y7/OwqI9cvPHryJt6qZjmfIFHn4SM8kE72KTdjOM9
RXo3l8lS0mj9MmcVCZWcsrl9vw5sKuQwPt96Ml6RzUH+lf5xL+xMT8OJvDzNEbXHqjapssXT2cC6
Ss+XLtey0JKnbhFzt6cPR793YJ2AuDiJeZTO21+2LvnQDJ3qv1heOS/iMxwy+EF4Diig+uzKNUmM
qo5Kvfvt7MTxQbb7qw4DrETs/kN1ilZbIWwLzFUt9WxYhd3Mv4vhhJ+KgSyittUwGOB/EeBdbjLF
JB4R0qrY2JiHHVl1joGqZFDUGHS9P0Os1stWVRyr2HozVD6Bsu8npUGpYxBpF6dmZuzEbpX+EqTf
AZT6FouCY0cQ2XSmG+VGCIYFv/NUhTfVUsgvT11DXfyr9VFcdooojQPkw1TnNh+WCp3VV3EQsXFo
8hVjX6OWqHRq1OmMO25CZn+pCpXOi/bRoXMmQTzTQlsAeXP4nxARaVehOryqfCHre6tJ+GOMOXvo
SE+38uLeSKT9e69UoNVnSKoqAqgD24+wl7qFcz2gxETH9AmWvWqHBM4Wcb0ky2map13IcZ+5J/ey
F+MNLVKkTQo5vuKmRvrJ81a/oQNmv9SiqAtChfFyEBUD1a7KFSiCAGwBjq4QWLUYO+kO4TaTyfm0
YPXUF2ljkWV9hCEROKewD9szklsGxaeOHnRqZbDOpVEKBK5ndWMiAg9oR8naoWxbIeHBhfu0wF1d
SmleyIX1P7NofWs/g5OHA0wXKejwrsukYQ40dt698SZpphpEmp8rgST2i6l7vHWsWvLcUkJ8BMUR
Ol4AVPj9pziidPgFpiY6dgZmSgmlQcMpVBESjvZUG2LNtjAMUCu1KnoYkrWZ2kzQMCYtcU9Iy35t
oGXQlOToNegVx7TV35SWywlgkFS0Ud9pqgL3nR0y6Ojn+qhgJ8rp0LSeANh45rnlRAKENmqKS3J/
VuA7a/1TX9K1Or9I1Wl9CS0kF6PNx/SoFf8Xf1qc0kzbvNsXWdzlATnkYLAMz4dg/2Pon3LmxZr5
t8bKsvnkWUdUeo9koW2ahD84WePJsRInAzD7HXZj5Ns6ScdrOpuVIX1PpCas5V+g7eLo7KsCCLUK
dglOtK0Y5pIUX5p/p/oW9yjNmHFA73eGNl6F/wo34/jpUkfICyoJm2PJx+0CKGPP7COPuynzVfjA
vyovKEDkWBEEozpiavtDpzcBWSfD94iYgxMbY1V9oWObySrXVQnuxUPPNLO9U8Ni/OksBk0J/JJa
taekDWAx8OAtkNFvArAaZzNF+KVdx4r0biWABmQfaM09+Dzjt3PHNVIOJAeIw2fKCgKoqxhagjX9
kC4dKEr7Vkuq1UKR4RChL1bHoj7npFDkDaHwZLo+tXgeT1VgRVfNsBqy8TEWF2NBwpr1Sa4+B6lZ
jQWiUsJI9F1BxuQRLosKnYXEqZ/AkMnDTT6JWItVo2DjW+FfRbCsN5j3m+yNFkyNt47BlQNNftRC
LHSzBVlkMoGCVcftMKWyuzBUamHC286ytOhdr9QMpor9ViDf/xQ/Za4jubhNitoo8YtNj4uP+lew
HDMnOsCUu3RawSxuFQs+HJUN6xu2TezcPXRs/DXeEe8L1+erJPS0WPou/eI7AIe30oeq/iiGBzgu
dFiDHejvqKgehT2UZFMrTyUXocMYWs/MaM/2/XkoioOd4TVH78mUqiEUZrecel4s0lgK3imIK6IY
wGDl5NumQ9R61dhSzp+DG8UJHaf0cVyCpPZReHviVzx0WG88oMlSpgEjHuPVq/6yHB9T4BtEzVvz
fIM0q4FnmJekwZmTy+ZYtulcBz/k65CqRh1cTMIt3S8I8VpoqKM8rkC57rX5Oig3FmNxywtyC3/v
gjsiJcvBwO+WViK6PaEq8yt+nQPYjloYg2i1uWxWjlIUcguHE8O+Dt1DU9nfjqw/rCLCMpqIuncg
tA3uSPm13f0U6HuOHBi+a8B+8FZBP0tnG2k5ddQxw1wZs7AXRMO5mPLnrwhxxeyynmsLgDr0xTce
qkUPtEHZGXklJAMwHC29Y31lU53SI+/FKiD8UHIrJDTYUQBE08OdTyqzKypBOrbOJ4uwyVF0GWBw
X/lpyVkNkpQaDd3f2jNghCSVSEMnFHd+3Gu32ep74FrTHl4+3uAf6yQAAT1vCMf3uXrDaTPkMnMv
Pb4PszN56K3GA70/mgc8UFyHckYth1mxlNMKV2rJzUFP0KfsjjHyUAmUc0p4klGgoKuwOL9Sdnou
3Awr62pBkleMzifZAY7WOXCbqIIltYBg0d34ZGglo91HRuTSbkhtn5v7vlRPHScrhujCWjfUkJ3S
3aph9TV/NgQsc47se+4ghBiby+uLvq3rgUMbZzyA8AtvAwJzE0eHzOqj+YCX1a1QH8NUQSg58nu1
Sy0+49KzW25kphZw5fWtOqA01RjUjmwLmCTdd6cywx28WKRsvVRen+jC1IXNH8CWgLz0uaaajlbf
2Y0Zx1IuIgQ1jPzfZG6rctCjnzqjAJ5tP+un0wU2AgscmewWv5Y8ISELrukw8xXB1LeZdpPukMOf
hMMDqCWXXft8U+eludiT6bgFmJcE7RR8bc5sVXg/4G7VpH+PVHMtNWPBAN9xsqygl0AaMPMEtVcY
h4ND++JP2WgGvfGTpSDZ28+bW9HE1PvWwYPe3EZLSohaOGGozmhO8XR7UfwIfNCKFv5M6Bk8bDN5
5u6/UkyGd9NKEuR7Up434US+uXglZDDw4kBub6Htn8ePRz8H/iNdFyk3ZqzFzo3vhAYSP5wvl5u8
COwevdpvuV4Lm+InCynLXIvaBrfQfoN33udVnnitiQu3V5P5TjL0POGWfUOUeHT0gpCYWBhRIZJt
Q1i1B8Rml4lnLiD/5QgQ6uH9DuMQNMX57u/iik/vNzlH1DYXY4s0WP16Py88GIVXvWp6rj1aD6FH
K2o6917rf7EOc4902/6XcySdtA04vsbRnT8HMYr1ABCmV7KO7P5BuC95kK9+SyK9wEl6GaWdmYQ5
GVmuwMrkd+1GsWjVMj05r70/2/GNZ7GFN2aJdBReAMSj73fOrq3XNBBnkVPhpQE2rI8vubgS0w/q
9RjUUM7VZJoeN2xWIhm8ZuT9XVIpLH/TM6CK1b4q+O3yaAf0PbD+EoiiQ84VKLGUBBaOnBAveaMk
uRzxviQL5xpMn7XeL4RB+MTCKu7lokWKkEgz5uPpuLtpZZW4T4w6S1VhsbY+D9xlZGlkTwDjXklK
JcAWoT+0uxm8cnf0iPGr+OiSfYDrMriRGxb6f+WMnimfvI+kgBlo5Q2lgHhwcZ9nR2dkpV0z36UR
kMk1w9YB767zMEgIqWfkZ5yGWBYttluBYCS439+u9IlI56ghQdlWMSfuLzrUQeIeQ690BSewHVLx
j+1+Lw8uxeqB0sOArYotjbq2JVT+e7Mg81OL94IQcDYjefCVE9IDvt4B13Vp7baNGb4gYOWI/S+R
0E6dnDJxEoNhKarIDTqSLgjBtSG303roKGsM1Dlj2hB1GtMlMC6mM6YkdPhzNzCgL3DeEj37vV7N
PjjbE+GcI44dsxXGhgotknfOofDv8n78NCCwvmslvl03akab/Wbx/hLwC90/y6C82iztkImoTjRg
tQrIFBztSz4vkhGc1uweD7/7ffN5M7J0u8LQQoRgeaP0qRDMHwOlJqeWbFq5SMxbBzekMd/BNtLo
//BOdTN6gSa1dvNHQ9c4g6WDnjPnqFLjyyWzq29bMQBiJEqJWeZb99nhgkA+h38k2pSQGZHJn86W
a3xzo4TX/eq9A4yIM6BKMMVimG5h+wmEZJ09fY/OOecs++Icc0O8yKw5MXXRIurUpU7ZeaPwzGfh
c5AS/dCVt2GaLx16qDxv2Gf0yn1TXBu/W169kS3GzAdqgTp1/gu43HzIRrxw7/kplnxIoC3P3Lc9
bUTmNl83Ynru+f8qcCfZc4CEArXEjVup4S7JAo9r3v8djg5fTwn8PPgi3224WJtq4InrE+UALw43
74CPl+V0fTgQCAAxnXAZWf/6NC6kB6cDWHcuk+fNdbTJtAFi/bzCZTag1lMeegPGMgAcw7omP19p
//DjKHZOv3XgECxacOlPnCACaDhQxcM4+K8Ymvt6hNJ7WaOeDwhKtJfs7vkF9LFSmdEp2QQic9Gd
GElycjUL2jAVTXg4pvmKLZUk9JYxbVV/N4DLAXSxCVwnqTReA90MsH7dnGUShHWHRFrsyEyZsVTL
LUJEXQL4d+6cypC1mTubUU//nKqjtxM7MgVFme7ekuYVc6F60Q9O3q3mg7SQEpgKeHVf+MPVcpCz
Cqn3JYIOcoG8l8+Ll31lzav+SOqV82sS6PgL0PDFfSSEPjYllhy+9N13bVEhktTc+BwGy2bq5enT
dX2W6bfNLafgnQJ+8wzkOWVePosF1lCHNHmXzKBhUYueOnJQJNeuyDm/GctlmZlyxMbFzEeXxnXz
P+Lwziqt94LUEcKmVJ31IGbvZ8M3Kv1xNtvRJVHWyMWPiufDNvRahsb6BsGunORQuL+9kKxleAL9
9NyllpkGhf7jGjoYSNSBWEfxmEKd7U7v5gVZyOJ1GmJjQc5/wncXdviMN8H/JZhohLB8sr6v4LOk
nWGJEIb+d7ngWYb2pBqLO22Hskb0SYOhtM3oGOTzgZnTfBcQfyYSZ+RNvdU52Qc3DmH3Pyjc44Js
C82lYjMC/x8i9iKtyAuY4iHKqZheLO6Hz7DeaiKqxXfXszwWxm+BjFS2pDCi46hTsICTZ5AqPD85
FarHABECWNhVJyFlVKp8G4W9rLB3SOxRW1AG703Y4OsirwXqm6AjeJn9gku4Yj2+aNrisCubO7qF
Zqmd6B10J6oIKJhGpwqHQfsdBtdvTWE1qc+7OyqAMvb2DfsVv+ncoF86RNcco8KhMVAWnwFNp9Uk
Wu/JNswtoJyxrByogs0sR6uHHtWNoIgq3eCi0IPmvaQztuTXa+sCT2xJ3WbboszhdYIiUYd7i7dq
jqmCGiFq6FYdIVjvFp8sZY9fT4Ckr0N9NvmYPJBzdg7KsKbNwgnaFQcM07CQDdwulDqMRE+yoI0a
E+I/Gx/nEus4Uk6DA2QX9d52e9eQFJfrDaHGzCzrKVWPE1kRlRt2SbdYIJtexmNgX+BbsNGEGEKY
rVlCaA5IqBcNpbDWcM5n2tqOtLoMkYaDvBEiAcgfveuhqjhiEmR94WGyM4wt0W1kZuj0PVsvptwW
PGt6OPXaGg5X4cm0w2pTanhmK1qF03P/+d98FiPTHLhR8KZqclzLI3wjD7lZfyBIv+0sxsFRIXuI
eg0w7PP/dmuh1Cqm997fmO/ORhl7cVAn0jJ1p+gG575qs8WXgbemTzH0qWJxbvOJrQliAZCxPqWH
1Qau6UcbwD2p1SPn7f3fgbGBcv5E1zqb2x+e4NpabO/lRECYgkqaOINBJfioaQERZel5uKlhoGlV
j9dFcfuxF5zNQEL1ijNhRcg1cvJ0jB/pO29doQ9qLwLXIGEy5ZQ5cbBztnbUA6jLhotyIqAHS9dR
deeAQ/UPSABxZWqVIdeF46Ob1W9gwHIkfD6zuBq/rK6P06nv0aOST+QBJq/4fdX1/89a67EntH4d
cAt7DGAK797CqnszKYaLbZo889sqdw0O2rQKh7/7dJRKG2/XqG/aAl7+8PQS4iufL/hk7mmfZEhx
n5L7hNbQU39fvXtrhOzxHb+hCgcKZtT9MySCpD3tP+gqo849NIxwtWtkrfv9v4XnJLiOt/Axgl/F
2gf9CK3Cfnatvi2WU76WYBMp5A5fATMeI/kIYtktRtYy4ZOyEGFnuG0LpYMkMCFPqBFdBzQISelg
Z8AttCXBMuj3r4r/e45MKOClBUIEYs9S+OKhg+b1hydr147+qXL+CggtvXtwMqAM1KvnYgOq9uB6
u0TDr+Xv04XntjyByELcgIZpTyur8V58grJVFger6wyY+/ce53sbMm6GV9IIiY2oK045M/KAwSE8
R4rgcgfqv66tJi8KxXn9fhvSn1DLTbpZA1syvd3fYeOVLgjfDQnbseTpvConuqanIRdgv7YEqrS6
RUi7d86Da1+u4Ypznmu/NcI1MPvsl3MOA2WG6QeeeR4HURaBkrAY2QhTSG7XYkn4Qzg5RpYdu1zO
oj5RjYdwm7ecP+Ypxuxpc52C8t8VTmVEWEufW+UQPtSNj7psBx8WJBHBO4LXh6aAmiisVM4MsTxA
U6UC+yaaYN27Oiz47oc54J6AqArkBf9g1jk9aYX3mhtvYPae/CrqvZJSCpWsVn07YnTxl9o1wYS9
m2rUfcNuyefL56bLGCLbQsaoJ3P97SiAjAZ2JjLli89zrRnmprfm70jnYUU0nAamU8+FjD2qAzHu
Z1CTqbB/bxpq3SWPcKySgYGIR8LGhsg9SOY+U/9PYk5F8zOEVTotN2MvCLA1MvZEWWO4ij3c6Kzc
ePzvX30P0lw51qKjfjUUSninaAmPKNj0RSCKCgqWMTpJ6HTzDmsr1vDPMbUu2j0SKScRWxwCjZAi
BVPHLKTxvwUey+FWUtOGJewizGE3Y79Rg/yuxpa9Lt4gV1Vx9oYajhJKUwEG8H32dIt4R40OQQP9
iol4h/I3sz6Y2tOSpr5vdSuASts55mnWLnWUB1piZpl3nOQ1QCvYsvlZSA4RH8a+EW3ExYnC2NGS
GNM+ELoQEBurCynqdH1vp+3REVcmGOiOdF75Dakvzgd+0Jox41BlxwngFMU1DyyoWt5s+G4VnRfw
tm452FdfFB9dgQW0ojOnHSo2QFnbVSsIhCZI//RT8qml+posA28iV/ERhbZow02TRaODtarYP6W5
VIgocxQ36X9yQ0ogAbem/c4dOSR0d4eB7W+dXF3aT98BDtveCpPdNCvggK5nou2TYSdPZVGksEi2
XHcBC4l6iLFkoTOxbzSFjq1vtiXZHrWetOG6gWulwPaNSAeGzOMgJz3tiPRN8n82OUUKHAIIIJ1y
DC3qPkHXgWWcqzdfG52iabv1p+VE3Ypjabcj2wVoiuWPOiNJ2FbGQmYY7KrqV1vMDCmgNP5OodAO
Uo3bEcKNsg1vjQojsC3I8foPulbqJqB6WHfwQSf+mbbEvkGd1g5p3FjrGyPeqzDybkadR+I0fYmy
sc0ImEKT4vlGBHHh1IBDsfpK1+0/aU9N5MiVbbLMN3vP+j6qopFr60X9wtM1BVrXCu33zrmVKkra
als3iC4yv/HXaS//2vTSX/1FZO4Xyt6llcsd0CdyztwRQ7QQRRJv6klSqgHTslWO7643Pba7Hrk8
QUpYRwJvZBZAm4qmKBSS1/orcD6ykp9igAJmwZIureoMN8ocIYQik9VeLkIXT0O17nOq7Dv8FgcL
Hq/hqI+1BgDABz+/hFQCA+TTwil389zj5wXhvgGg6F7JQ4mRTXyTBIqMERSl3FIzcsQS/WVxeI+W
0r25ND7uyCovsekhN3HuV9F2OMW8RC/puCEk7hX3PfVEuigZm4fKkrj8+ga5cho6216q1tixZxmR
p6UjWlQpVM+izs0bu53olkrPais8NY2Dv0outHsRKFhgLkE3RM6ft4HA0+aitCXJ2rrKXolNFINp
n5bAb5znx56UC+8zarSxOSlDyq/MPTxkxx4HbkU8t3vIX029aXksRN4QEEqqbDgo4hUtT/8uTfBo
sZS5iUpvk5Ai9WUytIAiMvm3NLc5/9n5pOLNOziQtk7jriIK92Gf1J5I4UJo7rD00n5+5M89jJtP
znJAqWMX2be8sf2Ht+A/8IW0fUC9T21e7Ho1eubyqGestt6h+Smgnv/CKFh/mFc3ejoVAYlrPwap
GSNXMHMv6nhVZ6IhxCf0JIU1NToLHOc0oL8nryo26k8EoaZCyo+KQ9W2LN+kmaTPLvvrLfD/E/5g
CcDQRG7xZcEyR3oRntOfjGy8t6R9oSv9WPMSLhQlJIN7QY7senFvKJIhiON8ioSEc7cJnlQr/X+3
VdzJckCirbCA9dGNFbdJ44snHm7oE2QAENsOyl/CaNjxFU7kBsaVm1LeLLXmkWwVY1hCj5acUECj
MIH9f+bABmd075HbpZLOkmuZgEhaj1FEkkBWMDqLuOS+zJs9Mge4lJJI28yVGkZOIE5u1h1VXftZ
w/mY8/orOg0HbKs5LDL2ukT7Mgoa1d3CUUQg5ArV9eoZFyUhH4mEpBAR/mbjLKV+VAh/PfhiHZbT
ql81MwX4IHVbQUh/2+SA9BE3OjlGek5B0SvE4zcLoh+c54TawYaw/pcl5/mD7xR67K44A8je4dLC
0+3ql0Id/TqtVublhFNo6a9GfjzeK8t6I8Fpf0uOWhhyn5csMUCZ3SPzHa2vY5XHrHwAn50cqRGh
OBSj2zy0YvYyv3rYMnqaZFGZdvkEsnknNHF0xmxEzmWAzd7ndqUzq/rF4mGg0T2J7AM2pdhXPOOu
EOO/D9NbNSJiMnOUrGVpRG2f+4R2ylm++GmTGxryPiwgjvDg2SMH4Oc8SQ8JXqWyFPyNni3q0QRF
8EC4grtiXm+S5xIwFsL3FRLfVJOJ7AdZI9nqUz+LdujFS8rErRcdn3DuK9gkQlshA4PPp8SsEAL3
6k5z+93FgYIDG00YXTlpiDG/UlBaks9p+EfRIHVWqWBflDT7DL9Tk3tr4if4RZtT4cZCqT4SzHvc
QNjcoqVN5EkN/B9fL//4DuovidTGHB2H+UsaARJjH6tbnewQWEZ19b8hWPsYXw/K6OUALNPY2BZ6
xZgmowJPnbV0aaMu37y0G2UcsYDD4lbTBZ9NlXeo+0hEcMdJXZRhzRXbxQlufBOF1O3zn7RnWMe1
VeQrmDvwOK1t9i2fhnRWYQJ2lIN25xvngh1TRSVjVuRmLyZIVhpGYzLTdU2yPnQYpjOqgXs4sn7N
RqbAdkUz2r8SrZVU0/Q5XZ575+y6YfG0JQI4hdnce4q+ZDpNH7iZM/ljuMgEvcmhE9t+FgNCMJhe
NydMY9CGD9qCWJMiWh3SZnNpAd02Uvz63AuCLdsqII4XP846jE/xLPz0D4hy1lRC4ooQkgI0nBH5
cCAv+AhyGzqj1zWkY9YKEjhcIc5T2UMFBm1mqlne5zxav6Pn1twhu5eELjygs+jMETdC+jw25KLw
X7n0ajS7maHri0Hf3nmrEJFujJMsxRcvbXFlHpPUfmTsJIkEMaZpNpXiaymXw4zkVI9lWc7cfEX1
TwhWevrL8MJ/Q4Ds/FKoaeNK/FznuBYTJqJ+laI5eFsVRtIibyKdskCdyMAJWCF96mKs4+3uN4Q9
Cjj8EPmwOYDM+Xa9tJ8V1yDYu+x0ygCuYY9Wgy7PqKuMTvin707AbUM0BehS2O7HKg4ZKFQepVwI
4pK5QmCE4VepO5rl/bIbZPxI04c6kHhigUC3Kfyw2s8BGCWyVjloNngh2KUKO4Msqtt7PjC3tQyw
pu2MRi1qlDgxKS6IHmyFgNelr7qg8FEENJzhz+DLFBbFmaKMHSgDe87x1vS9eFy2KbOqyLCqLrya
t8j9viGEHBQIoBNDRm99sI37wgFUiU3tW5phF9A+KwdOwRN8zQpRNwC2UMRnKbWfBQ28TtNIhMNB
ymETcwovXoCTn+YUEtS0TLoyroxrEpbWtsSE+qfZMaaoleG1huLta4WGi0gCAdPgGV4R/PBH1wSe
LBgJPlAEtvoyntvRF/bnHufr7nEITVaGxuhab4butugFa71YM64Kuo5bqCTdiTWTrA6kygr5SEbU
BOTSqo23CCkxWlGU4wlpy3FlDDCpr5FAk3BiLsBHufr6f1evQtNrr846IM+B5SAo8uboc5jqM3jk
PChSCFVZtkXJ5pQV/tE8CjlfxQqfviWP+0xf6id0XJ0H1l+rWAZaBszGWKQDQAp4o5g903r+zrJb
SZcdnzcCjzyOcerKvbeY0Pj0giAdYwjSKaZrJNYRwtRI3g1Gqxk5bdNKicrmmRcdJa2iTiB4tCIA
ISrKGx5oSYvvdWX+U1DyZvxOcw7TJjQPJQYDpZUqejAjQvak3iJozBOYXDO2hf9TEdCZvh8ZDNNx
FBzWukbwyRelOHsI+n06uhiQ9ae9uJGwrsLJe2+uagETH0qsSQ4Abo7P3ThWdcdEzz+X1gp5Yc9k
PHLdfNMClqTmymZLcgwCg30DhvSCGvYNUaY/IFhQM8zbugInGxWVQXgUnCpcde4jMMgVCssuylqM
KOtJ2nnujhs34ddZME+ll/nMjyPv+08xlceL9HhNWBohDmwySKupdaPqMALmLJFLS3JiO6yWsZyD
xzf/VFdbZwiubMFB8iRpUFALIgUc9hRS+B0G4Suo3k0T1Lsk+Q8Q+In40shMSSeoadNaocOUkm1m
+Exj8ymnvrGyBVztcbOh+5QcOnqZfDJ9mx2FLmUrUArMGvejHlBjILCWUOQ98s0GtiOOwBXIIPl+
ZZySfi7uJaB3cGc/cxCWwj44vs0QUvZbbv9Qzm280e3sqfKZ+IBYbvWWU9bgDvE/x085Qm89kqnb
eCnT+FwmCQGnW9DFrr7FWvFk4CC3/IWuMAY3z6xmz2OqIMq8tkj8BomdJpRBVDKr8XnXL78wFx26
+O7yh3F+SOQDXkZvA24MduttLWZPp//klVbdG+4U/SiZzD2FpNg4ICp4m3THDbLs+JExFiBgIWub
BTFKfc1Dp4v9VZnog40Li9kMTzrTSSTiMYTlXSqh+nFIWop4HwphvuTSHExbyBU+EiwALdXIMESU
gf+3G3PGx1GNKPnnKJ80GbmyMu0JGhGlCRYUAZBcN/GTobOvStWzA8MAzk4idzpQ7g0OXxn74RG2
5e7tClEu32bIqpjynLt0ljY6Vf23k3m2A9yihMX511g/sFp2giisPcjdT501KTLZoPxFMktSPus3
5KHsQmm8v+0V5WWgt0nAjql/PisI82UumiEhRQfAIhB4KLusQ5UzaBQAzkUjS3/NB+E5/GR1HTDo
upGYvMzjEnOs2fphpsIvkUJzlYGXvgV/OsH8BQHiRSsMwXHAJ597/ha6RyHZjGuDwugZVdorflPS
qoWtSYUtRgErYy3F8yx9BgEjatDXs2Rmpn4srxdgWc+EaNTRaLH5i+Z3aSdk4XkKxl0jAtHCrZwt
5MF4+McQ3AHsiv8Lcvs2On0DhnaBZC1G7moo1md749qMeP1Bs4/xpVm8wWX+ZTmQzyk62+PG46uL
Xl38qk5lRn2VCEdPwIFjWhi3+4d2sugtQSwOm7/jhOTQacGhlXq9S3WOLqJOHYdPqUIrfQFlg1E3
LXEkJUbQmffAdDz1uSrFkv/Z1jLpm6VuSEPVs124jWteZrmnZ1hUCTHeU5Dj7mB6QsXreLGMqK4X
TN153GUN7qnbgOCKytVrq4UHLIGyvMrh5iPcbl91vXLaYiAxBl99xx5kiRzuYKhOqPAfYuFd1m1K
QXp1gCqDutoipgwL9AernB7l2iIkhPDuOG5GMc0JJr5OG+VReRNxwrHWuYONOt5lX5rMmoPkmr8r
l1QWrMcFXQRu8mBhMl0CInGsm49Q6geFcHm5zURiwrECOzTTiCFMJh78cAL9m6pgKyFjqvz4N0UP
KLD+I4IHE9Mx60i3oob9bSj7VLqx7zoh4SqqCpSoTpgO9Qza4UeYc+OWhFLmVvK5SUAXn+FqLcXV
uJOMzktETtyBSVivzLJwXwzH+hsqln0MYjY/oRCcfWkYxo/rtBY0Re8WWN2Oi7tPYEuwBRJjmdsq
rR5q9qJxy0+nXeW4QF70RgLuDaLV0E9HgIa0dc1oK8ef/lTw/cD/zJwgwq9NPWQNhiz8Pfuq4qOI
/fNEc3FUmo6TWzFjbue+2nX99egJAYeCMAFLhIvm52flqYTOEfahe8LQ+/AkMAf/EAuSzk1qr/Lf
yfkU9WNCXUG2dUL5NmsumhDfMz8tIRToXV0NCU5J7Nh9NQ+y4iXO3XV/bQ0+tg/DJ6Pd+SlHQ5fr
yk/drioZipuMPtOuSads5rN0MQAH8p7PDBLEwuqjSz75hgoRYyXNKuacD+JsHr4uRfCPrNnM4405
leU7UGg4VKHKZoxYUDpF8GPiFGZpB5tuF6+wKp+KsBsZebsIpTfKg2yuYr70Xto24CC9PBzQww94
25+2DjBAw9rPUP+K9C/4kmwHz+g1SH3Git6iH/scImK6k6fneiRBuxbSdooF/smrMEmigUbm62or
Pdd8UUJN00rLD2RBOQcO+mVjTtf00QnJYPECFZXPMAFJkYRuyvdYolTRBCT0TU0UDljzf7nC4pVh
BDT+Dh+hToGJs73eXKHpfX/dejSwm4qJ0uD8TeW6FNJop19YDwaOf7B5V2aVJ8YRdyowzr7WKQxK
XM1cliUUsfqd2C7ATcZiIvh4XjM+SoiNV+a7Hqm1PzZG9PuDenQ5YH5nz3hLetLLMdhar1bddDNt
7sRIIIg2+vtXFK/1RKdtQzU/GtqitT677SKWr1SM3oqmR0cx7HLob7Ni4B7ggcynx5WMhbju0pJV
F/pbw9EyNimewb6SHD3K2ONM5jLktGs45FlLYBYgmINIe6vSXuKT1GhGCwlviztc4toZt+ATrsAX
e8EJdXUWyKWJYhoIna0paq35evyd0oeSYKPmq68GxRop5FNi9w9t4cD1PfY1vpPidVjPFm+yMuF1
sxM61XerWWljljPngXyosdLiO4wNEC7mBpQZbKdvKQW9b+foehmnvqLdvR6UjAnUtoC/gTgbHFrR
Sj1pSClDl/+gtjcSvGh3aC+x+0RHTWYmGXvM03UwJcbigkO7rBbXdWhg4HNBnOebxHEvJbJ8I7u4
Rkb0axvDJNspP9gSN6BV0TAJXiIcxjsnOTX3YuR7W8TPjo0ZEBclFF+lkzOu5pROgUBcKOxoIa7z
T+4VqsU77QaKwW60WOUEb+020mQKKXfAlO88/LYyino9UCMaLWBg6Zng924wVli+lbZED1eMngV+
Iq1yd50FgWB0XFa+a+Vi9l3bKFDnWYxrBwXouTTGSaLXuHMb49CARw12GbgUIrFjZqiSd5lrgjDE
/7UeAG4VTIGQRAoLWLwBCsO/oVGO6FXbY3QRCXpTKPitPfZfPScIRN9USgonbzxt03yOj5ztqRn4
JXNJog1tcuhdARNTZY6IsWpw53YuGZ42cLp66FnDPV4c5h7II8Kbf52dGJSGavyz9lWkP58fNdKM
RZafbRiOl8eA/lWHayU37LQRd6+OhpBEJi/JB3KLeH2TFfawRMAzoU6YX2Zza0Q/Qk13BWEiIGN+
JqKfZ0ORxOpWdgIePQ+j2NOHxaz4O5qoz46TI8JYpAsYNIpcSqFmz4pJssWDQkz1Gg0lt1qkFglL
hvYrOBtngBIfLvPfhA8ewkGP7dIwNK9ZzsyXbphVebVNSlqW4oDweqtjgO+YUuvv6CLc5iq+QxYi
qNtUVcehaTsIHVbZPiM2rthxTi74ulV4wtRl7d5SryEzWxeKbdDnuALjjhhmnI4ilyrDyBj3TUmm
iaNtRIMh7PL0LV61jHUM1xtmtapspaXnTV9ABnQ4IahXxXj7k5rWjPe5IdkI5o91pb0IW0usomLd
ZFmE8P9FULPPgTt+VmmB1btBPn6iwoWQCA/Wzy+Xb0JTx0YoUlvzG/fohQvbE6JGqY2P2fRg4bt8
w6gAx+pWKWXJwZEjWGhohFNV1MVIqnFYGR2iw4Ai0ZmIESs3UutLLuv/er0Iz+4qjifEBMh3qKsS
m526OQ1nxqgPywDFTTZ6Nofr1ouYjE6SauPkI1HfnEBStsQawtK/YmS3MPajeAGayX97CGpO9hXd
Ds97vyrxRe2F8TirI7f56XqZKs77oeD0qtdlpZUsceJCkRR080jsRRmyABIqgBI+8xnJJ+Tz3D/T
6nkVUVGeSxz+4GHX5CLSWgRwIDU4mHcoKpe8KdlWCLckQzwGmfXyT2BC3RVKNMyRv9ABf3Y3QXrw
Bzgy2xdFl2hXvGKBSio+cpJBwq6nXasqm6LmfV8D3BU43+LIb76EzwPo+FE86IWdYW3xGDtEQLxp
nEJNANT7DMvT279DAWZVBNN20sKedCa99/gjGnadeg2j9Z/Wbw5rhWUcHGVc7I4ed8n473P3j5lG
wH1HrfDKIiHpXyHw2bCZ1NnL9BGRW+wqovsT1uZq8incYj2ngulX+cf9zzqBXif1VgVpGvgCnpHS
IdkAGsqt5E6hfK9cvNAlQtZIC/7WFP8mPi9Ctzi8BKaXLKUP3qo1/JZE8ZE/oL9Jm+ph6YLgVxr2
/QJQTyf01ejJ3a/uqPdmjae4U5HMrtHR+wDvE+6nfnyhme79PGf131g4A8lC37+V87bLqLUUi0O4
qEAsHdWWtSENnF/zxe28DfeVPL5xbeFGHPBoY+q4lii9P7RGSKrEZm3qPYAnDirDwE9RZJqE68L9
fqwSjJxdoSF1Tdxc53RxrnuOFE+mqsfH+kwbTftrx8hJw4AqDUqDIqgkN+KBl7aFp2NWy6vWiScK
ne8ruc5RBDCd3sxbsFBKS7SjHB+FcKcwYBEGvtBYH+QpaxgK0gc/5wmnv60WdbPXUuGbtMzskAxh
jsBquA+Sjgw1H/SYs4EuoURB747UZv0CArvKlZXIdr0bW9ilZL5Zn9kIB1H+CW0LDTXS/YBP9jDZ
qmB4OCsCAI2uzdBMYdfcMCFoLX54Y/AhgsSu08RB5ytbEWm+dU3YKhhYTanL/BzwayUmgeDSVV4C
NeSTz0P6YY+wsDlx0o5QV/9EC3PfklOQrRhpmWJ8rpbNYZqscfL0TXOYQj2f7xACQCKDc025FYVt
myqH78iE6VD1V1cQYtSTYkTTwh0b/QxGNNPN6ytJX2CNtOkzpFO5zJ9Mux4dKJenRD3QYDozWiKO
74FdBrl8COrnhZq4EYIxZXJEoCxW8f3hxqlQbG/+IdFxg7CIMyi0HU/1D1HhHKaPbzhhUcgN/0u1
/WFsPqLcQ6l01KCfESW3DnThBIvkZTU/DBs+P14MJhmSA9fw6lKesGQIc/4ZLfTOD9C0wEAKV+nz
1Jh6Cn71YPssvOQ3J5FWcq0lgdca+xnYlGNb0t+M4sZWKMlKomTRVjBt06rhVUf854IIfIWPlRGa
tJaF24NjMsQKsOz4dLKBBvJ9eJ6ebqpbb4tpGugsG9AArBv3DLWTjfNygjHvWU37PV6Pl6N5JA5R
ui43/No/XthetS+RO2nMnWPmcNOceYFa/vdb9V+Oe+PfsP3jGRo/nNRXL76IoyAZnQktsf2p8OkM
Hf6Q0IYMxZOieO5Ce7yw6INueOvThWyxkkuK8D3bp6VCx0k+ia32z50cQ4tiBngZ19waBePSATWJ
mYeemiPrPwX3h4ZhdGOFl8fWvjv9u3sLmShmLR49+RV2TIuLkKdWcg1TXxJ2ruwbzEWrXr32pYZh
6PfgCDJDwujlSC4tlnF8NTo+hE5+r8ATNRxWm42J3NNsaOtwXYY+5J59gu5mOtO9t2OFc5KNd9Zq
RQphFlwpdJGP9hig3k+hJp7A1obWTB+rr7u051+OV2RkHuzc1IQE4EhrEdklPUwxe8CnHAt5RrxL
Q+wEAkf1U90vtd08OYFz2um3q1YLcwKwkYMMLwa1Xdmha1TKpMCCFNWxlSqk72BIFqYsYVVDfC21
d5C42jimuCUtHqutvQydOBEtW68Hmjd4+Ksg9VLfpEOejW+gnjAo/VRPAH+Skw3pXOPZGJsjXuIu
DgWUqed74tALoVUDBhBN6G4eyMr4HMJw1yx0TQVgmyzXWlsO/iFf5k4c/AA0QzhhewefCeWEfUhW
LUyi94+N6o/Lq+fHUaQk6kqhKXJQDrtfcZrdqPXFjVAQ4A+0yl0urYMiC5jxYuUkO6IHEUJaPdFh
Jc58uy7cFrqD4q7Cv6694MoB5WAochcUcMp0NF1i9Vt1k88OxWZUZEjcgCDJ1bkxTgdoAiIDTTE2
zracQ8hMe8ispeRx/tZwApqBpMrySoetQbiJYF1gyj2h5BzeWnZEx/UG2jVIWgXqi4RbxevJS/HG
lNryK2Z2xRhfykeDSm+MMawgDXuOIj5TdYun4wtassSb6Ps8P/C2LwuzZj0bfof0nFvBk19QV8w8
cJYB+bwqq6/nS642+Vi12Y5g5wzoMfiepZTaHBIQ5M0dg40SXrRSWFVA+Cn+SX8r3jamKiQUhh3I
UDO4l81y6TQoqMcKoZVCddQJJuJfkJyRzn9ldeejcxeWgN27QzTI0zKisyUQW9xxG+x22QY9j8Km
5YQU0aKTaNOCUfsa+YCEeGwY1/hpXieGGePYjoU4pfY+5E7Rvu24VLAHlL7e3iNM4qY6g8t5XVj4
PbbHTvZKL3yiFMca+8Bmea5HfUNwaeQK/LkRY1GLCcz5RBKiQWFIMMW9xl7Pbz69JJFeO80buYOs
QC31P6BK6Sm4t/2RcOSLydC2bXflC8Yxr0M64oFxq7FZyaq1ycOgqJKOeEV6DLpbXz56O4hq/9ns
lC93iS8WaIZyBr8r2xuvuQHa5UdAR8xtR1XIgJJlH72PMw+qoQuSE2SGT9ubrfw+Z66Pt1fw0NBU
IqGqY82qHHYBi54KTgNMQPpc4giwr+nLVf47fVNr3bHpqBSNPkeuELbhSm/xFVaSHyYaEGfLz2ha
a/bK541gyecJ3ey6wY8RkZ2Q9+bOHbZYK5nfdjA4VyRSiYztsNlN5sQ+YYhPIq4/4tUxo1QKw+yF
Alu2kznXBliNwk4LFrmwyyphJ28oAhfJfn8q60xn3OUqvxH2K6GwDd97GECoJjzObYR6bXFFbvSZ
FjdMcHQvvxj4Ti1wmPz3nWmuY9l07FHHldiG0c0eopLRP8kgbEP3gvYpfFU5tpJuCMj2JOId1Z5f
J5k7Kaybo0+R1oHNH6vcYPoixly4ENsha0O1VOPWme0qYuGLUugTf9bF/tHB4zLqzkW+X//RttTS
MGxiIBLnOtqVe8bGCwCXBVoHKJVBvVAgheaCXyNDSKKxtfVm39wh6rgORXjRUGGzgeAbPh3eSdb0
RtnJBWi2oNRKAzhqDMQ/HTpd+i4AGKzOfowkU6OVoGKrlstx4WGxvcVu+2t57c9oyinXi0OCfsJD
Fk3qgdqX7M6FgIhrTr1aPhn6zmoE8qoPoB+eFOGoWlm8MzV8PPVsa3NWouFGnNxV9VZfRPOSPtw4
O8moAbY2bXqZgccXaJLo+IHFb7XqiW0Q8qOI8Xjzp5IJtVomDPKDtqx3XEWGflRyvtm/x+wdwUlz
uQLGgoRg6oKMpfdQu1xpw8kwuRjdV9n8dIXHk8g4lp+5ujMS+b3ldFemPTujHgF4S9t+Ebkfp9H8
3MSTdT9qtOSTOCQ6SC5/RNzgBwwmNSErvcdNO4p6INkWruxN12piGyRUhYEUJqysyOlBKCxv0sB6
R6L0v4PZAtKOyEQBPPMKXfgyoQMm+LjSf17oEGNtyBslpp9YOc3AVJL6SJSf88znkIkjhVqtdun2
HULvRXE0vCQe97m8z2b+0RJr9vXNKDlUfDW4e9zymYbyuD0mFGyPREqZGYV1APbHPRDMxvS/QNtv
Dr6VYKC75WveuubX/sij5yqOiQmbgrzCJfXs9h+oGPjreTPOHzFC16Sj2ofOnWmvsErZzkzkOCfF
NLXLSUaZWW6j0jBWCZZtUnBj1fXw078kfb8RFvV0mZw99QyItOMiQ4GXXIkad0Kk6izPMEOAVq+5
O14NzDjfifBeE4m4oVAyIqIpIMPiq74iyqTCOs/O+mwLx+B8KptHQCYKpiEEVxTE5d3LdYfrSmbL
TqhyXTYON+rnflsinOuLFJ57/2t8gkEk0O2WPzUGP3YwLjGfqhq1kshE1uIkH6UBPzNpqe4ltRiv
hY4bGRfJg+sN0BOBMpaRU9wVvtQHYhmv6IoFAdgYvsxY/r5C0n553iLP2zT+Le0YiVhIzYLKkW8s
8de73GU/CjYiOcyQz7zN1NpXxPABudh8FrZQgnXcv1VMuVEjDDRwQEV3nLnEUbIXC4p8unOfjZQQ
HHAvHON2BBW1tE/H3eSM84XJPY8LpqPGA1gsc4BBkw/187dcW/zes+3Y58pRuLtMp8FGYIgpHGZU
GzU6lxpnRRbuqeuZ/cwNWQzaBy6Bj5S56MtQBogt4EFxRk8H77TgDP0NGeZyASJi6ozgTIWjKj5e
oZCJwuYTbtXSAYFDoGhmbWssfQUTaMoY40Ibh21r4zoH0uXYHOcmbIQoWQVGCccXVRp62RFZNHf9
ShtZm/KpnGDiI3WuCLXwtMfHFg7bK0qNWj88bwWGAXKvzJybMxoPZuCAFEwep0ol8WLkWCpLhvCl
h2E4MxHfQurc2ogkKUeJ5RXeDOf1Coa+eZPaWe1/xZdZcwMyY1uUmRcdrmoD7Cdp+tDd9BQ8x8lX
/LPs4zeI3YowJQYmFYomVS8NFUZwE/5JZ6NBiIv7uR3JtE45uD3OTRwpypv8txl96v2xjB3pbH9w
nSxyGEGXXKsy4IU23KXCfxI6+/jNxaYHuFuu2XJm0jyoXigvsTes3Dd13Iudct9s/5p5Ni5ewG7V
GW87hyyUJQ9y4w48bAOKbAu+1iI73cQACBcFhyqVTh/CW+GDJrMAL6EKefu/+zJ/3rJUw+JWC0gr
88JWt2cA6fMrzjGPQ8X65+wgdsHTmpfGT1/9uXa/8B+w/pu8HCE4ovkgKMcngZ0kiRTqqYgK4R/c
zpp2Xavp9QVwJWfxbiuYkQ83FwMSmMLH8vgTm1uyCr0wJwJGP+GCTQWF3auDBlUVXyFHbI6+HIAJ
AO9EzDz7oR3662JQxEaKqWYu4uASFw3d9mH87mKSIoXMBfxiarQHYls0DD+pxcVw8w8BXMrvybeS
ZVJapVof2ymv+D5ussp+BRVH4efD3rZzvpRpsQTfINmDMqK/ci4BwoSgGOl1+0VXCf1hBbJs6iF/
w1ftALcWjH51RXxSpde24C+msjWxUlc+51YqUgEWsnZV6RSty8l1yS6tdx6ixGSa8iKwVuwmWPst
k48gdn/6KSumo+8M5n30JlsLDP9QsW2rULrojNyH82GF+lHtW6MFwfxoNUQ4ZDKKWU3O37c5WAtO
QGUG4TOug9Qa4BxdaLnk1GmCxKXrhqw4aj90ROvyL/ognMU3WKXPAKIQx8KhNOBMDWze0JVFKC1Q
TZRsZhXJ4yO4DxP5WqhCemJxf12c0Bf6oJ1bkHJv/SYgjPS351Muo5TKD3CCFTfTUtdVxbSwY61a
ZC72i0vaIEw0PJi2yKW5PRDe6X9Jb9fl4IqJhkSDY5Wf/fc7uh9sOt9m50c4KQXN7En65VgN8Tyu
rIVWQap5pgWE5py0vsBQ6e2lipEjajMT7ef/CxXKbkBkj5lZU328s2VKEujVpHaeMUnR3qlvK+zk
fcz8365PP2q4HQt2tshK52cdVre3ArVmLZ0zl8JuLGHOP76wjjhW4lc9FBJa+1h3s8nVefdfAtpI
mEJ2LV91kKy3MrH87gHxstMnmJydfXxWMDdZeDn5e0b33UVXcuFw1xzDaNOZaJ5OrMEqmjf5iCBd
v2Fs7LHUIRWnJ/oleqApUS3XdM16EBM10hDBbj5m1jigZk5aDUmU/e5GsPw0xQ0hp18v1swNBfjo
pGOngGbTYHLGBt+iIRPQhWePJhTQGWvDRjz7WNng1nArzhluHTRoff/FzIo/e+hItgMG8celYfEq
G8ErjNWN6dnP9MJOlJAKHGP76ott4fCf3aII/FKLMqZVYD1UBvbX8k1eUaeERQYUDHL+DEv3fid3
w85gxdTUfRMEyNhw8fe1uHHEid/osPg4OxgxX+lHGM1i6pH40i49mYoeDkO9ZYiCS1xFb1MecUIZ
Wc2pGg5UCJTS6vT00bZcZ2dklicYd9H1jFQO44SnlMFTtEmbP96YkHjLd5ZRPbC3xBRQ2LQlFGtL
vByIk8jMQP9eH0aU3tUEQ1ScchU169FXAi79PBI1oUb5y+RNkwfHKPelFBCUJIkgBUoM82cO1yxx
x2k4JnoYjtMPKyU6AP2lrg++cdvyMD01XHwrdnyxKyB6wSXSJERzDS07HzekAyaDDs1USODCPD3p
aM4h/Qzup4EqQoGYQZmQqpt8kZFhWxvIi6p6rwRhv34MssCKhcMEQeiHcpfLQMgjwmR/vcSN0dqY
AXyRzkoIYFbhC3OWvxhsc+gldDqaEf3kDm3RVAD8lKLLBZVkUuLz1DCioyfAtEVM8jYUm96ucoei
v/xpmnh115j97CYfs+e5mLtWp3HTXBDcB+d7M/gqQKRDXOAUm78rIYpYB2VFafc3GrpPjYOfIVVT
s6VUW4RCETHXrn5VTcu4WsRYdwJChhw5qHbOwsbUPJC7BwSuCv8lR+OLdU22/VpLZuQfRHR/5p75
D5NtxRKUjseJw5YnWrMKVFYSm5EjKYxuB9z1NYQkKQ/qp0z5Karu9U6p1LnReg/UY4i/F3PhV1WJ
wEt3H0WZa7EiqkasAMoLxcxgbPnEdbQfoDlZsvCN0mTWVewjsb+xUR0WyYy9t7wFWM0//3rX/2ID
AHuNRrUJliwKMDEsb1EJDb5INRb/HZslSP1fmj6vbpXF4+F4XAxqMFdim0HWP7+Z5LDnM+RmZ9Va
1M1DhB6h2Y0a6eqsl50Rf/+vkvCTSNeF0CiG6BBIGNFN1YqcxXvGqLLfjfCpmQMSHCFg5Dib+WNV
tWknCloIekFSEB/6c6KUziaCSUeeYI8M4KQg2mjKpCnEV1HbfVg8oSxtDOsSzC3Rhx7DPZ6XoM0d
lJmR67SfaxEPTRnPuCPSJDfVQKeLGK8wEJLz7fCStfznAeamP8kEMNalJUtO8VF2mQ9CLppxi2+y
1EZV/O6BwLtyNuxIrFmaFxkxrffvTAnZfo/nLE4QIoOY/qqXhvbp0c91XF8RvuaGS+eVDY16sSGK
ONzJMVNS7mBXWwPrQv6/AR+L3My6qcc81q2uHd8ye5jdSOPe7HouH1pvyoGgcNoGb4wXV+kS5dmI
Ki1PMfKDrA1uf4MsevoBEMdIw4d++Ta2CRdMiSE1h2ntwHHdb7A/dif9nnWAaqmoWfbSYR+8Jsfd
W16Twred5N4Vm2GxzCsq/x4mHXw2mGxL18H8XQkOjzGPdKeVMX5t9DQGYOCESjNioYp3wSZaqmQV
JQnqJUG61D7Nng0CXpum+votqonXnxWL9ipeIwoLtJ3Fqm2T6mRt5rqTJHlJKFvcZPAON+mfElbH
GSuWl+2+KkQBQkp/8+gVY6QFvgpFuwUazzLKZOAgAayTkAaDcjTs7KUEGX1PIG7fIt0f8Ii3WksZ
U/En0bgZqybeiSTTqBvpEM+KTsZgbQD8Ah3FpWZQ9HFYCjGHI/F54cRL7TVuTt71Lyzxz6ZpCKyU
nXPZpTlgRkAwagAlJdbZ8fUqtXxvE2MGhra4sF7k+7Bx7YvuZMyKusI6o5eFQgg7iAtV9QwZXXg/
auVrcuXv2XNMsGy04XYlKieyp+c73fRPG4uyJl3V2ISM6+tkNkIwpF81UqB/9c30yr9W/yD4gQNz
tU3JEAbVT+Ob6tBoTRkUYDGPDmZwo17R0xDYXFGozattpt1jqQQvFokX8KNv0iNP+ZqAkANaIDyz
6ZDayTacWcrPVu0mJCsvGoQnoR65/kBlRKNrjUh7YQ+cNF7oXspscbujzynN1Tdbm9OAwL4hs34w
Yv++pBUNCZpkfurESWDxBvfDZ85a7Mjey5s1BfeaVpFC2sdrFXy1yiDiQ1MBlz25wtmLw0i9MmGI
0RBgbbbDmDcytE/xGBop7q6tvGa4qwUO0zuhXBCwtUy0fFuQtEF0LwpUdSDVGF31TvQkYc4Iwh0E
NY8rrtjES7cC8QaOo+UPvtHyVgB5oBwA49YJvjHuor6FMM1zYLSUvoRX7wpg+yBaERRtil5t2TsS
41K9Ea1TTaiE5Rl9YMMN3X5iiWVtJSejS87Ljsln/+KlddLK31YflXk32pk072eWj0ZMUDzetI4H
BBAmrKNSCUkU4qqgvjihF306sK+K+/fQzcmiWKUBTSoa2GLmtNXtiQKvt2glDi/uHA+iCVt5YXOH
j2ercKeBHZJ85j5zKVbqhlDuBWrb32hLptGsgIkYAbCFthKTKtzxNlg9BBpI2LcuhdaZtH1XnxWo
3lM+0qeuRlO0p4Km2TG+Q8RX0GV5/zDkiIMhlGmE/s4e6GurK6X7IedMayS2kAy/zwLWw/z/t8fM
wql5LOehOes5+cCsu3+2VgobziDZqrsVuAegn0N4FU1ueKAL0X+zrmb73NxoegQo+s7ctwFFn4yz
2606p+eWYjEvKMbg63ZFyJuG7xmhOHySXp52oMpceXUqxA9OYFmhpMFkw6CRECUAxhA02I39XU0T
5TUpaYA0eqHa0yiso+9eQIVyv6nuo6o8+BLE/zvxj+BNI+30OiW4cLdjg5+M9IIqugxde/ADXs+j
DG+1PvJe6qgLuNsqD4xkII4fK20OaQoASx7Os4fuAcD2H/KZplbOTXL8jMn7bU985xGJ8vVksvYO
yNYd052RvnCnBe58ERZgEJUNskzadkdnmBqiqOiI8oD9Yu9EWrdJnOzKPwSLiRVVj7xOm8zxSF2X
zcuihmxRMJlpI70ZwkBIybk0u/W0Y4AzHuyGm7NA+e+TXCkvgaEDRzbmEtvUDhdIAQtY54KTkKUn
6y1bcyLXg6bPS1UI94PZPMFiize7alJLSQq90cMRck10Zr7GwhzQJisf460LFj4biE+DC4O5rkBZ
cZVWgXDKUTFxtJ87t6g2BCtSwbJMKyySPVKgzh+IbGO4SrjNf6QLxmFg41PFYeWQbhlddmX7ewCy
dv44i3oK2ZjZXuAYKkUSq2lt8U/Ymjy+q/83rOfK4SWgje22Azf+1m5B2PixZXY9f7XdoNo9sePY
JC7uhcrT7DdY9P7ScBl5F+dBvUSE1/Mm3INerPfSNW6cpjo3uCbOnT09k418nSkqEByP5kjEvlcR
i3fgm6d80IWXYdkWj7Qprn2jkc6gC2b6hkQuP2dOWku0US+igsI/5EmScHaEerXTxuBVzLTeZWVr
pX3VGuwI5iZNBmFCbXVuttuVxid+JP0jz5expcsMPeAXGIIboa17uJc7rpwCO8KMXLFZnkvbWuLd
OqfZEF5KPELN4XwbKDmlu/5HZApwk1q/WlC5g2CVuvluFV/xnbxZjNWnFNc9Jkrt13b0NknRKC/l
qnCb4HfmPw/pEaL+XoxKRhyJD4cT/G3kFrapOebBF6sCAT5ZdGIDDqjS3i3heixU3Jaahr9qSCIi
V6tx8v+RWAL0EjAxoYBqJIgYv4l189hsH0+ZY4clBunbbUrOAgl4IPEhzTIPyLryPQEr1I4+KanT
jdUsCHaY4wJwIFjTtt+1Ih4IsLgZTUT+u5tbCY3HCLV+FSqsLwbT3BZQhwZ3l8V64gGjxMnF5t5V
KIdmXW+j41M6syhO+wqFiaHTVYK0LHH+wx4Ufy5ykV94s6kqrxrH5kU3JS/LevW2xToN/LBkxSFO
0IxLT2DpMWVCCTad7ymOn3AYzI2oH99CAOBZ87oUkvViBX4uvJKTJmDD74BKPCBpWoWzjFutApZ7
ZDDGCZuVSecJlztikHEuiB9WHj0bWmMpoLj2BlPWWL9nHgP7OhGLQ6ACrBCm7SHNwwBnl9tN5kBo
rtO31xMO51oNrXOFsSoLI+tcE6aC1JCQmi2da8v1C9zj/8hMiZ6iAd8BD5NinFjjythRAmoXfxO0
Le1N+L+mOEtK2iyzrhS8RAxBRXqhEMV9sYfowfHLvJgQelgU2ATxCN1xqq6x3cHDzd1DWdy4dZIs
T4Qzt9ryNhQ4zBm5BHv6DSLMux+maS+DrVYqxzbvmLEzmBX6aICt/1Wgza0b9upD5SG+DsY71A74
BhKgNam1Cl8ccZGZoyMR6WKIXy/JU6/ie1Y3BdSnV47BkPRj/GcVseWl5+qPe0Gvhz1nVQ9W4zOy
rHsqU1d3rNmq7jDaFakBTpHMN3vc02htGN+EFN4hSdJNDU7c8QbWnv4GKru7wDw6iya81tQjIB4C
8B397hr6x0KFGhPi4n10WawVGibHb7FffLxiGfnpDqrMQv6R9nb0OmS8croqlSgWGAXBzI1bLiLa
kPGSBPb6EUCoJgOtZ2pSEI4D+vDrpnJY7c81qnqmwho4DvEb9/q92InCzugYKzrqRDSR0rTyYHDx
KnHIZiIYSbWnChJqUwNm7tJu3Y1k0G/kmq3PVmYP8cYVspX4az0/4y9e+/0S31M8/hIUaJv84HBW
pC3JVBEIAPtXuGuW+q78GDblLmqX+/Tv2ZRWsHj96reXv88W46r4QY6TuGQCmUuTzbxM/MiuzSMJ
yLwEs5OTLSQtLRo80zgeOS9y3CCEKbmiS/UzW9V1KcSx6CGfjAufvon66q5DL4bSqNnS77N+iPA+
lFQ/gpQSeXX/5Csx2jmcoellP6ngwG381QJqq1tS3tEZ14GR2k9c+5gRB6+t9GBqfIL1vpTwSGaH
yzE4rwAJcUkSkPJGVUxgl5Qj29fVZMhbRaAuybCsfUGHhIONvD7fmziG6bOu5mSl2DWJT8STyBxu
8ajTs01znCrg6N1scXFTOQI16J+QsqOxTCkN7WwWWkNI/nmEPb1V+3/53TVDpLB6SNSk1DbqSOCT
jrKsthH019M4EwjtXFttCRPzRpQbFCTr5MY+39vKKsTA63Fd2lU0YXKYQTXVR7pNg82IAU2r0XMe
7+hyydjVllAjTLIr8jhMEfbRqQHyUDd0P/VkrgWWrySOTkfLYaCpenaHburbtodU0zlHIfoNVm4E
yCazsK5CP4SN+ZiWZxoD9jx9LoxWRagrrWlTJ45t39U9xLI7gZitbO0bz4DzDNBlhDxZj6bNot/M
rUBh6nTKyiXAPYmB8iMuhtSnYZDrZZhVhuKhEHqcYrsTIJ93KZDXYC1LQ7np+CoqjB4xEYgLu0Rs
PWXDDo+QK7XXJLMsbbw8AyhDBZjtd5CTI2GTUjdEn7UOQBrG3VgXw2FoLGaFpo9AxuFF+04gujsE
CR8ahgiGyZ4vk/8Tyvewbpw/aXJ8/ADOCNlcVMsKyWJXs0XaPfC7muW1+tO01RVjKwAlAj8chnoX
wfKzFi95/IdQpLdXQguDYcs1VrqEnImiQELaFAe0ZBIi0ypYq0tTZPa+Kc16IbueHmWHB7/loRkI
sW3zLWE2YlAOmY3Z0fSsJhTcELyJCEz/Z2Kipe1osxXglX63MJpRAjU7GephX91X2JB4VwCukIEF
5D1BiQwTVDLzrEQ6oJSWrd4aJl0AbZ+BSd3sRCFj14hl9uB7QxmNfhxK1XKrTWjYHEKffR9+wu1C
MGQPdzc05qLGyEmJ6kkfm7+Y6KxqS1v9w3BsK7hz7/C1xwQIn2UihQjVVD6yd4jJVRW9BgYi1Pbp
gLT1V/SdWpNp5ijK9Jeb5MZZKcTX2tHhI34uuhVWDjbfhcIgQlqQKoFbQEda13UashD/Cy+mOlUI
0NowhIHt77/OBgSICKJkU70mpGLdGDbOpwEAwWZHIKsIj2z75LpokJXCiUItnOqSHufNYZfNnNYc
zQnAuyIEI89mx1zaCuTgJT65dyaoDMZ2exyiCG1Mv5SsuUihz4b1si6ojF2L0SX9PptWxbiU0/LB
y+ZIaMjkrqbqXYfSxiq78BhwRP/hLKCj7zJ4KH3sKVjxbk7fNEvAVKibNFm4Z/aFuweqfN3jdNwN
gYK2M8UUtMJNaQAVdiGL57eMCYMKeOrnCxb6dSuhdUWTEVhCCAVPyqmSbC8FZiFD3eDLiVDzzrJw
iBEsRDO8fIfQ3E62gLKe13Qfl8Px2ZUYn4CRgWwwJInSl90Bxxa0yTE7hMhIZB2IYjaSerKre4bz
7TYm4V/S8UzzTRsI7KNV3/a1oNydXbrNX1cc6N7jODbkKT50HkcROQP/LGZRS+fQvoF1jySybwjy
9GnskqQbfacmlRMFFKtIGIEVYHB2P9+aYcIfUPhoGe7lmuqGmNGGOPQfG8ddn8CpGcLLXGJmMndW
R3P6TAk0nnK8t+KdiTcqHiJFWnxjlblsxnicKhaPTwIeXNK7aY4coB+hzPaFigGOoIldY/5DY/9L
2UsUZK8SpJK9yOI3pNeyxIhaua1sXJ0LP30OgrwslL8OKjKajgXTHgMI1VjgykjDL7c+OW/vrwPa
JxW3Wl3eXsofONetqP2Q7XhYuLNY52oJHvm1M0miDdVZQIczgPNYZvEOJWwRAjlbWYdTtJy3e5fW
mOQMYyZLbxKyiS/Q03q8s1zDgDnaJoiF5pqHDyEICyTF71GfPQvPilM5kztXsCcEeo9X7dAs1yfF
Ct2mk/kSqi4b3RQEFYdvvwhcE1zrWZSBJnlDSObUU+Btes579EAjZ6//LyNFxVpkX7+gPi/quhRB
E6yY58yhlQydxJrn2rZw9ve4IZrpjPERpzPqXv1+/j3DeGuOuRmQ30oXDT5bapeASsws5vy0Vakl
dYIX+OP6bmnR6KCoOYxzwS0+zYwiLAPvy0F+nMDX9pZULAxvcCzeKxRYhlI+27wQybqb56XYzhRm
VvHYt+QR59CqizttBY6Cr1zSWyDNMElysxJB1WCl0XVYrJn9MJ0hAGpxR4mCuBq6fww+tI19tJI4
3xl2Ka3NjIePvKT+HrjzyUxOZEk4aw4QCXCOmQ39my1TiZ58fxl8TSRbeFhDawmbWxBZFB8MvES7
5QVK6fqvgTBqyJo8bLC8tEjywUWwWFq5tid02Ux1yapdh/5o1CKT99445rOLuQaxAIxcUuQpSQQo
0WirFshqja9ZHMPKnb8H4J3ebfosl3X3VtQn02LduUJurVUi+Y1vX0IcriIAsai0aHyMg6kr0aJ6
WDtYghMwK1qyIdJqP5TewoE+hb+RjXgnL6nWhVOZzrUxoNn7+Uur8GbUSjrBMW3eOFjsTvvu7XQ0
BarqQkJFAH/OlIo13keVtpMbXCqSwRW0LPT4svlUKu289dRT1eye2E3bi0wy44X24gBpugey+tTv
ifXfuaWeiIUzL0Ge/RXIYrm25oX/rBeXn6IkP/Vwe/zqM+pMGoIcZ6yAGUCQhFo/ex8gcEyFaOnP
3tgaoF5MoeTVKQEeTflECmm+ZjIcte2gWbc/WfugqgmHaMSKEt5CrIDlrvVbiJBo2wmT6PYua5/d
V0yNlfwmp1JDVCKIv7CUnrkZ3wRWPAcGvmZYMy7LuRgdMOh9TaBU8z62XIji3K4NaokXKRLV6X8g
TRBlkLIU8tFabfSHCwCgk0oC7adrGaC5aMXCVrfLW888UTa7ijXtnJyIOTYOX+R4uH+eJDgNL5Zk
vSedfh2QKPdE2O6QJS11K8KNQY0dX3IOiZU7MvFr84bM8zxpe7IkgnCDlZXJbgprzFzGax8i+XK/
SEk090cafuday0AXNIz5xPO+IIuUFWyj2DkoesBSlYHGxIKryAmT+rp2YsEk/g/51dC2QhfV595g
9kivDBgyRrPzUDB1dfXFiYobbFIGc/fwLRYbweo8j8du9YkrLJKM3yByfwULLlDSok0LTIneHKEW
fDMvlpNG6VjXMJNatFMeWhdzmL3nD2b9FXrSUhC05fOXkWmfjVTiovCC1ipJAiEGSK05L/1eew+Q
CJrVKvE69ni4CukPPGlEOcQJQnrzrVaRmKIpf5jEBStdzQk8O38y/wmllE7t+hXOTbLtfqmBGXRB
1OKRfIUvm3Yqjug9ryHCAokIl2ZGI2FYY7OSpaEXdXTf+A0/yVnnYM0eRUyOlQ00WT56oXLHZh5+
YOOaoia+3OHRVOvhi7g3+Lr1+duiaVF5Gdb7vk5Ck/AqN3X+Np+U48SDajlxUY3fYkpLp1giHr+C
UXH0nBN75JUW/uiE6wrPueSLbzqmje7FaVXLunLutnkQvmSuTmRPRBHUmV4tXwQi8yr1pFXtxs7j
K8pmByiikPBHUbDI0b5tMiz0mD7heCjq9JSesvVMMfK9mcNRCOCHxmw+Sz6Y2Afge/VH6WT7pJnS
/lWRbE/bOMRuCG6OoX9a6UJT9cZhVK2sOFCUT/qd806vMxvexgOS6rsfFNSeNjR0tc+eIjCg6Iqc
GSjxeIbg4+jJCT5z7Dngn1ZyUgICxkInQs0EL/O9NQHyz6W9orrXJz0aY5i2aH/+3qPU2t+9Jvyp
yV1cpU4RvYLacUvLWON8b2tg2A5VYB6TNeTkP2kdc2H9ZK+9uesET+0RrsYK2xIC0N6SRgXE5DTq
3U2SGuljo9cw8vyOCBRHiSl/IDenZHIFStWXssjHd+GvpQF4MiCioU5brIPgup/THorcvI2pVm6K
ydRmv77KWMLWYAaJbR69NK/LYiwd1+0ubBSG8ZqX1XiPbTdyAorF88YCntC11BSx5iIWX16atRGd
uwrqrF1oruPuPleF04BJkBfQxEPvpaMJiGODap3HHegTXGF5CaAiIR9cm4WewlXjz3EAB4st6FDX
MXrZYQnsBQWA+BlOvUxfFAiapz6tNCXYm8FklJLr2xJxUHPU/mTVu9QHV8XSMNT17v9vQkRP7fde
xWbW7pJb5NLybmNXIcf0hN5PJZx57XR8ICrj7q6ClHzD0Q3bbXZ3HMKUT/MfCZkeV6i5nFrLFwqZ
y1kFXDezXld5HkNAhiBCOzhNbrXsWMkdEWDp+AqSooLuifHRSTLEWJsb70EmXBsXeUKjyLTxzlKb
TVdoYvxQ+kt+KgtfQVEB1qf0GVuR98Ill4FXBwB/tyjQSB2deTk4HgdgbDa/JVDlr48JwbBiUhaa
YSjFOVE+BHLoN7x+xT3N5OHFEJSQyRFfHk4hZsLS2Tu0pCC5owYFQ5Zg1wAu3iX1YvsDKWQX+p7U
QKwssIMIR0Fl+dX+LPlLG6RPCuuEBH6ZCRkwe4Uf5SKBuzWjo2nbDlylYwhGHFWoEt/B4gBySI6h
s4BKX1hsb+JEZSREC4fbaDUJez4tKrtGMaN/Mhmt5uhccnMumLxVuxXMYt6VLgIwQEc31gl2fr6R
lF6nZ4LY9YSZgsMgM/pc0XpKMhnUfqTp7zHnKCA36/7m9+Cim6LWMy/F+B8mDgoav3Q1gG8mXgMO
DpVlJYbUEzdmcfbLYRzORqGJj4yQRJxJDY49Iy76zIb+RUJsk493q63vLqGc6IHT3y6OxydnjWOq
OCqayD0gwqcgNqEwS214smJMC8vSfJUymvCP3LQZjeSLGjTP104bg3JpoYi5Un2xmvzWHqe/7vMz
ytg8nd8yj580DNvPccFdY99NP8k6L2tydRqeVv5XmaL102z7cArb82ChuXlRoK++nxtWwrEo9ANq
s385ILCSxh37ghcDGXYwi483YIvLH82i+SGnhDHMuCD15Td4N+45ljfYpPZhSlgewB3jcXgQtzAc
Id8FYc7WyaXidSx/Wy3za5xQiYCtyPijksz9RFsdddTLMRLZRLxROK3TbGLxUFpzswsW/2im37rh
zldx3fgKVai1L5JClwhlKm4rn5CTkgvvyPfBRc7hseArVcok33Kp74zOG2lAZ/bzcvPb7vI86cDl
Ax+AM+RdXqBtOi7W6aJSCfdBWEZwXjhqvtky3gVB/irGzIy9eUOfPSwiCEqRgPTP9jPEJ1kXYHi3
NmwA4P/TdSY2M25wkjN9B0vTafh3f04HIF8XDsS661FJenndG119k4/KyXJrCOqkQS6p0Ya3gY7a
VPlGsBBKRl19GTCwNzl1V1gv6rSZ+5j2EyXLTQeWUa4VWnunHzOZsCPQTe2TEMcm1O4YJT4kaY26
LlchYAR2ci3VGtscGM87nPz5/40cqMuz78QMMIvdTSSTLdIuzWX/u8invdLCKAw5HLUWJmL+dkwa
z/oSjwW5lI/OuV5+Siv2rBM192DnGPqGnwquaXUVIcIbK0Q818GC/M82hOs9ELywn/53uGAIzAEy
tCriZqn+gnYkAtjp0snLq8vP+PMf6af2vfMrIfsz5ZOcKKpuq7ePlGRF2xNiCXTWpJ+YU/D1SawP
cKfLgHBSdqiOn14zv/aTEPdev7PQYTfuSir4lhSJ1JYMryfvCrbXER6xyebSSaJ7Mfwix8dhJykl
RiV8NEWw32CCLLzM27LhO8OFMPS7sgQrZJ9pyNr+B30h61ETxaYvVwGCIb3lNvugIWDwGOSs4qh/
8U+OdK2qMTerolc+MoqFKAh8E+xa9jx9x7FzfcsutxZ0tHqwMmPWF1UvVE43uM5Q3jSo22MVEV5t
o/IDTbFy4cfW/KSXmgNCmfgJwnoeTtR6Yq36pFbwzkHSKqYGy2YeoJrkAgf06OsCLAckzX1icENk
cFFEqflklcAcMIFNtrfmAJWiemakY7NbB4dLa1upsPxZJ0ZRe7UBoYvTvlp+MxJUFY7/Z9K6C/dP
UZ2hY6ZVVlDK/RFI1RKJA0Q65WBTpYPCQeAZd+nILI9C73iD4RPY/A2QGu8V8xOV+5ryHL8fOAO2
fO6AKjWsGyz4FjGlBL8roNV9NYpBr7aF574NnGh2b7A5H593ZxvCIqOfjezXCD/4z4Ro1Uf5PVrN
RvYGowyREvB+6+f2LeaelZXIot2BSZWuUoKJKPVwNxslk5LUlWJtBFFi7zTNt0QeQx+7Z3x0Jn+h
OBaP47zfD4wgLVGpkA89dtcaYwDSWfhriT/4IyxpcrEaoiMznjFJg1ZEml8UcaG2OOgsl+VThiRs
KHeuvCNgNEYP4EIuinkBJ0xFFBh3fvIFL1aJeg0ZtRjkbnvVv5/Dt04Pkf/6ePBDj1EMfCtDG2P1
dfkGmqfNWVN9oxq/LG/LfELzL0IDxRrTWagSjbw2fKIYic4/L/hTjUKNrNjibspv75wZHS5FpjYk
qYYhCRlq32t/wYgBpJA3Q6ap6eyMUnD87ZQ0fBnQLvoUudUtB+Xk0Z6HyrxtFlLIbQFD5yNrTQWP
rbo2tFGRqvq/hGwMG8TuW5ui5Y+OW7SMo92FYcby556t2V4OuzYYeg/dzC6zqwFU29HlXarG1VoH
dWsK9G7nFIpwJSKZLawvHXPT8m3vUHJusEwoP4sTXpE14G5uR7zI77VftkqNKVfktbflS8DDhjPC
8jqmLfeGGnQWr/pZiJ7ToFEAJUQHVF9FcWr8iR5HmZcEU9133paYSaFBFH3DY7qccjDlpMkH7XRE
eU8zN32oPnoVW7em7ks0NfWQg08C1Jy92BJxuAQdC7/SFkcTfIGr8du6eaevUEp1y82GZfXLz2Xp
TUj1OcXye58qAGkdYh93lQJK4AmsH3EbNoCSmu/g0UyWmYH2OcRimS6k1IfGGbv1f2OAB4H160I1
6AA/OdE/mhQvP48OLDEqklEs7YwOLyRFb4IpxXDeu0dfGW2537nkbGE2HwLInBgtznvO2mV43DJj
TaKM4HvR4M3kVlA18p0fe2uYKRQpvv9Qq3Wsq6J6ZqEBQYKwmCYGrp1b2Hcp9ShdZGpwrK+hObtJ
6C2AXesN9JLcAqu6DljTJPukhn+WcXd6f7lmSnCAlGlg4UyusB8kw0wb9lcHXf7/9YJmDTq+hBvy
mPrtHvy39SbaebI5ZjK44do47sGdnonqjnyVzQBfZuMc+mF3o/bbyIPWgKADfPzVLlB9OeznwJ6o
x5f5NNGFW/CXC8aZn1EsADw2cjCO6WjLgtDsRMl7PhGrqw22ytOKHbjOfRCvrpiBcF2H7P13pV85
nlSazBhO7N1SOZ7Ay21YjxQUzxjFH+gpB4pARu7XXFAMjwJ5MmjmTZTfaORtQZ6Xa1VnATgTwUx3
Yzepd4lYV66usV19jV9CJsT2TEzBktgh3f3LYTKghGz6nml+fwcLD8SygQr5r8mqmELSo3cOwn8c
AHuBvUP0p8sKWa7u2Xs3iPpvJk3hWDB0VVYEfFR/CJD+/hoyxvjhF9ktKGV+wMkKxAbRiDD6Gz/V
L0sxCpnGaABSwLYG3mnA7KRR9TQAwYRkYpy77tundk4G9oYTbF7DIurosz3lSFcyE6j92uCTQcOx
YSPnn4ERvN8zWbKkAr+7fDfxqtiJAcXHHHvClZKQUMWqxJLdf5oH/vzZEfwHYdsytjC32z/GGSBk
ymF4aEEuGvMm67ws4yCPkSxegGqVrxQNjQE8gl0OnZovHNBcNd4FkP/F6Wbgg6DSrwCt8F1JNmeK
/euS670imhS8VdhStMeB+KIDJjEVjQo52yovJ46Em2626//+Xhrt95u1TSJ7JtbEcUgiI0ylc5fP
UbGPa4OS8LBdmozNL+UOC8ZQoiQ5olfO0f/mirIasMhdRlvaJdAJwwgf+a3HA1JcV8yPDYkcxQSM
8pBA6g+M/qXx5yzvaBu1mtpoU3T+5R1AhczhlR3KlVwB9XT16f5djAayUKfAb/Ub4iF/sdKimZHB
USGdOcgwNaawdIpWSiFkZTOEoB3gCKidpTsxeGBaklIN6dOMAM33Ekc4C60m3pNDwcws8ffB7WNt
h8uKX3FZee6To6IxRl3She15J9gfz1yQGfOQmYf0QstzVv6jJWMyV0pzAXMV/ILURTVbkzWHsGCI
FDnix0pQOe9gijlay6e6AcZvwwhTQFTREINliM01cWJaaPTuU6y1rQcU6Xo7u1F7hP9VGvDK2BKb
+4k/weCAXxECgagtk+wHMfeR+o87LpdVj91gO7oRkerGjBarKSLI+ReG8+35DJCXG/S3UttBIPSz
h30NPDuOW32LP9luwZF2eFBqD1j50MwjeE/52nYnO6n2zQB3UX58MmFxKDyZqvyFFN0nPHz0C8Ag
WJCn2y/acRloFZY9BAQ98L9V8828xEpHqDaO3ppFGOCWSwMCUPmMF3twAi6rlQuU2DSBUZeP70Ou
WqALj9aDP3p0qUK/RLZ4pm4kiUKO4HSn90R4h6TR3PWaP/w7RaBQF8QUS7F4kRPHocRwcGMVWR5V
yrzjeDXPWAVjQvrzttEahLnnyrEckB+7ly8Cvt2vfah7+Bppw0tCPI2Xb+LvAZOumWkyHY6hC1Hn
dfetElwJKnkyr1kP8uyKhGSIpXjfNJkfChXqst/m+aK9JhNAtP1ru8m8bo9Z1R7XI+3p0LvTsueP
W1zaygzZaW3LDMrP9ROulwQoV4Ee3WX9YoYDYyO4aHItKmKoeP9TkV9M2edKGMg1ZWMwpsxPQifb
cCv6vkMfZH32wAOxmFMhz3WOtTC2+oM3xDCNgypGTEIVGHkLAHxzzf0wj0jONKsULwPhqSaDEc7d
9BxZPLrJFLPKu/0z0KcZXDo8rLnsP6/kUtoj+YjYxQHTIIG58EYsDFzjvuX7xbOfoqTSqlyeRry8
NsNMAGgXQsZvMBNpzzNd91CAISA9D+X6/wUqX2SfOPY/bZESM0e+co2tFBSg/YVUCebjoaDjUxN4
JHPaWoRmILmjIFVHmhwuQVwSpIQkukH4x0KskCFE7AsnfAadkjE3MTiBoo1vTkQfmy5o7r5FjgXR
umDGXjG/rwpTjtqw6SDkDpyiWRfOIRYBMVqidoLIpNdwReOJG4sPoObLPvrAyV8jYT8q17e5ze08
kW82yHiKuM9o7P7PO4raY3quQO9INlyIfsG3niVkWlUNBFZVsmF1qkc4lF+M+S3Eo7YFlvXg6p+n
r4j6JKuXTzk2ZKxxadyHJiee35/729hhZWwDmj51EfWkoqb7xrWBkkKg6nWLgwqw9oUZvd+lWd5Y
BXDkycsBRWOobp0sqwUkXky2nc97/I6mq2VyppmtdtClE5aqruCHwHe7f4YezL1jfYnjEimabsaT
0RelcymLbCF8v958TgZloqDY2WyLP/ShafD7yxnchEIt8ylsOCSpwSVAa9QwEBsf8tT6AVFSwhc4
b6VzROMs/ieIhuO9EaDG90Dl+3JciuARy6BDVFFqHpFibJzcCoUv5hT8A7xd3cy2V8trDNhYaf13
jihPIJRpdDgEuOujtxjr/ZsWG9vhsY/Zj6qCIEnMc6dyrcQ/rN7jWD1MbW4C+vk8zEdyQLeMKEI7
SXwm7tMFmwYgft4lkP9sZAmYwCK0TcolOGFGsO4YQbuu3RbVOWICpOZtTQenbvmcB5v4BsebIN19
CeJWqTFp+uSWisLi+HSkZk+FS5HOHS2h/tm1KMpc2HYW08eZ0hAMhjhvTyTJJwHNwKAUmX0CvgRh
FyR8SiiXjMpUhrct1gn/q6T89QtqH/10BUNvlE108Nzshw+i135/3fIWIwVtV9Ge4MwGEcq0ng9j
86Twr8cDRJH8pZ3uIQhBmD829Im4jJ9Sn677AiPaG1+fh9Pfl6YHrzK6Ew4UlSzRbIZD096LlKOK
kJUONaFOCyFCoB1mnnlDYzBL8gMX4rBXRx0ZuCVUIFdtcQFssNuI6YMcc0RLAMWqUZ263RPngCZm
4DNwIiSC2I7Sq4D8uiDfJ7EKbIKaOrJpG0YA3c1Ve4woZZIYcVNCQAu3LuKsV+GoHFwC1+HT9pnD
xpsygilI3HyZXUMJNiPMuaJWz9aXy4IwLg1YxuYRN82QiwN4QKGKUX5GTRiv1z/jBYQOBrI7XWfU
gfh1goxRk4eE7c6uZIfTYp74mSPQcFFx3ITaIrw9j/Ks/G9aZxrhBy2bci0c4wCiDmF7JNH7Eg36
Sv3QGGW0JfuTv4f5r9frd4WXkPlrOpm8ZeBuo34tvILra6ftBsp7Tim5MGjLSZ22887Tw284sT4P
zy8dkKpOC0qdYvwvNpc29QP598JMEB+VairaiHHIEgpSgfWmTVA9tzg3mBIy80+JMXMEnwnhmNV+
vUAPrr8yXFcjwQKQL5r6ePLUzyV3qgThM6ZpKV9lNMFCyOddqC5E1hPfMz9rXX/ZO+W2oBt4B9xK
I+KlX5/VzeC8kGhkIdN06mBSsHDQhbzOixmBsKgJK2PM8J9qEVrrFA/K6tyg2tOc2jJ0ewZTOLVH
SaoVIu66fjK0SWjpnL6ekQhM0/nzY5YkU6TZagM3eWykioHRT6VXzHDnl078YaETf+0g6Q9Xqo1e
VcUvy2uYho5MwnP3GypnTUxTwDlYLI+tEssZc0VyPqycya45SOivsfS/F6M70XrEhStusE9RcmKo
kSuTHrbkg4Bv5vEliSZ4rpgiwVpl6S7BbaxhSzHaDaz5B8rwgptaNH6mLTI6NROhmHiJCp3k4eLu
IZPb89/VpJ8y7CV3DzuyqiR5+Js3uA/pve6YHl6Wv3YYx1n3Uio8KlGAwpLlQV5czf3fNu54uswN
yaQVVEd0dghHcvrDQREtZhPTUN6+fLqwvMxbEqCVYQTC3OPmccrAbeyXbGoOgxs6YmXMWsnm25vg
r5FWN+mPOt65n95U4dS+SqVDEqXlyJ8UW/yXD/0yTZkbeG40d3B1Yr24SAEMvezW75w/GEhSe5/Q
wP9lOSHm+uSfcbvLLCmqeJyhzAA+6x4CrO3Z+XyW05FGVK1zZzxOzGFRE3dlkHyzQYivf47E1Bzq
flWWzkVsAGF6Mwexj2/vwR0u5Q1Vd1tYRGAUPbA3qDqHWYh9mzj2bt5ft4EjxhXIqBzE/ZHhd0HY
PQGk8PPhoUDRMKOXmynUajpU60uyIJuMGtgf8pEI/WzmRXbOGbd5BHnE00KqqSURNR09SDsIyoD4
6UYlf5oG76eIjY5d+bYrGFx12oqvfF3TJsT2oAhc/YqlGEq424P1hJbPzWUxPiFgsUP1ImwNnse+
B2/1pvp3L7K/P7o43hYkD69rNFzwhCevQS7FHLeSCgB/BNGoG6QDGB8qKCGiFbpZGPBkSSlHrKzr
aERJyRsvW+SlvkPmQmuDcPmPCbHCYCSUnXp1uIQHcA12e9ThWVyAw3kwVmQNeEcDZNZUB7/1PgO+
gwFx0i7unhhi25B38oyqtPqbauVVnQSpbWxRygMzdj15XYzmjDrkg/ea/yNiG7TcSd6Bbp2Dbr63
rablrCDmPR3Ix3LbjQ4dIrhhgfvQINerIY23DpV2xKzmvhDdIpON0NswI9q/pdRwAvH8fa48YSFd
kUd+Msm0euUH5bWRGuY3mGu9nvew5OUJrJLFaQEfz+P4kogI8KwrDig48rqwRlMV/+r7kQFUNy5p
fa6ZrobUGIl0EayEMJZ3qN8Yq3Z89PVG5QTeb/GkrVwbfNvtuj0BboNonKaeQPByNNIZqkOgp7NP
L9VfqAos2DTsC69FcEr1kiku/rIHrJaaKkc0ltWrSx8q+qSnsxpST6sqqSEou3heBFCt6Duhb6w4
IsgUHQgTVelTukcJuHxDxNkJW63KSB4i3tb0Fbnzffq2FkTNGHiwSpeiAmrXOVkEzXhnahkdUUDR
btUgykx7RdZo7C7G41mqGz3FTP8d3ksDiKOkHCxlfCW3e0+jK84gr7sRDKDNS+2TMqHJmzY2yQVr
xaPsAr25l64nREfa/+HD+e2CgKLEfCkCQepQLb4K33YTylsWhiTxIj1p3gj5RjhjH9Cybwfq2Nhh
r/BTmO6m/lbcboqHsf6i39lCpLBE8fgnPaHD8t+lDbt68akIbskBU1CpJz1I+CRb4VrpMDQBcsTs
XCxt4HgViplOBfkPzvpCYZfL5HjBqZn/JPk0YHZSb1u1q0bC9idjgYnr9R0LqXf4C7W4o5jHd9Zh
TWzgAC8iYLXY4blbrx0P2SaVmwTpcjsC3gmZQrTtobbRpOlkHnmNXx5Ln8OJCF4m6Bzy2PXeUl8a
EDckJ9UBR5A9edt44Bd57EPLRej4rCuQHeQ08n9Fss6frMGOVCgLFdJcesR8UJ8nubJvjbzbPqya
xu91Z3+Ava33Yuqg3QDO4TBQXuqFssX4d5UfcsZ3XBLYZpGAYPj9ApaUFjaddohj7+AYAdbUAaWA
W8twcYh9rPw7c/8pWdsi8Hcu4YVFqm8Bg/Ty9kox2mKqP+Q5fYG40p0rcMuUCEEw5x64n84UYYfD
pHw3jfUdg3hTr+J7OBYRmJ692zBb0KD4hc83lkW84DZaN9iv+UCRs1gkjIRD0xnmtkjCM2+0U4L8
KDgnJ6FMju3Q+ndlRMgDHVvosDAtGPq0n0iz9+J8KiHXJHtWKXHn5XgxYEWOHeBcP3BAr/utfvob
LeXysxrOm8Rfpq9YukQl3x4919KC4oUICBtqigBuFM0C61PclV1u4c96jB6YtL3wKFBL4jUt+2HT
2F4ovo7kCPrAnkmrIBtGU/89tNzJsgAB6dr3ZbljFndI1AgxqE7WorkLs+U1D9wy2+aRwtaec2CL
7HVE54oSn7mFqIxgGt+gRidK8QKe73f3dEO1pxt2pHISH6PJD5RU3nbySSK4DnJV+Vt76/dxvDTD
i1i6jEGnMxgw5e+Z0Up0z6p9rIYJjg6atCWU3g+DTZD3baBP32zIn2x43xnW3J+z0Xlwyjx4IP4m
tl9mwonk4BxQwKhUdn7StNH59BMExPrAxmGghGX/+13VXFTHCIcRGDTV+TutfGhfDVlQrWU6OVgl
S75QxfuYTeX9iv8k8fFWT4TjGBEKpI8jXQuaiWsa4HyAW/KdhzMmkp6LlZtYiq23rgZ7zWoqGwgr
NPBSlULSRlGddVdccQS6F6OeKbgEQBt8WXYaBvjyXZaXjeLgKrkrdimz9Mn2LyZJ/nI32opoSaAX
qnG+b4Vy8kTnkXS36/rSfWfD3CEvG/2SulUm0YZI6gvANK/KZI1FdJJemJav+vAs87zH0eEbyH0X
G61hwdGAOh+yvBBZrQmaeuXimceTr65L3n1cKMpTEZY3axcLQ5liBTwJb8TaSilsbaKdmbqvNMT1
gvRgsKcLRmHAiv9rNpwtNfNDTHhP1An7Mz4sO4Y3uybRrpTKifRmHcfI1jFW/TCh8fxKT5+b4gIO
O3aJsbHc9iwFPSGbj7WVByq+JZ/RbC8Mb6dswJNgUm/GOkY87TQIri+5DLC+vWff67pPNnahNISQ
ASAysQlUZP+Nky/lUWOfnyU4Bus7nI5aMfA/rhzfO5UEzfd2OrsEZDcySyvMk1GjGF1nYn47Xe+u
k7SvPFwwEtz5fZNSsYpS+AFQGNMvzOIXilPd/6EzBLbEc2mrEslrf4JBfeLqjfjqkT+Km8BijQFq
lUBmt8alTHsHDv9n7Exdm4UkbRBCTH2r3tHxEHsCFxVT3gBT2nXT7NmZmbwX1/ggucnXsSxPI2Ch
DmBkHXLcfRwX+49Z+pR+vd0C/PTxOaK/fram0RDKJg6DylHKtSdetL36KqsjhOcJeA63X9zo6mKR
t2/olUEO73bYny+4Wsw8/77IBTDJMmdm1yPRmnSP6UEOGeHwXAGw17nOY/mDj9zHbBKJeuaGYkkT
uJLb+voWodcDzFxVvzMC4xUqT7Ujdk0HW7m2NKSFDuSq+H6PG0/db1z0BgHthGm8DcFkZylFxBrD
UlGM0X6FCDJJWnDAEc549qgsYfq1tbX2bPd8nssV1RdCERCr3FlliG9bcwHRv259C0CjNsCWd8Hc
jRKunKtrTibjkD/X7qZyuDivqDRoI7QeiuVCXTGB77V0l4zkazWxRG1geAwD+cj59OPDpIy3BX/4
RGx4l1ZIydiNQpXh5RIfTA8xs4BIGIse7e6P+b95dXlSJEi9c8+cLodkS2hAeJ7Ps7w1kPIebSCJ
EAngUodvFgFUpp6TTDJuFINegNIwPtJuqc1BTlq75Ysgmc1zKmKcJAb4uvcNAU2TQ+Km3GPSV5RI
WQ9znfgh1nPykl2wTx22/mkzYMzcj3xCczlyOH5hDz9lT9SzSOobt3IEvZM2O7YIPVe7YWUOmD2S
d1jrMpdyjbk3wmjJy5OxGDrgz1ox96VxaSsjdbLeq3dncXOaat1kX4jmkr4WueLYN+xUb7FqOECq
Y4cZxJAH3ad0qyaY9UICG08Pk3ghzzsdyiFlG18H7GV3zPnNNZf8rYvGRMrRgxN+e4NHBz4xF88N
FytsBruF6mvTIJ8XfYHTusa145nmf02cy3OCbw4LVW6DJ1nPA5OLYblvTL6JOrLUpD8u4IZUAgzd
hnhH2KeVr1mjO57WmSKwLntoVbYuJCX+B8USbm9zaqX1tCtev54jfmnPGqJ7a9ZeDLicTKE54iZ8
RdR1Xe8QLynIAenEOpKXk6mQT6ZDAQY9WXvz4Lamr9a5mWmpLxDU8w4AvIwkJyTXDWbD0oTEeXlm
Q/WF2XKfl/YwPRUGCzdeGC6Jbifi4xyBM4fwmKwA0sn62eR1yHhcLHTeoyM4FCesKixtmDhhqT5y
FipkHQq3lSE83u/akm2IwMEGKq3uJzyYT+0ldlMwMVQE0M2I/kjUBxjX+ra/41CML7Mbq4HxOgmW
xEbteYipZxb6kZ359QbpgTISsHyJQuJLD3qqNlUc6FdIHWrAOymzZnBMr986g65rzJuxoAyxlUff
Ft0KCH6DJ/NX7XmVsM+4aYY5uPiNUBajrEyqzwJYSx70x9QN9IuKU2+gSfkPXDAGmSvxv2qhSKj5
n36CrqqaFlhdE5PW6Mt2HVuEwUqPX6G/c9ptYS1oQDHjPYPEe/zyB3/kOaUWrqsUiw4acMeiK41C
cH7ZvAfUUGZdTlXRX1yWuI0xJyKtwbAie+hX1Z6430sNw4wDQUDfOtbsA9lj3uJwKu4aWEGpF0Gg
3IMSNvkfzeNkFf44NppCS7MpsNEX5Fx22TL9O+HSJ1Vdlpkow/IodI+I0CA5jWf+Zg/ddmSEy6/8
TupWZl8rnu1hhbThRDX5ZkXbjUKwx52lJwqeFZVcfquzSnqnscKp2ZEq4as53sdHM0J3a/BtgFXb
NTbebUJuLfYHr4B8qk2NDWthAf2Wjb2Jrrh11Uvaz9vYqFibubsrPo8hywMDYxqRF7ZwwUKTCO4g
qm4o9aMFZaD/NBBGJvhsKZAFRLLfl+q5Xa/XJ285VCcQXMh34NqOetrVAClMmlB0GK0In/UPlwwj
PR6o2nFG1rnebVUkpBjMs25bPejZ5XUOlbHib3n7uDwjfXh11f2Pi3++QDP4FwsT9Cpe7la9k3hJ
rzp9jUwVx4Kz5a+Z6nFHKc0HQc0Sj4SZCpsvNrSw1KBsCLvxIhmRF0ZfSgQKDSYdmthNJ40Aqpgb
jJXHnbdcZ+1JMfCKpg+grXBMKv3Go06y0YEpnBTTLzigtvzdNXJlMg+f5hO4W8U/mOmyZntB6bfo
2jnwOJHTzbf92St9APzjwY7fZjpB2dSSKYligQQ0Z8KXO8sMgRyqYIzbbEAJdbmzRCM1oLOcv35X
iSoIC2kCdBakEe44KaHQHzmcqcVoF3rU1mquZJd6XBRlGeoQ/7mY45YrQi6qrXy/R9ho/5YjAwxi
TTkNiIiODVsDZD14vTe2F70Jt67wQcDDJPnS0gWbvn2nu2zHshGBWJbwq5Y98EcSMu5jLA7xpoqd
EQDW9dmkyfPt91J/b8RhmWh9mF0wcIFOATjU/kpSDAWOEq56AbEMtk80UulVRWb2Wq/5KxoYnPIQ
x0pK/LQzE7Mt2Glratwaj8lyZb9oi+ak8zjzJZDkrrU6exMsFSw1EhkOVPfVxXklHz+Vq4z+C/jD
a9vui25ptgB4AHvEYG5mEyVSPbSVXJdvlf+1pVoAt1pyj10zHpCvUGSJXvjj/dJjcTGgdb23vuPy
4oGhVMY3WHFy7WP837gF/LDOEDhfdw5bJ2qJuWIFvbi1pVzUAHr27bmYpGWbYexBvqWYmbeF7Xve
iZNL3CzIfIYEYz7j71ww0XPfaqEaCYzJzNYgHzJ7Ygc2O+A+EySWHME80mDech6h8/9Pp9ybGls+
94GVkcqYdLym2f1bbJvfJ/inipbIM1zX3HfvsN/7fWK0iXRjtToSZEeRjaoieFK46yk+kcVNPqLg
DrQ0KGOGYiRUfcT8XjPNPzMO/o9UHN5vtnt51nyhFEcg/mpOfdKZoYGfMnvYSxUMfVzo5dBw+T1W
E9MGQrXkmlFAucEAxT0rQr8HZyTYEMMB5tPAD4ajjV8SeHPaFFF5U4QnHe/Y3DVoJwE8i3PG+2GE
5DqvzV7+ICttEoHE4zn3b1d1X3PXHgvAGln6BzgN1Uz/erMGRA5noT4pmfYNBa36kQNXwHuhiumO
4ZIQyFFxC2y0qvmAgVnpT+jzsfSG/hu58rwQFwtmYzA4a31cdHtARqIZR/ipETO+qyOEK3gLA0V7
Wnaex5g07be1Ea2/u8IxvVvKhNoscGfRLhCAiSNbXM+ccptLEo3TFRd9x2we9b7IgVTkGcv0132O
9DmdsATyFkgYB2sfRbKvW2G0mS8ZF/Le8wKNz2YtJg9jkdWq5MQnqRS5KE0T1s83qOm/VY4bP5LZ
6MDiJPuNLNBAi1VRkf7k3nn8qtWdrmQAXVFrTA/C+KIseZHh6RxURxoyVP7dw3TpB4PeK/XAo8db
MrIqfZMVMEGXv3V35fNMiaBAVHV/aAqDy4gkuSyYVDFCfHMws+UDGXx0+6MYoBC++vD76RBNezQX
QbRlhULDg7zvQFGA7yIDD/8vJIlyClx9zKDVQhyTCwjvjAVasUMtcZiOBwWmK0gfuFRcvymjsd2E
M0HVSUjyTGqJ7xP33bRtoBicRfZvV8zu/4FihvVWQbqddZtRgL21P+z5vXnczZUq1x8kmfwApSHJ
3jLac+9SCq77TlVCvGmyO2GOyKnxk+pYteiknm2PqYDgMOwr8CAuuComkMlou6uCuiUJrSlTnZbI
HybotMxw9FeQp1xUaJFDA5DzVR1ZXVs/6jm8+v46D4ikwS3mbAGjJeOiZYK8F55rIUt2aTkapbns
dgKXy629TnAzhEnJkXRF7ODAPj42gF9OwtD7KperBoY+DHfByhzHeDLRdx/Gl7HKgy5cIAQRmdzr
Mbi3oeFeppS9NomC7Lfd+HUa5LO8t7KrkJVc6SrlT30Oq1HNIR2lQp6E31JTK4qLFQwYUhurHL46
UjcbTpxr7TfzEoSD1TY8YH96fXTfwIpXYWx31YUdxnap5aZTLpw6Teqpu34Aswz7fmLuKTwMziYy
8Re/eyB1JtOBz5DiVlSpVHvpzwEEAAMBNwa/2xpUq3Eg2ThkA5WPZrCB70lHT+OJ9sZnsS5/IwkC
pjkuqx3/nmSj8Wf6JaAPe8hZoBqBI2T77DwpAlR6lMgnTEVnd5E9Dp4okBr6sms6du5mH2TlVdk4
1Wp7QG+BpRFiCba27E2yHvKYrHNWVRyq6HNWl/sr447UI7eTyzdRayoPN+Ejyb2l6qS9SlNYxVXF
1GbFTpcjtdjaRbkfu9pxROaOAJXswkhEfx4mo+J/JpnPGSlyaLbjH2tdCtJac0aWouI581q4bqmr
YmmmzfjuxxF2XIJc6LSrO6JEyu+HsdVzdqjlGPCi7nLpBSdh+EtTNbNGbjXIJemHjdBxp9SdMAPh
zNhfZQXp0KqRFRCfAKqB1n4TIQ/rk7kdhFnUudHpzdyiyHPGis2hGv85ksNQxgNeXv7aReJGa5LX
uidWA7ivEE5ipk1IipJy+Omv4njPmMky1JDZ8BHR7QTaLzeQJ5/LOzEFMmyaX/z5ZPdOA3S4VvXR
VI74XgGqPnC5XEJjL8/YxP/tu7FlWtUTs/meQt2CkHIICcHfarw+7nZZ0o7LJuvMPpUB33GLxMO+
LwcAnxKw0IDyW/GIYTtxPaDMGpZW2abAdUhMfDwpAyWaxbGlN0QBQ/pzs2n52LSb38pJ2aqnmpvJ
GooTxnABVKbixAHNvcRLntopFH/rjPFsz7G39KdvEnY1c7Tc/zXZRcv53w2LNJAiD2XG1xi7gpAI
McnNHZHDrt//jzFfprmMu6uB5J1EfI9laq8G5gFzVtXWiMwyxB95epNZ1huRKk9G7JTFmIUNNlTI
JvKIODwl409S2LKyfqVCZvQPGnfaJ0hjzlV4bh3kF5wSNMW6TdvNVsRvxFKL31TxPt6d5iv/gWf8
EAFWThqG8SdYSFXRbhnnfYvxdfbHkADBqzwj2ukeJzDTVItafoILpyWpG6feP5M1alAOUTa4tJ+2
JRDcy3gfu5f5Yz/GNbAzLEEQHg2W0ca2LylEPBfwbEjWIYuRiKr8gQbJa3X+GEdhYA/DpmOoYitJ
THP0BPe6lGRp20Ym7qbOd7LXbGR8gddIJa1UWIcpFs7ELp2pYzgnirxMcLDk54194zLZfQKU4PXR
iE/VYRCqIYRL3/UZusAl5sthhqv5lPOJ5ANxU26lR8VVhFhr15qBtvwgAfoLOzOpUwuTnGw4SfgR
JLl14sw5A56Q/I9l2xDWkm9eONAZtZg9Zxe8EHzjgO+VnqERci3hFAFZKNMvAQW/psM7F8DvLcFI
ZscLXjXz1EHeetdt88j0GTUwto5Y3LGWnRbr+emLrZ/HrRH4jZPAPXp8CGx1IgPrqeWiD/MZTt85
DxSHWPSgFSJGcwPrVXRQc76HB+u3m5QY4T0kAnWml6+Is3eqYQp9dMhGBOLHe3a8mH8jjNMRUiYP
NIMeqaCLciIn9l0p9YdoZsl+/sVzi4FbeUzRmtNp2l3xcKSwjU++h+OS+E5lVeZb0J11I1GFRIHG
1ypVgwTlFxuIcTz1DiEZLC9Yd/Q8q9dj7FhQUr4wESLU48dlwsueV2y1otlR6yk+lm75oEN14JWe
UPw4Q0OpR+Ez8/+kpUe1ud2IDqn5mUvs3phALVZicwIXOZtXsazskitLOLXOYLco7dM6sMOMX4rK
0IhaCgzoHizHJ/5Z9CTC2kW1M6DEZqApURfkVk09ixkzmq078Tg9T0Jo0FsWXh8EF5HmCW7DRrSM
eIITqGCy5rgP6MfJqqCNuLALcI5IDuv1wl4ZB0RM6j28NYzkEA1Cosrk+KzY5Chc8YQt0C/F32CV
UoUEZcIVgcjFUOSafLt4WrEguixqAYQmxBR9r6ldyKZIZz9NLRwgX0EUxkXLHyDE+raAjLfu1TFu
mQ/8NdGXbDsipmGba4El8y4cvF6sYhQu5Ykt18TMKdrAiLsOvtGmMaoy8DwyVBhU3fgr0lfRDTzQ
Ph8qTmt2uxykwEl8w+2UQVKbkm6Wy0bRECBZ4/r0xKAC9RQ8XFWoT2QbRUnrkOY1xNA8EPM6rDDz
1T6pXfX4VjRKL65YlgFiNFiFvmF19ilGkW/KoSXFy1pAioloXtLGzIU1x79Ae14+JS4di17WjQLq
LqAGsBUY4+z3W2ygVM82iMBkCKQUdHFE5vLfP1syEXxGAPDuKNb7BCA7IY8grL7Tj6AKwB1OLXP+
Z9kSPmLrCTbt7KxSxPWQRL65Eqeln+/hZsSaWs/Yt24TEONe6GrK6vBO6EujCVjtB5TAkripjrBw
9cSu7Eoa/J4aVsv7iHJIlYUqsBYT7Wn/2XdgbNWHj/PsdUeulPVv8i09xNrwPKmGPxh4fx/HtcZ6
c6v/zFL0VgOctT1PUrVepFy0gbRaWw1+L9/6A8yaBJK0G/QJW1totmoXOmQNoHZbF7q3fKR5nXp4
IT8kS9LmlhYnamYDy4QnhpEtKeg5pdqsmzDxx35185luPYsw+uCz1QrVMd7IWr3hQijgnJgXuSNU
0UTkL33vm+YSNyYmJhvTpm2e7jcU3JdxVcMZlWm/SMIiGWJBZ2Av19Pl7MKIHawPLa9jjfQF8xId
zD2LpVYArZ871LaoOjO6vwbgKLlUEErgbVKilZNcnXaVsjSV2Q5sS6o6EUVuKAwyWF/vp0zWeYjU
ITBCJgKUWlKrVjzX4+Ni95+T45y1LxuCQjCJNA60qDMB5Bj4H+ELV/E/9mvOTB5h+1U1BieHKK/5
Zv3IRoT6AeQClyFnS37ItbpAUr7NwXopXJyW/Bn+snBmHZrRI4ln/X1iDFIcqXqF2KmunvkGRoEf
+N1zs50t5QsbJ/ida800g/bAfDJ0Oqvak0Md7pZsPKsNoWNIriU1/iYf92NMDh1GIxeeL90YsTny
qRUy/AdisaxJ5wr4CO68uPVhUR8Ivb60BGjW2zc0G6MyCxkmV4ZpkduylQyfFiis6q+Ka/K3xsXq
GM05O8PnR/gLFRrxmwKMBda+tF8FJmL21wdzB+8Gm8KD1zZBnWV6lLxBmDrQhYMJUr9sCFkci5V2
Agxrz+fuX3jGXD9abnc3dlGB9/+XywsHoUmJZF5dSxXiipA7jvdDmjcW2bn460t4BjiTefwxOZnw
Q5ttRLZpZHZlyXxlx1yorqYZQ1vclhZt6ejNZ734JCzRpfInmpn2t6FLbKP7EwZy/694DPbdwuSO
aV2g+IqqnNuQirYGWEmtA+wBUyrqsOu8jpEwNWzFU7Q9jcuBTmrY/Z/2v7DR7HVEKmQi6FItKTjc
7TI+N1kBQa0/QU0BNm14z64O34UBgSqS6+pqEza7ec0yjuKTfTusp4lz0WNYgNpIy8uDVzwDoN3T
CrFE3auK27c2MMEkKmFc4/SlrimJzlvUms3NRlYRBh2d8HWApjWXys8/n2G2x10WsiPX+GKaZ5ZH
EWJGbTmzEcHyhi8lSYgJPpR5GbP4zokG9CTiklamAB6H15UAAay9m1cgX8DVa9Ch96AXZcq3IDyU
GleZgsvsXtExHe/bdc9XkUvwZbmlpwOGz3P9XJfMpomE1KMtNBxzfd4yGmuNuQDv0FSwCltACXC9
cdYj4yAX9moVoMfgrGVDC3Ver+3DN44DlV4Z2TPSK0smkfnPdzqNppVV15lCbFFnX8QTzdmiRv5o
jq3mBsNdyoUFVzvRT8JY+QYNJ9A2auZoDsqAi4IP7GXIrlg32CGXEr+fbjOwZiK9g7aBfNpstbWg
3erFFyaXS5FoFxT4gjYABBlSxCMnJ24hBgbTog7Y9DLMfZdbPAjRH21/2UUwc6SB7Xjd60X+OFM6
X0RYoyjPOO+fR6se0y57kcGdhV7IO8r2cp+stKavQ3QZkCeStgrMhh31pacn/BTCkkdzN1QX5//p
lsELKrnZz0takDRJZhe5Crjal7AGb+XV9k5wLYDRVsTLTXpKM0bs1Gjaih19FsgLtold+aWVWgaH
HmfMlr90Xk+UngLiYyhLOjVkSvHJ4i5ajQTTBnw5LodhCcNB9s9KHvCYRuABtUjzSnGL8305eBmB
E7zM2rXglg8irmKv3ptnbJ2MHTKtKSM3kGpHpit1aNd6PCnG0VU6RyGtqGtElzlWzLOe7Kcg5Rf0
yNr8SRCL/3agFtkMA1uZc3Vt3pImr7gfx4p3zp6mQV8M5fUsFPFM+wV/wvdmZHQlL6cioXQBWLSO
Ss0ofzzDFCgKQcqAI1d5r0XcvuXgjAAmzyxvCz5v6+kAzS6Q9WGEvzFNpMgiXorzyX/GCQ1kmCO+
DPGZ0pZrdqNJKODurHyVVBnNDWhxX8Sa/734dWB1SEgSXVE190YzQiBRqPM0qbI/SpB4grbJaQEB
m8g4Pl9b/k1hu95i0E0Shbx5UwchtLMFWu0krv2ruapHn5rXBdoITQ40N8mjxPtGvWidrI5IVT9o
03DN6LpVElygy5VnUVeT50yNFy6KL/19iVJqymy1gKiWhCovVRjxonHrSl7/ievhnRAwxfaCCF+F
GfZ1y7XMjnBuzT9WTydvBhza+5omeUxsXMyyRUYtYocap2iKcjsHyzuU48A6f9i7/aOL07VQg7c+
H84XK4Nv77YTQm/AI+3wphYRTBHnuZMAbkgZTglnVoEURZ7swJYQgAXtbP5L38J9sGemKCRx/q3L
/qbIplj5Z8IhEgNvJvHtetUs55bUBUAZS5qJgccviPzU8fMh3b3zvhu7eCbzIQI5KNec2bFsX+Ta
L3mN4OWSQr4Ef2L5wWIaARtz5nN5Wz8229lQam0UBXbJrJv7b2BflJSKBQTyzVT6KkqGKdZRfXv9
71HngkAfeQp2flgQkP4hKbMtaQvjpUHN65LYehhvoM2wQkXh10CxC4knKkV7AQ9siMdEqt5Oc0Z2
fwgRlAIwSQkPVzXX/uZKCtAMgWSjzrBfl8R3o5d+qXZBSWfMbaECbTxquZj46Z2lKOYC70wl14ql
Z8r5t78pCpx2QgSfhfuo0iSDCEc6Ke0CdNV8fFSDlN77swX5ZY74DuB/G1bUDaLkAt34NOAiLiD4
4EwWjj1pfbCBhQJ/PKfas8m/iYv9e2ROoOl+gn/TsqEPJBYP7vA+e50g313TULiVio6Erog3bcz3
4NX/wkZzsI7OniCseS9sdpi2L2FixiC1z8xngck0j6oIu4ZqQ2Bo7py6a4W9t1HN0GCEeMNKXF+2
bNmMy773ySM22UKQIpu5apVcLw1ek8A0sGEtDIZsdS4QkDhfT4djNENfof9Hg7ETtG64J2BpA5Ip
4yo2FuuCQScgY+82nNfeiRp46pxqZzy5Q9VDCTDdVK1rO2lTQ9XdSq2MPQzx16FhwTVm4kBxxBpq
pvqHduRBxbniGU2WovkzbaL+EkxFUntbMoxkzCjcref+QkrZ1FBKZDJxuJK9X0ex0x7xMsXIn+qr
MYXqitoyXWS+LRLe8/uP0p9b0IvBTP6gJWpLAnAWRuXnfPLFfTq3xbMafHq/TVv9RIcdfdnb2eZn
NaXsb5Fx0ForVYVjKvJu6JSPmpfyWeVFpkwzhoY8TCa3CDnJxL1mdOa397d4xkdSzJGXlRtVaM/b
6YU2k9o8d2y+COvuFr+P6LJIL2kOIcUom6L0zdaU/b/XMxA9+eXJx5sUckwZ8CKZGavValqncm4Y
UtUy6ku+17iE6BI9OD7rXw3ZrXqODcEeiXZZNaqvGIlWQA5clNhpGVnHu467zUNrF1q2EZisQ5Ch
QjVr3bBViCxdBF/v3UR39GYUkGJDM8P/xDOjZF4Fg3g0kjOOubXveo7m2kQlLwN6EesE97rowkcf
c53rmgzZcUCIIdKPq4SeGZc3ZAku1QGA8oEY+5WpxX/iwpoL6a/ij58MBs5QxAwXWPQiPPj/8Gy9
x2euOJikdr+4D6ex2pJaSN8tW8Ow2vy8eQZKdmsmm3oA1IgQ6xhRsotKsKYHHe5/Kx0fO/4XshgM
SRunj61gioJKT5Q+22CWW3hx+cuG2t6wk9zHJoi3y6JykyhlDiVnCwfTcaZrlux7BP/D3kh1LxAG
69eyum4/QyPQamFygecqh4TRZuuWGi3IKL/UZSNRdTyIvxgmnYWqWPYXMavrXro2QO9iKo/p3Bsi
oibDYTnbeT7sJx6ZDzmO2LXEi255JYvRnsFg/ubOIr/qefco4UsxgmUTfWtDXOn1SrmKea8bo+o6
2yJ/djXXJriNbLZbbV0P1qbKQCaXdcd3zWil++7weoQGgSlIjJCAEd3od3tkMK+G6ch5BHLdqDIH
L3wOirX/xeVG70lW/1ol+x3radgY8za93PttGwfiIO1CHmxijo2d5QtheNNYjQ5gkMNzratFtlYY
X0HFyQjfRiyiYzRh+L8XwGjEB5Ys+csfPJFgfVo3h1DqDf2Nfms14WInYss3VYax/XjxJr8kct/I
ws3HrNxZ2Gh0rMEdIwOm/MDNN+Al59pXVzdS7bms1gxWKoNBRACHJOT7A3GKNHwpEA6/q5wvN7Ix
erm+UWldFPnxVBE0g7AbhguivhqWwRSvZ2GzkeA3KCe5iO/RVWRsQz+j8eW4SvrTTQRLJqUEuEv2
zx3dHLD/aRUr8wmNlNzLPmofCUDgKpIBs9MfOSJle1hshVueTMAwQ9IZZCWbpMDPIltO3h+c/v6u
3/+czdnTxZga9mCdjoZBZMNbdg8XK9uHIFgGRVb04G19ElirbLOJgPItDuW1Xz1YCDoLWT5ff7oj
CXpl9HfAr3mDcwWCzx6owK0eK7K94LpezM/h7uyUBKEleV6BAMr+Ab3i+ntogYAkNDQ/+RzSlBCX
pXDbcCsIEE1IyWSKNt0uQJdU+83WjxyDg102AmnhnERShH6HvhMUR6lwVoqFGzWhcvLf8GdaJLtN
WPO585RNMN3QenFLzys+x6AAGI/7EZLDhOmmVatfOjg2glBvB1YPHIsmx+e6UENt2icgjQKfdotV
jyguEvn1Ec5NXbS+dismaIzzfPr/JeS3P+BHE8XEJAGNPCcu6LWdrfAE1ocNT0jyW0moJkJV1gzj
LXh6Yxn62ikB1Inh1x+VeA15XgvZQwzwzqrLm6oliSfvimn9/9/3wlHGGJ8VDLURGCdrnjeM6dBL
wOm95iSek9yuVQVBteplilROXZA4c531bLzvrNwfuqCuTrn8EgT07gRgcKJE3PWCbnhAR3h0cv4P
VWSgyPkIs7PoXb58q3ds8tAs7XhT4X+z6PvXftmaNF63/evG/CHayXrdBBoHLaZh1A7SayYjd9EG
dca590Ekvs9MDyZ/yFTX1TOz+BYei2FwgJPTgZ9c/UwGo36VSDzF4e4veG95j3Fod78jwdBceoSl
zZoydhKgLouJz0jqLuarkNJ6Q94YrQ3dwr9zIqbVbPTCqQUxh+DfXfkfDmPlm9pr8uB4cHr2oZjp
2HuvIibYeJ+V7BnX0lJzNpyRzOeLBrHZPPbg/7BNCdCkwU6ad3tGR7KUHbFufzymaBZ9OCTK7vXr
dPhdlmJmt+0M+KyXSG8ukHD/X1tpOAD7TqUpLqkqiLgcnATC6cJd7lOqXZPYHFzL/ZvoJvLd2ylq
ylraLcHsXCSX1zyrUANX5a2zgzcn+Fi8MvxsDtt5QHYPRXxngoznc4HZ8Z3MGbf3a5u0jdAVPi2o
qzLzJXpw2C8NlL/XvMeqQXcfbbLGCE+95FshY7DsP0SmVhzHChvZgM4A21MZ57FzotPtvqELIk1q
DSJF81GR1h+/dTYTvadWHAMbwqXTknIb+Rs5aHqpmBeWIdrAjAXbRYWZtmNREfYdlNdiiunjoAIn
L6eoga1GrJuf79sFXAWRcF7vw8hTY2oGgvQC/czvFIvrEaT1iRPXPEsMqsO1PHsL8rF8I/G9PpvH
TAumSMJ/UVlpK4jMOpDI2kOhxgCEOlNKnVHLGzXuEEeWORD86+EdcnC57YDVHoEdpNMi1p/Jt2ez
dw/NLA7I8ihthKbBZchYMfE+7pShx9y3sa4UQBPD3jaQAtng6BrPvp0vRZJ7sawyg2TtLH61Lnfy
bPQMF1eSQPsafMvPSXfzziDwoccRWrqp83Sp7xupcytMPDjB+JlssQzeZ9qBN1N73nhKIYN4IQWF
kk7ve4dHYB3/fQzHPqOF30WKVZp0sKE8zWDtn8hiKa7Te6oydNDTnGK1b3BKvjr/W60fBRB0eLV/
XivUB9rCXvMDCkOFsbkM4c3yCdXfBh2TAmv1pz+suqewi8q7Bjji4aavGCf3gu20VaBP+Z3wESqB
uKdzzhJF5mrBfj8zadrND7UbJCJIlkqricousqVxFxH0RbqzhhUzZA0ajiQM13ZCbBqguG96CxI1
uePNNoaJ/yT0O040G2vTP2s8PfgqKc+CHcDHhcUfxlKouhSGbzz64TuyiNK6uzc5CP3BppLLJ9un
RCurgJD+dy7IA7VuyWrJQiIF18z6p63IoY3VFe0BIchl+ICskjzeEDfoGQxiQE+9N3yPBaWj72gz
FeJH7aQyKqf2225I89cn05Ey0i8FY5EIEyYySKP5fg3zSxGZ3mpPjgxbqPh8etTIVxrbo2gjwOXb
W8pOtQ49Vbt/ZWhufFcyzDzlLVlhqtX6r/I/syKtl58z2J8+0u6MXaPb0Uin46qS4F58Dgq1h/yt
ffdtiSSUlAHVsnihRi1qDrKrn2+Uor5TxXTkFe1gLVOeaH7JmbYczH6XSG+ryAD3RKexhidW9UvN
I23mXK1nv8of7wqnfouut6v+I7Tmc3//ZRuD9L35RmHS+65iL9svdGl6WJwFWsQ9F93gwfE4pxEs
3HCSzK5y/rbZhUz2qjW3k+Y5UoSN+frvwdX2izseIbda6dzUjNfoBops99u9YAOzvWO5r2AMXMzZ
JUMStZFSgSiFXWYhymgTYaUQgVUY4A43jM7pPjNmBnRiZo76Iy5HyF71N3yhYPtUzErrOxyUeHr/
D5XPCmp7RJru7ZjOIAI6z2wOyBfMvWQOurHdHDZrJeVsuIdpmaIK//PfcMETA9mECkGBgp3ut4D/
TZheTgUyXlGc0Uqqufzbjx5dzohjkI9vo7q42cZ+uRA8yRndTsA7v8QsX+L8CfFxCe4Qp0hVSCLX
PjqlDTMTuFHCZmf1l7wNOWhiZh5yQ3TIZ9XqgE0yUVvB4aJPPz9sEoCqZLkVX1+KKMriqr8yUL0b
Uyvmoyy+f7YViXzWtb4UfQnJmYxk8ucxtTCXEws6wuCnJ3XKDNjEkru1e+YYw2j8pTXzs7AZjcX0
CdKnZw44xIaPBdYkXTdPCKRWNJlYiw7Tud2/OU1CJc6d0kEiN2RgcDZO0cAqmOGEovLsMquRCynp
sYUILEQiN6ltwPfa+/hLecRRF0KN1prPK12cKTxreZxIW+Epo8odHxbSDo5S3TTKtRqEkkMExa/0
fPeemIRBQ9JXzVeMp5Rveo5b5qXW+eVeMZSVa8w8YYAAMtGwFSXLTKom3g05mtn+AQgnf1lBS+CL
4NV1NMj1ud66Yk4/g8DynEBPMRa5URmKwipbgd+k08JUYSxms6hpMoIcgfBgFb693bd0XFKps1fW
O0YADptALL/6Ou1+nm9bGddQwzmipw7EtX5G38Q9fu7PZXrbSw+HJR9v+wNUH3CxWtOxe7+On/Ld
lHcq9toqZetXmRpxWI71yByIBEvfRzQWmYy366Zmvi9aIy56O++nWiWMrTI/m6ElUOiNP2WCAixH
44CilH+Rxazy5Bi2ZWMJ3CF8Px4taGil8GCbLL7XhLzOmLegMNz2PC0k6dL2Mwk42C6jc630sjBh
+F0MxsgFdhpiJEBuDAmOnGL9TwJwmSokFsi8aT4QiuC4hGw7YN2lU6QoYg3IqZH+On+VxL1wRMsq
+n+bd4Us09G8DJoFoFyiZK1uxXst5GhKAXBkmBiL5oG2Fkm804e4bAsylDmxMRRbG0Jbvdy2618S
NCKwxyWTJ/vGQLeq+ScB/DEUAz0dD468Zg7AqGkhwuTZQvRxzheWWWo88p5O+oHT2VQTebNKHwfk
PtkTI4m7hSfxEDzH/W0Xp3VcwgjswytfATSDEDIS9ZlOsxAcBJtTAbjl+MC+RuNbV3WBBE5EGAEs
OvlTKNz00otYXQLVyKBqiuaYFG7dnxrroHm6570fY/iprbeDMvmLjk8YeE9VZ+pcwj19I3t0Gy0O
glXTa1OVYpfiotMT+0gbo++jCO3/1iiLAiUbNhi3bOHN4PSux8dPR4P6AI6ePZH2/CK30bIBwF4x
PsP7LKIKZVBrisRXn1SWGsk0OSMEDS5au+rcre0MtH/uVvUvC5e6IINwtsrwHxnU9aE05dSW8bjn
axOAH5M/I/Ev/spcdgNgt9o+NTdNzqVzjGYAlrBMCmbJkIRknXGC+Ya0sPgEEgZYwAh8H45UtPKS
kTtvZId/nLXCw0AKkTSfVB9WPjMzv0wuN0NUmXhs6tVgRxVK9gvdVFRaRzUUl4k1fUJGmS5UB5nO
ddM/VcUfMItudA8ZpMeL/Ur/EVPCciyO+t3wCehSWx52jTYRDTKe1hqU6HXJrbxzqXY9qmpGK4P4
YcNCrBMm61WW0eXdx40yp4MdJ0o2OObaCIcgEnAljdGeeO/YGIm6EH+TxPm09RKQMs94em+3VVNG
kw825zq4X+XfODg19R9Mmfcwnjo5KDzG2UII/ZeilinwvuBobjNC5L+GgSalITvr3ClIAIIU/ul3
m/o0gm6fJcoJajsasmFjnmQMkm4UssPfE6jA2QTZwC8ENz2XaEyYFBjMguDVdXwyYC4n+JqI3wtk
w5aqflBidAeiM5Oe6HuWxWax2w0ZefDKAJvi3WY7p+/kw2RSpubEzGzDVRme4jaztQZgNNoaIFsB
B9eStzupdknsxvW70pct6cjjSfpTmhi7fTmI5AtNrMztlCtUGyu4ZHtNkADKokdANTcr+Gko3/vE
zd/xefdSj2y0ke9OvWIno8t8EBGNcvsOH5P1lHZ5z2DRPH/zhP/jv7TiEqRKu7x4nhDzJIXni4wz
uQvKHCbpeY+q3Eo1tVz3WuFUXUA8ir4ECIGOOHdzoSQSLzd5xLBmN7e+okq9ITwDYxa4FLmYf3NW
++aOZFw6dyDkXLHijFXW35xhLdULBcND/aw+FYrTBnOy83HOsU+D4f0PPzDljtEHyeBb+lieq5CL
oXUyScR4ZPEPsgCkpfkUVEgJYGImZ2bGIiUgXCYcaVCxmZM353hWM693yOwAvqo1ntRG2Pr/llLP
hPlAnOjzl0JDhToe6sJJCrMSdhyR3O5BtNvi1JtlVWuFrtNL02wTYO/Px8HtQEuZXF6YExQG5JY8
UA1XcIkhIErM8FyhVKjsgsDWvtOrajZeU0U7KAUWWVVD7daHZSSy3gslf70WFnJb2YCxrElV3rUh
xC6WJ0SUYSMAibBTDp0qwGqM9iQL6QTlgW90b6hXtdcv1bD5skSzxrD7zaK2m4nxsm8S4/sSd+n4
WFCXKzSdd/oxt3+XzvUf182KQ6Hn1a3WTZL63EXdzifLot/xuB/vnYxETSBhpWIgPBXJlQKE0ewz
cYlxilPgfg/CPgGGcTHc50z8FWGbInZKXiym0ogWFZSDbAykG9ZfCg7+sTpMkcy5qpSc3hCW9gMv
kyKYnaaUusJ2ce2uFoNKo4hV9ofTfPrg/NlaqWW3in3ti2nV/vgUJsjkqHPrHSgUU7h+Xb1aDTLI
V2AwKFAm2wgfxxFYqoWI170zA8WDu7RZUb9Uqargvn4QXIA7zM/C44yO/yMdWpmL/KPsxxLS2H0U
VYnoNsIcU8vFRa/tyZn4TKCFT1ZAH6w7maQB7QPQLouTWr7qzgYGOJ4jbe4QVya4Z11CiWaSBQxt
O1vzhcHkZh7mIQWGoBcj6X6pLwF7n5rxW2pLeoyjJe0NqWOBkvkFCizOVQHhyPKgedqXf5ed1KvR
sTd/5YprmOjB9xnRJM0qs6P2g9YiZkwwB4XrTpiREUr8CAfiJOAr7pwQN+RGpGevYrKe4aEkUYXl
NU0rYWyMMXl263lDN4WLbIzRbt61BHO+ZSmEpQ7qg4euAH+A+VKhcTdYZm8HJdmF4/3IYfqiPHQa
m+sN3TzgQmSSvozW4DjUG5fZS1fHclX99kKf7Bjk8fz52BwPEY3su2GZJQ1oxdQfLEkDlTzE/kKh
6PCwk/Q3cDoi8JXz2cHnePEnN5kFJFFoHxojPA+sKuTjafaGXFcqukAg+/bbTRf3n+oqrQj6HOzV
KkdTJRtPLeYbS+1MuVB8KLmo3slNhvAOMvvgQ94NaGIKPalQoLPYIC5wQzsV3NKCB4iq3yvXlNU8
xK7QyJInzJwzfrjqoGjzugRzuHdQVGf/1eUTK1dtfpKSPcEoTcpw+sNGZKwtUerMP+0bYXQbF/nR
P91QTJald0Vq4YWPAY36J7+1D2QT8reNS4l659WiRvvCLpSJGtHKoUmE4eCZZtjNRkSYXuxQfz6w
+mZpM059ZF0aZffpHnsxl14ImrT4SDvEsMSMELlQ6ek546QZ06iEKWtqSI7ZRamO0x0SKn5jhKob
i3cozRV6u8waevP4vkca3aWcOVb48VGvEtRr9vYNZQHvZ8pLeHwODoI40Yw8yEwzAUpk0o3zFYSa
NedhqweuLb8z5PuYHH18J5Q3QEw8x4eHfhn0fk9uS+ca3qJk78yWF3hzhBoZUC8zRvJv4RNVszO+
69kv/ueLunF99juBJMFUf++Zv7gFHO3W0lNYg8veFUYcqjHWol8XDE7w7Zpjb2oiJWiSSlKr9/7V
1D5AYk8uYVMBN9czZnMvRASJiADPvA4mZ6eZ2cxZIdt6SQgUSeGkcZv1yueUS6hm3bx/R27rZW1S
exeGFzkYa+ArE4efPmeblZkNclv2NNuUZawtRRNzxnJwtmxuShDQ4oQEL4Au+48Ebb3ECNJjFd0r
N0lzsGQwqvi0uX8+E9NlH50xuM4gGMOowtepCPCzDw+U8Ycej55tqIOkL4pj+x9GTGROYGp2YPBR
tyJypn3zfmb5Rs7p0i8Iztvmu8JbJ+ik9ADxw54BVi6F84mdzt8HCF5ZIzwlXrkyQLtF4LfvlpP/
XGX/3fyrsxDS8/yn7GyQymbTUxFl79JhpChXTOFh4VUq7QEf389VHcnt7Jb41iWUSU1NUVvr8H5d
43rAciNHxgAmK0ubfV/Xh7fmmFtVYUxyzHk/yf8FkKMq4yDwDd0bXopoDV+P/IQDYG+5btLRnUeA
IW3yG60oAHi6kFjkj4GQy3jQsdlzbqVt8f28sAzESwh9gpuaSkiPjlvAxSDuFo4KdLrFowzdMibH
4pTMDKnVboVUrSXIOGG65whBstjOUAHvWBi5bnDvxrM82duyzK/uuj6zdjvUA4Srg30rWxLigmPP
jCWc8jvnK8F2ZfdF3cgDnsL0loP+t9NLm3YcrUsGrCzBhOUR9rLCI4YoBiPiOdMNPsJGf3gYGGch
DAeCCWGN9XdYpJ9dZs8EC5DFoC+bFFw2DdXKgHyJzb/Q4nbxJM9K/ASyMqGhDCjk1VRwNaT8iGUU
kD0dxsfLmRE8HxNmyLLuufZS1vGkr/Bp5DBpyiU92WXt7q5Fmb/csW8T/m+EY5QWjwD/Rd8oepCq
cAMn1oXSnOvmSSlAGwUeWxGNwmHm7rvJwMP2qGBFCvRXBYO1t+9wGZIIdVGtnVdPW0BBxd+2grj9
+NZhMTJJrKjSyLeTSxHkaIwZJ4LzCtNTldGzXkJQWZg4rEL8g3ajQnd07HUDoryinAEKq7zWbnFb
OTNY+A8wOe3h0ygLlMcvuuAwpLtBVMK86WdIXGB/uIBZozQvFTUOHsY4qVHsd5I8i9ObwVjGxoOn
TA+YHcKFP6KU+cNj0U9lRHQtWU7NkbLQqlFPvQyvqujuoyzZ8P3fI59OfBsP0ugWKORrfqK7jKkp
uN/gARbkjruE6+6eHkKTPbZTP90eNuKnxfIekOHHuWYPny3KRzNH/Ftl9ausQcoK8HWxMUz6sm/N
4Ml8ZRs+W5Y1b/2lp87e2jWwKMBFsHZNiGv4ajDstYYViZNJATbv6FncsKrtBh9f+UBTfc6LoW7v
vZJchyBabBagSCUPnI4IFO9WqsAMxXgUyhxtNSaB8pUA9zzis/xGAxLuWvNTq2pLBqsBVQuC6UMV
EsUnKy7lWHFdQBEbOhmn8361gvXI0NEMW0w9bYmPZyUJFDCN29sIzv6kUeV4AKnNjxJkygEFuyUy
b5dUc9LW6+YIx9qtojyTTfG7M4O0gt187GSnU0jkV4WYA8doQe0Ht8z486gGIswpKLzRM0ZlTkgo
4TzXCzFWvI7eYtJlz9NcLo7i7YDqq2cschlDD1FK4fCav3aqpKpgWMJ5iD0xmaxd1839rlPSfenb
XjhU66jgtckaMFk5+L51MT/3viJE/J0XldMUmIsRLYU6LRRYd9qjpzaqLNGpEoWhRAuL/ioNDcxQ
rIgzsh0WS88ks0d+nHmt7BrC3c+sY4vC3zOsxz8SIRBJVMz0bdHByqrx4d/8jEzLDuUcpd6XCDE0
ZtmBFYb2yGDoDyECuxgIGtTLh7eHT3d5nOyh1exlY/Mwpj1cMnJ/1F6DXUrDsP04XFeVNceo8FM5
yXCvCGQhV1cgBXbvPWGIslV96+rPd0aiba44NXD6ibQDvLv99RvpWVXwk84Uh/oRuVffDuAHJ3Jh
UYsFBwDKxfklSv8ddMdzpD5/tCg+O/UIJqfC+zoNtN7/4uwG8cLBzrzM8+zXdLQYdkvKdYk69MMt
ODRMwpRH+c8mDLENkRQyT7hlQDULiioFzyWkVTQRPP3YAJ16yVvMQLMdRxIRL1QJOf1pkj6Eja0s
8SPJYkkZYCWl52PzyI2AEx5CtJaJkzw3O8WAgy3ubjBWKfDmA3cG9AZe+fZG3SfgU7OKjrWLLt+E
3+C8b9ystcVDgfkvu9Ssq+aMzWRCRaCFMTF4lceysLGmaQlFVtjAhApOVYmvna5MxnSO004ph0cc
CnGrDR/esERByEHhmrwv7rAZPiKsGug3MC0ZiFXzXgelmkVGczP8JzC39Adsm1+DOUNOwHdAuGqg
HWA7tY0+NAWAuEMC5CHLDdftRexGcBEGLbNIkxNeA6W7K1vWxDSc6F7ZjpHiuktV7EN2fhMorAUW
XL7Amzse6opIyggYiUYI+8WzjzihMvf4rAWXC+NY5m49DhmHDY8Nzziw5Be2V51VOGY1IVxp/A4d
GXdXO0EIQ1A0a0s1Go5ATGu8uz8Iag91nAItUcAQEaDeeHhFaXH1DdRP8bGXfaL2pY565lrTVJCn
Yvse0iR1k/a1+dczNxBbIl3SvHhHWDWI9ENI6gfXZucvXH0FbgNEiFTJ7i+I3sz0d03lzy1rXvvz
wu7H/l5LrasgmZk8Yv/jg9GcwmqQ18yokpICH0KWXaxZo5gYkThkVsg96eW/oAKZG7QAgrqVzB93
GCsCfC+7FKEY9XoAZAk0/5CTnQxqqdZZL304IrlkwOkN8eceH2c54RVth1fW5JPrrJhKXcTFHWmk
gUMxnVpCt8V9umoqWT7gtZrf9Iw6ReplZoLZVgaLGcVhZU6YoOndrVMRsOGxuan9G9Z8uBbIZ5Dj
DiGI9yabLbycL+BDo3/SDUQKyU/Urjnqh2awK7E7ELsrDq9W1tYHrWQanpJCJILb+9PvV/aY5r1Z
tm8KymjjV8wmsXWJAswVnXTTp+sze/Y/mVnNXQ/HHwbMXMuIHuLbyhm5Y+s6skv+tHxNkUxs6Qbx
rahfhFLIPLLjjnyoZNWyeQierPR0D9ynCGCagJxsV0WemwwyvBMwNwyBdjS7JPDayCQe8re+Pq0P
daDbW/iSUafEoD2CnciJK59234XQwUG/+9rluzUWnzPwleb5GoqW1fQgwLAmnZjLARc+9K1zK3wm
4/HMAlXKEHCU6hO47301LunJQ8jUJSEZsKM4tmq+v/pmmPbzyV24NVKhAyatbhb2Vka24nRgvEgj
uB0QHPqqHMf4AYj2pDJq1qVyFRykTRqWAn7hrEflSRGXGqlhYFgNXvuT+yT13tR+aUkCN32U7hLS
7XQZspU+KYG16InzVVthZ+xwKZ/aTNN63pUP23a9CM/LI+ITkKF7oYmmp/YQQIq1OUT58ZUa4tb1
Qop4XUmR/RbOWgNLAyAdWqUrIn/cki3H5moKwi0jhHnEdewis/jdQXH0lHLGRIlAkP7+CuDKHUSI
Ev01/2a222zweDuh318nnphiu+6RwY9L0lbyuaxb42gfkAKJJ0+DTlTxfEWeIiE4C1erCorCX4/s
QWVTA/+OQBrBP94pp1b93+MgP4g/4fgBoKAhtaUKusYmDO4VLsqgG+vAY52CkQrJxMFfCZzfpptJ
FrCv9hrSqpYwqSFy7StlTcottVYpat0Dvsb3Pn0KFwBx8Nh6x0CyXm3XXJ7UYGpMjJV2Yue1GvLM
DHtZA6t1IQqtQPlNuYtQ9XmGZ7P8JSAWrdw/jO0sAKm+NUkOV1ZQsZ7jFoKOjKuoYRgvYIfgz5Bl
/8LHZDWJgLZmugAgZHMdvXo3jzX1ISX49MiN2KspfxwalVSSFskrTvXZbJE3rXJzuC31QeBp7ItK
hP1kQH7PtTbKAzSH5KmwDERrCLu5dzadAGJWW5qerJVRoTKDCgmx9NYIXuFnXvjhV/PzFYGK+vbc
TTUd1fQ6V55xYeicBGRX0TxoJwWo58+qaWWcfAm6QU876gA0ovCLriBvm+BAm4u077d7xcW2wUhT
zP8a2nvk74fUSd4xzYPVK83Cv5pHL/IgzU5QP9kBEuaskVR6YZVHDlkGA/GqIljd87/GZ4FkM78M
0x5BEiu7Qrb36ET/ICXuoVpobpnvTa2vk4HKrqpzW5vqao17SPYGOTC0xwFDHChTQiS2RApKKuxA
hRXzH6flWkp79G0NFZw06SxeJBFC+AzLAeS/rzWmNtM1UoDgLxDdzKQnXd8wqhzQFaWvkZK+1brc
O1B17AhpoPs1tJn21BLVlctXOfGKjR7vL9oNQQ6IgRyasUEg5j1cMJK79UcCE+IWkuVH2hcIrvch
gkSywjz1/NZEO+c/0jEeAYenmVPbPFU+M5b8FUEJMCt1H7FJ25FH03Pff69fa0puqSoATFCTZ/yI
xVzoRGzO4zpgo386fbPGb0pK2IUqVc2XrISpjWOzXu1lAsvHwJ5DuYJL1CuBtFn69nnVQBh6cDm8
KKb4qZhVRVjabXXj1ttWyOZ3PRkCTtspiposD/6/9ooeuYIbah0VgsjWWFjJ6AX1GA/RqgPdPN+P
FHP/bFdLoC5SFoG08k6A2RX2urx7dx9jQ2XOQvy/NiHnqwKzzUl7DJm6ayETkdZ09LGWdd2xJTDy
6RTzMhe27fQg1TaI+KQ5/zxxfFQaePS2KufngcHAmBn6cB9+aFnKRshKxYaif+JpLVvn4EjnI1Dq
vSdpxwcLtVM/ReWqQKoSr/svBELiOJRiVNvgORkMJlzuBE48dz/sko9XonncAHCGkO0aP3jmefq5
J0WjK/8h0tQfThEMc/Dbesp5glLwOt+Ticp47YlrBHVEamAW+eJlmauCZNW0bdHizpQLArmbsIJ2
wEUmsOWNeKjfE+eXxmYNmNuqlxJyiEyU62GGW6fNxXx/o1L6Zq0WLARSLjBc8IH2nPOYFWkLSz+j
9XARipbLMaPdKxXVMr22chM4tVbtwdjmh7/EogCmls9w9aZnSzDQp+T7BFtYbm54ngXGRfm8nDyn
jVU8L5UCc6owu+SMkpQPodO66swfJYpIk58M7as34X6t4MjPSuuNAqnwoPtszPyzoeiy4nTkIQmz
tcrS39YKEmgNGUjNDYJUlbUS1jfS7/Ui5fRDTzKi2YqokbrbQ20Y3PTtOwy0y7pj9GbhJm/S0teU
/0Njmit6nXbIbwNikZ2af+B+VUGMsvLweSkfw29iwliqmPwIWcSOrLo6HtQh/qOAK81UWqcp1uB4
Xu1+M0Gc8hWD0R3Rx+s2WIdcEMkxzM2p2tUxGLbC8NJEBXXgkfzjcXd6WlHm2ObkztuI6BKSrsmc
MLStXjGQhPPzJnYGewLkxWHCkcLnvt0qP78KsCoGGAjSJi2DVS1IMnE5hWZgnFopuSL+47VxboY9
lQcqnT6HfpFEp2ALRFRBORMqb0jNJI/zxHCeq0cuh0B36gva3OnSx8AIFA7p5jXxR888Zn2Zojzg
6+K9sXlz5+sN//iVp1xqqnD0xyqQ30CBG61z6+F7SPZ5GCS94XjW1aAO1YSfxD0AgBNFhZM1UjSf
PVcIxgZc3j3agcfBIx6SsPyPq2l1a31Lup+C25D0bxXp8ZG7HmcwT5dnjcPRQK1e0A5A3F9ISs6I
hI4u8g2hkvBZ3nmAWuPuWt6JaOEywbv9rYt7vjMTWtA8Xd04+kmVqfyqpc+2C+S4VTo+dp1cFOfw
xe2vNXHFPqXUU1xTQahlqFc+Zldp5FFOUL32ztnbk57/tuXbSkbZkdepbFDCzQZ6TGASyRDjD485
N4gTwFp5g0ZvJkQmUotloDDYYhPIAqfGs94J/6HOBgBHQwi/pTRPlBXSJ6yEmjf3SVMo4ehNgSeK
aXd14Ek0g5QRcztIBbS33Ru6BaLRdYKTzgCi08RNHoFPXucB8DQY6BKIue9swCot4ah0Ym2DUJXG
mbsbU8yv92/zIDSmIdlm6xMVVDo7bmrQpxVeXz0S6lD1YvZUEbBTXSuoz8ozjkDLAz8vDliIqKHp
rhiQEGskR+rPtlfh7/B5K03YCDG7oUymuzRHnVbpV67gKkmAw5m1gTSVRAzsosINa5SjQWtwljbI
CMGjDLGPmrVHzYwt9JnwP7daeGdRNyN1rbefJwjFhHggoPx9D605jtTGgkhY7QsPLw2EGlqYOK2r
yNab4W5IUNqPvSNrJA93yI1AIVyiWkeZPxxmDppFKDliCRn8W+fICtFfFBD3/NBKaBXdOjW8Y2Dj
BXD+Elk/D25xhkGnn+qS0xCgsjBCsW8R4HJTDu1eHA6EXGM7FbeDRTL33gSq+rlIcoe0fteKHFLz
sQ5ceCiAShUesJ1QlRFMEbF9aAjgDH1bJY429TbsKe8ACFxuNpIyGoIhU2WIYhSAXXQ/XCISoCSx
bT3UiloSF+9c6/f2pjvkmkJug55zqEwsEB+s6yoyrDK+0t343p+jZlXcVUOtxWhGwNllEfRH3azX
Gg/vgo3a9VomI9/4P7G9UBaY6S8oIXONQH32Y3L6U8fJ1Bzvt5254bN+u3QWnQ7nG1kDQy1b/F4n
7Iqm+h0pcCjDNgIERsgriWscznjU1fpK88SE1Hhg1srmItSvygCddiMyLSbE/PkwFJWhuK0OQ1x3
MgTTKl6g20TjnPwhMdKvltISrkfR+nwLjCBQK5sLe90OTChN/Z5txIFikIo4X6HHERS8a1I7CXLV
JNu5UFAp/kwrE1zXItr1yGZvihv9eEYc0I/VuF9PVv6Lg9GmPq9Bs0seIZnMP7iEkXjJuSm7QoIN
VdDi+G//0etSC9Fp2cpdx7YJMt2n09RIf78RNtQ8c77khE7/74ARkhPVEsIUtHw2TMhN/asJxkH9
iQCrYqJYrCVSkK4CoYM2d/H5cAWF5V+loYXn6gom7S9hhoCGMbg+YmfaPWMqNJAPinb5aoT/UcL4
Sifcr1/dU0yZ5xjre5agME31RPX8W6xcGtWv3NBy2WsS72PDQWQKVz8i51nk+6jqqlrlayF9sg46
5bt3HphGkZ5qh1OM/5XXkFcGXooUpwUVcH92jIiZGuGcf2nwc0BTZfzlH4FEVQH9tbSm+zGxgkYB
cJ5O6sLxHvfkjiW5xSEtWXfBQ7i0+roginEhRFFSZIXscExALI/VBB9BGVhV/H3p/oL1ZhEgoLef
p8Vy1lAOOLjMB/8lkEvUgWHKhhS9aaHPmdVWhuOb8C+TiCETcL217lTw0/Xnt79xSs050OLJxgii
vJVGbtshcmmMHTOZcvQhdfRaV211EWH9DnnRyAOtXKqoEy727kDLvwttDcb8hq1R6pU6e54SbKxo
w34o0TXyXNtYjxFnfTyfRxDSlMmivhtdUczI+34IQet0Ar0v56z4yYilNk8v8MlU3nydFmWho6To
LGFgTmr+N4LgWNKE9j97L4sdDFZ2mQ4g+mPIW0iBvvaQKzFdAyGR71l3wx8c4adUsDG3cnMtDtZd
UjjPXv2MJ+LT8yBEQkyESXYzSmv2WzoqTNBp4ijAUyFDdNxHyWkT2VTowoMKN+6B6dXJG2iygKCE
qda/NgCGLfB6N/QrtnatD4x3heGiOC4KntyYjRlwO3JWs2IKTKyC6TOa5Sc9FmgsZpKkAjzplGQl
OyCrLcdMLu96NzH26M9vFsruy22mpD5VWO+lNg7XFEcdrvXTYr6TvEk8JqXyTbLV1bsQVX9s4/lD
DMj/3YaZ7MQNu2+hQJZfsupvp8ulA61M+2R19zoz0LsM0Cele6GnBMhZ0a7rT8CmtviIzF6CxW0f
7HtE6xVbuhxWsHcQE2GqQHt/6GO7MKLIniekASXWo3MIGGDTGw8URKKEKg83746HI7n3cW4ZtEtT
YR/dZQ6s6O+6uxi4WcVlr67vzvHi+Q28+q9qvirKygcy/gcQ3LHxAM4AhsKqvCCxcGUd+ePp/45g
wTOwEJDVvEcQzbAeHP7Li9LZ73De40tdPTS8KM7w7u4CGzGSsldI4w0psPoFlTkymoYYSFML8qA7
Vqc9fy043ySLqETmCw4uMPEFOASlRfTtx2xvWAfY7Zdq4A5Ivwzien4745hoM4tyl3/CSaNyvkio
r0wfgxmSRo9X+Hqcb7tUniA1XTYrHTReuuFsZFi6dJ6xXSi+wfmlwLMPZwAN8TVCa1eHJSs9heFX
c2l1MLw9z7Qz6pz+UoRRksfC/V1SQpwkYPhCflBaV6FBNyeLlDcaw6EKwCjRb/TuTjl4Q0NmW70f
BT1D03E5Pt6r07iZ+7n8kTT4oD50P3+pwq22n2gG+wLzgwU7m5pA/9cdzEMBMHLaWZzpxC8mAyAX
wWQUbz+wdL9B388oZDsAyucMnVNTTPWkoKrIbdWkBJxCW5EwADn+TXVZXC9TrwgNG+2jW2c0RGvS
DnQS5KXppIpFubXmbf3SboVV0+QO7EuCA/uMUw6nlfRKUwmdSUNR+rhlpZE2pX+a9nvYhPEBaHyF
PaQ96QSZuJROZ2YF4D04LObHiJU9gH0z5b84c4BnwvkPZ1DQ6WKtTpCdFL7ux+h4vNsrH/Vwtrex
ORzTA10jGF4aC+0ZMhZcsvh8HydZlm5bDBvCfvzAUFBc/TsARhX1rID1MxAm4Y3GkZR0nnjobSHv
Ny67tuM2m8TzKHN5c5LICdUk2CzZl2Rk1VseVXN08HYfITZgwkae/XKakkIxp/kmHjqaT2Vd8+L7
jpCA5FgoefgudjtrGIUBv3Or4kjuPs9HMSWEB8J2eEMPwdez+rsA18lbvekozrn0m4S+YF+AUg2v
fxy6I7f9BNBQsfxhx0YckRbqsjEIFocfTqhhSLJTas+J4T2sawV37jqjy4jQKjfvQSeG+0EH3bRf
v/zT47Q3ESFHTfdt46YfDXAo/MwhraZds1RW2jrpxtJeuG/9z9UfenJiBnnha9D1r9MAIZHP7xSZ
c+UyRVB+2Lm4SrEGlMz+YEi9RoJVtK5zuQ2kMeE0sZxBFvi1AP/vE3F0mBU9fBymaojfO74lsRlr
X6lBqa5xNdupSGak/QWbecsD++w74Dq9Yshq0VB1EL6ye1qy2T1yrYqKBHFT97L5WCndeRl6NcOH
U1yRyk9vwtJtGA9BMU4/L8AnI0v4jKIWkHgoJcO5B0A635mWc6WCN+3MXGxaORhjDjR90GtKO50K
Rg89fodksOibDWiiWGvtTSUGOeC9wRIPxKvoRjzAimqhOYzvg3kfedj5PXcnmb8F9rPiktQsIBk8
DH5Uyeboa4YewCuhd1KU2lLY3YHgaTfSHyH3hCPx30cKelN9PM4AWOaCWXZ2PvlNTHDeBaek6ppb
XxjmrHszL1P5oh2tcsqKMAiwmuhycJ3v+FjVGAMF+7nZBvgiGEofbKd1DrSqR4aBF6gUKxeAv+SF
g4NhFn1Adyzb89FaAfzFF82vYmW+gqmcnr+JTxmluyxf0puOd2rMPtB7H71LqKdEMFAhuEg6NbjD
3Ops7K4r9QBgKnjId6U/Zy/FpDJPlkMQ5+8YMQ4F9gY3Ip4J7FM2gonYaW80GccYbqkwzeCm9Ylf
07t0HtKcBFQbkeOVeDhhzsr1b8KU4GqFAs76kmxRzlif6Rytuzg4MM11j5agS84Nm8ZSuNNA+fpY
Tus+ktVPvyd7TKA/gEYbb0kt7y5sBp804f/X37E+XbK8MeQ3N561Ioy0AUt+hLrZtXZberqQEsdI
oj47ce2cDkaVBqoST95rvCGuJ76nYkfMm5tiJAcl2Owg41DGivVWDrYYsRPK6wLRITdUa3E4Ib/X
YyYae0ag+Hb6+5U3nmbgns76/Qh8mAA76Jqp1QJ4R/eYt56KEqbWkV1rEAbz08TeKZF+M5TCDCA+
nZslVAl08o0ahKv1nONPoWarDVPLb3J6c/29Ws6hx09dCsMlW6LbEyfnABa6nWMCpfF7JB1U/vmo
/tN8xUx4VfcvdOIPKErw6EBn5v/qeRf3py7mSsBxH9bbxlQH4NPi46C4SKnC8qtR8WsodoywGyK9
44NCvyEr7Ix4FVTxnnPqkDJHxe2xBjcPftrZuSaCwqNoMcvAKAzLRVzUrfDmbWv8VA+avIEAwz2H
FQYSVlJb73PUAqdNUZsJT0zAFCp6z7wNkTmHbW/hr4uFtdi8R0sOYyGmNTVFK2pZhKXMnuNjOUFT
o6JxmNoR4wwDweKJJf/9EgGNeHJaiuCQref9bvbT/da4QqOOd8MRjXoerlDbosR+ecO2wbTZ5rvM
Q4Hpx0sHlulER0BbvPvp/1Pg47EpaN0SVboROqNPAS94S7pnBDRvoaBiSg30iXeQ9FnWadLWc0vd
YebCvwwqc0hoJpN6ypSvj9dHvQmGnFbiCpQRyHx1wEkpwvv8YxNdzo7KGym5PORbfK6qgD9W7Jur
Q65+vP7x1oZaqAhl6kE6QMiKw2ux9fzBfyHArG821KDDka/G3mWKP85C7p2W5gLLHviM1uhJWwpt
4JPh8oJU/0fNaRyO8QZeWe7BvLtiVSRYkx89ZgR5AI6I3xOHv3lDBcvq1pIdSrSnsXJwqeh0qkYn
TYYmOg8iYCZ93iYaKZCoocVvZPPEZJAxx5ukIghUZ8wtM42RIsmwfoc61tfvnOT6Ao5dqcw71wU2
f19KCmiwoRJz/5xT0WzFXAkjEbu306YkcOf+IaMjYg02Om33aQYWWt/aPIJ41rznKqnp5x/qEjLU
8cZGRHhz69aPnI13M/eXRdblniMQFZJapiEOEh51j0BMI/LseB+meVlQIhNtm6nbCqPf+ss+fOdp
QEAcgaww25fiu1yUj+fL09G+L17uf0z+lISjXsN8HYRnqJjT/FYzsRIU6vB8EFhSWvQPDSgFZPyM
aRBdCtPucEsA8VgGmZ9IDJqpz+uyblpvO85sp1NMgdJfQOGaVUGsbE4wlqZmlQA3X1kO1B52RehE
bTA8fk+lAvqQFYc2XGTD+gdUYStjgzkz23RFcI7TyKLLXcY57OipACfiGoJlpSBKMybA2tB0lngk
RjyH+xe/5AWm6NQsG6OL4EojXOFMSoi5EIwzlnRwt5hIaoUtnIy0KOJ//AGyMa6WHVGDyQhtnqjW
/g0gmRT4VfYqqsnKAilbCe1qSiXeAn4CGlPQi+w82wneMYNzLsxXZ9aqlelpF25dqqihuQ2FCAiH
gy8SuYqZwV9ZD6nUL1hBj8IZ0yJIromoHpd0/xvDiEi3wo8hNLazNiclqxmGMIjU8byDpIIJEK9+
us3ICpBVbQy9kRnd4fTix80ENTQvA+hZ5QSXEbE0Z3NZdHR31xEKdZ2zE+Tn4jbwQoTFTi2GPpkO
O3U/XX9xSQXWTBgbH7RWA8Fsun55UDEdH4lCG/hykYx/EOA/1kDAOOBMRBWK73vRQ65jHM7eMT7N
xk9dcEne+IvdRBfVznUthiZwcUK4dJr9dlNZ3Eg7dzSxgpWkAPrjf/m72k+mNMI/mJWAd/JR6Rxy
vXLdnhbmMOJR3QdQGgABDQW+/FUawN0ZBl8MXUrQjXAHP0AFA6dMm4j5B+wQKuLhHndclDA+jN7B
5UVPkmyrPzrsjyrs1ks2vp3geuXjYcrWR/BjfoqExww+B+wtyoApd52nH80fPZThLqUX7EiSRhCJ
8F1pk05qBV3ufePPAIw2TmUUtIJI4kLyxrIQSNZxH9alz1ld8muN35qaLtKYHoPky2gQ3q+q0sYz
gI90PMUdPwU9i/zC4dHQ4TqfX+Ef+ZsCcSDXMjuzzeDujJcM3Ellamw6qmXzEIsJvanJFurGkJEd
7sEgolBdGV28IK49H9/f0UsuQJWzlmyWz2JJbkTE60CC94owUCdNR0wqzJyd83F5KvXAK/TMQnuC
gKcJPGveFK8dkYhJlkOQ3MF10vBCs8KEuumT4hZuYoin9YAjawZoLVMr65C2yO21v4cI2eq4YKH0
3gIhVSbQ/KQvvycQ5LTQUMnKk5shMlp58E0o4R5YhdJYqpZzuL54iQXLIhIK/nbvqM3Qhvbj5iOU
F6d6SM/7ADraQ11cVjCOS5iFg4h3DNVI9z5tKVBK8aTFpYCCgRy+Q82SXz9MmxsYoeNcyXH2JkkY
NIk/Lf+nz9B8tUoxHpiYKMaL0hOjOzbWhRiCh4upBhBUzEowPaYBZAbdieKKDzRBlbsi8wOGzmRJ
z1HyOMBEjCmTLxrj/sF8ggnh7YaB5aH67QdYjxUvk68DIvK8skRUzCgyMkLaKWi2VbT3TMzAQV52
BAhkNSzn/FKE3yud2CbySo0m6PfygS2tYdeilorA6sulIJeDPadNcyEwa52TAmUFQnJ+wCSUMgRT
Nu1sKpZrZUIb4oWmIGpkVcOfUIYvTyuu9yHtZZD/UshRK5077HfhIafy4yzpS8Xt/qDw2wm5TpO0
9+e9L2W9tmOzWWNPIK5r8/27QP+dzveoZ1LE6VWDtyjbxMW15gKKVWNVvlbwm7cnF9HBZ/PfzZK7
loXRlZ/JDEN/GxzcVpqxuNfdPBO5thZ+1xfS1ufsLBfSN0B6si4yr1zz41fw/M9UFWCKZCBNOJbf
6RMqGYnh/lOQ5Kh9b612epFHTLL4CIsqz1Qcuzyul9GGysfB0ZsAZWRS+kuBvfGZ3n7WogPsFV81
cPSTuBxjBZP1yWsRb4rbP80H0An2zmIz5ZV0BTG3xvwM+DUCsbvdn4LNYvFqQzGPrCI0mASNDhZ0
BtWpn7yoKRhLUayI9orYb7bPx2LHS4HcTDvjn8dJi56r0X7inr0WUmnxLzqKdNcskESvc0G8KvwX
vo48vA+NdRZFlRhnT39qOLMiljd13t2wL7FhlxnNM15+IFZv81XdVN8SI2i7cNahMr/2tlkw3D3A
5IKKm4szHVfhyWt2cVfkcvX7usIkf+QztVsn1drO4T2HA7Gh5TXbR+AM+hnRZi1OoahkBGiIkl+i
EwnZp42FEaDhwSluDSCN4q1i59OLSuEgnTzk8XuidPwS3yarInLoO2cyBn3rbDFpr6oYY+ZfcsfH
q/T1RfftzMCGdMmFpY6JIzIrXghkbRNLpgqntVe3k1c2xZDiEdS739BpMM3blvrbaP4Vpq+hlZOd
tJeaIlsGaD3r6VUglFkHdbM0fNEqTL/L1RBYP36kWF9UDbzEsT1NBCaw8Nt//LOArSrACQUWphjF
skePv48VQcpFeNPowmXUS/w8HTw4xD3n9lhyLdocxYTz5IvX9PDD3mFrlH6mvF0ruMCwyDZt/tyW
EdVc7bMnpSUfFxyVziD5Xpx13P2ZVS/32p6qcM40ltylzqNIbpQD18m4UpGXsfFwTGBCf8OZuRez
ylH5Yn+YJ6+cQhakcJe4N1v+MQj0zgxWMC9qkYfquLbrTgIFIrff5+6YYfQK/C8vlC3VPvWIb9q7
CXrzlrAXwUaLfUIIark2baisNNrXMfalgSk8NobjfUWdJWguh6EcdRtd2OkRwz/wkOnlg+TRmvcP
Qe25rFWrzjQcWIkjCEvPbXtR+7gu/9Flvj3zkE8TPPxcScAtnj6v6+IRGxnQsxDinSi/v6fUgCjV
1kvPDY93MfeoReXRqiiaQDV51LGda19kGMJFDUStihoSKS3KKXnZ7e2qqAhIMECUvRhTbivKo8j2
uCaCsggXBGb1ppzKeJHQvjMmks7YK8p2KrCBZtIfd0WOXILe6suLYVeeUd+iWTzP9k54ZWas0K28
KSSnHcKBxbtb5miEaJDdChSBxcy5dqnbS79E1+qNTvVcAAVKrh2Tr0ZNUbmYN/oejffM92F5YcmP
nZl1slDjD+6ZNWfZ/03haSciWfsxgK02uwoDtmvIlnaCkeCST5EJ3/64jSqAkxUA0p10zrXtH23m
genku0oTgWWDTCFT1XfXmFKzLXblKR2bR1LGppnETmuzo32UGqfzoSHWFip6uoevXKO1j7qgIJtl
q4laCPY8XBwA77UtYJHRIPfyttgXAaccBm0aBwVNVOImmWvqVfXEgXz04Jyo9JtOMOt/N4zdwOYt
vJnTra5p6ZmGW1U2x0z1PpT2sHzYeq4086Rxx/BM6zQoVN6/dwZBa+CTqcamUhO1XymwC9eeiCl2
ttTR1OC02tdiN7mFNEuNnMNoqVG+vWMuaNf3Sikj/aFOUHtPzTmqctGwESySRE2UFWIcCGOeaqPg
Oq3bFcQSlM9zP06plJUW9I1s+4FgXhpClzMlME5fmNVnbSVwd8h+MiT6euqi0NR4OUlaE//RBEst
VJLstBzN0HC22q56YjmqH+UWjy0cjZXEG6nguN05bLH8DRl/gRABOosDPjngUJKNUegtKjQM+Tw4
Kvpg3bYiXjuQlmY1A7CmgZjvYiavg7nTp3M26G7Qo00PVEpzk7bL83rY3M9N4Li3XTrJ4avNRRYt
++puiThbjsmwpqzH1fyBcuMQ25qjUiypgQPrTEDfIhUHv0K3q5lTgWiNiG5DxIeKPpnyWwuZ/VUj
uYxlXRUr1ssK7MW0d+0Nl/Dl9ueigqm3PbnP16iq4ON7NwLzmkWFrqCK50aj4vQdggqW2fckfnHy
VC4yfFbPX71ty0JKXkppAQwOZdhZO400iIiopYx0B3uUS/37ocUwyQw3Ym8XqRyfbcks4sPPfITT
YeHN868EkSUVHf6i9TauXIP0ug7gDL+dEdMYRF2cEsr7YsHOGhMTaXgmu2VQva1i8/qiMunTkGwl
RRSKxDstDaDlq8pfzYhTAJXemsJ+fi9q6aCA3vgsEnRMTxKq2Fc7Pblek44RKKMQ6ZwBzzJj/gDT
6mKE7lceg5Muc3wcJacuOT2ZLokn/RA5ruHV7Gp00ygKG8xWyL2119+cYfOJ91Rf+o86g7MxqGDe
WnWnv7bDYVqBavrJ5Rt7LCUcIkJL8k18xTE72r6SEhhKbtBWg6zzempjO9VDQ3S8k9QxOoHtNdSE
zQj728v0ISzcD37sB0uoGrYKg8+saYXGFJFnKN/NMfAZfUBNyx9h3gt6MklFxSWnHhRMDkx47KPX
+Hvh5txXq2yDlKUBj8dIAw+sTIKjRRyKxrda7FtJA1roCpflfp8skFhJd9dLxuRp0Ze2NMm2smgI
qYQmN15Qd0+GGa2KjUx2nttJDo2jgB2eBheYKSQftO9YJixXwizTlKi0UQA9oE4RCVQpX8r6hdAw
Kykp1eLBxUuDbyCM2uDtdKhZR02DP0Cc+boNxLu0B0d3AisCIpayMyknkV75Btl3nmM2pUlCuNpg
/BQZNvBaFokKzHqPJp+imsZEw9wGmU747YmQSPIM1NQ3uGmIfVYeMWeKF8WSPLdWxUmBm1L+TxOE
Eh63RVPrzQ0FS4XMJqbuS61lsjERd7AYEXmdozs3kc/siOCtTDHXhvdGRcvke9bY0KVje/AOWwhZ
lrzyLKdLuuk8CAsWdsmqmG0vSvQoCyDQkni/7bFKH8tOaAjXnGBMnPwXSjlmIRQb+J5KgIJOChUu
aDHIF5zXS5qnzOkhXMBU2jW2cYzPrgU9scfaARHe2g9BMBSqlWRHG8c0DC5ZN0z95u6OZ7zVfx+/
zgyqLDP0esUt/cF9ROzfaxRvCwUKCbXIJFHo9IBwzF6cujM6Py6PXFTrDWg1LTQLHKBAgBTqOiwB
nL8O441D+Nhs/bjga/R/FWkg6YUiWyNYtgC3heXkjQNlt1VKkieOvfeyltm4t2b8mb0ZrHZAxTcg
fRKxjer9OzXwXr7AvyXV23D7H3zElmfiVcnfhdsWxrdjY9yqKZEpY6khbguj7UyFKm44LZHh8BBg
AAiCsi7KLKpfLlTaNZHywBt8Gslmq1F+z1AJL43wvxnDh5P+a3uIbiJG+I38bO1NFIQHGRPNVedZ
ylIU7a6Sz8LMcf34rPOFb7HYNjrOa56zpHgjwbDFWvziCDGd4VBsTkolugPdC6PSKgikpRXbxEHh
A54gkqU43+/IGPeuWG43YpMhEK2hZCCZH8pxsKcDU0fYlc28XuMPx4Z8Sl8BN3urtEN3BJ7DDXlJ
96f84Dbw9TUNrOXK1F5s9K/qw9xJboFtKA49KmUSYtb1CWFzLi++yHk3ZILq08CSNYfOMKVP6K+8
vzCVl65pV9IgTjp4tnQJOa/YrxjRZVqtl33Ps5a6/eNXhUZBsctylHmbJ//cdLerUtrwetZvfM6q
eOju6J9JaS/+KHh0Z1RKIIi4Img2cbpMmZ8v/Q5gvNZ3L7jOPNJF5gILnvwSoeiamhtKPpaIn6Ay
06I1p0u01cdN0Vyia/gpxgj661H9g7SPj/8gHHA7Xxy/a740npshtkQ3KVvmrRb9Jb8ayjE2UzPK
g8NGGeEJ/CQvfSVrBHCSFKW8XzeYqRR7T7a7BgGdz/Y/pfbq1O9cNdiiuIGSpj5asUcSC7FL/GF0
AHYtVS2xZ4hZ7kgG34ndwNi8kIcUz1FrknylrAeII4yQdvGZBCVvc5M1lj29CeXThNX3+iShjGEC
mpY07GNhuYyKFtFAOyySvI7mmu+FimDUexMBo3ihpQkMmuCXV1Osk8u2wyG4whJHnk7V1m3bM8qc
37Qrlfaw7Gt4Kq9A5SvM/KjFr4732c5FU5OoZGQxWMI4h6/Tp+9jFovcP048Q0KKdVobu1IQPM1K
qj9vo/oSczmA64MELloh9QSIsto3cNR5GYqndH5UvRPuZ7sAYXIiPgfsLiY5aj1mj/PgSmN62FBe
+LiMkE6tS96y0J24+YroauRkHljD5e8S+Y3K4DPJJ1D6A8MeEV1wJd9HDasEDAX0HppFGhGu7maB
vwHCbaeHsTASiYfAlULWm26XBG8ha56P43khnLah5hbPe0Sp+dJXZruJc8eBc6qpvT+lf4fIHkVi
25bASRBM8EFRywhwOx2RA7/hW3fj2+bDCZhQeOa50U9Kai3S05BLyCEP8xOMmC+9VFL5n0WCq/Pr
1YOYSIITlxpuP+uI89sNLWogLKS1z5jnJmshnKF9tQ6CkdoIH9w7j1LZtPEa1uCCkBCp/+WqzUat
+DfPmYUAovRlc20Sh+yVMG79RUolKAgAf7xWaY0RppdCrLY5z2Wc/v+TuZLSQBFpG9SiieVsrX+r
b+bnuniuMMoL/Ci1hp8pt6d4uZy4XW0OQd6gO9vjy61KLiLAndKTWKQEZOxZ6ZJtoGjzzGNN5PIB
iJJalwhhD/jss4vevwPE7wZcMO9m6GsIrTpBdoB4ag+jVZ+O7yMYG9dGoYUO5kpLRUUePRMI+Vl3
C6TE14KNZOL394abTypMow3QAUuPVs2n5krP1XE0wz137TQVICFPMgkKAGPjT3aKiLpI3WC4dnOr
mdf2MYTUlvFEOUAk1cIKq2NTHJY16DfOPR28apN8hVfhJ/E4iaCt9+pZ2gctkeAdu0FdC73+BZYt
T3EW4k5VQEw8O3zY73gNMOXVe/RMfV078VFSIJ69DiPd6mMzek18c+8UpWu6pVsOjQPmZawx0iuH
5c1CaKZg6bW1t4oXSQaiuSA7564j0WxxpVLr7uas2Jgsipc6Fw+OScsgz2tImVX1XNf01Wi7ZjsT
NiJ8X08SowPZp7AunxEzhAusB7CQQy7OK5OmZOBm/eoAVWfF4Hr87byD+hhGG6qnSd3gPCAt5KoK
/ME8/slgx3L0JKgkx9YGITXRBSIZvE+fatC2lAT3tIgagd564JWo4hGjXTQmDpCmJuKr/fX/w6W9
RzQfT8X3XXR0uNbv2Zwx9dCJpLoJW9ktAq8rxJtVTG11qhrcz4oYrg1qyTofyUI382oGqJJ/7erc
/f2gC1hHwbHqsC57gbczkOOimOb0TGpgePhV6xtzQLPNXQzSpdO0jlTw+576xABdFyWj4zkJ6ufI
dcwEVdojlUWJy+/KSbeYIae4V+QHtKzhQn3WW4HEjlw8d7LmpsJL8B2HQjjCKuZFlVK71nHOz0Da
ekyBFs6cjXKUjE03Lj7+eHdYWulOwdYQErP09jLKZu+WlQcTqrhaRa9o2Y+mkf2YM9rL7Lh+hEii
bSgcYIELDWNUKreHqbNByTEeUBmRR68vGcACdIyZE+zsI8jXN746qz70QIhfcfPV0GkzcqVL2nHg
1deX+oGZizDhz7JxcurFeypacQ3F2u4S18yMrUNgCJhdJDlNdaxaH8ISho5SWouXujQGtntLBkrk
ZjzLryOZycf24Qu+2K4ABZcAiCOTFtE809W3xgQtO8yLCwjTb5652OA2KOZIvil1Jupkdm9D1dP1
HIIpKC8mOObARsgwUUdwVCiLd+qvP5ZHMcqA//mWNvZ+y17BDrc/5fHoiXZ68Ykia8gRUc9p1cE/
Wq538aDqTfvRAepVdrOc3fKiPotTgj+DLZQy+7/+/7dA+YXXSFoBrkZa+4sx3FZFzaitKUMycfil
t9TI+tmq2Vnf4tPkrIJe9TAu4S5EmZUNqpWEMWQoqjy0lUn8080G8wih51YNZm+W5DfvdgxB9Lj8
w/np8S5lsVHymmfxGFoslNh/nlqS1o4pOOWQtYmXDaFhFSNpI/MoFWse8EymCpDPSMraSDUMXh9w
LF0J0G/UnHM0ThM4jOs8/yb4lLr/YAJT1aJDNpB7kfsxvvQFIAFGs4BStXeHCnXkIsm0Thw0qSCL
1sDLX11g8b6IQhQp5MrapZdL6T0g2C/QTTRaeQFpQB5AnWvBP1ITUmiCoFQE4knS8y9T7iaG44xT
UQ/TQ0VjDkGY4PQPvkgcNQapv9TQPwplU75G7wotv5jQN9UKOXbT6cIkUVOWB//CW4GFGKZXa1+z
lcmzM5iSP4k20Iojd1K1crZ4S/dwRGFR9bBcD/plTIUVxRL3SCIiK3WPBqoXGn6Qm5DHzgQHhmgn
FOVfvUokKjA16AdTA1pukTf7WL8hO4LN6kkHfoQupPdcQ2RxL75v2zl2WJbVBCzHI2J5VuUIyrSm
XaR4X2QVwHeP7iNEzB5CMXaNnhkl0rZQSj8B35ROBBZM+TnFFI4aSt4W4IV0iruBiOoWTFWsMslI
3l+qZ5TOWAmZ5rc72+sfUW+TUIrCQJ/QNpyErg2yslakosdid0GLUHj6tU5tEeqBOgCNcfqFThzc
BoXNBNEkTdoFRnV/4WJ3j7fn6W/KAxvIHdh5NeBfyWrgprJz8u+yv82MYm8ghwrPJy0snmRyomM7
hJrk9pEwFasaXjk6PDM/W0PvUjhrpCsUXgV53NJeXEYQ2vzMQyGgMmvUHmGBuzoKSgXmZCmtlBef
es8GOutWRaLmE+m6sWgoREcuza0S5FHDGc92Pz0dwTPOXTntF/tPORDFUkdFHQWOVYF5sLoFQkSj
uhE6i+zeBYOXqe+EFZfp/ie3e1o6X9vNurPExEkjtp0iXgRaj7VYK9VfvKtfNgyyM4r2+xv6E/Uj
wG1dHj693k4/qpbvPJHAyiChUmnkEwryr2KnImXkUxdsUN7fadX6ZUHcBcMGrX4TbPibkd3pLfd3
w5/eJ3KWtuL/QcBtBMAoAqtVTYY0h5YS1IFiQRch66FZHEXiqNYn+2Qx7bD9Jp4aa3fG5nCTdB4D
jdtXj2zQLivvt7DIiuoQjRDiJ0PuwA71+fxZRBMMFp65r67rKVxP50lp5ZOltPwSfDsPCLMjcIZG
kpQYT/sAuou6j3KDzbwGR319sVUNzEAPfehVopVevE3W4ycCx7nXTBQOeuiyRpsuScmTj+x2m/7W
fdA0R/DerdlGXeYx86vrsq26InxudbjumiLo2O/xHHbtjqp/mPlQCYUzczqw67d/sxf+JIbJ/MIg
/gsRhKWHFIIXCPUZVKlvVgUI7V+ZYIcqp21In8aWihsYVQD4ci1qU7Co+x+LXMKsHQwB0RNbc9/f
tMUxuG3E91Hdw0s5hoTn5mTunBgmp7GWgtRrW7blzAWlhg6V0ObWZr6zPGxEl4xOUFlWtYwHbruT
//dsKcUla4kXpp4jv//v4t7RrTsTvjbMuLG0ZRUkMZMIDylwDvZSek+zsMvRQi1HuXwkFJpo9WEV
dvP6EpLlXhi9TZp1OPqlmHVYJI49jTUb678zvaS2xSwFXeAw6dEaRg9y84Bk9B/gKtMivf/Zgw1h
Ms2GrocHTEs+6caP+x7khOetVwQiA+gimGJAf9/20q7v9rja5sfg4W0NGpPbumoQS/7PJtQPQGGq
w55FdYOXyFQfu1B7X2PkUwLdzyEtPa61A6dPQ+fZlSH82pKRKydA6L/OJrwNtQhZryuMP2HRkOQm
OFDCgvZQMPTmGQai2nq5H7M8wy1KZsnNBKG0v8QQHHgiaClnIZRzzJ5cHzGaecOxZZVz8JrFLr0Y
jTN4MLRWSSdJh2tsaovENNZ2d4IytsBolZGPaZYODfNnPUg0eSGetlKyB7WFOq2eeVjfnMJI/SqY
4W8qeClJZ7D68WzQs7YtzzG5SQKFccdxQDRPnu/F+Zq25noSaLk41y9jklkL32OC+bR50nL50JA9
xhXEBhNTjg5YzzsFS1aXQFl0CamEmVMbXHt+7ACFidFSVV8l+ehdgbcfXwPO1r6XgUtLhFvrTKzQ
1ROn9Z5OjMm/kpkXCKywN5tZwOM5eIBcEGLjZdOPcT+ir0/3RtfI7dZ1HXNdcjCJV2feUraJRDgT
ynJoUBWzsvKltTaUHL2Nu1PV+7Gzy+d0cYZW+ULPWccUHSqZeOxIW2d7D7xa3uLppC4RKatXadFg
cTH8F9mJiEX7GfkB1/DE4d3jCYt0cACfIsmxoFmhGKjPZzOnzOIc0aZRWNXnOVHsGU9fwBl/+Yr9
VH4sDZkq49CJQX4lo+75yQvprgeu6M/3svyf3lfcwjkBhhyAtgwUfP+6y2naTw5bTfnz+DOit+jP
jjBxu2/bmQbaldS7Slwo0pomTP3yrEuug+AwpEBYVHuOYJl/QJyhIwGDogOJF5ype4/37Dji8Fu7
RZI1yQ27Gd7Ucq9LEgfiKxvlf2zmRP+OPRe2ie13H0f7GceeXfbi4Qf6hozc8SAP4Fsp93v7/DAg
wk31KGVXNpAiagvwqhD10icruaSRU4cgxXZ8RR2/VC0wkl2nr3dqX+d68ravTwrJ4JJHPqeWy1et
/wtofV6SkEyBla52MITNcJJlhNdXkJ9z/G5yaR/NM/Ztek0l1FYhLJhQ2FC+2aNXtRGl6DwNXIrx
zAm7o5rhzk26c81saV1EPIzClUzk7SNWYmauLF4AEEXq+qoRmBwPgxiqsp4qVS5v+UyWvODrY2QV
FfMGgVfIImiCsqpQcafATrnBCl/BE/Ps94CPkrPdX6fwSzn8yyraf6qcj3IlIsf86m4IB/dT5eu0
HdkNi8SFY+vzp6r/t1AaVcfMVGjwIrbhphXhCy3++7nzdF7PgCq7/RSZI0yFEoDovLWVPdVwXczH
+c4Nb8+UWzoP28ObgfRL++qnesPFOvdV+/TXgeSIY4UVGF5noYVCCOEmoqSpcNYPB7AVqaXUXT1b
pUoARwbkVvxTV5BN8oCjfTCgOIzWia+M3N9uhWPer04vFkqlc592wPn8MIUTxkUh6OsH1VRbQj4x
49694+UWnG2p6bLYK7uL/R2MTFFI/GkoUSawTrkulYCOMiQPfM23hJ46i2yDVU3VjKo3sTO3Zokq
BJ0+or2lLqamQMN+DZFDXbUIcYW9OLFejCx99ApV2+eFRWso19s8Bv/fgugvp8rT6swYaaiF8x1h
prQ6vMHUwjmN0H1JlEsVOyr1ayzvfcbYIERzLXnVGlfqGL+j0OMczReBKfApR5Cy7LRNezYO4Gzw
St5E/YEwcQ04Vny7Benx0ooMOOjZKjAvnkiDG6NVOzX9OVi7oV8LphOeSLCIh2FzXDv7u3qfnIYy
BB/c8L0DPK0qH4RkXGsPj3lqh6uox96Tk0ICZdaVld7Ml0iYVJOQ/a+fYh4a4u4XFjBvIe7sANcP
0a8OS2M57NAi04mRGbCc62A5Jk0BRmNfQaRwSY0TPBspMTxfohveG28dulB8wP8Ggi2IjMj1j1+f
jNXi2dmE7DLMHZdvKDxQ4FaDheduthtSsmj7bznLi7MBs2tnZgEaTi9p8AgNIZX1UMqXQcItV7JH
f3VHqFfxhZyqWIoK0bAc3m28EE0oT8qqLqLhuc7PrMVYXH/LPPfpV5vMAER/O1394JIoSwU+J1XC
oYF48GM4gMdvN7Y6++4tcdiKK3UlxQPPw9Ea4DIVYTq8oR4EFIsKJawSgzVJjq4obDUe1fqqrBY1
8M8d6Is9JB/rBGva4m+AfTbtZh7nfeyEhQt9jujat3Nw0Y+NR6NQSQ6my1w1n9GBgLjvYo2fWR/l
UrKoshZOZ4wV5rrZBVIHWLyUCrErab+whNnC/4WsFOXEh3godocm35xXErZKWqd4qoIoDRiXynjA
mL4zjUMgG0EGtYuPeUBiZNbiE4ZOORkKwIiyylh71h/bj0Q2XnkFOugpyB7EmNkBaEdp/yar6M0d
w4s5kUljlXqiuXzSIVxClaljkoEEy+oBuSiVE6Nhx580klg4ZI2fhYrashKupBphBje2bmzSyrYb
I3vzC3qwm1ZPYWclEo2Zsjce6V0r/a4JRFSuuMD6y2n3XLQrXT8sfPoQghAHZ5lvGyEmHlWHlIvw
mwCTaZwd+8xsfEzi76ewjXCuV/GHGQhlgX3yauRZM6hVwyIWNi3pn+2uUXNvs21spwUoeIihDxbt
xajqVpnibtqEWR7mw0O2Iw9lrG8sRQBAwkeVxz6djyiUxhbX1qlP52D4LpPqStB4OdjmODMCZIXR
6aNZS4rI+z0R+UOnf5ni5jHX7M/L32SX7tuIcL22WgjDDWfUOfqBfp1rv9qG1efJBevSEbYDexWP
oAYgiHXas0a26JG8f8f768a+weoPidxza/YkvOOzqU6/ZP7xfci+FKeAYqSwmsumQEmp/Vtyl2xq
wahuFrNrnlinIrYG5YV0HaQTT3En+r+xpXNG3B5tosEAe21n02An5wcMGzZ+OIZhReECyB4EqxJs
0Nzj/k/4IkxocvHQel8PkWD2WgXr9UgE7sXnnUaveuG9zwZTMUZxGxQvcYRaMAC0pgdZN9AoEabu
nRmS8t6L2MX0RaJZYWHvwbNAFeYGzm7PBcLS3IkX+vrVEDxz2qpzOY+d02bwxterV8ITQbhxix7u
S5RyPF/dcq0AK1wgpMG980Esdw+A3e682y8C/4LYTdLyViomxMn6OHNXo6Y+7l+eTNA3JvUzE2r7
1ck4jML9Nt489UNQFPXoWumDyqlW65ZbIyc5XIssMiFGu5GrqwtPQUB2zkrLoR0wbD3cIujJMmM/
0LUakvywxJjYJJibjAuZrZk/a/hHJE5Fvh5zMGVPPB7lGSfHS3d5cmCHX0YnfIwOKShGDiPUYlU+
b5CTzYHLgsOFsqlTq8gy5qf2AWq8ixAvAO472/jiQm8oyP9qJkS7PcWmsm0myLZXIz/XW4Zg6doI
TIxS8I3NvPTguRdJ6xObcIswmYcn4BPYm9j+dZGKj9h+5BgSaGc3b3K99CPL+SZ2JFG4OkJdryyA
lkK8fh8DOzoBHgQXOPFJ4iSvUL62AYp7Ze9WFhvuzyA+p8j/FcGBiVB0ePEFVXOFyNXXivg2Mcy6
DrxJmJ4TC5ieh6yIzRN5V2cc9ZEguSrhY16masVb5A1XSGKwypTGlPnYCzpoBvi82qlOMKnYJ70d
fi687XrNHkSMTApMMOha8Bot5B0amI0m9wbW4p8ZfC+hMXv0q+SkBe3uuw66WIhZFUH761vvMK9Z
UrECimqjX/qG204F8Roe4viimARBP8dQmk0r6YHQTAswjCSo35mrLYuQrVRiQe+t8LUGmqlknJIG
keYs23XhmMt4jZSfwHNjp2z7QmeBfQuhP4BdxLxQMjyoURGOpP7SI0qqi5q5womvjut09s7i9z3n
VngQPfe/8YvJ+KEKreqdErEuGmuzacxQGhfdrelrsPObmz0dkRG/X9aXdoFJvWu3OnodETTikPem
qAuttbo/ohds0rzmbDDkwofECQa0s8N0c3PEpFltgW0G1A40fIbP1URDA3qYOVGdiSgZJKr7ow6U
M/0fMAqbIu4DAUq4Um93Z0ktEmWuKMUzeWrMPxTesBxQ55NLSMrC3vQD9jhNsV0W3Se0Xc1QTVqp
nWml8jCBpK4XgbJYwFiybk60/x6pnTxL1nil3ayM7ELD+Sxsn512Pk1Kv1pJsHuuK2/117l3xRE8
KXCcl05xmuxKtxNX0woYJbOqx8W2OySsBEbOpRWCzHPMz8pPIeb7vc0tMQZxI4yFnXvHCohiDk9e
l17zpyRiMd9k+vgYzKoFos94CLgRmqnNwLwwgpaOES7oepONWjcm/BfDdS4IDQqVQG2fvv3L1e3E
p1e1pia6mNHc44/xkNjadDK98o6kNDd4mTRZ7vg5zsoVTk79z7T9PTwLc3AnG62IHjVx4VNmdSn1
oMY73R+2Ceu0+1o0CXFmA5CWohTjsSU17y8swrzCcPX1sKyBXaN4tvsibwvoSqUfGhO/nwdhnih/
9yCo7AdeNmVGUfGoYhXyLT2YOq6pJtYX5prvyYOj/QmpQrqL+RsdOKiysJkmI4u8Iy0TkSeREa/z
WPxbQpgwE+39lMnAkO4FMvlknv7pcn8NZvg3nZH0ciV3DFEJhRrcU3epA4WQx0V6t/8YOzhxzFO5
SIjuF0STdQzuvZySgZlyO05J2UYQm2lC76lWW6Hw34+kRqjXXwTISZnkV4WqN0WJXYJjttIircB7
uw2SBr2YXbHXIQ6c+KxdFiH356EQI2izJUX6K/wwXrk8qKmZuxvAbWqrRZ4LDpF1byPWa18n2UQN
VmsojzNC0JRZ8SiczngpCxxK35f1En6hXaxLR6BdEC23w51Xp4+7ZG5cebqez5cU8bTItEUhbchY
T2bMeHk4WbMia01jBG0PkC+cwrc6DZNpy+V9I2CJzCCpSkTiCeD1muia5wXrMTTctYMbtVjUUwio
VEMgzIO40/VOQPd+dawGi+/A4Gg7PJCF0foApkMwB7M3pFz8yxPTSMurNVup1vKW1cXUoLbj/r3k
tpFJJTIpUwvjkBNj3nq1A4uKeeCPyxoZexluRH/jjEgbRZVF2wsbypd4xOR6GMUKmW3VhI4lwAat
sSqh4M4dMoJBLFG9E4Vm3D6ywV62iLSHwVAplXP7Oml9yOyh/HKdiLaZL/FzEwCVcmu1hxx/Cgs1
+H7ruTP3FmuAIs2q3ZAS+vw4KTo7WJKlb7Y3NMMih0HBfFfAdflA4vJ3v/ROyp5TSDnUT8f24wIc
IjqAhvqq0XlJ/KZEDhpiaYTCvNifrOWUJBUkOZkrwNmp8W/pBf/3EpIRXYnJg7cTxc7yyYs+c+UE
UWs6McoO0vR9p9oLOtK6UpaZAfc96bAyF4hlm/L+AKKwuyV3UttbevP6dwIgiE/YT7siI26ziQg1
C85VLV4dnwpVSGw2Ei5INjau40x4DJ7Agzclvh2d006XEC1TR5uvCoy0sUZHAHA5QctDyfUHom2q
gBoGiPpnZXDTnbE9rcTFs0W3cxhA8CHegleekA1irQ35mCH08FDPDh1zB/XQn1/B4tmNNT/FV5Ox
lKiPruQaJ64G/R7vHyEZ4AU45Zk21RP2r1ES5CQXTHg91yKmxp6fZJAmPooD9hun4Uo4S/pqn95V
4sMQlqPcAJVDHiJr2CEY658dxyrMunCF3Ae4NWB7VqYaPVEMSc8e1LLoz0amot8kDKGsIZL5aheb
fQ34Upc5YjQh3LzmrJ/u2zHsyG2bQS6eZqrB/iw2yUTsHDtpg8uiurydX5XUrGMgg7imEDvgX2af
gvDW4eUuzFrJ2Z1AZJDEfijgsPlLlzEzQ3KyaUyWo4ZNRjMInloTPTZs4RPkAfK5bhYP+wgj4fIO
kIaKtLMmgE0tY5Riy57SUX39CIEFtGuH0h60jZnxLGZFUb1wJz3+QJl5Spi4XrSEJeWEQ/cAWzCR
LheHLHgRBojGUONeBPvu7ncMwk9APjFlG89jSWwHWSQcy/6KhcHApBtFjP/WM2iFnu/ITJwezgOA
VTFKtIc18lrNj/jBDa/D+jYqoV8RDJx4F19ChOD2o6PKrG8b+Qqyffpuga8shdZfC+tdvDWZZK8E
XULnXcpZE7vv4XJTHpEAb+7Q31XKhHjO2hab15Q1Pu00k5TF9xarFbznaoh8uG6eKQSZcvj12RNd
VgnNHZ/nHqJL/FtCrdAoB3jdq7xRjlEAi6HTH6vY7L/w6Pb2PDqPCFglM/+m6ENc+k3uVUlfqVVp
Yu6Zp13cr2WbOKKNvI0SMOdl9CNq40F6YOiT2duLbypwlLJ7NR108o/PcBX4fxUpPXdi7WRwcnpA
P3EGQV7Y3unoC9yQru0lvTA4JIyZffeSsB4AhRTUH0neE3qSK+66lCld3jB/xhoLjmQaDYQ5spXU
jIgvPhP5ge2Xz+LGP9QMVoveax/w4xyZwo9QiZlwmzZcgWKmOwcgJzdRPMUM9R6UtwhkO5fvr4Q1
RCvA22ILBL4HxGstgKHzxmGm2npVO5A0bfUMd6St8nbZFxgEwYkKXtnF/TKVZkkDUqf9yYU8k6JK
c6CqRgQaJ8FZy0xHqHUk0agGs8Vpx+3p8mWMQpTP4QkqsOIA0ZQS3O/xvREpZjbIsNPXc3Roo8bX
rFinXjhwjniQQcXvlz9yjvyU4nlCCxzvHDlzwIAe4g8lkQALkttbyAVjfQxhkfHaXoiAVeUc0iXp
1WfIc1skxzblHl2vQ2NHw8kiGjC88C12hYYSDtoTXyOIkYvFhxSLqfhdlGw7+CNVevdUF5jPH1SD
SdBwOnXY/tPalRRaWC/89prNDKxUcF+diiBlH3/N58R+edDt+ZhtdEfSuF84PASNcL14mePwEybn
ZMNhwbE/SaLF/DhsuZZqg0F7bXwmdv0YOBRVdPNIRKHXHMHTdCu94SVrpzjdo8YUE6NOUh7BFi+J
g3J4oVocTLgrj9f77dW9Q14hS0LuIuiVCt4Oi84Oh0CVlFqkyaiqYqUKK+hLLxmmHTNfwXcUb4Dt
s4cTtR8TXtSgsiSHOs8AmqNJrojxEKOXaBJmcgIdKzx9XlH8Xonosxwopr5y/QyO+URWe3Xyj76j
J2Hiw2Z0zNAtBs6IiMGNEaVf++3YesKwm9AKgnC7/xhqpdJAzgU1Tow5uKQ9EeKEwRaNuN/4rhug
HgWPSzZ52/A7SmxMGo9Ee24Vwfbhcc4KqJjr7dAohZYgRA2WuZboUvEWNSC3zm4+VcL8VJnXKSQv
ACL+TnowYGhyi3JqE4JnxQciWlJN8pAPePdLT7Nu4c4LJl3/zG95t4+i92npmskpfbDEHUFMKIkw
p53kvcTODMIGNlnZLSIzPzWuKKrp3NE+XkbXJgF3RUUtj7i/ZLD4o9jglEDYcUew0RHJKn3Ejy/K
guKw69fEhcu4hPNypj66jC3uQgjHfB23WmLCeNh5gBPb9RDnzqX6YlaQTwv///4lDAQILcDa6BTm
zoJdioYEXz8x4/iGvcnj8rGT40+LVkZzHf3Rq92Jx8TKteq5GiOxTNSMOMDG193LhyJ/YzLrweUF
bIgyAHkG/ZjIidLFVDh5c16q1hMUFi26itdKpKVQSQW0WB+m9K53QfLn9UMqLGlTIsUXynUmeH6K
Eim+b+RoRHhOrYO3YeAQf6mc1UQhLpwn//bFLj9i6FWzM/tsLIYR0tL8u+94FPl0ubnPaEum83OB
U+T+cW3LDscxNm0NldUtdUgwVChryhnuTHqm/uYQuJwgdqM0SXESoQ8MrZui7Eml7s43wmJgDpsO
4iILMr8cfaJlPaX6d3Gll3EkVUNpZHG0xh75JdrLIu8h5YEr4hGbN2lI7x5wXZRi+lWDsYXeYErI
mm8EtDgKsU/WbHebwV/GjT/D2uTZXt6ajpxkOsBNMla6ES3PfpSxnTM+OUkG6skYglTiWVcSk+Yt
I4o+Ypnzd48sf2kMQtupQYTSZ9LCYEyaWcOKBZaJOBmhfrle6XnKAtwR/NqreK3tmthnKxMD/DBm
t4Hi2KXE94aACTli5zN71J4GmOQ6VZhqAXZLXoBKXBl/NLuXADE1ae+EtUYpoi7HnkukeUEy3wCG
vLnxJklDWPdJShZllgDWmWPwSjRdlos9gRYALPlnig3qmRLvvTWs14SonyOqymyKftpaD7y3r3vh
XrdJfOt6Z/3aWBTyOXsTfVbN0G4lwYAuSaDU8u+h2kFCuOJZ7fQcMbZLs0ZjBnuEsklOmChsqXAD
a6CuuDWsDYi9TrvxgR/46naii2sziH31vR58wPj2Ma7S47oNojEHbZKDlhUVDhiaazgFApjK93oR
Ia7K667wf53RWIZssSzVPB102tfsY5cTyYSfjwkLkvJj/U8tBgxEHgxEAZijEtcwNvpAlqloaZe3
wqYSFoFM/i+kcc4mmaTwPXeeJ/vH0BM5bIgpYzDC6pBcsAckoKL4tlVvMnGHzqbUu8bxjx4oIaOI
BN+HYYwm5IjPeNvHl86iOUi5QgwLCinbdzhvHhkJfcxxKCLzCES3CXr55zpb88y55veuv1rEBjXY
79lBrTXMeQQWOtV8EQz2kjmBDm0GNlqHzknEHJ5VqSRV+wSTlIvxXAloCgs2prmU8Pt1I0RBrzCa
8ui+QZxEzUaVn559jfoHvHpHnbUPLbcOoQ+lGUDqFSlPR3xGK2cNMgRcSduSpXs2tFGGDsoynFTZ
K/X8H9ONnfbu/Ce2+HJ+0PCxzvVZwiyZsKKGfx2VFt/WoDldTXDvfbfyYTbX4zdYrkNK1+YMxzGM
lx1Y4d3PXtyLQ5duE/axNXdrUFZySWlZRVzhOdGH0no3Jvr2BohsNIGn+9qMLLCzp6l+Kmg0bbR8
DKr3hDdhsHwVyK+51X1NCiADpMhXShs0mXroh7SG4nvjyG9Nd1CPbDnRjt4+5XWO9cwYYg/CLVMd
g+4lihsgOlCiOYEWW1TdVjDArnLeirnJzGBUKoTsdTCyByf+/sE8VwpGRzXfi9xyll41lB1lMVAO
6kVwjEQHvAhWuArZtKjNdK2vy28ZZ7QdxGRC+5xvDC98GkVvTfCKTSSZWf/ccwmCU+77JH6QqI8x
2UUg/N67ProzdGIFaH1et3qaom3mzayUpG5BeRnWf3JR0GAhr3Hd4E6cgBcBUVR8wHqN/B6pzv4w
jYlL1cdQjOVCgBdWwKsk2R0wS60Xhpc818UNUN41LX8SJ3z0MVMvL6Bnl12o6jcYuDvDO6fusXCn
epW5rB40VRgtVY6D0Ausp67vp3j282JkDtDl1poo+HJB6tzy5Bn4Jc39QTytKofUt8StYZwIyQHh
B6v3h66psGdo2TtqqQ6/lApkergWWL/mhBmndONDxiWQHPNbu83gQycuAK2i+kt6Hhv6seQDbyxW
zgbjaR+h93/onNJa3Ra2K2h4CUezLeU2dzgz2qVuowICTltgggeJ1XNvc+UD8A5SOPPkv1XhLnNy
eU3FgUFMvxbzcFqxYyq8sfDtDbu+SGyQRS7ZIPFjncvQPrLH/pKX/cVRkHPtNdMgG60yyJJtpswN
TWf1RAGwzP3XtRym/9vJUjRjeTwwNQ+TMmTvyHyohrhaoBAHF7U0urMu5UGL933qyRxPtevoWf6N
DyDv2OtY8W0ezEnDN3zP9aIWjYyq6EMHihOd4GEMRjx9KatCy2BihNbMECk8jHqy5CWQXM4fMQIw
jqhjPh8HwT/TTUOJJdhcg3JqvIBsDIbZKxHOmLRTVc/lTZF4QK66WBZRbxBgRgoiWjFbF5S3W34R
Nu5Si+FA8wNN6AU7LXnMK7S5C6YncwhZDzlA1hk/mHTHprRNJeElyR+m3+8lZ8EBNNBArI+niv2x
8HG9bVp6bILYpLJ9rXjI/Frhi1SxvWYsgKnEtJ4ihlRwfLYz6zvy58cv7NwNbaUsuaD8D1lVWu8X
+3uWLPW5v6bZ7XQU0EKrPiCvea9zekepX3tZ2gyArYCxibhM8hZtslCFy0VasdXY9xPdBqtgmoNd
+ThtIuzh/WGj9LTNq0aKlCgdFZb4tMsawEae+PDHZArW4I6DH0V8TD14Dhc/bJAuTqPXUsmrhvNs
L91u8lXzn3GRxWyR+qdS6utMZx0rpgtXAAqZSx/icE3N9eAoRQBzpzQumIl78F2mkiQcRtfHuI+c
gCtTR4PwQGYlpjQWRTa1K9nQtLU9NkrNNYqQLRR/HpyS0cpRrcHuZUANIRYoo7ssDJCxrU2QDxFW
QBaTtqJbwCyyXKOb5a4nNX1aTSwYprrGk839ImJFoHy2Z4rvsOn8zERNQ5MIGhcTZsqoa0ZjSCWo
b1e29Jyq3l+7YfKMQdGliZSLhFP7HCuCuiCV9c0gu/9PErP38m2cfjZXKn6F9MXg9BVy8cmf9qn3
gjmM4yvQ7F9mFCax9HK8FMSZ0K+ANFUdSMva7rKroctXjDLd7F+MD3nOfJLe3xhYJJuEYq031JeT
gQwgOW0r8TPf4KqCNKi7JjowhM9rk+JYRT964BI6WjLyILaNsmpai/zJ7ARtNHVUxCPyRIJn+8Eb
JYzns/7zmJlWmv460fcdABLChomFGM09pEIHxltNEUrNU0C5g7yXpgoAfrs52DsCDHCLTagoKVb6
DD7Ozjh25GuuuoYOCCvZTFpUrmKTf72qkxmbbtnWKFXnJLPEk0P64MOHSPpPlX/7R8TFr9Pz4E4c
62OsA8affCwVXMBQAnV/czFUX/9w1ThtWdLxgajrKMYJ/q9PXFYJG0TXP47NO/0cmuKF8Lq6uxal
VxCXUB2mv3XNASSVeCYVUBhHev/fQnk2NciEEQictzXoqqrSvaalVWeWqBJtWAEQY7baWfdIRoHs
ySjYf3K/CmbpN1zZzmrukDgwvxH/zBL1y2DGanJa6jiMe9cTBok3wXuQ0dtPr0zS+UsWg3YSjg1T
6V+d6qJ5kHwFXNzJBns0M9+r/nLBANoYdw4AVzfHc4dW9cuTDCIdBnp4Ji6MvBwuHwi7apmW8E/Y
P9G9pytQJsYEbaYgrGpWpHXDcLQIhnqWrT5e+Dwllny+nsmggLrWb8RcC9vvnpr/fGU/vUbuYtdT
nvfsh54YHOEfURTxe/jVZftBf8FKNG1sRbCnNYQXgkU+bx+ByVoKBaHccqRzGbTYcU5ggFafx1Dx
DsUCOb2wKkG5ks/ds8nguQuNEQ01UYvXvJ4PmdPLkHNj8pg/3OtrHQ/14jSQIVd5/eAET+FqB50R
D15i5oYwt4f1JIsl2vQXc5Ui6mCAWCKYwCkXtB7L/OjaWWN0P5zLtqur3X1p5SzNfgye7Wf0qotu
WmwWfqKHM1bbn9Flmf65sOdF4ZwSogP+iOREeyptQgYhqanOmkQRcSCCSNRuL4HaAHc0w+JjbfVl
maYFyzwWYAxS2ruoLBhk4opo5ApMbj/hpCPU0fgjC99uCZFhhJ9CTVdQvoF1slQIqNcVxxpey/8f
ntXcwi3AA+xWl2ZYI49YZYS5NoFa6efAOXOUGoEC5PSFFarAO9YntPBKtDRjuZx1L7P3WWZKPbPE
jUEcqO6Z0qo6AZXNhd4joFVWMMcRiNw2havHNzojHhubNnEO+ASW7vcSFmLJAeEOSFg4y2XVMuRw
5BCqtufqR+IgyJ44w9mG8ZEvJr41OCL43dhzh80etk0yKNsI2d9W6lU816CNiUjsNWbyu3U+Hnbq
lli+N1T2H1wxUKCCYDL0m2SS8km9iETujQqqPVIvCn698216vPYxxpfmcr30XwhsuCkMwzeX3EE5
NNLiDciOiO6K0cUWuCqUngV8e9RQJG6dcmfkU3E2rtiyVdmtSzxs15KKSCZ9nA0RkG6rmkIEttWH
2Mk3lBwAfzOaG9A4G8PoIdNKP4q6YfXRByY8+t43yDuz01dIxWN4E4RmpsGtZQKeoUUJzItoBakZ
z20U2OkvCww+m6DyjX/V9mZcdvrUeAHrE6xurlCxFEtL1TsCsgor7CzUsUdwesDB1q43uzECgLst
iMKfv5Jhv81e1ZvlyYLNj2l/dOHMx7kZiXeDYgNZLOqwrAG7W5bgS7mZGyfI7k/WXr4bX6FA1771
B2gGBW5//U+9I/GeWHXCVMMZ/ad3GHyfzKz/s8dVb/Zo207CKc1MtNr0l8aHTRPIIKC/KlIKwsow
cg8VI1fdzSMcn9sWZFBfp0e3mdJFppH0I2E2Xlrfkl10Wb72u7XAT4VdRnQlCUpru0SakO/2rWKF
ix+F/GbCg/phEryCI5FlTjevr8dYPFKHOA06fH8uj2ZA9/YCergmaXIoLnSGo+dKKh/8pt9ODrHe
ep02IrUOwoKF/vEQ3mK4dFvL9CnVaIabfE3ii5Cw9IK3eF1XGMlQycz5JE971fncnVIqg1fs/D9S
aFrz55ydyElboX6IRdULNS8zAtOmppvfT5PXdO9Q5gCL7h1lEDnicSSUSmpdIA/ScFmeQQ4CL5W1
gS3L8rcOZMcophMFLP6jpIXz7vLv38Qj3jg5lS1R4uBnCDWF11yRHb9Rolcv0O75Bja/Lk/tIn2+
jYgNfdwROqEacf8KsanidnwC08icCP1mJlmD3x4zMmrSHbTYHwVFqShSGXlZLLvfxCg7hxoA979o
onjZsTT2JSQUF2SKTkPU0lJxRvod7KAhiBGC2nhtwTTktgTpKMT7mwX6h7nCb7eVlnDmsbXaTaHy
YGuGCmJKtUBSe3dM1mILeCKygW8rDQsc3zBwVKH/oZHYZpdJ9Hrd+8tVl380HQecyVPU2VPujhzL
B1srftr/fMqLa/aiYjYdWB+AwAFNvBV0Jh2u2i/PSCAOnWtEDHstMYqSAFaKYHJVzUtlH95g0+go
Axr+hnlKPjmDBwZVQaMl/YpkJE/4rQNLKbZpoYYcxITWFBcYvuui8UbhQOnSlUcLTjCgd0urGGyg
b1sqBgij3Ilha39pjKqPe6LsYrHNeS+U5rWG0Sq3OGGio/RxrJz44iJcxrcvS3LUhOZfytSL7dxR
Fy9TFIV9JBOFUmvWwZt9QDgTJrbL4mBkMsgJD+7rm+Os9Dv0Ilyf4kzUE7w3YIQmi4MBoR/N0Jyw
mPkg9ioBEpCZuyTFCAuUBh9rcWzUcRIykt2/C6k/J1NXXS+gWcUHQdESx3r7LAqOV3OTr0YB3JuR
vhJHa7hkCslsWroFsE+ghXTEVdagtB5/YrBQEfo/zxgcDUJ2Rx4ibVR4kkfMm05r+p38GPXVm8a6
N3OPyyH0iaEbWazWBI7oCWVjBbdgiqWrB/V/TErO7rO7S1A1Ry33WDwfPwv8rHmKnIqlrYD+u5hC
PuPL5ah0e3p9li8D28jTWiBIB9ZmGU10Rg468g/OQmSLhdENzhJsfNvN3Gja8Jsg5aQfoijyjobk
1aaW+Ti8V5mFc5LRlEcxpfjdTLcWgcZdL69ZbmixYAruS0WNGWyzexRdZwZG3/tyec34VFs8CQgp
Lf1TpcYZjp9FHpAm9/uf5f8vKpjp07ioQa8S0YEW9m0QiK87V4qzdBcFZ1a3CTx9vi/hmWNSMevp
PkUAHf0kKUumKHzQRKXNoqyXhtzYUx7QClFUA/7iyHHL1vCR7B3R13pkwTM/uPyoqAXyC/Q03dmG
e6QcIqau/NzBJxxgd+2PdRyca0wgmukRPoEAq5YyNqD0w1TCwq5OdVmNzfuBmsvpUxN4EosUD8hN
H5JXDk221gZQuqtJ9UqQjY0PaaKG2+L1tO24dWkmyqNTKGvus34tDfE7EEKNWzpL1VWSzswqt2/U
Vba6dbmrcxlM0W37gfbDzR9Lw1119O9dXKN3KHY71JL/eYDsFnTChEN6vXGiu2yjbN0Pm+0MTgG4
CPJgboSdrlRU+H9fBwYxAXexeAgvVHshR22YObIcQWxS49cWejRKTpSOWUw0mfcBWcrf7k3bgpzI
xZSIxxNBKZ74D95Qjp6jzQYI6j0/bP7Zmp2uDffWy7vFyoQj6g5KnkwLNJjodSiULnUwH3a1GOV7
7gtltlSfVV+kxYS8RJQBk7qfVtqMcZMcvQ0oqVAFHJj+EgdfVurW7josMutMoomhuh/y24zY/M+O
EKTzWMkeNTo2D7bpi7kaA5CS4BB+2BJzbK9ZvtcpYzdKkSrodLeltaG6yOEA7PVOq65KrToq+ECc
8kQ1d1pTCVoYrhOBzpdJfy5DlP6Ag1Lq8XIINcsTqg7S6dbSzUIM39897aB50TfYfCIUoL2ck6Ep
Ir+wR2u6p/uKTwY/gLD90n4Z3HcXCu5TczPKe6Oi1Z7v4UJLQpXSnqEufRDoqo2gMLs9fc9b7ynX
XlVroutA5R5NGFA1hROX+JWA1Cmx1Lfchz3dhf0lcarma3LlD7VEMebz+vpPsy4480Lu9muVrle3
xDeKspqerskQCISUYwci+SSXy8r5M8IFAmdcCz6Yhv12tAMGcehLxJcnFuCafEN2gWM5Gwuo24Q3
1AdQB8n0T23cXBseV2UXMXJG4oGYCUc5HQBnJFwc5gJGuPRuLLf2ND3jATYaRJjw8z94VesRK68k
M0G5nJBX1D10+mypuUFlus18AyuBfm81i1SNrz/nvKSobhxaylLO3GXMqsMEulGRADb5dNMV7VlV
XgLXLScJsfAobMR+3Lwq14PtI2CZeAOV4haTscCcByanHljUZqaXbw7rkGZDlhDGfD4hY/vpnA0E
zSHxM8RYS1Rn5txW6Lw9Acs8lURKp6FBM8Ky8NfA06KqY5BEYY8cOI673i6h09SJc4KLcT4itFSE
4PGVtLK5lccErqFySllI/WXPt37PpW6rD2IHwTAJDySo4txOScfbQjHcd4hMdFIqiol7IxgKecqy
uH5AFg4yGV9N+sZuSwTS6RfnxXDoBPpgiP55LbZugIY2nDZHICDjTStMPsxncGaGPOnr0yufV/lf
kYQZcgXAdCbMMjr8GwPLS5lU3OS9OQOrtplDko1XKiw2xY9y0ANptOds9Cn1yGqS3o0T9pvRan60
l9zlx2gSZdqwPX0cDuYwm6g4d+EM7KeCck76LP7R6zN/dN+4kmMfql2XAPVqC/RMhq8OwzNPqtOG
3rh+q0JDFuwbhVPOi+KFu5DpOfDJDxtsE7D7c4UmIH2+1VxR3C7vnFZif2Ymo4Rm28u6NdxYJg/r
3WTmCeyadzxJXQcSeYhRg0UpMCwP3qRgrnCjjsv9u0+/e0xDmMonWcE6l9qG505fjFp8U69CXAXQ
ki9kL6gxwClhfuQi8oGP1D7Cuf6WJPjCxfFlxbIbC0V5xWnQdRb1Ailjau2RjH1ZmKosFOH6H1Ux
ykBjOFh/lVt2lvOXaH911Q3UbwEa9zsaZ4+dXg5E01tK7NxQ52ld9v7FtTU2PNZSG22rGShIcyAD
m8bKM13SagZ3j8yagaxtJtOOzx/megmBxmurZKL8Ky6IJ8FP7PiNLWKX8PdxsSTjR5nU8HqO5hH5
65K9J3e7t6ja4Cf66M08RswDHLXa9Hecw6ImerrBx+cSqzc+FSpUVY+n9EaYJNLqIRvBaJ2E70vc
2L3FU+vX4aShsVPghtlDoxgPhS9YMkRDbgpgt2ox/EqzQfxqoPckrqd/Er3zUvmzY4AlttK53Kd2
kcUEgnNxzfTMvtpm/ta3vDC2cytJwqm4YDcc+hA9JyEihlk/c/kBt1kxA31DEQdyjY9nf4ywxpYs
llj0Q9LCKNc8dgA0Vhekp96mMDaVyXL4M7xweWKXntsgGufuUpujs35NANO40XjVgx7MnVyD5/oF
mxXs9HMwQAt5pzWKgPO1HpE+G8vbMAYdS22hBSh+kAZnjcK1/F5Bou7JOClsrmMjguS4t1Fqsm3s
84svtpi70zT9utqznEYhk+p3UdoBtxG3j2xmObe+rmV/rocJ6gj166uLMkFxkwOKr2ZoLtS5ZeV3
Mix02im1ySPHx08PzxIN6ZirAKHVNNoQQhwDbw0Jd/7kT+ksfso/seIDrYVsQvtZJYgCG5FO6gIi
A27Oke/6Z9wz3xCEWYO1aGDEJ4D8UDptvfOTtUqZUZdcGMa/Ghp08AdJrXEw1otEpz9Nata6bfJh
RNYZX2FrFWKL0Ejp3WiglCDdDvB7CctLilDMlFqFhvzmxOl1NzW+U9AGubn3WjANBkrrCuwFbPpg
5TZKppTrGmmY0yK1V7AL+PRvWc9hP38AYMouaevm+GXCqXcTcBM9Xn6mz0FdIJsryTsOzHIWekyt
1TvKGTLL3SikSkuWaN8q/0h+13iEgUdRqfDqV/SFouw7mDNtTNULWKODltPw16TLX0Ja6PAFOS+/
oemgWuK/OeE33jd9pDuvuJ1xvqRuw3ekMLQTI0TKo32o1oBfuJ7N367/vR/6v+/PI+hl92QZeREA
rSfN5VeiVp4EIJ7uHOtP+B8IxIUmH/miq7d6QIcJTe/txE4USSr03Yntk6S1FxrBBhFzPIbGTPjx
RxK4Y0gjHG0J+JvE0u93GxPlWoEafl5nnWQJKuCX47/EbGjWAdb05/HBT3j/JnIolQGRm4texast
tx4nGeDNhvVRIQ9TFhQ9xT8pkeQ+HKQNPJSGjS1hjNyfJeo/+uhN6pF3u9sQdmgJh90nKLbw9GfU
kWOmuMpV7l/FjdSOpGlgG/G5aQ2yoT50eEK/J7U4ys6lAVnHSD/nUgwXzNNyxyug8fwqOGTzZ1Em
vNOlqGnXMkRuoULpYVtKsbiTGafRSkaG1ZqMw7sAFJ06PQ//cZ+hmiCBTqcBqBGEPJ55GVcPAQQb
zup0kd4pY+lrkDEG7qbnTfVk8s82+UKyKBBtnTfkoEb41U6+AXixJbmaK5oz4gultIIlHJZMkytO
QNVUcK8J7x/pmbDOT3OuOpP0JtekZhGSNVtigsTnzadfbOt154GNcLToniPj+YjsZgtuILgXf5fa
2rrpp9R22PJCQ+rqo3GdnLmc9HcP1qly50tVkEglA3vFAlbpEoE5orkL5Q+NgRVqIxBmrsyyDWdg
X8jst44D/QiZT0h6oXLUEQrM9AmK4tYxJAFAOKoaJJeaWPRF6s1v7jkJqjanIHgc+iB0t3LplvuX
OGZuOKJ4A7Ca13Z7hO4Nngz9JMnZKi/UPRDouysZqg77c+ZfRHJ4i88tktwSEP3NtXQ2Zxl6KPuw
Y+H+cELVwoTBqvs57FLMZx4I9hAuG+i/+A0A5JaB6wlDx9kqCiK4G8v1ZZ5IrCvhNOygnlfEpklV
fAgv6hEPPt+s+dZZUw0UePsmk3Wjoegz1jkSpqANwsd5Mryt5o5RUhuts9w8zVTf40hvA6hsEwGf
HMHZaaVGtFYk0a3CFeSILf6v6yH2LJsx8iEX+04UGnwkTQb3Da2haKJ4lKFhxQ7Y4jzcsUpcSsJ1
6OWJbbvd7hNp9h/78dOoIrA4PeZpuOZF0JtClNAFNz9NVXyRJ1Lu+S6nBrC0aFP9zE1P0ymS8blp
xuCH62WKhmgjW+buMDxiYu4osUK8QuqFuM/S/pMkKc2/U4CHvmkwOGK/Ppbzlk4S4qCBAmLwctrs
sMiTg7ZjvLGHkc/EvN+2EV1BAeRD+3o7P7ZiSgh7DX3LQ8RxOotE45T2nU48ccaVJ1lFZ/5EF2Gw
2Ahe/VkhNGx/20BKVHcfAqui3cI2RGRKZr2NbN6+r0HzrrEtCsdX0G1cvFDV4qEFWMpZKCGnyPAk
lmmPMyS1sLcCSmuoTvWVfKTg1Xq18YX9ccBFdmM0zt/6mPRppX87EnNBLhpqIW88yFrGeNFMvWgA
BkVkZxcz6wXpf3k6kQ8MJjBBGQUcVOLL6o9q2RVwVYsjYbRp2+F5/tvhYhNu2hPK+R8uPsqbFUj5
aKXokjiQ1KusFusZJTztOJ+rYOp/If1tEgq1kjpsPgJWC1YR3GJhwqTmwDTQ1jrVaVuTUP8/buns
vHe80lmhNvVbBh3SJTQI3074TVvLrEIFVGuZOSbjKJ+qOQa3M1izPJ/rYpjpL2lc+9d26VZYh3sE
DOD2BXHwFlHJc6cupeAiv76mkppSULcWgmgaTg7OqI2muYIYZrDx8b1LKDmwhU13Jrm3IKhyMVh4
ufCuICSjBN42KjYgeWUyKgssz0bpXhyIVFjOFi61PgjHjfRkkOuXxGMFhaYnVtMrVYkpBPPipOwy
A7UB1dq36HYHlVWEGHjWUHBXrZih5QKwqlv3UZfXvXwJCb/sldCmfpBvdgYglE+wNV9DlxS7sELq
VgWAtQVcEoFEGMO7r4jCU5Ktosgg4ZW5ntSNLxiidhhZhkKnChc8UYV9dfoh7T9W8CpT/D9+Bu+n
Xy0Tgr0Y7D+xexdzNlyRKZR9HmLkuilsl7UBrk13Vvl+reiVKJ91VumuoB0BE/eagnUf54UicutY
kYR6bDeDp/7GtFmZz8leI16B7BXmL25zcgn9aYDwp9rTKF184p5cFICrOWx5pF/oDZwjLIdiO3ZY
nSnNDfu/BJ7dImz/8GcJXbZ8K1ITzhKy/96jp30YQdz+kK4fcZJzcH0w03f/tc9ICGjC7vYgHBNR
aDcAtIfQKbCwnKnqugQHYo1MoONFtNtZEO16ko8I2/6A5euKefIU54SSUPf5bd2SltYNi9E56qbA
8rTwS66u3Bdt8ILV3SxRICJD8DzC3CVegj80PyowIv/9pJKYOxOS4qUHh4AoS/UK4l1xE2VImmZz
t+mwwfYvpg8hnJznY5A4lWRAODGEXe3cZPwKMUjYRs9dNp+1O61OLqvc9/SjVJMjdWbeVUKnGjpW
2jkUsFgq9KW5HkyY4HQdhXixTbUJCmFXLolm+fJo0xxdxUwl+Ta6CtZ3KZ7zyMxMwi8tMwBp/KgI
cV6dkgowfnMARd7Ja23EGsMVRgr1iPtDumdXaqAJx7ytpcyhLYKb/RGJ7TRjro97/T0hWL2AufNE
+RehgMiWLwbg97uk9Pq8f4kHEqGSJ+1Jo6k3jK0JaK7yN5D+9IDy4n34FJxBmD3WFqTa7M/3/k+K
vdCbefdw/Yw1/nnjWvmy27COzVzFoM6Jg/uN2GQZHwKkA5G79vtr1vYOhTIJZjbfsasXiQSdAPtH
CS7YB+b5+bm53IK7lICst3xRtKu3sQfKopBXzIpL/wW7Rnbe9jq+edfqy02bnRdTIiOFUBitR/Rh
IbHJ5PyQhGQJ1hdBGrtD3rcb9Zipcdy99cHemN42NN6uqHZaZ80pmxTrnHpKKk0808UHwXIVO+Of
sShOp+LBE5s3BnupvZZiFTrnxgTkMKuygER2d1x6ZJYpKTqmTc66k+XU6oDXMFAbb9Kxc92BFYE1
usKUz1KomULuB/7+BXIyieohnrxVWzJ8uxCrYSdGBSNZaN16q0kAX1XofproiY/gRomEdFGlXrvw
GfIwu4oNcvx5d0daWd8A0hYAIu8uaA3xzPhEv8PMZ6fRJNuYdSdjx7/ndsK5SXP/S/0fDaJiNVNd
GV86AxzazjJjngYibkFNN26kQDWEPN6e6jxBmbHWTATxSmpEOVEI0HVCa6nxiBocV/NMyR1b9x26
8BrBPdXjo9BGbDWN2Gr3bfhCf+i6faumsr6Pv8QGTQz95aLXFECsF/4odEYkooOkN5yDpCK0v+Fk
g/6DXPiqv8QFrq0g46dfmCm2lEJOyi5mP54zKUPzFz1hURzOufftNGoBE/uTcr20DJItXxfLrXMF
GWKK2ElvY8vdnsZ1ycSkoG2zuMwGsyvjA7QGv7dajCrTZpGn+wvFcH7OodyAr7HqFW3/K8+EpGYL
pGWw83jPWrbCh7lT8R0+Mk+SjnlOomTsWExxWtS6DTZBeTWwo4RbGwtXaICQBYJKBzb5Jhq9aNOd
N4D5hvd2D7Gb4sfPT6Dh/dvEIcBhTBXNWDA9Ktcvyr/7QA7elhpxqUZ0z93zXpBl9eMFy1Alv00D
nxKIb7qLxS2ipNhgXpUvJQAMfdvwjBwqOphEY0UwHalf5QjS/AA/d0R1HQDA53bZBuPQgt93zRoj
NVkS5n/0iAoUzQIrGnXR33+7lorD1GrLuiDj6Nj8bOqNHfBTosP48Jd4V8kpqmuaTe5LU5oNQsDO
5D7Wd5Evu20GPztM/PYrGCurcM61u32+GliOT2vS2q7f1VKwMXcFeO1xGn8bVdcXWk0rNdkqqEbl
yLaE2Oe5dlZNXjqcImV5lZaOmjJYMfpxwluPPmiWPqh2g+UGpaBVAhi6arX3vem9gUvpleDozuZi
EP8Sdb9vzqATbBq19LlmK66xcB7yRyxqBYfu1lcWbcM9Om8cQTzjuhB0sxVXcd/X8AQrZQ5yjJan
OiFqbPAUTypCug0umcTV8DWPR6lyfGDgXO0nHuoK90LRAcDOzRAKAO4EuAfcXT1aJ81ZwPZiX2MX
jiFoIV70766GrjIaYExTjgBA6f7d3wRvjVjVNxdzjCsAypaxoLzEPEDXcxPppbedyyCTsi2AqMkq
FopWVZZnpRW/iNjSwo/IueQ7sjdfIuq/QML3i4ilsla08WDV0+Y2227CLaKBHUHKcMqYUiaqI9SE
4Eq0CVyBt9gkG+Gy0VIxIdxR7Vn4qvOiSiXOzNXSbiYS51zQ3KFGxF3AhZafeDz9TIQBWAuDkk1g
HW/W0xKYlYCNQoR0ekS629AtlSvdOipUwpt0wqygemY6lv9KNXZm6kNhlxia2dPrmSvf3H+tu00A
vV7LpWFA9dJ+vr5vDSrVHiz3mT+7ng2gN75N5gyMQwboly5eO45oECwiCwj2/v1rqer1kSKX9klD
dCDl61O6HT9GK3DciQD5hHu89e2/uvPjKp+pzd1+TX0/3hYqNZFgFXkx6xla6LLNcHvQaV92uL1D
h83FIQuh/jd8Acg42aP6xX+45eUCbmDzCh/UZ8F4PgG5/XKvB8VfXAn6ZC6e4FWW0Eru9gy+8216
K7dbbjNGwMfO86v2ZIgpirGVzlLSaNneVGqzrUm/KWfk7rL8kjfrB35G8r/PmHCH4UK/OCXbFyEt
ufsnFqjkW/Rx7BJ8U7gbJsggpylo3AA7K1EWQ+qIGJqPPptzI6mX4v2tsyn4m04O2dn0FCiMImvR
ymAHhDG2l+xV2nX2WK4VuiJN5B7cQLqGQerR0K1eMvD3ct/TfoUNp7xsO80eJoa03uXTGs7F7tRe
RW4ZPgKUmZO1GcjG2DzCyNzH58pOhsuTa5XAAYisktnD6u9EKc4ARRPmof66KWp+AdzR6CJv7ti/
LbW/GjEGEPnZHiO+RkexFZiAq7NajwPDvLRpHgUd9urr669HJYzM0upExE4meDys3oMsxZLSMxkT
Vzsj+X8xDLpst+VPtiJv4rsaZAxNc3aMP9jxup1fZtOcDaweOzumKMieu3gAgjTTEQhs7K9W6V0o
UNJqAqUbEWat5M6yByq5YdLi9GnlWCDbBhaju9PVNEo4DHBaDbIFbQPvdFEPnYiYa4ciLL1F6I9U
ZTYgZK9Y639nNXVWZKaGtGmlI5PHO/arQt0OzN3Kc25WDUOY9+PAkvH7c8Dgxx1IxTvrMZLDUExk
HljmIj0BvYpQnNv+0yZi3vnzjBb/DXdaEo2j+cpN/4zY1E4IE9vYsPcOhcmr+jmDFhZFFL/lMuiG
GBodJQS5ykI4v8btg/tLrOINRaUfPjTKl+MVk2ofVPXxy+5L5CgpTFFIiDw7hCYRfzxcMhCYvKfB
1BbanQXfCSFmcxBVfCfblmXtlmaEPZo6woa9MipZMz87x90y/90C0Xxqgbt9VE+ckeNwWXmaU6rr
izPEstQBjowALOaZbwWY12hCTpEplRBIcEFEjpdwp3FEJU9h1ca6+vvquud+pwmEgZSu5pF7wXoW
WIQXMPeGLPrErU2LTm20lHhs0VaVx7oe7ca8SSgeAxDjkEeeHR3Hms6om/8DPApjNHG5FbDESDGt
49Cvlt80wDHrhdW3lWc4O3E/E+/H2MdtzRi/d6P/bpPT2o+R+32u6ULBK/WCe0TKxTqOO5tma0sK
awoEgGrvRWqEauJi+BknwjbQMvpN3GEV2PJxoCnBgc0mY5GKCf9w+NiVmxia+LaWgkSshyBhE1rb
QrKKJ4dEY0vYhZ6oxKx8Y9PfHsM4QpVWhZIAWg4l56Fxh/0lfS7KBkmO5iDpCho7U1ns28FbnarF
75Ed3LyQDJW+z4BP72FZB4dfiBFxz3pGjkddUb9rKpLZ6mP/FVwkDutA1xYd3WsNbCCVJ2odfyAG
7X/fhOWl7gBA0dcbgkqtlsdowgMJ2VBhHVcA+HRlTKJ585r/QM6T/AKnmDi1Do7LvXQDt9pjLDT8
x1e88edj2L8cBFsrAzMAiExDJBkVRVTxIDi4RU8csNKohBJCFhcvyO0QIJ9iioCEITbS5CviTv3r
qeXlGdR0imTimj4i1dLK7d7dvIe2DWj2UvkyMhC9swOpXRLFvEjz7IMO2smm8gfgBveRGdryQKGf
f+PTiCOHm7T4jtu9ucUjggG00Ghfk6BvuAV68FdkEkUY0Xpjrer4LwE+5k/FF/7vzNwjD4I/Zasu
BlEDHiJQM/+Q5nKB6dVsCkHr5tKnN/PRJ/mD2o3yxXCzePK7FAVZd4I4HJE33SKHO8+bk4H3jaHn
1MzsUtI/7+6OLCWpp2Da2aEkkNVkwWz0MY8FDIMZX77Z7iMjcZKrLqgGuX4wGOrttTzkTekCam+r
LKVrEXiI/YsQMJoUr1jvOaxyZem+4hYhtUbVFTS7V2Y8zWioR+cmh8IVXTDlmztNI0qTEi7iQGjQ
u2/KJSZqOrQ0LFI+PAcC3GfrPy9ZgbH0ynb42GoDe31IKN8pkCE7nCYIClTtQlUc7yvBE4rP2GpK
7QKP7hxhvzV7XHrcj1obBz6xZzHhUJ+90+Er+6iyMUJ8r7HVzZ6RZt+fVC39i5bd4k+N+Z0xOMhQ
oOZnZhxz3WPpEnwrlaPx2RSZNF9ukQgXxyYagpwXxm0KH4qD1rE5/uOFGY347H1WH+n9R0FUMtuK
q6FVXC4E0TPTzshuXoLjXGFTm7cjXGHvLdFse7+KFJdtxdJCv3J8WwOTiR93whYYT2t75Y9tc7co
cCS4NO5GTywc4wl2GexemNuqFwDyq4Htzu3ik93X12mD0ORbTBO7zINpmR26najIpgioHJ+FaCWG
ZBvTDawEwk+hKtq6nvt8IVCySJmUe25wY82fSxpY7Z549yZOMPUVMbbJ5vyf/9PPkizrw262unie
H2vOPe3k2QeFuNquG8Pw1WNK59mfpqwASiPHlQlms3x65clKmeQ75SfoNaTKTPmE/23QmCwJTFFQ
RpQG7B1uwIQ4OPTyZL2rPZd/ME7wP9l0Gfj0v8FdhlPHiAR/IJBn+1wKvaFSD1ZSLYS9+Qe8jAy1
mI9UAY32PvA6u8xUrl8qA3SRjt7nDR3KxBihR3cyk0Lwjlf1A8Qa5PGBGxHhJ539QDpU7cZzh9Xg
jYBDppDM7f0eDEQQzbqK72GtU8S5+ZdgcATbwbBZM0yto8Kly9+VDsUSEzrhJQtRQQt6YHfc4tTL
lF3LvbXZ+SlaMAL7FsqEoOjlSil5G1c1BG7sRrGOP4OF+uYn0EJK6vbO21sD4nEgYmQ32af/cRux
EkpSnbVLwCSgIgj1ll1Ceg8jOTcFXL+qp03plJ+xoQpGVn6W36/z9ffIVC/cW8AnNGZ+5+TR0rQ4
gUuLZaZEiRVIXYh53sCy5Kxi/po+gpLOFMSIvnU03iGcRB9PBcA3HrFfCYc8XDuhrBXA6uytKysO
jEpvdRv3jfQU9FFdaLhXXGgwZbX1HJjxUppbsXYeq3suP127Zk169e4ELySOtFFlaotb4OGb3A7o
PgJqdKZ5S6lprjR2j3qp0r9kkPYMvoxIo8HintgoE6FLqkq00WqC38Oq2GsZLViPx81o3S1pnFoG
lTyF1MZQ7iSFEnymdn+RXUY5+AifQ05uqfZrcYXfHSqWYRwo+Qp1iBl/JTh4dNbqyz8Z4DEtwoh+
nOM1vGLArWqX6Ps7OOfAhtBFKo3iwKoPN1OXs0/Qlr4tHJUJFVfFRKCO+/vpuywMLb4zD2tZVyjx
0JQ1I3Gnb/6xwlNBt69MTFrpUJIC3fOmR7YIoPFdrdWHg6i6POYVfk9rEbglbu0maWPvCLJ52M9i
LlWo7L3EcaCBTpBQpI1rQR5RxOwSSsB5m/JVKK7uizYoFZqpO0iYVjdfDr/wkn4C39OEaVa+2DVK
JdX/xKMU3qG85nk+83iTNIeTohxBniVYWTdJyDzfvYJOPJaixBM8fJPPshfKmFkfhFDThiycHT5a
dMldiMLyDGk4ydmWxm6gy1uuXi1P1LQ635wVJdoDWBVoSFoJGMA1XxhX9oNH5q0DN//RQHqbE+Z7
w9olj65tRELWNfYE9le4crQ4QI/kDCUxA09EPAKUIYoKK3XhwM1JqOp/Qh3aBnFjJCNNdVtQ/HHA
Fo/CLxhcXnggm8u9R0otqzi3048oBZDSg+KgLPqh1C6CcnV2BUln9e8OvNfoKGf64kovEal8FYyY
M+Qg7LXEGnAnq4WP0GlSb9H9FgGapFpRZRKdpc1Ns8Ps7qWfuCa6/3vcNJB8FMGNme/iuzcuiUhl
BsSMmIKFgfKG9P/ufhR6/TtuyS02hRhiZE1kYcnW1MIs//uFi9wEwNlkYVD5Ag5ixC3ah9RnYmF6
IEv2j4ZJYK89Bus/AmHZ+sdNDVuyHGL+LueJiNoL00as8I3sSWYVaj/CUsn22a7+ONfaS6IMjzY/
xuSZv8YRuYLL6QWbfjvAuZbN4yyFrit7n1DxHhkrp3G0K1OEt1P7inNitkhEDDewjYRUpojmjDX5
VprnJ5A0sJw/yRdLjL40l1rgkqrTOrxX38+Dt9mZQsUAXgeDOKaiBKEXePhqVPmaFd0MEKRpz/wA
B+Mt73QpcjyQMNHYhSeyPTqrbEDlU0odvfNil9vZhY2UvG1egQZ1aEeNBOv6bEFi+iQ4szgqeycG
aAc9DIv62og+J8w9yQwKKr5ul6s8bdkugDgvP4SEhY1ZGk2obbF3Jjf62b+7Y3ZsYnzf67cobIAu
a25ihfSYoH/xmk4xR6W/SelKDm4qYpfiX7oVUYOlktFyvzQB7+qjqRIFvd6ldjGFUBTTAZTFd5Cu
6hs4atwCygXtedEOZDg++3Awo7Gy8x6HFxmzfXFX80Ay9VlnM1/4DV278X61DlkIs5uuBNAVYkFm
6SCP/7ubOa5Ek9QsHT1sXeB+s2g/s3NnKIAUCDmE3LBdx1tGcBBB8JhINjiGU0366cYSEe0u+wZS
gfVOeJdCAIVG7O+LSZZt5uI/17vAjzmpCr60qHg/gDy6cQvtwTfGNVYIHy7Ol+EEkC3SbXtmJMxS
bOLWLzB/BdzG/q/YF4p3FSvIth8CnZT94X+szpv2uEjmfbR0k+By/uj55v80mZywYjewWmlNh4hZ
kxdvisZP18/FsRhXTfkGcGjfZd2dXbDJn7fgGS98qdLCpyyobCyK6UuK6kIjWSx7VUIjU5wSL4Fn
V7NHAU1mBKPNHgdAOimP0tNs6h256oSl2VPZjNUWzP8U19dg1BUPhd07puBiwvnmNrTDcr0s45Kt
t+7FmacsRO3IBjp/TS3LaWAw97rfDku+QDDTVupc6C06VrYhpVUNcXYXdfcTvvAZcrFrxbgb0rBv
PH3AhlmykTWTgf6AcfyK8HmnG0VZ8KCeL+3Z8VIg/FhpANUuXfctTv6sOSZ4HvJf7nT/8/DUIRY3
v1iCitejPGYxZKf7UUpWRMJ0UMv08GaMY19BrCvAQCzauMTV0x8AVvpIbMNI7uS+ihwru/yF9kQt
QLQYeY865y9ZrAGf2OtdS3FylOoI7rYx1nvqY1JePhrz8ojQsy+nMsuc7Wn0QUhSNT2EbAALLyQE
0z56eyu6Z7+9vpKY93N5e/l649564+I5BSK/er6B5coVVGKTKGA2cBpR7lxNTv+YhIfxYG7tjRrI
7Fikbr8Bs3C5GLT2uh+L0kudKrmBBAa8RCifuFOrjGXDA9zGlh1Wx67oHX+c6vJRa2DUf3V1bRfb
VwjBzFOp7gBQpSOKOIoGtZlcy/pEWzBEJtlnDs8xkoW11RdNiNFHPskiucxlhebtxHC7iyhqi7Jr
k85veR9gcOXFHYwqqJg178CMZna1jCuVYGQixKWqcreR4zgQr9qiLHDdiQizWjB9tqK2qeDryLRz
M0Ux2Y5q8vW1NXYPwLcEPqHb9FrmCi8OMKg7IwTKB9Nqu3aB0LyQeSaIFYM9ItlrfMm0qnEjSmkb
Oo/bWR5IClhDmcnd2bWDk/wmwQtVyMLTtc044JoX3Xoz5a+6xjonK1Kx9aVHQdJUJX6/NeJqzYL9
eH9lxAN3rEnQO0e1j2pMoxny+0TXi4r+Xoiz4iVnPcpQ9uudAooak9OSnX48qdibaAiY2RSbBgkc
plnh1p/rHs7Bxd4N8mTLi05TnK4KBGgMD25doTx6aC0rVruuLKU49sPxBsNPG+X8f5tTL6V3psqw
qJwhLCqlHR25Uk8hE4USzZy8y6Dk5qMeAVPVtC0glHn1prGVUG1h3XTZtL75ECaS5KUdolQ4JQg0
aNmGP1BMNbBrMBEd4yKCM6caW5FB+g3KvOgi79ZXn7VzctUg62jq45sZuxir75w1CB4QFBgtscm0
wO5s+wvdodJx2JiVYLoMyG1a5dvoAtkINoVd3K4Rho9MdbFGXSLOiq2xYiBkSwnJFgqTUiXdfmr1
HKeRgB8lL2nj3DLtAPqr+oGWdkwkj2gjNlebKQ0pmxFOBwlAOaGirnASvKaKsPd3/5YuimyEMG3Z
lpkqT7/jjvvSH4UslW+TRVtviwaHOoUqqeesbbNDTWGwW1+wm2uUglKnQSffGCx617FNCVgI7EWm
n5YyCqe7W7kaYALXt0X3PLuEylVuVgfLfIcB15qjWZuyrUWNwMAd8J1l9j5w2oRGP90TAkl0uU7b
1csgF9/+hhK0POE6b0aMiAMu4GIeAuwCER//27my/uqluE0r9Xp8xNFaFoEfbXGQ1uMrnblcx0Gh
tVkz6eArBfXtDPL/MAMe01/BVY2F737G627PtL/hn+ZX530XdLROBthw4Yo0CLe78pNwwkjahiaZ
LEEQZZVYkh30Q/WJ51WHBrZUqXyo9msKnJsRjGml8B3zdNGNpT/T5Tk6dhET6wotHNanUdskYeox
avXEVQFTdZlZJ0fG0q4D9xl/QinqdOwwL9RltTuVkN47WLOvTDchIEAuOgJSJIhQ5vlaAZRDMpUR
rR/OyXFf8uJ8oTOg/Jh/QD1ZIlPARzD61vmo8yKsfMSr2JAXtCvD+Iqz027AEeAGhmqtlPA5rcG1
cFqPgIAK12oDOedkcScOoOCgep5DgJOKNHYB3W037+fGvKBlKFekOMxyyk8puv8my4vBbILFhFzU
ourXLPf30cfkiLC7m7SdXDwSxXEUHH/Js35g6Bji7qd34tbch+Qyw2KM0QDN1zBm9jsqMM/xgSTM
uVE/OR1eJcY2zwRIjYnlxtU0KNcckwU/QKqIj9oQ0Rn1lQ/xjcef8Nbc3FqDQnLGUmAECdBkuwnq
8Bh5dQqQJG3hTgKlJ4XNc3u3uwEQTlbftJ+E8wF1EhXVXLq78I9d6BP7RiOBudIYgZWJu6GLIZhu
NS7uMO++LtXeEc26KzVmVHhnbQ2+OfsDrm0/VmhTGfJxrkyMgrKZcpHZ6MctZJcJfxrPKWomCqsQ
Tyn4FGdBMfC/4NhIuh5WBbKNPrlF1cjn2uJw16f2pZWn8BxJVSwGy3Fi0z6S68gpRP/Ko9GOxiV+
xM2TbOp/X9Y1aCR3FIVv08Q/14jsCVB+Dk6PCaIf2OHOsDmq5qvWaGZTbQsV1YW+oVihArrdLsoF
4YEV+N0Tuc6areY3eQ4LHUddjXLBl8DUWtSr5FpcKls2Nn/vz5WnBzzjui57ncHvi/ywF/Lj47av
Y98OeN3QZoVgrJAqfCGN5Covmuatmd3058qTBM91dF/Jbnm+geatECiA/7frMgV5igd+7q9eXSUE
haFsLEugAvyh2N/8XoEcwaLY2o0U+8HbJeNhmsK1Lu/YN5xVXc0dWL6RDGp8DBp8m3MbTIF7vut0
z+FobGOrAM2emVzRXRReIxsaZhQ7l3nUxM6gjYaOmLafTwnWbtcJyA7SrQdBx0Vv643VeNih+nJ1
wLvsG5KwpSoTMTASto+YDVzr+z/07Kd2u93pH9oN4sPo9sd9g9lb6XQWk4LLObHkBtMTSUBvA6zf
78mbjXRe9B03UIDfvS5SMNHkzJT8TWyvsiAvWrnCkI32xXtzFHCb3EBSqpobog+rdB0b926LmM6/
SZq+upxk2msNXOvLpVG4UxIfL2k1NeRv0xMep2vYEi3/ObgiqetlCiIJnen9PjmQxpTNoHztOS6/
9HAt0gmpQSVujAk5ODYBh8BxKzr1e6oy1KBW9MxqIvDBG64DxphDdQ0xezzJVuk3qsdyhXJipTN1
TtkFeJ/v5OBn26fhQsY9abGx+FyQLuiaw5RLCx0KGFYp35ptEuXXQXIL7VIY11jvcMlhfyvAQjwt
ZcQ7/9aG4C3j/mJ8Wy/oPpyRArtlL09Oh4E1VrSUDM0Ka06xhVCVd1xjZhch2QDkIttcbjhrqTFW
JF4ppUJ4JyizISFODf4dmzas/bkzrV/tstaVFS4GbcHDEhy8b/R5lK8ztmBFgyMnPxP3hZriq08+
QGwpqOtJiS7bNoNMKhs6THpncMkktfb6COKsesaO8j20gtoxAVK2giEJ5LFHECBgOzsfY1QgGEwP
PEOrF20n7yk+XgKPmwK1e3YuKpfnMfOrDS026yAbas49LeehQlc8lrCdqhb5zB2Nt3gQOxgA1IRp
x57AYtu1EQcyGDlmqwTWeRNACJMkVulRbk8qfOyZPl120ifizpCkBR7LvfdWv3ZU0NoTUk86KfuE
tA8HXM+tDFp7qvjmVpDgTtGkL7KgFbOwkd8vlUeOx65iGv1gvmgj+m2fm2Hlp3TqKb5HXj2kTqYq
KHQr2NlecpX31v1/Euwm0D9k9WLBHwmTnpRRRmMLCMkc2hJJmP7Q5odeQkQx6/fNlG7IOy4o+aDL
AV6aND4t7kLvV7AnlI/jAUDbEGI69IdVozmjkcW6/QrgzIWf6UySy2TkljBsixIrmv9t6Wq81Kpk
XsVTBrciCT8Lp5Kfh0KpZdRUIoTQx690h14vTOWOvzCwI/z74g8LrTuhNpsHDnAIzARjxDXqbeP2
eaZhB3MzIicQc0cR3uz5hMn4fjvP1r6WQJN1BCfX1HJgw713dmK23rY8DDD1U162o77LhlgKpQjb
mOJEgaNKrWZRwJXJufWP0B6ugDoW6A8Y8SzfMWE15tz60CQpQojawnMrgpXspvY6K38KuFnilxfO
r3qK3F0cVSb2Oo9YoQ5cXwCCnFY80P6Y/NSkHSqDSF9WWlhZ9Ici6br+w7HSm0Cny+GjFJMG1bmK
DI5APbDWtsdFK3CgSkNWXRTiYsahvIKTQFJcPnLx+EUFTLjmLvM8B+jabnrvi/AT6JnFtPkGlQhK
dh3tutqFrZQ+wF73bpxyyCouYwoQb8XrwU04KL/n+7DeAbT+U7l5pHe3xiflfDZ6rEuqOWJ06cnz
RB7o9eZGEBGV3Uu7GpD7K68kUznbUcVlWvisR/s9xMMTyszZfxmWKDZ+fWFjd3zH7r3rNc13sAYo
XeDomhbPNBHr6Jro/X1/o3eCqmKDIqhEs5eYjGX7gIj+ZNtgEhj2CyhFYGNLBML/HklvbnESHkvK
ht4I8CR6AoCMBGjiUqnfEGYhWATkzyJ0kSuWqqgBwToCFosl4Ed53e61atnSxDLFSK80zgCFUL7b
C74eak5NHFjXwqsNEuNppsPMKKeJ91E4E9YHhlXlRbYUEfVza6Z54EEHXr9QOPYiVlsQ/DQvDNBY
iOcEojAUtcso07uDRlVUjOVD2nkwZBmB07ruV7Jy3AhVxSWFYZvjvqP9osVfnQN7YH96i/wWYHNM
MyqZYriRE20FwzOhWyFxqg8Ku+NwQ+GW82M1kfHbV/cd6TazKyHNJImVAyo9dp1ZDYVIRZl/QseY
z58SuQB/zZVw76p4u/UNkCNz8PhX7CsmqeUjol6F/2A6ATkK2m4JKAe2VK/x8zOliuXo1XXUgCLf
0bfyuKzlzZElVCApUA35fXot758gruVB1qumwJZxx7Kd/KXUvpnQRMd6+34vvEFy+llVemwX09ID
H46KXGXt0efGe2c/TRRhMSjwtv0IX9VqaGGjHFZyI3d24wgESJKvtj7AzDCiPqQ9pAzVxy0z3LcF
FcoESItZ99sSAr5ovjjKhZDHtFKAQHPo/m43oX2xEh7m3KPwqto7vLCOSpHK5GZuVSOywE3A2M8u
pJvwwmbNZSqb3M5pNpTrpGYFwCPcH7Q+i6cQHELZHHptNHglU6/XoP9QIlzEVuYRLcdOFaH2LAKS
qeMHA6b7rxdhbVignsf6vGmv93Efn24Pj4UGWsT4hsmZhtMbNvqJGBhZ1n9SqyMPjCxPIs2EXdoP
uclBrZWG3XV57af+g+wUKI8ln9Xjv+0T4Rs/eWsoczrCcgomlmUM9r/GhnbqLg/6fvqz0f2UYG2V
zXNiVHin2qSfQ5Qq3RUFb9Kx4R+dvmfYdlEcVzSdVHE1/GTh98whvqLzzfQWlxq8vf5pshY9fEnd
BlZBNXKUzUZr2170rPg8e2DOxKCpacETVR5X+tiYR2winE9kIy/i8Qn3c4VdQcaeyMrNTZBQoBZ/
SdRs15wnvUYqfvA0OxQHmX18tYZH61oMEWgwkfmNhXvHFjxao7R+B5/3dJfL2TdDR9oByoyhbE/n
iqAUrMnRW2rG0oOCh2tOeiUkzuWrnXHjE32FrIprn3WP6lLZ5j9XLgC9K11kQEhFsXoxWJv01Qdf
stE22w14oeTfGZORSTYxExKQzAAMVFvV4UNBg312Tb3YMwqKPZu1K4oTewBI14oIR+MYxHJDH9XD
tdYt5mNhX+LRAhM1Fl0NZm/SsfS3u8zLpd9Pa6ptweAlU9dQjXlOcX00kAHnRCA5AkisVF0ssj8h
OjHNe5AyQb/nAtFyDI/9MtUN1OSeRsVEd3z7CHq9m735CQaOh+BGJsAEVpjAfuXk6Z9hpqKfXXuW
xmNE4AE4qOHcZ51k9/nT9tTsTl/gNhSEme337Z0mr7AsRBTiFJWwP9U5OBfPqCqTaz0t+JU4T43+
2QLprxh5WYlLx0G/bisDsElwW/b9fbV1Z3XSP5xw5YGb0fEIPGsP4ueTBwI9EHWd85jfcMmQFwFQ
7HdVrgS3ehE90tjkpKPqfLCtPypzT4lB2uuzWJTDBdEwykysnp3WnaCqHrjUZqOQ0Pq6doXwCNL7
ReRPAer5eQiqBRKRRVz1ykW7PdKJLpVHjANPJNtvwXyQAA3dQSIc2kK6h3gQwvKbX7bqlAHgiKjj
jacJcoez8TP1/ceMfr1md5oY7VHPxzcHBJpQkWxfPULsTbBf94TzVkCCLGnrD6nUus5lPgTbjk27
ywI3loMT/8nRgGbxJ1hy9PXhje2VMe4F+AysjfCFHx4hZVhhvdsl1YlEbJojNurDp2Eeri9hUkXg
o9/X2+AisRhFQk3KmA2FZGTPsIzGeKAufIkn6+kvN50kwHZCtSZd6DnE+tutRNSCcJSdcl69R5UY
PttvWPdWT1rX09ajRpixooZbtVf1ul57qsPnBPZ2bBr7SLlvssv/BiO8CNvHBNZWWPNUNS2RKMnP
dshYn6cJG2cNCYDbWHlQOSrxsPXSgK0YVMPIgcgaHXbh6MJhrHNefBwlGAqkmtYIJQSv9njYojAJ
GSLXXx900YjESD1t5kCVhQF1h1nRcFhSKVZDdzwYihs2TYIMCYBf6VkzJBycy2OKikPzU4vP42OK
zFYpNHuoEX4UfLCXXedZD4Tuajdvll2z1P/+9KXIuDxDA9NfktkDPovgg3BiwgWK8+kX8+Tp9jgE
icHaCaaLTUPBSeIR5Jejwm8/2sJxV8par3tImZpVR6jyefu7bbW1RaWNfZjXHlmYiisBY5k4H+PE
U9GlZ9piMWlXA748K3HaZ2IY+KOU94ZmrpiOmCBBXzpc7CPzkS9rXvrZ8UHUmGDud1F8mibWZJjP
2p+CZEmemEGOOacYFf+x8WnIKltfu0iy0RB2B/ABD948FEBqULcD9iiHAJp3tEWt/zkdwa0C6uLn
58Xnls5aHF7KTE1iJQHNYXbjfjQtcsfyshSRlbF8v5bPFWL6kmfX8u81jYKDVvGba6uPVaAx1EBh
fzVvSyy2xWXwwCLV/p4L6S8tH5S9vs6G3zs6FjQI6ivtR0Eb8YfViBwHtd8p2oQFp8fdsG5GgkxA
Ighp7cOFBu69O7xMKFQjFgjynMrxIA8I7FGUQl7oGDKEgbnpYDDJm2TVAZTtbfqInxqxE7JPYePK
1ulANZSZIxztlKqKow4aG4nESh3krWAKEip0zwZyZq73iRd671jk1teBHYrUcloR0e/j8clX5GOu
xLG+4BKFkmSg4vZyT8uRv9aJ9k2zNZzuQ7mvRIoOtvvTYzFNMp1NOn40Mw3cuUC6vSVaaze+8aG8
yNma5Xdp/pqgorFUswhlC6QiDSCMnuKYfF7XNr+vdQ9LyKX8VDbwnAvVnENxV02vtC8/eZgZquv+
v5o4zRPD49HP+HXwSt/2TgsKssMf7xrGu5GGlP2gcyXO4+Jlzsy6HNocIW1vXyT8dhtJijsQToJ0
/o4GNEXSJ5d3W75jn47tRoQ+CHDPQ/CpdVWq+QHF9HHNFgKEpAJXAgIuMiQniEuNbHi+WRfJpLjn
5hC2jWUTTdrEH2MQMSgBbU3r58dgyeDbtWip1oArUDTEtUKeaEI6yvvWr+Lh7uy2Un7j5V0P+pez
ApXCTtj+nCuTHjStJ8hu1G2H5NF+DOLOjg0755oeTM5mktoXhJAa0RPeklHpDhidWVQ/XsSdxNMn
q//1H4+5X4vVEU5t++4ZmhkVtLQAwmhzZjSIQ+0/a6y6RVWLwkL5mhlkGAgxFjzFjmyn5Kabpt+3
SJhsvFJ7SqvD0yOGiQrBX4xlNM4MSkYstUx74vcfPB4WovNO2OFI9Bil4Km8rtPKRyP7fPiUYR7I
2gV1wTaRNo+ocXQQIicKd/B9+ciMqmig6A18EVNPdktps1g8QItxtNJG/kUvdoayBepgCYfETsCb
ZYSF8S7Kke9IM+yw4PmeA8838Ve63UowPjyGy6EPqUIiIkCS0rlfoLbInVay9cVYzVthsUDutByC
/8n7sl4UbA3RjJlg01Z3tOCMcoCVj+1khZB5QlnVrf0V3CW5TMpU8QZQ4LRUWNSmZ94LlzwMBmAh
Rw6MWv4kE/3oiCQlKBGYsmV98tgSU+QM4iKHtOuk/qB5GCCOt4eJPJEqnzTJxbkvBYT4PlMpctIE
YiLtxuU6AsnJvIc7pLDiJt7B5wnbsRxxiSntBlbZpXpx5UVVKoVoRbtDlHELuEbtC1dHYTlIJFo6
IQw+Ja3nPfBdAjxCadjZvZbes0be8mmrOZl8smCoLre4LkpNUtL75GfFpI32wymVgu104fIUcU9O
MQICzCnCAFMj8LLcoie4lqptJnNTz/69UoiC5SsQGivLe6b6vKyHGF2+pHaw1Am+vuhLuVk2Xmjq
H6gQXaqXVxkQ361bHPSJB8fzcgDIGZUkUco30qGLGz5dbhdGOI83GNhNLwIhaMIDZFEKv/WC9eas
ulf/B/Cj3hDPNlj0R6GEGjlnZpVHuJSP6OU4WdaRhLotlKxriT5Laa6PpkvQp4btP8DqcUFhWcaT
0wPJ5cYagDpOhWa2BRlgTZ4zAKwrmaRI513FxD+VY8do3mbtX71h6CQlfmvvuoYjI1ONkJsc6Yvc
t9Y7III3vc4DXBK8Y+lp2Iwt5Wu3yiZYtvy2ziNDTB4W9WTZw5YK1nwVT5e9RSFGp9640iqQXa1E
3RgBa1937IjrxYhBKttsetehGSj6iJ8pHTBHsBcg09PYKFM7kE1zRjYywVQuNPbBGiy9aOSXQyOa
+qnGEqIC62j6msOAkjhOnxcV2/pcw7Vii/w1Eu/CxUqmhkbGXzuERJvXPqD5eCWlcygiX+MU+omZ
imCpxsTPq9bz9C+Aajye3XRgvyKVPQVsYq92yEYL0cjJJNBv2skABOU7V9DkML4t1pRdwXisdn8P
7mP2L6u7Ibiv6+n8jLWYl26c2MRwn6BigFoQ3W6zPLUmLPGLio9s11Gy+r3we0tDjYoHUVbszVMA
pyyAcbA29IId8n2b/+D3SfJNw/Sep5iploUYC5U/N/sJlCcOwn6Xcla8JeWhkNYaxlOpmDURcoL3
XzZ9Bh2m/m/iDTRtz7gzSXJgE/vIy7KvYMvhRWLcGiYjqRu6N6vob9EiM1yuMC0EAIg+zTD262rS
Q5kA/3IAdyo9cg2wQHOlX0SnTWiUSdsDvUaZGBFEjngPfkbgKAamt0CUKDHEAH7HQyzuW5dB0d+k
y/vkVYGJLL/92CJNNkOEVZzPTM0R5IF9KgbBQKPlPXqH7m0NKTq8ha168hkMRVSPkDfi04v2MNiF
9slisD6L8hDSkoBqZAWL9Nu0WaCk/O7euP/nIPf1fAHPacv7+JvnJVhU3VsuKs5I9IOcQ+5kSm5Q
TE+YwjfPoVI9wgOqDHkNfwE7Z8+Erk2YDNMHfhmf8zNXFThrj8a/RM7MOos4ai20NWk0mZKn4eY+
+FAf/u/fVN5VvJO79xCq28szFqs6Naq/M9tr9GkCUWW/WGHKAsPmL14pPPltwNbVttQvXr7lIxrV
oimfW/70Yz1VZa05WLML9lNGXfPQ93l7o9/MEz8KHUgCtVAVm/oW9K6afvb3fbEGgktv/F/RpjsT
H/7eKp6+EQ5QpolGD5JN1womVPll8GQKvijcCo86O6PKYNDSZPq+VeraPGh1zZOyDHzb8NFixVyE
BrTo1SqNaZh/9eiX2akzFF3egI0Jkm7hfMFCCmElMGlfSBqpcBggqhXoCeQCaEpwebvb54tuSbXO
7wsTgIdLUMiZx3deIZTuqFOh5q+xaETLw/E2q0OLR+p7nz63Mk52YvE7wWpVQlhWhHGzd841j5Dz
VJUGo6kc5WFF3cJ8SKm5UsHMM+hdaJOboMCPOWpbzSepLDtQ6uci9noDOuFsDHLr5r5wz364l9+4
YbgGkD1VZYjzw95QBIDTB/JaPSmZTpxsyXePTNA6BDEFGXB5irBFKzPN5CuVE2V3+hoQWpEg37xz
QMOJ4H9fayxhXInt/gY8ni5zNloEjTCEl6+EZ/uYSWyU91cvM/b4HOkROC+fAZ0fXLlz+sTdspbS
4xEF9/mTofPnh4dmMo3jVqfwwXDlrUiv9RceIcd3Uloy16Xx6iJrs4nO/aN+H5k2Z774aJJjUp3z
nx748b30DdSp//eeNg9GOniomAOxsBbt1IYi1rj4dOjF69if6pexW8BXftfk63qGyBZV9gOPK83W
Y+MlDwTJYw8lrQi6tFDmPZ8+7Ax+pxwqKnLbl94y+pfbZBs2jdNL6oBQsrdEyQEqyjWj3iQUkn2G
fJ7kd8CTXMzxeurD/Xl8lBLayIBsi/PCIu3NwLulERa4PoLycEiINb/fx68s6jcUZrtEvcLkMnUH
s3Pp3yiQIKySLDOo4n48OzRpuU/7uNrJhdtH92p2bHO7y6NvGov375ccTTGQWgZX0k8Is8AyRg2M
WBTAG7XRL1tLf7W27ahqiLqqtmxT+SlLMX25iLSaft0iJlj+vd+iUP9jOzwWgPl0N2zB/2lArJzA
3JzMI/IdAdT+8aHjXyCRyXqs/8iKwxWHSAWwevPP25bD2Uq63VrZFmwUf0jqTEkPrcjwrWpXjWR+
O8Pj8ltt7eLmoVrq6ZSWYHFuR4M5wtq1YxlXsFmqXqY/2c/DilsxeeQ2uynXZdJgu/YOaY8GtxTH
EmtjUWP57/cl3/YmOjCLZxNFb0CnKkkndnJPXAduQDgnhgVr6JAVqI3Ia+twwVljfY/tX0PwFTWD
umdvz48gJofCtS2FbQoNOj+fnIEbO3nmQhykQhpYMQrFJIqI4iEkZOL7aFWvUAzS6iJ4AWRtNf+O
9J3kyaoDogXDev+qUMw7aew+MKVl4wgRd/FaDDylsqmBRUYmjVrqcIid1MTErBDIYK0735i9D4P/
CFC/H6tu9srvc6dS93GCOOXJKf8618ygUhrMghjInSumtqRFTTqBsAL6aTsvRq0YfiEoauXujTPj
/2utjz/OFGF812Cy9AgF22URb7ggre/05lvC8aUCrsLGpKaL0SvSg2Pp//hWtYff9ZGwPlughoVA
76jUoNE2UNsWb3rnZP36/fFs3TekX3ztR5naO4kv2jpfejxZGMDBJXF0I0P//2jMyX5c3xKVmMSO
8Ip5ypIsKSknUjLmjD/19TLDFL0yNEhdzqP3QcDyoNgl6NS/lWDzmeDgtkJ3biBt1RmzIuFwixvJ
E3DSitY3q0dye6GO9On8cyFyce4ZgBoZvmptMSPQMM/wE6QiStTF1SNFpMY4FIQxEZFMy+aHJu9X
vU6g6MyBWnflY98mQGt13PALelZNWQp1wZUfIkaIzlUtodBGnEqQJh7PUkvNsL8SnMu0bR/0f0UB
Lgry1etA6NkNAKHo7bT97r1bTq7qBOH557DFhYTBBwtML6EIR4zcnctmLU0bMxpVekedDbsuZI42
w+b3sfzR0zY9BU2KtB5WNM16qo3xuxeOSXa8Q0t5QTvFo5Z7UuAg6LIVdSAYD723ZuOGDRfbQhms
ygv4dWz8/QnW02p6KzumwagY7w0hGOXNdz9MAVfMF+qHxwfk97fmk5eRjvRVSVj1Rim+Wz7jmeL+
EnXtfGU+n5yzouLElKitcecPJJtehaLwescOPIAG2bR3kgdPHKQM6TtMQzGMSqWGmQ0obI/8D/32
An4phvSasNXnTebo3YE15KphiT7UIMADkTJy0x8XG4EaXd6u9eu59s8gf7APjiev1zS7YUcQcjmC
kiVXuXs8sIDEcpiwkLOLdLLr6Uh/Bnca7YHK5VP/6tAdU6FelR+AOrpHOyL6OeHyoNjC08v8tB0D
BCjihe7tx7wrcU4AWD/Lq/c/DdiBAYdFUBGKtzRq+WzBuzb5MrdHqRMyW3EcJufhOp1mI1qR7STw
J/BuVWmZzGy9g85pn7O3SanUHjPFTavsanzWLeC++xq+oPKJYAKaa0DSxPdi5Ri3l26EveeKdsdI
7JQnYsLtvRlSMjnLG1hN03emB6w6QSINSJYzYhamkr3x/O5/WMS+Cvvdc2W3Oz8PQi0DTTgQx/6e
KPfCiijaeSuSN5zhxd0CEVpcUxHIGogQtuYtchL/TAsBPQNeNlJvocnK+TpXVFZDN1AfNoRwRccm
TEsb3IbavIRlV1R4oiCyOevhtuR2+iPchUQSGJwOibn1ZAhEaNJGY8FW6tJVB/tqVlC+cCHmE35O
ElAWj5775X2Kni7vuBceoHC4PRhkOJq+rX4MJm3ZCj9DR23USudTAL5dPgMtdQmfU3jGYGp/bdeB
ZcgV7NtUyyr1qaTQbb+vF0yw2Z339t+eg2Wx1L3eXScX/tjm92sNFBvDtKfEbswVXxaF8ctZOq6f
lnYS07mOeOrmxhnR7rCH7cAJ+MJSNevMWTHPa8dsqo2YtWcdIMV8os8mXMXg5EcRzpAgUyOZbmmO
2lMa31dNbgNFmiEDtLQjQhrJ7EpWLBSjpDMtx16HGBiPrsGTixXVgYHm+Ql3eRYA3xQ6P+N2Y+gk
cpAAxelOBMgROeqtbNK6CVQm+L4rJPNgYxTAhIM5ggIl3ujB4e0SbUx4cQ2wZNfTACWPt859KQ5v
DqOVSm7hAKSeRAWPIrAfV9LxKEgOrNriYxweG6rKAewWMi5pwtOxAznSA5rsw1Dfjrj4/U5qkQHg
RhtUqhbmZT2ZG8huwKTP9j0OGZuWjJXcdW2SNHKRzRwdKk8GT26LEDIFor3jgoQ2TTf48dU2nVum
uI+RVjFL0VfVWZago29qm0pUK9WdcXJHi+jeZVJhIZf+ASpip2w/wKAmtxcWJIE73hrM8uluUYjX
f8B+2P6xlJwQAoVLh61RZU20KF86lV3+jbvQpH4IBAwCfFBClVk0j+hOQPQcjQKqAMG1keo4ZtOV
VkBZMCzDHUEiy6qjM9S7i4Ir8S8o7wd8CupvWJHC2nUOzvJb8P2R+wKXmUuwo0YIPsntWoT4WCyp
zqftxWRm35uAgG77TfzVX/3vkEh4nx+FUbpu8grDLXvd7iHlWCDLO9jekl1PyyEgc07r5ukgJ3Ws
Bqw1W+87jVzMoUiIqMu1rVMEVJIKf0jEoYzMyW8Ij+vLthEWQp0EH9fjphwb+3iz2wJgqoUgDnZ7
JwetKhkLrR4U/d96w5J0ByhXLNh52DKHUR1kuRQnkWAsnL6JH9H+63i9Y91LRWkyUjPKwl2tLbzD
0t01eylzhGT5IaLc8whJKL+QR5s2MDJV74X6+UblfJw8Z+r6i8gAcG1wURPUF++f5a7fP3hOJnSo
gpydSsSzGVAxBQBFRBDKJm0NlTyB0e8eOi2pcWApAsHj/a+hfezxP3dja3ItIPAqF3Lx5STK9SqS
8L5XEy+ZXLN43MiqpIwj4kZ4aoBOdCFULgubBRGBSTiOcQ9LB0heMHwuKzAXS/k3cm8Qy3Z4UeXv
++wJ2uN1nCTxartpommWzsUIfGpTko2wQRKNfcRfIa+c+N1k4LOlTA9pjSwo/0JK36HWwPSedhYT
Esh0KZuX4MJle3OKTaZpeR/RrKA5bweMdh8c6/qF5euUXeMo4yDL6Cluy+wU1+c2SDgo2sia/Fdu
9jminM8AaDCKZ+Vag8CQCwoHtS0LnEmO7NrZvGQ/vZzVPDtCsoX7lqSPVagfH8k7Lymz5KjW/Xmh
dlmT/LXUAuWamRw3vyHhJFAnvIM22u5CA03k/jsAF32TX4qqTIYM5udQ3iuEuDndX9zzjltUka5p
7gaLjeJIcOWLEqaWsSU5KwhwxJptAd10YPXLzEP44/7KPpbVMxvCyRxkIl96M/41UTGuwPGiERN5
3VHmg8klNTsVZ8tM4Rjwrlrdnh8U96vrQwtpsYogghnLkFFO/YphrmOf3EwLLsadCyyErGXJ4BeQ
9sXSX8/SLidch2FAX2FMxXhnU99YIQsuHZVN0NnRvsUeteV8gHM+S2UD1loFeAQ4ng4tmBIRPx36
+paMHMp02rPNtvglfTxz62WtYmOJ6DMAcEuWd1Dwe4wyAB5/PxLfPdFJ59xdTgble9ERg6mUlw56
lul4nQCzhT6YjnhpWgSq3WVAZmCnbYXKAD43UnRoVbKMqUAUQMJm7NfLyKfW0jY7YlUst7maldzR
FY9h0RXHKjCKCwIoaMoGkwULY15h5uP2024BWDurAw04aWrlZOG28Ufj+K7bYtFtiWDIB2J6dJaS
zg1+SzQFzExuT8DAzZMlwrPBbs+wPTlgETAQoOZSgoSeKNJqpHMebBra5JN1oX9fi+1aem8s/9B7
4sNc8wwIv3G2laGbogEZO26AGGh7K5FDP4pGAsP7aQi4TfcuKnvO5+8fcP+tiuSSrC6i67hNSibv
4kbaqP2kjwQT7JjPMqC41cpBOf2y0lMU0eDrGO5Wi8Odfp5/37qlPosfchmMn15/3OXlYBfn6d/O
zBUUc5R7VSQYpUBK1hVBGLNXU2CTKp83l1oBOoSRFyqJUxczECc9tPv0cHg25VqnwXJosLBGjyDn
qKOONf1r4eQwQidDhr+RZQi31JY3VWQ5EVYf3ET2X+GLveNrGe+J0WPM/o9SXJoJa5veGVwTK6uJ
eNdStVUa5zWTV++qs+4oZwUkduo+sJkrUJPilgbOucTfJOxXQ3j+3dAafW0EjX1sBcimUuN5q81c
ZbGpv/LOm1ikW2A7z30QdAsRq0nv+4H8f5GFfTU2ph1ZfiwUArUAnUy4Jq6qG1lZyuZCqJ8gl+tk
wBLwzw+ofFhsXu1jZO8sVtrOOPOthPr9EwljIL7ylNSvbpXooo+r5pgjZo7C1F8O+Ce3ERTimvlF
x6xAcEGAjtRPhRY6Pc/4NLir1luhyWWR77tNPIenELOmqrzCLZuzq+HV5ysc4BLXYc8NwqHKHsDN
Q00GrSyNbWibi/NAl7JtL4ao/2T+k4VafP6+pYRnuBWAYF7yCYWLCoI29q7gPqsq51QwzkGi/jW9
+FTtd2XCCHc9jPAaBBYfj6UF/0y4YLOhsU58yxu5LqjEDm2rg749So2RbhiefzgEtWhzVHdXW3Jw
B3TRpc41lbGee6bfI9aIyajzfIDZWrGkiZjTsGfvyVjfvEFoODXvS8R2Dqjzuv1jJobMNDeZ0mVA
zOPoTu0LHAwIo/jS1Jqnh/CJX4JrIeVzpf306wIwOI0E0OxdfKzDnhWHieaNlLNkDPlUGkyIzEcE
8nia7t/HbfBX41Wp3Itfq2H4haMN8J9F9c1ansm2JWqRT7mUei22OMxVQrKvwg9c3A2z/wScQUvJ
EE0uIKe51uFMZceh0Y7LGmozLsUiq9zpM2Fi0Q/eVhfJg5Sdtcu2LbcHYmFh+IcYH6eT8N5Db0l1
18+cmNBye0Xo21lrMCUUDm4Z1dSB4G1sOb9NShHlWFX0N7WV3Zhd3ZV+oTPXaMss0Hzzof9FFjsh
M1gZynC0AOseC0JhgHK/k/eiYQWAz6OqfaJPrHvA7xp5ZOB/U7twlPVgbYPDhlfUcZD2zsRjGnyk
v7ILAD2lIkus0oSeCo8mK2UsSLIR6c8xVha/Pw+rlpdcoNukVs9OPtAkINnV6rIwhprYW0z029aV
6gPbsqBfYXuN2Bgarjcmt6GtDR6SHoTqGqXoihb+f1sAxHooITjS3o/uBS3lqu1nsc96m6vLsJRa
OvS+8Qab+uTpbCLrtY1MhO+pJKzZZ8M4wORlA+WL0yzE6TZ4WQ4mAEcMaOXUejmy22i4UP1eLv+I
Sh+1t4JBxfLn7kSyDTJa+yhv/beVOw//xpb79MZ9u21Mg5ksBC34DE6yWifuJdexveR8puIfQjdc
tyii1QiQg8jhmoP8Nr6fp2pMXVHR9C1l8U6xRxUPMke2tWPtW5mxbl4G5G8a/pQKVkbLimi9+LNg
o3bPTNyMFQttRtnO/nUPlhcBdAKKcfL1XNqUG1RXy/PW0XhLIHZ9qlW/UFXFA5HuxY0a+NhfztXL
QONtSjgdSjmwrRghu9IkKSTWQcSmqzo/JO5AEppQUTKZjXe3jqTvtCgpLUxYBejff02PvSdXKY/x
qm/7jdHvZmJXNgfz/Tc8JDealmpy2ftDgl035QIsMQuOGuuBfeo9GTFYHEWqlrQYBvl8rokCoRs2
0DaVrGuYwvcB++GueGSjrdLrL+MoKMmtx5f2dIfzFlgQaBhm1zDbRiflGSLmns/RNOwbQzL4b4vu
TDEaO939m4lH0AgnIR0791Tconlqux/U1DRODM5q9E1sLPY2HujtQJ7Eq84RcTaT/S9CKmc/aQPE
d8rQHH2k56IvC1mg9O3j3pWOG80M9sH/FF8ojfrl9NBtHmgMml04dmJyq01UbxOigEnfaIi+PGZJ
QK2gIYe/TqSK7LhvKhFN0hZXdy0zW9qZ5kJN1ojYojv4F+bqMD9/sNFHkgZn7dV5LFfl9ECsZU+i
buPVUI6d7q20r401w4MYXPo5P0fYAf+6fv7YolrW/8ni2Pp9J99MSCHYUF8DuziAJycX8R5JEvRl
mvgHwtbD/diR4QjP2Jje5EQVIkEQB/F3bJnsf3dh27yjVjcGxZk7UqawyBB2FnTeT4QQ2vedOl0q
G57eqR0Df6xbZsh+yj3FNVIazz7PFKpCce6QJbLsPLPCBJ6WIHusnGrCCvGg29Bx4LeqM5QhozQ9
klLUnomxumztVz1YGGCK57bBDC20BkXXxeT0QN01/a3jYiCSTqfmQTUwns2HvTWOHGaTPeQunOXz
tb0vkdK/4zRXNR/kITLLe/Lmk3fcDFp7iypzGKCtsiXQgWezCOXryKQCR6UhgwVH35O2WaKmHELG
tWzoA5EBRPrptRMFX9+hqP1Z3AS5YRRjNCld0nu1UI1P546TPNrZnlQOqJSW6jTBTH+03H8q1bqI
HDchezZROnSx02wt7NLyFiFstjrNRuyBqQzxb5LWi5IE0NmAJNEaEBA2Q5WOVsF7xNjrZwLh2o7b
8WqNcydfjbC2TMJgdERBzI3ayUWBpC71iYpqZyud+VBQH3qyqM2mOW5YyhUSZZykNGvo2/tkpt2u
Ovbvb752hW6y0gYQarPEhPTxa1wQJaP847QrPwmMjGstjUq/a3B9J50j0u71kdzAOqpn83ETgDfD
w7AqBD3Rpos6HIAANzGc13B+xJpguBhprm+PwyNYsdvPQohGwRjuGZ2QMdlXv08YyFVL7UPqOOY0
G/bKhb2LrQtWuMkl7hEmQ9MOUqAcFd7cpmtK6acj3PecySJDcxeS0qK+YKBIUXbWRPwgyPlHAJ6v
lCMGInyzOCzptHJny9WMzsqSJE5AuY2eynzTQv24ibvOzZBilcQBT4n2ChbYUHa/9JUqWmnfNEFJ
mzAL6R5e7rcJjR7Q0jxlez5Tmul7HmWrfeuUAn8UZS6DjhACAHwCXla8QdjPAqfAMnyPa+7xYeL4
4xn0Rhq0AqYK8DB35TRCyra9X0XPrPGEt1VLY0jJzCEMrJrRrPNsTV4j2PHfiSPm1t46Vut01j9b
mIRDmgMrf6e9zLQzgSGdg9ewdSLSL179VSZNYouSb85bppHIj8HUDUACPtnvab33+sv5Yi/vSNcT
8ZaQ/QRYHkb1RIwZHjmgrwsoB0ib+6Lp6s8+mmeAy70aYvddeCJOmpzujLyv0I/LZMn78O4ekEex
OjwRBMPRiRB6VCIHxlEcctfr383jDY9bclIH6bqXWgFKjB8sRGdh/Yr1G2N6T3wig0C0fhGShLs7
is3V+PSjzYMmqnE/y4JycDhmtK6fFJUnM25JOMx9IQ6gn1caJoknacJk5Udx+lhhB0eKiNQ7wmQZ
aBbD4sthUW5K1iv6e9NRFosp4pAUq11xQI0ptvJkwEKn8/ezq4BqjdCb6xZZf+vGuCRu2GEsD1XO
I+UwBV3u67DcTblUSms951dx37nOh96aMBriUXdfgCwcB86mMcyDfK1eIqo1hU1lNEG/9Tsg2ZFO
orqILM04mnhKa0sUPC5NnUa2HFI/lDSrxVBnwsu07taGny1oQi/19oGFAIHI3q5MfDblDO7+s/o0
fbz48Qf2C0JB8ZxchL42LOS47tpBTddqzX6qrFqeeGfHmiD4a3vRpMzfd81Y0s36rZk4UvcuiMUQ
lJSyMiBPqEs617SBndFpqwGNIAGywF49/kUWr4iMexppTNfZmo5nGwN/OUr6TNPMciJhYhzoGlPW
IUWGb3PpZzEr1kVTT6VtxgrSB/+EaxFsnSMMzxFBkQjSx8G48j+3T5iWBbTgpAGInqSdkb2cGGdU
gpA3MXf26CTmXSS2a/bDctThaENHp6x+afTJJUUy7+hRsTqVODZg8KBTfkDOsA+9IBvHv5zZDvSO
2le//gX/DtfaniNGIqUlCdOu2Whm4NaPa9HyIi7S8s8Pye22ZlLanwDwIEhA3NyUMGXTlzDyqhdW
fuJ2wzH5lAM1kTaiY3yXfaECD5L16wRG3vPhtZgi2zgamBV4s56CjxRPAme9avLizfJjrNWr7E8O
Fs+iixH9YvuUpKu/1VGaxJ/msd3TxaHb4YSVPOzPLHISSN549OooC5b69KcEpSjkAwzMrIoh0arQ
Ok1DPw6ftWEf1YUEQ6xsl5aNFrkCJfPTGjag2ZwB/tHhIeAdMZnQAdHtfXyaYW1cI8en60iriolv
ws4fB2G66naffbk6hRBueG6liZkMHEsNyY1LJjJhClnJoevp3ogt4dkduLm6pTeHCZLWM4Soq2Qr
fmCtdnkwhB1QLQ1LD9Ek1DseaGC6TDa0o0j9XGebYz7F/RVydOtb77aRWpPJgFDam62/KevxldCZ
j7l77VTOJXVHAn3j1G1ItgJTeaMWMTTmEIHcxyjnlyIk4MCu4Gdj7lKDG6lXTm7cNvx6YxfbNQ1C
HDdwIIRvohfwY/MchxsUjq7OdnLxVibzxHj98Uwv1IEbUV9QPznUSDy37qtsu5dXMkISLKsFQq26
hAQLDFV6vfKqaqp8DWJ1Lt6vmO0FvU/Tb5n/QXizEEQSySp8u7rePYW2Bs04fkx/BnQtsWBSNWoI
CF5NfEqZSNcukPS+GW6Tz8U2c6ygUkFUihqzPJltSl/LLFlzUEanYRspXUnb06Zf1n8OoPz4Ti/X
wLJ2BDmiUQqTspWkMjMz6HhzUcKjOelKMaYdtcjiDUx4cLhn1Vb6nMh9LKD8h1d9NyxrgduYGs64
BV890cCa7XnPAHq6Mv88MxhOhUM8e7lMd9+pv7Cb6NVj/j422c0mPSGfTjh5WNZBiwRvN6dHSZnK
iZhx8w6njlPoB0tS/62CLqv1tG+ZHQBKtcjMeB5eMdZjKcPu0VPHCCwlyv2iG7eZdBhiNSWO9UQC
4RA+sjgYY3xDqmbBXBC5YF9fkbTOFH0u/lDmYIqtY7GpKMT1/Z0goGFWYh0bjg5aEsO9py9W3ZMo
fwf0ksij25kvD94lgwX4BHVwcAIrzE3cHnrPHS9w837IcnMpXXkL2KJCMaUR2aT8HqmMz5V1fAxE
dYrsbR9Wo09iFGPNNee1NaA9b1hPb4nGfcwbVUxyYDj26zJAXtgI1Vj0VTsLo0iPo8aeQK+TVB2m
jYLDLonTip6tT3/F0dfdqpIK/RKS3T5eUfVZTpDEpKc3DTeimIb2megtpfv5pLtvU+jlipiSmK5T
AsTxuUhRj4DhHaHbcu2H+95l9G4zDqfL6szK29bQIQIbROdWE9ndND+eTEe5YoL+BWfsN2+OGLRU
h4tyZRFtU5d5IRJEGXylrnZZ3Xaf1BTM8oU2qkBn77fSuxsj4mjTjXSamNbayMaivsmSHsUq8vsP
YFwCz1da8YsxvCeUW/2sCe01T35xP2WEPe5hidhRITMuFPLge7jwpqPeXu8h8YSJP0zM2ilO7F6T
bOq/4a2KwzXBE+NGQHXXTzQCQV+zEtYqfC4lrfRWg1Udmz5QUaBNR7U1ta25QZKRetXLgjdbRwle
901YTao6yAR67ZjmH99jGPazaJCgnUHq6+TW+nEoVLckTS+mNM3BXPKv5SzSn5/Q8QO35qpfFAYB
07heQLyUR9A/32fPURYgdCYYAyvILxJK6t6/rRPVYnoOq9sk7npjrOav/f0xsZSUsVLDV8zmbUZu
e/F7gsB9ttipMIfxPMGeazO1KRcFF4pXh0fMgFz0SoQa2SGBvlVuocTYQKjhJSaTiT+nujbaqnNY
hNkhRpxBC47fbh5tusFGQw0xEXahFOtRyIKCFLgIds2r9MoMBSCc6F90sIcBC8aKBG33uYlS21Q/
OmLEuH4l4pKqvMBOvxj/WOPPPh7Y7CtLAARhK7uPpAW7GKf5icqYOYeQacjXd+bUb2G1d+lM81zP
qrYZ6c74E/Selnghk0uuLTG+VSLepoEWokCdC0Jqmn17uQGCrikWeCZ1T8Rcd7M590QTOAnLv06W
Jl/my6NKV4bJaiwQ07RfRa37zb/3kWYqT4SPulWP60bHgAEPb540YzViaOPJkA85dbXWvX72yelM
zu5f2DJYmkQd5WjQejwmTkSAU9Dbi8UdvH0Yp0eHCamxv+zFcAaQc2Jt2Pb1xrxOUULxL94JpF9s
LW51CgFFgCYBPQxE6xbmARJy6DiAPE2lk3g8OjAlLxRlDRhTuS3sTnxGAIg4Y9ArKF9D2ovPXB1i
tCQtDfI5QR2KmFhpm2ESOITEcb8n+SQL8ul5pqaUg5Q4sfHBgkYVreT0kGnKju6BnqdIphHCRl0G
+dFwAQQzrjzu+JuVz2JEXzi2qtrAm0U33A8sOLaVPqOuoOozkB6Z1W1e80DOSwPglJOvjC+jo/RV
mFt+APntS5Oc836O6NMv2vbRo81fnWMrj4ytLys/3uorkAgtVWcoLiCz9yl7QdpttL1Eqanx0rhe
5BSeczDc4ReKV140IlKr/mvacQM/58dA7kG+eCmO7wVCeGdahZPwr5oZUiGhX38RAby+bg0mV7Sr
3FHUmIXBQXOUAE4fjihNNy6DVA7iUNh1CrmLE7WMpPiHmKIxE1FPckeD8ieUCSzgO8kd4gAKrzCx
fyHV0GFHJUzDKGYQpcD1t2c0nKAJxRqbXkASPVCzrtZCJXoskij+DzCezKs81cBkF3OldCGAmAs/
RqpQR8Rlg+3hvGdPyKPbGvqzKsrw/D1wRICX9sN9rmBAFXIiLlwKwXA6tmc6uOkYRW2vQAMGCs+0
m7iFWVXFFk+OK9uz2g5nj4zolHzVE0RdCqDQTl2Bf0EMyVToJNKnnOGEqBEX2pBqwm8Lp/h/UJ34
Hj9wUy895uLnZ+4I4/1680S+bNtMaIzZG0SCY2GoGmcXoCB6IAP7tG5YMO+lJ8kCf6jCop/tfZ8+
sPxc9FGi/AeKLnJkSwBOu6vnAxj0q4/PDZ4pOExwQtFIw1uRkOyKcN+DjgTLQO6Pq37L1LMqmOj+
mUCf153WjAHEahxqa77kWvltSDaNEJPBneZ5xuJXiA4Gy2hQ5WyRKMXEhddGV/fE3zYnuciAGiLo
foP+9vKVd7StAIsRNBCgrF5hhS3llXiTd85oKcAO31UpitMFUvnILi3uLhf3piYHu1dFqf6fAmFw
COFguZG+eF8tu0WNX+0SMQBCbCTTa1y84wTA3VqLcgsX3+59TX9CYoim+vWzIZysC2Opa8iGnXw4
Gd6AyWCGs44OR9P11kAjn2BO4YEsisW01/CoUomRjQfo0kD9YBK7kyD4Xr1kGqADyZqevyM7kZxy
xTh+1NQYGlS4UZBhs8qLadidOIdYJz8EW4WXiH/4zZpXlQ9C3LHlzxQOIasuFfaJZ6jbBj6VsNhK
k34/ouuyAyKTnjwZlF1yjvu86FoTmshjK8eonagNj51aR++42N7WayxVAnYeh7pwOfAXd48dBMPj
KyxqRKhoOsVDhIz04a8eVWnWWd/zv9ftbPhCLTAyn8rkPm3PVm20UiXqs/yNueI1P8LEYRQ0yjY0
82yU7TcTMEFOYS4WH1zoplXXuSJj7apoec+OgeBH4fr/U+yKZXTmXF3bIP8hcVbfUiUGG/wobhBB
Ius4HWUrxeHx8rQS/QHUqzszIs/6oRdWCUOF91ohwgKI4n8s8+xtxKcPXEqPDcuGS+/F1qJPlbhc
wt4enFc1ltM300wQOzpXW0Rfo2utyKoRe+M4UFXGMpEJUOlLbYpVQv6wOD3jLaJiKw+XM2QSaLj8
tLvi++lCCFghxvw3uj0c4XjKrzZcut+0cvq0E39xwHXRqp0loCzfthEB6y61Ds3wn+fifi6PpXYN
eVUDjfNUODsk4JVDAiP15yuTRbWyv6YvcpCE1exm22y1tcLxUYun/2iiHILNqk/kruURxG6AqSLO
IkL8WsMYerG0oEQVS4pLYn2bKxo9t16GQ3S31pzOttdut7Kd27j4oS1LRgvfJVX7WKVtr/z08wSH
uHfw3TuPfSL5i5CxVi4c2rHktk9ZCKLkP3Mc0Rt8JKQB6ggSDM8/RNcT27nhLGq1XgwRJeTGy7qK
Kug7qTKa9Uopd8zbRsnfn3EHFG7EJ8ly+0hb6rIyBpUzsqrhsoyTGYi4eyZb/jGvIu4zrvqg4F2N
GAID8/V345LeR2UTrjxTkuQi4hAqhe6AHUbfkk8OdcSH8nJf4ndnau/h8G9Avha8AiHXDvrOZMJM
V1+GaQKZ9rIvRxKeGs7RiCnWTKwVhiMQcrtH2k+FoW9wWb158rzhVd2BmDgu08Sm77ItGAR0PpVd
7QshCBFRfFBwCgauVdJucdqi8zlHLf7k1HXRtFpiPT+pTgrtVxGLJnwBlrFnDIIAdbfmE1pfmz/A
ZRrmcSPTbxfwU3CvvWJIyIPfAPbCZzVBG5u6TrfAjWRm6PkS1eAPnf5BAZb0FWDSP2x+ITzuk/HX
IOhJ1no5YiKpi50c/z+WRu150qiz/xp83vyLBYn+xvrm0KZtpTVUuuOxN2h5xo8ZUQ/sEX/6bjrL
4GHSdaStaBqeg8Hu59KeT52xzHBsXlSJYESZ9N2l8iRvB7n6nAAegiwIvOIsBYFesOpZ4XXyPpFN
qn0jUBzk9xtGWfbeZWfCxlmWMxOdh8wkDjyO70sw/FSEiSXbXAQ1zuv9ouc6pMZ7dAZ/ldFJ7kv0
QnkNoWTFCn6ZvTOhwq9MSniEqPeqpkcuxcK2dHRe7EQizgAeTmOmGNKVJ17DRuR9UAs36m4n6nv2
DiiT0S55h0odAQKz507KhcoIWD2lIaPCSuGuJ2fHBOG6b/BDmP//08ybKk7uAFt5/6jtcIYP1x/t
SpybHtGLyBnNDFoLIdicJXgqKmOMU8NEjir4KVTN95+z59C/Qnr5+E1TYUfpJSScGEughDaxSfR2
tAbYxURNlR5H7ofmeKJE04xFVR46q36JZDyss6APdG3la5ezXqlZnKzWCJlOW3Q0k0Nv0cokxWx+
Jcw0dfV9XAPKl1QH2koFvqG1yVmAoLmiMrNkl7im9kjFPPerk1SSFQhg+38XTD+AL0qm1CQgjjnE
I4lKRcxIsNGRkI7SJnazUXEoijMsJxDyw1WtTOLWi7k3lK3mvpzD/6zwCKk+N4lGtimSE4wNTTdr
sNh+p08INWPpGi0vwCeV+gJqDISBZKufkJCj/cM/hWEhwdJgQYm2Ui11xc8Gisv4yqpDk0eWhCwr
WoafeinGvBHT5cFK1n7ZHXkPKeW72fP2wW2C/yHZcol/ICVagmFzpCOGlQ1OZGP2psAttcOwLNYS
opie9M4RYp1FN98FdcMSVOqxwcDh2znZHWm2FeDNSDiD9pkfT2DZEdDaPUy+ah6hf2LcCC+oQPLa
UoxT4Hd3WZ88T5JJfAgbUow1JY7N45si+TYAshtPwlP3/9oxkDS8YXcej+87n2zB3nIC/B1Jesgj
srcIjCIEzmxjWOqSFtHEgg+0eRGvveilZtW+llU3FIBnimFH0E4gksHSQQvQOLDWGjzR3PkDwxxy
3NRNt2T4LiXdZa3p5L3L3i3vzmjelVz4x6D11OfVZcWcZm80t0tysYtJChazR9/b9FmmeyMi3NUS
D53Pu8KfWjz/QebhGjlwefxze0dZpY1tk/QTu8dR8uINzmbL0HWpLiGRu7Tfm59c44hpJyefbW9s
en+YFdHqxo2aX6Kkk3DxaGBFWU7n8EQt/DdOiRk5U2vOyfEzfU2QJK3+cIdBwj2MvQotUugUMs/D
Ge8xyzBRsUPkO184VYsPbOB5d0Y9JTsN/6vSPJ0VAe0+WGjnCm+YOBK7KKYs9HYohxi0G7j9tJNl
A+127x2uUSL6uJOnhbTwnLwWxMTgopdOR488knQDLwsu6DuxLAT70XFzmCENQN+FMQF94arpxTu8
ZkjMVItf4LRyOaqZ/T+LfqAZ4BW5mbqFup4GMMhZ2fEmvVZB72FS1IR9FXTcAam6gVhQXFn4dvwK
XO4/w2NFHU3jwWGkiDT9XadojiAED/l0sZI7AgNz2xqWgzczIegPOxLyyS8kcA2GPPNsvWVIyWA1
OknkAxWVkyuni+qK4Hn1kH4IVcsfIFakWVuwej6X2+iP0piumarTkVeiTOur0+Tr+LY/6X2Kuzsw
xEaw48fHwRV9KnsprfnJKH83U1b2OCqz2R1ZN3aRlMh1r+TG5Wr55btJ9HtIEVmTXo6AgH1+20el
V21R+nouF8TLxkkA9usrOzfyQMTQa0wl+WO7QXDHcWwczu9+IRNU8RoLvTURjB9x7TxQYNYgqufU
XOH4RIJHIYDNdX918yWQcafelNoYKeFT/MrIP+YF2wdxLQ3Ot2vaHqSrkeD0seDHTki5ITosh/9N
R9JktVxvpxCr02Bat43gLimaNgwCCKdetUgjaAEQf6tgSqkL14Vc64SL8EYFs3jzymQr3QRpHjZM
QZb4m+QVSHQSJBW5MwS4p0KYPx988dJ868KMsKGQNuF4IvEdHZ7KYo/l/oNB1LZ+L7+1QO2FisO9
eqgS0/iGLkdsx5nFBtc+ZWeGIuoGeXnF7C8gp359RJY+sK43zIHmHImlTPtq3unWnG7ykapnrDOC
YyqB2eYxG1r94/PcJ9VgSeRqwt7lKioRLR/mHP5OG/cHfvjFHfRmcD/xxiPNv1GjDtFhPTv1qNiN
/PTPlUzim0efyGETkUBjO5vMb5FG0ROwgXz8BdLN5hx9hN/eTe/vlygix4Vh9o0Z2cFcRs0lXXoN
fS4ahkbfwwWlFw70oJ9FxvrYsrE/E48Fz0NjDep2eS2CCc628o4dKdB1hOehEVZ3h2DDH2ZCJAtd
K1+9RwDAU0b1xlC94WRUIZmZMaDh4N6gX8dM1R5WRjr4HNt3r8fBu2Srm0UfH/KRyD1D9/96W2Cr
H4zWiqFmMN8D/JAuusnxQ4kRVgzRZFPHY+ou0dqiJB7ZBJGl+TICbZrYfhOl8hMuE2OR1PnCUjcT
v1gy+buMQ00ajwhyDXk0uts9ybdxC0x43FzPDPakl/85nw4DyNnDunfmQ7GTo16+zPvaqg/oSzGt
MkNNHpYfD7SWjEFTNVBIqumRPcrFm13/AU+8NqXyeOSFFcgz+/gKv21S4JkPpUMyLfY4JZEdKJY/
01RkMAM/7Fs9ZQBDlgd9oZFJgUogK0Pp78QWDYYFoG1Mecdv9yfn9cTUDAciUgoUBvdCU0aPbgE2
HHTt0mHe0LBb61/HyjPbzi9P7izhLBnE/p1Qj/NQS9hDFLyXOqqakbB17slN+6tqUjVH2jSlL8x2
H0GGvsCsH2Sb0SM5AIDbz2eH0aph9KY/cJ0exMvSkK8dDUHIPg/yKOdEiVZEklAhgBUEy3eD4OrC
KvYBcdIGyO3onqZ37K9fV4yeEKbjmRGqiDJ0eOitIccF8ZdsLH4PU5yFRsrb7ywar4FC5RXlqTi4
3KBgklvn7Q/KIUIKUqL+ZMMeUOp4x1EzXmo6aPD0nWJ6VldvAeAlGZWc1Nt/EIzX4IhXeAQ+TnxR
l8zbEjkxe/qCIE/4GvdNJXx7YWicuxBr2eEwpUmYLjCXHLIxMRgsuVGReTdVdsd/QCNUZFORhIuL
b2Ts/fdFlzD8Q1trzvSNqxfpRbsNJA9NWXDGkQXGs2XDYxY1HUfwq+6TW8+iz87+SeT7CrwRMXGb
f7qEoOnUSg/oo9sAsUMSzLKIp7BxJMSi66ZSz6wTa+ROd3ayzoFAsWjefFkJ7X6R50LVPFGnSfdt
K65ben+JV21Hr8d9+s5FBDPDXkUQ3Z08GEQFk2vIbwQQgk+Af000zSQ500F36d9OEXtlHTRRhu4E
PfxfSPOMux9nADJ6V1XgRo7vrGMqZJzVPuX1IDrPq6ZOsrSvxqpHJqGh76F5uLxeQExRYV9thIaz
T8JzE8gOUlD0U/JOf3fYWI3KVd5mpJko5tfkoAFioFapS95Ce/qE5RygOKTTd3NYdVYMHTvchHts
/6a01mj5Vd+5Ra50VjQ+NCrChB1iSaEnl0yI6VYcxrv24mGfoaea+8andCWByt5ptx5RtTF07VXX
YSRfMgL+AVNjzHAzHzRAfpPixJnJHGCpDucn38YDjUfRMb4Wm1A6KykLCopEcySddZPhmXJ5T4dH
UerFXDeQ0q4A/m+aeA2NSW6l+sfbNL2rcxERzYa8lDFCcOsQzwqOr+haix+2nLQFXwihymlrmNhz
XMn5JCouS6gWhYcvMJIObOFcxlpom5yAC7YHgQQsEXKTwF0whpz0E+xn3lIS3eeHMfsbB0pFyT/b
QKiD9xf3bbMBWk9Awp8dMlNzFTSuc3yiFw/rVt259RwOmfyXIHf61iXcujXJU40cfNWDdWf0wRtG
kbAR1E/kI1cmQhGBSnT8xQ2SwH7r/ay9c0Cx1nNhLMAd+FP/IjHxjC5wLXVdJWy1auhsTPzg756k
CsiEH4Rmj9P50wknYYJ7OQzJPyO+9Q3+zS9depVB409Nuop/XZxuvE9cyqNPU7FwIeBNo8T6dUP0
z5661sfqTM84ml5a/IQ+etKam088IX9NElUta/2VEptZnBbzwRNsfW+ZQcgElCoAIj50mYKk1Jdz
vI02KuuHl5FqYTBqYgL+3VH0+5uG/RP7m4m0WTFljPaI2/tFtnRoamgyriAgXdZtH1P6cYcFY2nY
kdyjiiXdTAgYmoM24HKLQDFgYkCZGGSNnwZ/OBmty0JE94QpiRWIx7a9Ayg9cZHxgytf988t68Op
CmDGQf+D/dizTCI/E+picZ+s3qoikKrP1lUoqD4qtUdpDx2duJSKgcj7NB7JJdUEUT+zZzpXjjcI
QqXEXSwaE9LBhr+K3Q2p6LZmJIbtIVqiDBo4g5vK/xK9PuD2Insy1UDvxHTIyoCEYj3i8kviOpel
Vrjcm3mAOcB7X6HaYwlzhPOT9ctJ8Mjj1lRTM6dryDA4Zn8tFYhIg/g+wZBd3RpJ8GFLRMAtQczi
8s+8B+OVl9AgA4ZXVsjmHPofaymcrR0OWvm5Ug9cTc//qpzgyHaAj1ysejF4hAOiWsMmXdEKCX1o
Rc4hx9bRTkWOHBwJr/z4gcYynJBXwGu6HkhOK4pjM3BeQPKJeH3vIZIH02DUL8a3RtD1d6PSeYSz
nn1WCk2bUfC+6L1o4lNljFqsu/BfPycilQLOZJ7KLgiolUPwGAEn5sDu+5d20dTZFzj9xQsTGWaW
9Ti0lh2jHKWjZBASpUsD5EO9AqJho9KXdjAnEzXJFMnAjYdAOoxw/o1kXHLL5/Qgun9FjTYfUWZ6
+t2tSk8VIP3q4deUWh7ONQsKAOXEw4smdTwjZureea7b/lEgUr8GKcPru1SkCBsY5qSlH1iH99Vf
pI768Je36nKk4gvE+sV2Cun13BKuiUNJNZT91RKOIvLV7JfKtkXdaw9By5PMk/BH45dhlr2BlbDC
2eGUgOpdh+UsTXzW2bN4Nt/3oItheh4pBbJv5rSfPBYRsdKMp8e60yflSsbFM9w/fy+jStKSuq45
QVlxK+fL5PXTLsDDmv3dI3gSHg9L0qxZ8P1S6To9lR2N63FDjN93d24QOqzgsWQwdRsu3LLdKlNG
Y8O3sjA7eZTi50MrT/wnQp8Doq93ZL+jZp5b7oyLgeFfbZY8i/q/4vN6Or6bbKpzmBxoJTeyswVv
JeFynsWa5x5RSIie5+Li7z7ONTO8xA/dhe/ZJaL5fI/Dm1YYjvCzMR2aZlQ7GpEOpdtA11fHOZuK
2zG3tJhyx6l9DCQhXQmm8qimoeM7T5/6Ky8stkzjFQ1WdTTBFlkzzbHYisSUmI1iAGDBxwMe4HQl
TMy9vNVuMLMgd2RRTQjgF2K721FlXiC+uaggbMVNuodGByDFD49UcIcCMZDnil+4RxOh9CnpR38Q
df6BY6Li8c0VSFh3lE0rDTKoKIG4SsaUd/z1J1xpkX0HmLGpB0rNbZHnL9MQ+wM4EsJ/iI1xMJwd
XuumK/vca2sSe91itp2mZC3pa5Aqmuasd2SCbIiC4Im8JAFkRUpsW7J0fNuAyVvTTlGnbfLKzCq4
hjAoluZ0ccYgp9bLMSX/6QiiuTVKp/2lzg5w9KoBmLTjGFYAy24RgDO/eiZCBZ7VnjA4DKRvNIn7
VsIiDYcy4sQMzvegLJduU8MRBdAJAg+vRs+pHLJX2kgfEMO7RkhZFKj1ncih9HcvOnGqRCLobCqV
Iij+4XesJmUsnRDB1kG+C6HV3F8KX2/Z4lreuovRzn5/vjFCrxyj78b4d/tbqKQf+2JMAYj6cOA4
S2UJV/vTZoOo+KgBKbHmmHD52rKIQkn8dbEGB2hOs7pchl3NQkYo/9sk6OJO59mG72ecuBKXRDZm
Q73HbQGWRQlvGHW6YVSZShLFGdxSUTjy2B3Y5otCWSA3QM/h0TjwpH1iiED/wOY9ZbKB6RqAG8kQ
+/W6/YHymX2A908Vv5aAxO/cWej1oabQJmPXWsJPDBT9hlgYGFGkvCv21conPWbkNrJvPrIBRJPn
RaOsGPIVE8H7NCttzjfpeQdziTbBIqq/smGSpp+dk+Fj7J1xc9J3sj6vMx+NCmgcsyVK09ADKmqx
JiZp9ujZ6D9WfpQcLuUDkRrsSI/uukBJvnLZtQ3yvAAbVlLer/JrxEnCZr2IZTwM7Kf1sbZqLkF/
lNuDxcKrLqf3M/OTvNltE1f5Q2zHsAUI4MVFlRisQjREPkcWqN9aZLqAhtQBvifjc7Ok/0c6zHSz
98PS0OykbBYXRTKbdZJyFQdaudEIYGQLZJ9I9CZIkHFlb2x6TQLtANTTcUwYS5i+rr1pABGi42q5
pO8zM5u/gFbFIQHTKAADhYss3O0n4R5a2h0ILK3sT9gIyWf7WxeIx4supIUkOKyrHW+w3QZdq2/f
H9LY72P7BxVnpMMD0GMbaJCb1pI6p9jFGTUty6F94LH0FrkU68q4Y1GSHnWeAdVHeyz8VpfpWBYz
dK9gXaYQGlIydK5HLzC0KcHicTr8nf7vOBt5tXBmHM+H0JS4RPUGZkxaSnlfdzZResCel1X8crkT
gdn9ZsHXhXTnUUrix0DOYknH4jVnfJ0TGKwJDHa2DcjPTwrJgrNym/cGoI2Y/hdNJErnNUfOGWcn
lXjDx9dU4ex2kbqrBzgltqeLLuz7rcFTxrGVeIqfpEMKh4T0V90RX0mIiX0PqFbgemH6gtMTDkFf
uqs6TlY1YWu4FxxN2jRYsxSZpzXh/NNWnkEa5F5A1+byU87vFmeCc/hlS5Zltbvm/APU7s6W+fNJ
+zLexMyE75tbVTFl/w9MemDxo7oto+6cikzd3aVsJZvVmCReqakweCJbBhnxeB54dDAVDbgCKOnV
8+YOQYgBTOCYvahLMnYgjGyPWT/Wp10WQkNjhRB8sI8ri2QO9qgt4tDG17SREOM2v4dWwbDxXUNQ
qIHLg3NV4tryWTlxyiLYwEKpYO2q4kebJBIRTOCQa+dvHrC8PLNNj24NrlAjDkiw6WDWJEx1v2ym
WTRalILkd1UlzjC9E21RFR0kRZJbIwmUKbsBqbVBuEDvko4yP2ZNhnXmP7utvNnw1zmj8tENot4V
lfBrFdg3k/d5CyJj2GwqUoMn+xB1yDhqh2ToyJpbTzHLDj1yFV+WpinhkeaBnOR+L+9iZ13DAVj0
in1QIpUeX6yIUlfiuIyCpwHpgx5qPYHdUE7x2WogvBxfkztY0+ltedJl/MLXoP4mfHcsT8q5jhtm
VX88EWwZ38NflQ40QvjO/VVbmr/gNGdiXnTI7d5HVFjX2FszJK4BYYMDGM50s21D7JnwCPFwGWeR
QqJ31+DZOY0PHSjpNV0NEKUURSI/VPpEs/FSNSzy5CqA8oxSR6ARTS4CxpgdGi2RkhEuLGE9mkzJ
Fu9pnuESpb8MlyTx7mCPK3glfBv0zvOn5qYb3Vxge1WXqPeEyDupAWoyADgSTTYIrnACzIaZIOtu
6yxQLRKTcF/HO+r/lXqPH1xjnYxx2GENw5lOae7c9+f3VQ5o95PFF/JbGi+L0n64nD7+RZ/D1Dec
djB4K4JLjwPwM1t6yhppeWhXy3xbc1KUiKlbQZ7EVdICH2W9eLo5WrHUsJrgCakuRQ522Bu8/nHy
Bxcm4/K2Qp0Wo4y3zB1MLf+qFcaOURTpB9XLUZ3IU5+8EJ3Zf8388JoX9xCQMzSPkAq3Vu5Rvp+L
QnjqVHMwSehPaZ9uFbRXXXG+MsXq6igG3ic/CfgV4eiCxUih+D7GB08duc5hMk4knbrL1Yw+zl25
tHSZ+SbE98xuTMD90EgGPYHT4GUrdjvljtMH9io/JPSdFyfoVKqB4ApJemg/0M2zZnzDM+tfiirQ
GJ/x7XM3jC5ynSnSZdk99E7JSAPrhCq1/2T+iZPTrACsbX0xnpO/h2Pxco8wyfZ9wGZAL7ITI8WA
6i1bdyAOvyGWMC4Qpju9uAX2HOKQDtrWwk8Cnh1hDU1k7a68fqLeYfImxNj1wegK6KvzYTOKUyaK
9Vjai8qdxjerszTYoaItjwm9UYrxMIMBuGjTXKVd+wHLLtM0ZpJzLCTIgq4Heeo+0EwCcdf6s6mF
fL0DL8v8HVGuBRS8RMHUWlnPjblubxX7OOYlAZU9+oWdmISaGCvL8RNxa/tD1PuroybxfRmwxRH3
KtBbPTiQqXsyuCvhATjBD5eMWD3QcDoAK82Sb9ZqMhcJ+juKvAfERBa6jrTFFrb+savyW+i3uO5F
ouAUBTdvkFbZC0Dc2XFeG6aYF1dlpUknvO4Nau7iqce9plc0HmXpISJOpeCsT4nuTcMKr1b5umC8
vYyEpsTJmVsevPuCwClrtdFPuEFLjMutCDtBxkvvsc2A9gRpvofb/Cd3PyJEDwMXBarQXaihIXjb
FDV7v5vVgqm6Yw0ntucJO8c68bEx0e2FAuAqC5aJ9DkFbND12vGkKE++jbRUbARI7nf0oylTj7MV
GLD3kCpOl4gDhRLByPlIvAFZYhoDvqplfxRWjH+lszWcCXl7L/Tk6A3unmWoNO6707qd/12W/H1x
AjenCwQ/p5RVQ02uWm1gWlEEnVzKI+Xmcu8fOgapJeQ22moOIB6r4mU41SIoVPitjACGYhBzrEm+
m8n0XrUpeZGsi5al5eJOpPOj0V39LlbsDBZqJ3O6ukHZJcWnj+IGtZekNIFHzSiHJTWe6NDCNEje
xdjzP6utfXOSdVwKPUtjMJBzqwu7EbVvAVbUDqiKJr39eeP0qijGcnxSdVdfW9wJ/p6bfLEKXviB
EH6jWvYY8B/4PWUTwUEuaCuVx1Nh83ukJS/O2QImaFsGgU0wvgCH8Y1xnfRAfDGv/N8f8U33bikE
6SRrfWJpHvOv1rF3N+mCSYpbeSkMTttgKgWgA8iZpljYlFgPeDe1uJWHDqFySi3u8WGbSp2+bVES
zcP60Endduj6V74O2xOfGeqyDFUG/x7hteC5ATht23v3/q1xMFOb8X0xAZBKaUaU6eTx7gxq+bWR
zrOXv08Omaa/YzKPGbs5MZ+XVvsBOEPKg5nn8iY0OX40lIGNMtrrwIy0gh7C5eGnz+hJstzfKTWZ
GBDccBj8HPtge06U0F8JpnL3Llwl3+ainyNxMdERL7/zG5D33AWM7LkhvhRuCjtMl7iDmlkJb/OG
aaFPl9z6eE78qfX40Yh4DofnzSSsf8UFsVVnsi2c7yUQub/yD/4Re2JN7QwF/asm/FJxzjL3z0A9
IyEFGgj6aJXyybcYkhoSrSKN1c4vyjOBiABoOdN7ikrzuwsOFE32Yef0a7DVJUHy3bVhAl0UB4OJ
DuwkWInZXhAQrS4GPC89a4+4tPIZcHpUW6wpj3J73xkHlXhUuqrMS39lKrBWUcYyFHdVfltI8zkz
tsKBhdemr/mrqEE+3qBOhujxtcPP4IYhnA37bTb/VVkPd9KabS6yHExBbx8byEajGOw52N7U+cU7
Pbjo3oP0mHQjKytOXzwbMzJ89yFEthqgBYEQhFn712myJk+E+/wEdJwLa93UwAaEZT3xTMwpC01D
JAtVNfnJCFBggx+a+fCjggPm+SvAkIITrMp7e+WUAIgb8siNJjD4wW8Rt0YoS0fV9Mnv7YvGqTkG
u9Vz6KMEM0dQIqodPq0EZNBaxiHpJuKFS7CdHnq2VfLyPIRu0pzN/zpxOpj86nM+cg2O5Mmibosa
WH9orFJGXc/V4Sr0qsJpRweNHehAzRIZGE/E4wQ5M+4SXyvX5yLTqUva7HlbKB1997Q+zKAU2YjO
2EpDtDJRz6Xz5p54HafbgHqU3Ne0ocZKwyEhmGcaBspsz7dNj9Bup/0r4oIZVGiO9V8ULnXAsRcG
kw5YeELwXG6R87A58zXubbRQxUEnIDsmnD5gfL4VDSvPrLvBWAO9e48VQZn2EaMFLaCzLg4EA1b0
ZBC5orX1YhLpiSEaiFHg3nZOc4buHfsIP4Y7CCl/fsFXW4wckYdHMmaGTZqMUvxsgZQ0X619Xfmk
i0SSRmnp03gQJyUbY622S6xyyCbOnj8EOxCyfBGAYYQgzFZOa1sZhIUZsfBhduV5HzDBuGgubUNJ
XtLdREhmm1fz9M5FHViF+KLCzqG5k6x9LSnJsziM/pH4tAxUQsj95LtPCimG6YZHmOoq5z6mZVJr
Tln4p5DkPcRCk73YcPx3s7e/qHbcC+RpysxuF1NUvs/D6zOp4uHZvasD28C4k9y33azkNJaKE2Ac
xepKSwKNCCdlSQi03oxTT/uO2c+Ld9qZUekMlpTMacBwh0keHkj3F5umek6N2ycmnLJqmjWwRXn9
60Of+2VNpc/UHlaK/na9aQdxrkfZNqqXGKVW0u7jz9uGFg996TqSfjdtM1ynxKvs9cdNn+V+7e26
eVWBIywJtWVBhZTNotywijkS4TZLZF4/hWsQx/frpaJiTfGI+fe902UiLEjC2AfZlKjPRisuv7KP
Rz7lBsj9lL1BQsghmAbvlmfy4zOHux5hmTC7qOE0r2E/OQ3UbiOaS/hzPNk+xzjKSNae+wv6WpWT
1Opuzpw2cyeNemIccjw6B8C4R5ezNthFdoU6/5nRqL5p+/te/Uhp5OAuH7LCWPxbiyju7GpBydWb
9Y9pXA7J0dfBESRrKZw7bLcGefAJCUoao6HWzqJiOg9UpjNUX20Y6zHJQe61oXWDNgtLKeRa3bWT
F8S6I/ArcjyMpRteA615pWgfhFCMmNg7uiVfxuRwx/U1+Zb9p6oktdRmH2y0FxKk51XiDJIFE+KO
VfLk07SYssmcMX4Dr0EAmz60kVvaZwgbzwuqQegLcK7NpYkQ3IF+HdEd7CI0sinuy5gIDKk62s3z
Nnk+PkaKN/krZ32YnHbOscNAaUpjMOWKGs5gnUSCno1NQRBKg9BAqKdmM+EaaDkzvHeDCrdoBETm
qCVL1VAB1GwYBbWRv/9k/QVF5r58Y9My4OJdm1IWW5qHwpouZ03hcbD4zNc8xOjtgTyirBZglZBB
Lk4TzB/irehN9KZli2zctSj1UeX1DMR756+j5SDVpR52Ne3/M4ADUh+7iVZqMkARGKLz1zzzi0Dz
QkYTwkb+P5qSvvA7d1ppO4FKUP7iCuxpAzCJAnE++SibQxcXOaRb3P7ctdXplnWE3Yl8fVsdqgak
49EA1WXQHxSJhiUgOiflMXAVC/nt5cz20VLAH9wCU4MLNnZUuiNae9FA+Jfg17U/qM8bdsJZg27P
rzfWl8KhFjlkeFi0mBR99HGmqHoF8mfJd/COd7s1NuZOZiqiNpN+y7UIK3et+lrLsN5+Oo4HtY5e
rvyzKiQqvqGL5kEx41yCE9REj347btFkYMthXRWw6EmYqglOrCc7dcCm8xP7K0RvJquRJwUpCNde
odlQScBfKjs10xCcsGUQkQpoo0EmGGCFYzlQB9rSRSZMNKtfaEmDkU0VR/jfwt+Z7oGyp0nwBqQ7
MWNqAVYLR9HfhyaNRHfPDp0Yj4YDgWn8wDR/dziAeI1I/Bi7lL+ObUAuiapdZ6aFU3BJkAGE2TZu
iq9mgb+b47Z14/dTVTGw1OdLFsAYnjWfXJsirVcu1p6tdLtn7gbGeQnVbFDjIoTqQVm93anQSomB
rdATwG5DOow00hnLospz8TSYzXb9Jy9x46Sb1Gu8GqeS1QSwAHTjPhoyBNZLATt3ymrLDykWf2XJ
ddA23gVtr6BrdCRDrqIRVBp3ivDcv4tZ1WFHHcTquS34r4fZEEF0gDGbRZjEo7kv7CYKI870pJQb
RD5pinawMOr+8rYP85+DIapQQ4z9Lm6y0B0U5s9ExVgZD7KQF5VuOTnnIXlYXQoEzvV1FL1bn+sJ
yyKRMkWOiYIvlBlU7Bz4nUGNBGEZYXglqVyi8hf3ptyr55fCPVdTM3vvBoMgFqSpN6gKmxsWFHDZ
lsRwGHPeS8LXI5AfmsgNiINp2WvbOO7QVnCI90GdtQwzzh7EuUgQv3oTugkBlnBYi3FCihyKsESh
DEb88eSmcY4jGWjvCSPIwwmRMhgb1lDPmRDAiG9foALXC0Dqj5J3bopX25aTbnOjDhoDJkm1GSLA
OlIpnyp6mDSllWTiIu+eM8+fdqKG8ZSHxLJmd+MDCTnHeCn6G+0RT+OLK0ykrRfeVPdAnFOEDnHo
MwYC7d7yoSQ2lK0oSuTPxpON5EMqJqdNNlVYq2PjXG431Z7ZsROyKKHw0SHd0C/vOdM7MWhs5Mxk
mlPsyNOUPoBeOLW0ZY1q5hwjSnuTXKAsTgbG+lmoIqx/JsOH8onu+UwNfIvBDRq9eI4258UBkL16
n9FJDOibELfAyQq25/2zOJv1u4PB+YFAXZcJ1v+RvmPRFyQowsidEL/cBR/qzyBAm7H96FRwTUEI
0iCruRmlXiVpAUSnJd50+3QMP3Aolt1T0yuFffPkt7SX3SIRWFvqu9fVHbCp2KCU+cZiN/2Qmkgg
slRO7cPR/Mhq7u9tJqRW07JY0jXMVDopVjckSkhD+Wk+9kTX+Oa2n2tAqXk2TepwKpYN/2ZLcLcy
VUpJ5ptFag3vSPusczzhUCiAX9snAD6nta5u10RLisiSSHVYdRTpGKc1/S03+tflaS59DHNT9s3A
6yfvJDCubdYthQC7/1Jbuw+Ut308vqEYb6ZmYHcJ+Ain5QUMErXENS6KJxLtPkcn6cU9mxD6Netd
z2YFG9M7Fa3k5AOM2qt12DAGoImExCbDmSFx7m0RyzlcnYjzNFP9Tfhl8rPSuRo+5mrSdNsg8EOb
afICIojGUu2zQS/zrqgo2eGmxexWD5TPrcu1Bsazkp3uUx6H14OalgRYKXJX6eQixGE8FR4s9xRh
5GTPdgUHi86PBM/rLLUMQM6y+Cjoi2uWzBfqymwIU3AO31IU1M6WgltaNEyA8E52ZabPoE7dZ1tD
l6JW0cjtLy+ZFe6JinEAEpHIworb1vZ34f1toZv227LamQMfzTJz2wHUMlNTEtjac9lOkPvCPgIO
usmTo4lDgxYG17pN80OSagYbBgc1oCviLny5VHHAFVPhOs3ME7tZityN937pUArR11G9lMaAa3fG
2oBxzvjHALzNhf7xAuVgbLaZvpht/pYNFUSAx4yLF1YHBcab3nAstwWg3ZcE+Gle19RAAU7IZsIt
eFAoBlTBUmuj0BpRF3ybgzJqwtJZ+/yPcUy/XJZPDUNcMAKZ1jpfwRv8fOloH8vMJ1Jbey4ZgTPH
juUNxu3mtYFfsxNUWpiR02wgnGt2cTu7ORQNkQQF2hWhJ6HIn7cNTSkldMRhgE6HN+pz6Ia2kbBs
zClxgUViLm6xnDGXUkyBtciHYw1PbiKDsJ3X+wkpNnEkoXgW6sNQvOjHK1HU/UKMEBFMt5Gm25lq
+9R8oLcHPuwL1iwpPMWVZ8qaJgkQNn8Jn6aM/DizYKzWOMvQ5i1pCdPlqRS8VKLKrflHYoD1QK+i
zKfnb+OHFVrtMeRT/9mhktzlutwQb2tQphZQ8qMFBcadv817GlNwx4GqCBNPC29FXNWgAImDquHZ
KpaUiM05xcYSg/y32OohGL+FGuasDUVH94a2NMwFQqQAOTBv1rV8dWT+ywxWJgQK/l/DQDVi1IOM
6mVVAYPvGhxYxw6m57bMvbRvBiACT7RBtUDtG3wPMrn2J27G5dkvE34k0nRsnUvgv5WJVoOGK9w3
szmJEsfVefNrwSigIXheCUQgucxgXcBkpLQ63vX9hzyiexkEZgvm0CF06D9Iii1wUZELhV9m4/FU
n7xUWwXNfnKUwYKMUZJoLMfmKk/+hL0OCl8kN8zNfXOTVMHvCy1JbJKARX22WqPV8+Wch9GCj4C+
12aou4ADQuQFpwQGpJ3eUOz0eOsAvjFV7q1czwEfC+uf+X1nY7Xbq55RekUOwHzBJWLP2Sf/wPWJ
XodVzBJHuSEc/jxGBx6YgJWoMu8QQxaNgaD5/bfNmU5ZG0DDggzt13UGI4UGm8UL2SRvrYqp1wJV
54TsJbR0Neyi6QkQPGiCDAcEO7K8d9QNfm4RuVoSlBkrv6pISAiUUkGfCeGfLVzJRYLv4+S2e747
pMEkI8IN9oFIz0k1EYGXW0uo3BMUo56q0vC4qx+bGsB6ixAk0/Lp5E6yUaxyzDThkW6b9KDfEuku
5QTiqnmCDn6Nf6KZYJZMFuAYhlFxAJqWWWHaqGGfllHNTvOs+zuMXP6Gg9zRjpKy0gRGFc19DRky
ug8ewyvtvF2CkvY8RgmohdOGOsA8Nhi9UBQNThQavqAOJQGtRs/OltXFC6bGO6EMTVbKXRl41xGE
LhVzi4iv6k4LZbIDYO615OiR6h9d+rJ/AdAd+NF8fAy8hPE2DTOvDyeNFwjCccrTD+W62K3HChyO
uQWbA44v4CC5JaxbQnk+w5cLUvEpklm++MwqH+pkPbagVSlt/OL0CLXu5PDstsjYLfTOObjNevC8
kUlqsbnEm2+nFHlQdBMRz8i5C+4yQRFi4/+3aRKf0BBw17FhBDvnwjkvJUzsVItrZgWXUOQAKrTS
wgDPLY6s6BSVKFWsyyiqgBOx9iG6PiTBYtS5iThBI+88FtfpJ0f+6GEnqK5+hywwmOAxK4KSzGgy
v6VLX0iETRidhjxj5H2dmWZ0WCNG9AXlleMsascQZdiurzGb8L9AVUcQRpEXGCdZBXe7yVCFw8Ne
7zvcyol3V5iQCKwQsW4txPGR+2QXEQhiNxMNZo0BCeqjHUUt31Y7W/9ZKwFae+zgnUMxenUeajuV
K3NQDq3za1R0K2qHvlH06EryRRrg0VixOjSntHoU2XCsvfZ/s71NDrY1USK8A/WQhX3eAJHOJHNw
jvsngNpBc8i/oMDQF0FO57h17EL+7nSeTDzPY+8Hh/Arac+nzAk2OxcFhkOMmam8B56qINg+8swu
v1c+BMh/KJprDOgeZzDipdWnao5NXRYs+rFldJpbzP7DB+OMIVRdVyW26hVErK4sQvs2qT+uJLcP
CdA6/SNQFLN6RyI48Th5lvt0AemCwTfe92ZJQNKT7bsk5Xoxa6Hf8EihU9XpZq9phw8FyxUziRE6
UHM/hmCUnQGpdVWUKs6GpowBLoe1ePFaE6R+1JGzhIP3KwFOotI3go1+AFLiusXOdH95yzKjFjyV
H1ru9jRpEF6zaNdKcKjagZnPvw/E1VbbZ5dMlKQbPf5IodSao8hk+g6SkGslOFlSXsT3XwQRrQON
LNuz4lhto4w9As0UStD7R0d3JLYnFvi8KgMuSINt2R5L6IuRyXnuHr+z8v+c9RHUNtPBLSxqLm5F
7eaAF6/dTm0TA6RFbTuWk2M7PuZf21dK+DpvN6ucTa1lw+7NrxP3CSPCD4BVKgDVFqbTpqSe6eBe
ZSBh6orlCPvMag0odKw5O5eJrtMCrgkpT+otXUxpCgIaNC/mOcWFhFod5IQvXsgAgi2L059wFXsX
SR1EI4HMienZZFJFebYokAN2Nffnf/7U72jLe/Wpox1pJMvi4ZPnO8QqC9je00On9PUQz2BANtD9
tZR2cm+VetiII1wA/sldlxQT5KYMOl0LI9j0SznWPlTyqhtKxs5WJwb4l/h4ZJ/L1axA6TEJDKch
gHmdFaZr1O67H7Jbut5b6FYUOofyaNLjqP62aRXO7l1oAt+EoV7nwNfytDUxrZ1p10dIc5RTQkmt
S4dJwa4Eefps8C1lPBlbg6aL1lVxHscbdqzIqbiDZIrr7TKmSJ5W/rzvnloTrna0LDQevVXhHeom
kxkZW0VJ53QS1qHyP2nv34ej1VqGt+E0sdWbXBY1wHXtOQpJ7/5DLtVGjMgHni8Cm9cvOlUGSiFq
RbwL8ThF/8j3ptsqsDzj5cpMsAqrDYUyRowH3Ad0Big+6FAvgRfiaAtKakOERMOnE8pO2+8FFI07
+GGHYQIoddAMon/PteJShAfi8+epp+FmTFHUeYC0VUnVP4mnN1oLBpUPGbWGy2eV4oX77iaKcjny
IxpwLZNh8x3I1/8wOgosAOwvFKCfGCVx6/ETirObodiFo+xzJW7plJfyTOHvP+oE0xhLMOy9voM4
MN4AlJeR7d3y+Un/ypIQmhl7qO+8NtTEMKElDGkh5Qc5u73A4vik48gv4hfU4Gl0pKOjlXEK86Mt
c/Ca5w9OluZ4I8F58IoJPqrh68HqHnlTTlSRT4WqACMTovPW+UAKWjCOpR3w1u0OBdJkeY5N06Ed
CzDC/SYXu7jF0MxAQ4pLfPSE1cc+8CTPEO/zboBH8F6H0dZvoTNUj7bhZl0AW4Vf0wuWSKJTUjTH
OaPP0ktIHSMt+SSWls+OhNwtmG/hdQqY3JWWRFer1xPBv/++fpOm8jJ2yFdYQiXiNFU7Z9Lp+9+l
u0Kgff5gEw83k3doPEwyri07BjKOURFOWmdcyzamPWjzcZMS0aK0jmKLa09/7hKzTe7suh4S8j2J
R4SbPPMd41gG1CByzYQKaIuNO+5B+zcWOq6x29swD7ZZkeAifJc9lESdzQ0ON2CEDx6VHJus+xlA
akEHRSDE/CqGiy7iZsJfS9H3LZHoGWVqVC5ShMcmoYwVyox34d2dwyTryxSzZvlm5CTyy8CSMmUG
xsh47owge9gMmUYDlvC5aByUm0NnPpxzRcWQpS5vBobfDIoEkfx/Rl4cGzEv7jT0WrwZZ8bVCISg
4MwCEUH0KYA76np1Vh4T69nNtZwFa/sh5GrJaGKebMH5PEDS91tlNG3V7WOTggc3jhNrDmF87vdP
GoFN0X1EQwXigj9RIW+U0ELF1IdIiC8zosM2riyn22vJJ2uvNgpl3pflxWWOnEmWOcH9bcpEdnq3
bjM9qVih/+JwCdZq3yASJG4rCCg4N9TlNuDZofcSn3X/U9TlqGr4HNckWSMtBjFYyi4wkilc5Svy
toOoZONnWJVwECcz5y1LDkF+TQkGK5sYmdnRKFyZuIBB+jbRFQt7nyoOkeEkJfEtLrVmokAeY/++
irAnZGrcQRkHdQuidgIV+zpIeuBcr1KuJ4juwaoHQrn4PE0P+YfzCizOmsId6Ws4mGmjLVhyoYSj
/E+BKpy5Y/B5K6ASd5fwnyM5ZYl1cGUvpUVurOo9IxZC5GY6jqNolVfT2z+LnilkzhO5SJ+eyeTu
X2fJattbT3PV6bf6YQOg09ApLfmVN8kydWI04b5Bq8YBDwj/8IfH2njkrNPi0sgoHMoazad+ZLI7
x87vvdjBCV8+MfM9CYOvSawmQSeluxHuG5juFPjlMzpTKo3DWOE2S51ImnhYw8Ot27olWrof5WxL
aFPQZwmQdl1yXePWXCiNRLl/OaTzR/OWgTcujDLV/6CxWb87kpRojb6jC32ij1nfNQ84DBAPngmK
66IHMcrtmB08IkEOEVhIq1DokRM1lTeaCH/4Mzo069dDI5oDHGtjQZJF7eSfHOz/PHTa9BZ4apJ9
YSsZ9rTYlqjeGQVS8ZPTdXTMXmNaASCbqikvYPpBm8rCfol4Q6ofJRoXNdonq62zf78hGD3egpjl
balBGo5I6/zTpyt3BfF7hNlWGKuOyywQftMiqSpoWnL1ZJkFsNYoWqcenEqBMCvGblMfsgIsESEO
yz8rIuLM6XNND03SkFAkZxbSKRb1zJJxxn/R/c5PTx4fQeIjuNU6G+wcT3sS/ZTSdt9Ki7Bz53uR
ek0e/i0fa9NKmfGPaTByox/M/nrnZUNrK/LqgYQm/0qKtF8yT3FCtcNleWw3psGlXX19eeRCtTkz
aegiRrZORhyfx27a8IqgdAwNeQRnxj2suiQWIyp6nUlw273sCG0FGbE2aK50o4ovv/mhMpKkGB17
tllU6Cv0d573Qzgj213Iv60H1QIZSaDeN/00IeqhTwWdMgOQqXaKMpq3+9cBybIlsV5HMKKLu3BO
SARLXqZlFg07tCQ/pxLKXmLQgHbliUvVPnRoNspSIoA8Lazu1lwLQai6xDvawHBAjHfwBv0SY42c
MXYIcI7ug3l81U2KGP4SnPZfjiavLcp0Ce7Qpvu58JW2JF1FtEOMZ4eh7e00GLpADU/2HoUxU7ra
lyVVpPS6evjx369kV9jZ6Y3UVWMGwzOJoE/G5DFlrAFNgSwwsn2fCaN9wa0aB4JWRQdEs8oq/vVO
HtAiu4Pcdjr3JTuSREaJfmOiWYyy6aCHDRMGGEyJQzlzX9RyN1dYx39mlyEJaJseVlY4gwTCviUO
xJxfT4PP3bVBrY6jbnIBtg9w2wtjqbq8+AXsjBv6VgBruF6Nt7dMTqzQOxmnckJeEweJdaC2M6CC
k9rRRG5A8yl7uMG7lIKKRQa3HF6W0h129POdMHqPAotfLdIpwhQBrTj0aFxoDgcGFJGI0IISmHpL
ibhhVHTZHRo/8qQg9Mc7Wl3tXPZ8bn7YhB9FgF2SW1N4OIrsE1NstfFYLasitQkP2S1idaAAPsLK
Q6o5YtniDhFipR90JGfZl3wM9pNedaBsKTcLQSNJepvJJ4VODj4AYqxW8nJaSKWpjhjj/JwN2hD0
QKFDDjZSmgz3rveDJrazoGsBjb4cSMNVVwYFHaGoQmDUBrCgdFV5ssquEDwrDIveu2khRwQaAymK
BQFS5perKYuGZV4N6ZrMhrHwdurbmQBZRWXM2o/LOSacrjsbLAtOifrszHSzI54qGmWxsHO7pfMq
Yp7GjooqcikZyI9EmOnM1gwavlV5kuv/nCbUuzaTZa/IkNAAwRaNwKzXcYp9Gmun2qdlOcfluS7N
sV8/aUB+ndMiIgbirb5FbXG4icuT09IOOvVhZJlm4Qv8XUw38VYY9xFmuVrXtdwvqF6siIQNrMXR
MI75WILLD8s64+g0uBSuR5cf76f3i+mla9QJhUT8jCzBGzBOAy7Jel1XXqFC27TuRaOSRn5AKhUZ
YVpgzI5MCD9yKs85Wailgy0bAWNDz9AsnKk4D17LBsQ3Mcetsj3GnrYiUFA2+pq8jCrlVy988/rK
C1YkAxWw6Fq9c8a/0CBDZKtOZ3R7tEYgSVW+6so2jNJsrq9+XKQbbPq/RSc6hgKYgeQcZKa4OuhD
joJm5tvQM56jxJG6jJfVl1bbs5VT7l4zGMXxL/HFaFUNoZjwyESQuFBWjgTsNekz5+KxpEGJiY1C
lRM00ZRunI7GzWlje7vHW2JDnagyJNrr38IEOWf4i2LuiWqPH9LLrrH0kWBe0inkzhsehEdmnrcy
sSctmq3otztdR9eZ7XLK8NvGGJAzdcJMU+f70iAsENdSFVPAWmQxBk/mBg1fNjhpg1+Ly+fUorZ1
TtYwra2HarMq07XPP3XPXkKDzoSmtBxeuwzAniJe8jBMpFDO9L/UxOzU6ISgI0ftt9JlAWpnJaGN
ZibZ1mkBahowkbGehG3QdF8vJxcnaO4N4PoJDCws0usZUtegkDfjsdbcNvvE5BCZnAzDUKMFYsmL
mW74Z2BcLcCFsACbbV1BNA1H96R3QqrXRE24OiF1/cAHTJSI4vFxqtWxINow5z0wI1tBOg/Z8VE+
W0Selti2jnbB0+OU4mXm9weR56Qd70Wyxm+MYTcIBL1nr5kvDgpltCpCgoUtnoQ5ChhEFa5JIrJh
GK8FllcCPhXCMYx+s/Y/lAixpsartpCFP7hn4KgNGZ0Og4wZCb7woKwU2k3ptWoZHOeF2HTUo1lb
Mzimj3gVk+ksBAJ9QyJBdhMkJ+nOZmatEFJEd0AnUxOVNUgt8OUyfLMYnqoP4aq4e7MZSQl3+FGe
BV+CncR1LPAh05F0M4N77lNNxig0iG1m7GPZhXEu7DB+sU/Hg0kh5nI1oSac2uzyIkiSzgS3V9Gn
mJESLLSItCezAHlqtU3xx1h+lIhQz5pnyNaSsyFGXcG4ArepwOybl8yt0aDClCasTDMc82j2z7wm
rSahEuuejMOavqpfuze6y+Xjqgu92gOl2jCMPcINT9JDxHB6Cj+qe0YumcfaGlklr0rInIrrudyC
BDSsSquDrZTi6OKJ7jHF6epN3Skb6DT92Tnf2POcXZm5xWo9zqQ4HUNuDU2QZP7/RWoGVbNYgay7
NEfIko5QNs3UeUSkLcZMij4kkTVXY9VTmeTCVrkXoDbCgX7pQERvRZWtMh0pumGP090UoeEuasgs
UFOtbuB1QRatl0AKMzF5MmOlNVcxTeNOy0x7AOxk6E7JGr/q/cEnthd/e6ZILRCBUDijQ/ZCU4m/
BwWVYhX9I0q22RXJbwjW2Bkap6sO1XEwMi1tNBbPH4e0Nr//wpEtvFL/0HoSV3TyI2c9lpTTCcXg
8LRipRkLztCzGNco4NUWr52ZlJbotOg5WnRyP3/NR/RbNrw0yfwLuQHRfKVM2HmcRAhU7UYWmGWZ
wSoSsotYloKtaxYXu0vpqLDQb1AlKmyCygIJApdcv/IvmYs0uO10/WTBThD7ZJv9/pI0zMA6BO6M
eJunKBSfpsbSjAn2CDxZulcueVvoTEjtN36Hb8pQQpZ4+D2Z5Dmx7gjxuNetE9gb2hgDEdFvr42A
4dobmb5FwDgcIsibtMOEyskryS+ZCEg7lsD4GsjDDJMTnMLn7p6z35LHcXuSvn++clNCLXOZxdON
MhJHKoYB5X5HAQGGB+26CKQxkvZYIFG/2JzBAlouxD3d5uDIE5FzBEgBv8WPq4MYoLChhhx7ZofM
oUc/KWopPT/SEm0YljN6BLPoxdu+eqUQqdzldAVRw6aoKS9JUUxvhoxRV8VRxAIoqmxQ4ifsn+Ke
cyWXA200gxyxyEHuIzO/dUPJDYshCOS8GjzsAo3Bq5FnJUMZsEDuLUEcMXa9CwDGtBRMk4kx5QE1
dtGBYDfzDqWeXAt0mxFQ33Wx87Ixqijw5j1B//OFZTMZ/gBV+TB3WLULpa0UAHpXTnTJ1q7QPizJ
xpJm35k6mh11DSZZMwqrDrCjsrXCKzT84nGjj3F+pLv8NeHUfsIj+/dgUKdChKQ5O38PQkty1kma
9Myahyu8/y8+e2GWfcpkIwGQjPTJP/u6bJe3mtk7Bkoqlipm7N1q/q+EpaJDL0TexLhI0aXO1QLp
walkPWtlyNcoCLeFoOTU/NA8q0YvIjuv2jou97H9MuY+Nv+nEQ2pmheBJTEO3+jNHCz1eZvZzgJl
NrnuQ4PEBt3Qol2JOiJ3zz4GOa7rcUNApR+AwB96jDLQciLMe06T3zj2VGibnvew+B/uC1Pp2wGI
TE0obo38fKKQ0NLDBUAtXNCVvS/5WL9IPwGDvib4dFTHqLi64e1jTqPvimH7G84SDERVL3tSJPGM
Jrb2uKaQY1T5ryZaEIJfPg5yTOYc2D1kjM6nODXagrkP95ebKM37Yg4mX4QVPnb6+Y2yfoGHkL4V
16rq5d9gUaplYYa1jwKLtqIfstRmmXoweqBSn5hxYeAZAtlFuZg+x3VZyxsUFI7qh/ZC8lPMPJTP
/YpNeJRMm3K1sRVv4HNRObv7byOxgd5c3upGCkCQr2+8OTKM77lOU/qlSZv+11WHfJPKLAckZVdM
VH8apFHZJOPx4KfpwniNiJoXST01u2EgKCnImH0Hn67KcqriArxetjsaBsTxXQLWRchYyCh/Kg8F
jz0Q1JJGTCv4TJEZEEUajG55x2A3gF3T/Gydi1NHwVlMNnLF9mGMzTvevhLEYIN9UEe48wqBrIG8
yGIK3XXQAnFvAB88kc/YZIrkA7lWBZpEjXVhfVGAlaG9XX6KFO9TuAPfJlw4xRBmDPoT1Mq+52RH
3nP9echN6WOu4gnJTUAXbJbRFuDtoty9jrAxkU3UIBXKjhbcLMXM25p1SVM0Q6osvNvgN9Azih7X
6IQTwphxZiCklTAD5R/O3vV8bb4UX+Nc+fw0Mb6Xmzr9mfSEY4iki+1huEjn9z42D8obZuLBH42u
jIUyyprAmWJwI5/4FZyDJ/jX0WhRdI9soXkAdPZVHqxVxAZyI4Wj1sbiDuOenewAfbh1i6oUnsDH
+7jdBgtRe4FIXgetSL49B3bM0En16BvsmdZyNc3062Bqe2sCxNLerQv7c7HMjDi423CYlBKv6AEc
EBUxCmQe+BT/Xu/sVvm3LvtFGGBT2zXhfrpp08D7lYnK9JiAD4Yc30SCIlPutBjEvd9MSa6INyvX
vn0hDXftnO0apdHNo/HdLvxwpfvbTJQM+IVYmoUG/hFsDcvRsXGHBkY+3JTDSAIdWiM0TnjEeocF
m7D4sIRMdtlSNEWrM3kdP5zb1ctxfa061sEwmDARD/QnsnUkxLsqdcAVZjzsSc7lc4ImYVFYtniu
JLBDuBGhQ2k+OBNoRtg/pb+1heWLW+HkJzr9FGUKJivn6Yrv9flSay7rPDmAWUR8oULhedrjUQnd
6zJZeJ/m2P9xHtdRB+rgqmaDeT21+UCnkoE7B2ymApRz/z2dBiQxQHhOjqBeA2OMSo+YOjPD+JSt
MHMBkb83kzNDF1oCW4P0SBhWY0zxDsvuMtp2GWxkOn9G4dTmA+9YMOkFn6kyzeUC8Ea2Ea4wxLH4
DFF7crmLw/t/AKwCQ2NLbdVfhvmOzsDv8t07rCldMH59wqZiNZdyArfQ88VnodJW+EJ7p5UNpPZE
z6bkAyo9GvheuMiLNzkfnRzngP2PdcJMB9SqAejGF7YBqDjqQ5pti3Vr9UcmJqoe0ahUUr7NZlJA
BWRFFsETKZUP3FG9BiwgK6T7BsIzFWh6ORFYs+LY+HI5qQ3PAg2Lr4OBTSRZyj81+etwfP77oZEe
4zLru6zgR8KV/2CarQl0Km20UgkuCSM9BJwJrYXi20a5x+rejp4WdWPEkAgNh6l5wbqmtbSCzF8a
+SVv0O1iIYoUTcb1WM8k++9+YgFNcMKwLPZQELR2iuu7stR4vj5xgMPfZcA0tH59YYROgoZF32hR
DQ+oiPecQdgJVPk8bFPIboRvyAp+z5kSsPKxlp70A+13GdZ26wY8MTzUgcaij7YCyINnIlQBWUBO
C4wvo0KmCiv4BIeI6Aes4Xm0i960kI4mNDvjUZGpHtZxIcVMl5boS/a+PEL2xgtMwj9q8GrdAoAl
66ylc4rpHxzwDgivs6qL9fjROlLMHcZWCo5qvwt3Nboxh1JWxLqDUEyoQ/hwALXYOEmXeaGlhKkB
gGkizFsqEfm9GWRmstH661YrY4tQWHLtF/PdOH5wSuHXI9pNEdTULQFdIKWpVisKSgcKC7fY6C34
+tigs1kUEXcxDBv0ChfzG8O9yNPei030gf8NGkCNLcB3zPoOrubWmjB+DN22+ZM7u20JyMaI6i0f
VBeDMT3kIBRQP3rmougl7e08XC3wURptxD3D2egi87cHo5o/L9dq2rMeGyJLEDSBmGyVD/FTzqW7
n/FAx5L0FhW/Bh4jvfmdyf5antcQqfkTwWFr4Q+Ds0Xp+rnJIeDd3OBfoi3X0/JzQl0TLTPF8J7W
Km1nfqPyC/P7wds1q8bzngUiqT8sGTwrD4FIcDx97otKOpng4572BMSSQRODdaSMCjRXRFEWrXWj
zxV2j+62sUBjtapt63Z/uaiatUpmGQ5Sjs+q9k/9tKQ9gsXLqy6jok9XMnfD018LfWoZCEh4Q1wF
bsIBG3EGVwmeH9nEG55c8QUFCQ2z0kkujagxNwrSK+gHAxEFo4ODeH2RHztvf3Ha7GxL5pW1fLiP
dhSLfMOhnmmUnZZ9CkEdM7/N2UVIW+fSc50zihZg8CBNpQv0jyfZcl3yFUMfUmCn8JoUArzTy3Zd
KVf6NtEArLerhxZd1SI3+h/JtN9QckvPj8nTdvqKL41+SZpqymxgWJUZCXobz32Dh8MQcWobDwqX
AVwePArlvn15NQ02aN6iVAZylT+84FQwmH4shfn13X/55sIkBXcZSNTLApM7GFtLsj5Ll68vx005
J3cjFR0Mq7SW+c4fjHr5/tPuH7BxUIzlybjIhTDDCvVgMmq2PREWtHKSib8ydRRPI+OTiJeWSqGb
f2oCLKyvImsRTSdgAJBdcm9mzh8IyrD3BocQNfXtnIAlzhT0ht2SHr2JRsEuQXTdgjtMudIrp3DM
Ml8jsJRPctSENXwmYXiZi8jn96aKdib5D26VVTiyR71AbFdQmbEjSZNkq3CVuZFbsqfHenJmKDAQ
IrFMjcD0lcFGNRo7LW7gJmUS3zm7JN57UkVf2VsebQgaPmLO/3MTPIl+8cBbPkijJJ6IvBTzzeR/
xvZkSgvYn5wskxsNF9Nl/LAup3DAaV5Y+9xstFqKsfH0HfN838LfSzxZ5vPF5e/2i+wNS7sMb/jf
pKgUm7trpRzhBF6x0sel04yc1ABiRxHsUFj5823dcMDMq9poB//vs4OMifYn9tGjd8a+efOdXzbg
dmLjYwoJu4wA+1DKcJXq6N/jyUrrEd92RkbEC08FamR7PepABPuZzCeLccDS9IHt7j5z1umpYHKq
xbFigXjggUfOrhF80N1BvkGKHF7koMTsU9Q33sy2DHP0QH++yJ6qpEWa74rYFgVhEfnMQ6rmhEFR
wb4ybp5gCw2sLtogtT5ronAZOCK3bUNLWycrz31J7KNdsv1xGruWQ0O2sWx6OBHXfoypKw21qjem
9+t6NkV4juQD61MQ7nMoY09FRTihhS0WUuauid8X3mcjxDIv+fpovjgmUdvcmwV9/ldkdBfjU/wB
v0AXnVLnJdedR1S+GUX7mIusyDPg6dyZlD75hF4VpVZI9Ym9rhcyWuNYyBOesCiWtUtfysgXnk8T
AbQIQRpIFMdSATYo1jN3n5rJynqkkYUlohW0lkbIMUqbRwcjqY/ApnW52/u9H9e9XfB9TxU/yWq7
nkjyZQK4iOIlHhxck0LCiHdaWOCvHMZtm4c96GVwRuBbe5arSTGx8SSrdCsDhTvvQ2KJX6X9cbHX
5ULYQ/n02kSGHe55u3YpGBKaukk8unKSizE3sQ05OQKm4K9sUUvW7H96jD+0n85/yAjOm//yKdP4
0/1FQIsf5ahvy93qAeej1iq/ogaZWEYfpE5UgIGQpVSihbjM5RGn95yGZZV1fR2gFywQdFkBU4Ys
fR0zziHLtEWUgOep/uER2jJDAsUWKMTEe2BtmVLpkaKtl2BeEer1ns6jVFVHOVuFWavyTbKUqbSd
rnmNLXcZ/VZu4qLXfPDz8s2eZXQFzpQlwN/C4Dc/MdXGRkaODYZkEwS9+0xxmFDtwZKAyoVqiwyz
QtdXaK8rYPs+7C3dHr2JcQW+FsN+fUhwMJVi4dW0nrDTvGhg4fPbqeLyy145lkcU62ks7+7t+NWT
1Q+HqA5aSmjrcd8ljnHsg7pJWYseNsbtaX4SXh7XhvfX8J8ZdLjXb4y80ZOt1pS7QkqgiANxOOZs
Vcmi5JNcRPnSd/Ri9vhCexmWBeXzGxaoeLAnGCLoRJVVnbIWkuwkiLtNEGHBl9uLsHZkTjjKvhnQ
ChFfYmFbLAEt7eFJqSORhKMdzHkbhySGeJEyXAg80WEafrbNEje47FrU1jQ8rycm7dRHI44RODob
jBKUYhU3KCwxlkfzMvOcItgvne2Z9oPTZM+t1UPbONNVJapm4sn6Gnxnfvk3XepfkG7bMQYo6rtx
Z78Mw8ykSQQDXVNjOw6sqdNwDEWMW2Idlj9ytcqH0XU2avtaUzfaVfsurhUKyIJZVhaDJWTqossI
braRhUyytmqy7qoz274PGCo66/qBJ19Qs2zcSLIklhI4vUWJyozY/XDeUTIAZ0Bv/yNiqMRHNmMc
b0VMcH3wRCFv9Nmrq0vzhRSiN8ADaEC+y3u6wSUmepvgLWUswdP9cADwSRrshw43+22AFmPbYiqG
QknjWgLLRG7HdhKwTExAkd8KlokZoaiLkkNg80DswJ/JUjIB0/a6ASkZ5ylMoTpg4QtVoZtJAYvb
t0650SM2QJz117E6a0JqtQifN234qsn2dPHgZn4cqwriIYEJy7MGRaU2iL6cuj2cPCpwUuj/YE8h
aw1y3Zd6160C1IDVkn+JCkqEKrWOz7c/HlDoKTpJ57BHiMzOSEZiFR1OAEF5xiKCEIvq/t7/tknn
ekBgtcbooLLicPQH2DEbY9TiUENlD6iSxTz2Y5iSUHkVspCVHv2Pjg4taf/nlk01FwCA2VQFtkUm
c5+7RSEcelfr0VPZVTlmOaBScR1xIoMYCci3nSy77KTlg1VNvyM4qNrHjMW2Nl/B6FiQe/ukp2o4
ERoG0GSAvaxoyy2SIACrwWv7UTM4UIOUlwpOO+xWEWKKN0BhFzQvIpAY6bHT863Xin8gffDuUuuW
Y+xB69TyxYmxHjToTZXYmm01mD/5nahwdx+PdwI47X2N8d2AxNIVz7l5mPYsJwbN+Ty31ioy8P7l
XD5jbEKN0sHoOwzdZ7Wpi5gCfgZoQzEnexMTogxUksr7ol9Pymk6h4PoHrBE4wekwi+F7zsRcRZn
PdLXjhmYeBDyokqEWx11MamUr2OIa4dNFARrhj8STFA0MS76Ce7X+KNUZw0KjsQwrO0DyYG8bq5f
oZCC+SBJUOrucDOdo8Mwe5n9b/80hq3hZVkNiUpD5ieyR74RLcATtnVqW1hfpWGVP89pWryeI/3P
o5gZuNMLGhnCSO0+VBTn+bZZ6m105d+qlAcXVMN6A6pP5FsWGZsu+WcU/GDZVGeHBKrSQ1ZDBD6j
+REr+/iJRqzpksj/VjNqWau6nux/QkKcC0jSVAmgDahwIzRVyPD2Ol2E6tMxouPTpQJgd2nRyWzn
kzhP1/aPltm35ZuZR+Hmc3v4Nqb4vUnOt40LEzaou29hrAPxubVF+7wneBS/3DH22L5Bt4OiL9Kh
yEiFZT3xUghTvaL1NGZVStHgrWS1WLZcRPWX86813RFsJQT1PWlKObOmEDSKz4g2pkVFq8fniiTj
7nUzdN0eMm+npR83GiVnSI+NEeFRaX2yPYyek4hvOYmMGIs90LllH7340NB1Euir5Ksya1QB1hyw
0Q0Uyvtrr++I2ApCzsHd2TNB6WPqff4zMuXKhnRSKCFg8I9ruIK5dUstF3eHI4zdL8HzHnLc0uVu
5QMfuEXV/YeLRKjPKWfjIws1/rbPHiOR2lR7Iyy5pNgiTqBem1FtKZnBO8fOo159MKX5dABr6S+b
PqCwqEwk+55chGUmaRpMd/DMGe+1GXdLWxbeBj3fwspdqRVkWsGZemHEw+8SFJtV3sqOLH38OBq7
5XWbCuls0ZRe0xuo5WiP+1mcwZmhMmyz47Ad5eT7kzRBtsmSr+zOExnKBU8Hq2uA/I0k0DdW21ND
i/q26rHD8lilrc5a5+kztrGYFcXeyUYd9VZMhui6506dVsAqaGlFitGnRI916wHXb9NJhnmqfMSI
ktYdi5X8jSgSwc0IVtTdo0Jeq16OTYYG390vcVwf6gAIVJOJqwpzMlbZ6T0E/jYz3ea1tN1SXLs5
31GSmYBZukbjkMKxkt2rl1fYnk4TRszPKG0fwKbHZd2hnI/ew39tCiNFDknOKHIh8T+fMpbY2wbW
YFGJve9yPT3NFpcKZurIyAQf6rlUxC0Q6/4uWYWQCFi/8c/t/zktCWrxrhKmr3AaP7R1TCTWohVZ
o/MnRazgn7pcGidsL9kbtDCjKDD6L0s3/ag50dpXnZOvu2OzLRaNGcV3ZqoEtToCqcpnbsE05Tbq
sftFVwMlJX/Lh3ihXnMntE40vaEgCVSoAsXn8p+q9vjbxhRrW7QAZAPBtFXYEDpuPdtevGGzjMwe
Jhj+bX8QaTGaGEJbXjV5MRMEwKKNUJS7SoU09Bq5JB97COow/pnXaSbZvxdRAlCrWplEsAJe9zRt
ZVtpz4qd3vU58fMbHF5V7Cn6L4DZ9TQXTUmVohUeneqCLgpOyxbt5AXGNm1bgOoNTlG+nw+Ymqv7
qe1tZxpECQLxv8WcNLT0ur+XsccjKtLfYV/+f5gW4maLYt+025K7nU5CXalM+xCvKKItt4pT5+F0
peA4XPkri2dWnZaQ5e3NyXQDz8HNd7IZMAeiE4kZ/DUl8MEVuY2fXtMjEWWJoQJSzaEbxgJcC3iO
m0dyhgcj42svt6LeBwd759fFaJxWJMSltShNXvefSzxLrg1M1FlA0KWXGPxBoWZ3ja4YyIxYLj4H
90++WAlxHIMdDsCZ3bfkOz+RpXWgw2WKjaIaiD2HCDk4PhKC/O7Ei7xjPnit7GrxYVXV6x8/uiqm
wCpEM4l8ftXjAP5FsJNMiJ5tm9SAa9GviSNC6fK3zz/PS7j9uvybXhSGk0fpT4JqF+fo0Y9Xr9R2
nXxMLiRYsTsoseVDWzvdtmyZZeAD4mod7iZ5bZvEWZOwcq2SQ0G3l+Cl6HOb5kgaorDSfUAvp63q
QfiQNbsb1Nyebw9Qx+wWZvvHnrOvhIx8m7c4ONDj96llS0iq93EM7Ccg61lsOfCoFMvulgrw0HEc
EdeqPlzTaMHXyO+nay9qjTUTacwvfWOMGl+EeLy0lMcaOeeUSPYP3u3EyE7fB2uLeeZFMkBPN/07
RYOvKW3Ik+mafXKriG5IInO5inhB2swv9HySfpG2E++rr0yz88MODD8+6yb7L/zylHi4p7c+XBEH
6zj9bWIzOWVxCsgC+cPxsQbjKF+rXw5UBLAmGZ2Ta89k6HfojmVNtZ8rl1sqmUO/QGKAjnvBe4LK
LYACaaSSs/4QSufQs44NISQ3++2pqQPNDy5FEWBsUxP613OkPuIEQX3yjpn+Mo+65oluv5013+1r
1PSIC7aui8FyqbKOOT/vOA0wtRIrLyPT1NUBM+X9lPYRypM5JEykfzBuPwv7siMrWtcXiqPwWl/x
zBgX16BmwJoqlcVexgKpA9VeKYZbVPKdYHzBsLeun0pPWByRn5FGTYzk4ufNIF6tk+vbxaYPh0Si
68pZw5uE73Qpt4iK2mB71Nvr43zPXZZMWzhIKVURgEWYOXTAbAFQ4ofYn/C6PRZ0KIjX6gQWHBOS
mwDAY6lVrZpupAEV/LUYL4xqm79Rnt/qnWbeV2APX1ilsXXWR4LYymndZ8/PQYq4hOHjZz2WobuC
oQXmsoJYbL6oboapS/1khe7Qa9yQZ62FPJTC5m5M0/MyKaL5xkCJCmiTKvcKHNBDMV0OjVc+wH+3
fCZ8OslqpKEyYRNBYKRXyMpg7dz0Gnmw7/O9WS9Ychu6ONuVxA63+BCBcKd34V3EgQ8Ej7vOif66
sS5GZUBLkAoM2c+Tqxo97MqHWgUwnrysPUPNCyCOKLCPj9ttwybCTzeYehJZtGcwOuaz43FkfQje
SDGOjW7EVwVckA7nKtshyE3GZtwwpawP9e2W2cWv9P0pDkkCu+7QKEif57Q7CbpPkF3UTyOypX+X
Vj4Fa4ODvpQUbc5/tk+oJ5Umap7lPJ7MK98m7ggfMqtTUkhf7VIBLbv6yDeIx3gv7tIK3JF94SVs
qd1Jf8olcDzAfvXobhWco3/6GRJmOqUQ7RWBQRmhY/Z9URt7GR6HuZBebDvlPjuqm1iD8RxDLtfT
/2PAtQuOYPHlQP/eP9kK1YNAm7sV4E3Whb8gDFP/Ue39uwlrRKUyOQqyDcTuf26CJgD0JQRG2XD1
MWIN2dZ/5l9GMNYi4sw+L944pFAm4ig++HaZL8BjM9n0UcrCrKf4Mz3+JX8KzD1+fkWXT9n+BGPj
NfazW8dFB6j9N0Mg/V2J8G7UN65wkUv7vGr1PxXcB7B5gsp4fYusMQYkVsB5PLsU/tsnhs/9EE+t
jPpPw2hWGPgnRAl2xLq9DvkOPtaaEobROvMMrkNXxKBr1Mu+Lpqpl8wfMb3EpWT1LioAanTQ0WEj
nJs3jAhN247KVstKUUvpAS4jJhA9xuSh7KM3PWydLOIZY9KDwb8yBn6XffW+FGl/YgIAUIHMfNw6
ip2JELNaE4fLhHyptr07XF00zhF5jOss1QJ3cRFRjgUu0mB+TBnPlHNdOlPA4rDUGJzhb5JBbipw
Gh16dg+NcJJvWTh8I0YK6y4kK/b/h1z5Neg3AVK57qg9YXxrg99sj2u6rmXPUVRnQFQ/TiiP1fQi
r1T0D975GZRk8bLLhAsOJIAwlDUrwmwTO9QasgEpCSz+0gWlozHGsVLi17W4qfxhCE7WjEXEOpxs
3addGS0rsLDQcpH6Jf9nYxAOLfxW6inTPmeCLeVgnDwivKByNh06psFyw9X6ptw6GUTquOZSWlUh
OYB33m1hpj5bDPJqRWkbK2b3hkKW5egtgVwKaxt9pBQxACwOnqy6WOsOC0Ze+7tsYwo3Q/NH6Wkb
nxExYYpHcSdym5S+SkjzjKKIntiZJNUl9N699m+Pxgh17BF3ec4yALtsexPOvJ/7Vf6k+CXFsxog
lsiWP6QoiPjxxeo46UjVqBRC0jrj3rQpcCB6NCVyOfYggbhlXiAgpkgBk8diu83+J/PZQBCuz0OP
e20CelMvTWwbB5PAX5HYxOnaM196UeujSPM7W9bYMPCmFSxe0yBb3xwmBJCdmDaLfZdsaJP2QoGB
Tp07M9oHXN8pO1ktt4HimhalEh9ymHUWX8a9NITZp1gUcZr7oixT+LPLtgtrfWFrE93bslWhI3px
SjNqJ0ATnl7b2KFDkZ4/dRi4z68Kx34/OjtMGDUMDKFDvEXo3uPa/CXJXwBm8c7wtT87EzJkBF81
idT36OJJ5ckebnCDhm7rJwRXDuBrtWOJt7bc673bE9d6km5u7JMsALezfX7UULi6dNVcLDPmwcYB
8ZBvJ4NMXuqM1b8cspN2OP4HW8MoSvEnv08O96p2cyjSZ7fH1a3B4uHwK1jinTFRetD4i5t23lz4
YgdppaAkfaIoCdON07FmcM9j716xkCW/JaHgsSRUS857pPa4ICHEcosLavIsdYRkEn7yvL1nhH2A
OsQB098jdUmTx8ws86n8swD5AJQaaV/YhWays1A9oy+My0r5jsfw/eByHJlx8Q4PHHUpY0xeMCxG
FWwQNMhl9fxh8H5nFdqtXxse+hxIMco2aIvdh7nlncEF4VCul5uxficUOZyPWZENWvRhfKvK8ywW
PjFxLxDtCU69dmP/a1SnyKvCM7Wg24V4mXrJGYd9ly1bfuliKraAhSTUhevpIgQ/3fDPhfWwRQSR
NyF/cYhvTf6IpetcELh31utNEU3JD6dALYoLbm/YL5xY2rdh5CR0Hy8OSzL+0ESoVKjWx8S2vquX
ic3NLYE7Nhv2dShy+WiSQsrg66aYJvi+L3Yt9DRHKR6pONo5EypvS2UASh2ih8B6gYnaQ35ba6pP
uEnEcRUxII1Wnw+33HWJLZFOmxFOVqtdNOPf7TtYei1T0p26CFj4UwuTm6+PZxLEY8u2c9J+mnot
H0p/r32sq3EtpJAJFyj7CyMQLLXzovjoqGauitb6l6qY4hrMWV3hbrhCn4PsYaC8pUmPbq95Tzp2
99EdkKXvFAXrYn2G/RP7mx1AvAoRx+knd/2lw+TQXTeVUjkgoLFF1YRn8WxoL2S9d6siwY461TB0
+XvzIBWdaJove26DPhE2tLRLpJTKdbOFvYLoNuL05Ld7I6oCTTs8+safMStwGVZTiwgt+6PYRnvT
LollBDRzcvSOJ8ic3eJNsIUIeUfq+4Jw8SSFqShJNsrhVOlk1ffFwWxxFMLbNO50tzpMugZqQTHQ
gIBVI77meuicgGmRuvOqhtctOXPX0cIE9SOT3t81m/urlz4rHf6rQvcEiRteGY7W3o59en4DjFPx
LbYBxBqXWH4FIO1Z5yFOnMCYrPPjNo5BT1cms9Dsu7Msh+Lx9hRdrYIhKfNIDve8JgIsFIVet1dJ
wZD7tOUUZ8ua5c5gb58+lNpNp0DLUbfhEEFyecU2VSbmuEiefVgIYXinNu/cNBIwArrTjSh2WmFJ
L/O7w6608pT7696uIed/vjf5aiWznSx+LZqE4QIXKT00Og3sENUr+DC+fGuJC4pqu4WmedWszRI5
53JiMbLtaCLXcjxEXGjBj+YRiUxwekAJPq9wvPSF0TF2/eGEs6ZWWu8py0dLXM0wva9OMtc2G3UW
349GpOFf4YaQWtvp2aJyovBC3P2BSDGlufpIDOYQoLP4/W1qs3svhGLItvT/KDHKNSgs9/iaYr8J
m/CO6DY+Y+jJ/7uMZGpkMRfzPhcojhQ36qg3w/UPnD4bXj8hs4k1BO/tJ69HbQ/ns7HpsB5aemEy
OyOlM9Rllav66nnchWjc3aaG2TztUxplHSAbDivRGIaRXOpC5ICRalr1DUg9w30CP+aSs8dSbaJx
vK9LCKLr04ns2KyVELjPPi0g6heKa2lfCLzkdxhBLiHz/cDDaKxa2sg46a8JMOtcimsOMjh/PF5V
53gJYk4TXaFuwVjVzPkhkmBz/pZlNo/2rkmFrfKwl6FX1Ph63R0xsDA63qGcUtGekTLlraEt56+G
ybrQKnCqSFY7XFfFB1vWmPjRRelZToE5fIYsUnVmLuMR7aqydwM8W7ZJsXmhva4bvf3AB/Z/TIHA
6DFK3TZhNtv3MgTSGydnFsr8oS5G/qfjGKFUT6J8JGCL93Ckv2BCGqbVXKsJLFzGWD7fghdXNSdY
S+Ray4uIXFter4M1hlBeL+rw8z5ShVri0fA7uJ9q8SOpdvlQVWVNEAvhyz/S1J27iRaBra/JYER+
Jy27edADy4l6QV/f3dRJIA+F4cxtX4AyCRH4E/MkMXEFfg1ZUS9QDAZlI3BNpLPH2W5JRnddPSMn
9f4o4ycYZAy9vYGpS2SHg6pTlV++7QvkPqvN+015is3jQ+Nr682NI3cii7tXw9G2TgoHJtWaMKiq
87/1hBcX141ciRnKbVXTUkqwtlvq6aoSupvUdG3I95TA9pjVuvvRsTV5q4FKiL+IaAmZiIlFdwnJ
95S8+u/qF2Hxr2mCiVf8EIEqXULByXFLE9h2cBmwcU3yCoXjXiwpWIXdAl8O5DNNB96K1Or33g8u
5LScGGMs6zqYgzTFL72R9UR2b4dSeCLw/XXGj4ta+fU5pgj7sbaZ/PbDC+IwHES44JioSVi6+gGC
Tkacw8qlF+5Fc3vStrDL3X+78rfR9GhNKpIsPGwcVQ8kwPpgqMBnb1J4BuiyEaoh0z7VFHvoqAkv
FQbcBokHoAuDVvtU8IJLbDP9E0+t5UJe5f9Us1LQjoidefjfK6S+TI0AVB8gRsmo6GES0CGbFSn9
G+OI9+Weuo1bi6ym7QGWrKL3Yf/W6UJsnY+Kx6kosbmbTNRlL5Qt0y/dd6Pyjgbd1AaIzbBHdZLF
j1+x1KzSOX/xeI42psoi3C/+SHHgQGf9gVLh7PwHwwbQD3HQ+AZM3MnmWKplZlq/Svk+c0Wvd7ge
rltDLDZcg3MzfsSKCQfyADUMszf0YXa5rBi4Wr1xd3iPyK/vL6Wao+xvVxdRf2DTF6JfH6PZV5Cy
op+3ad+drzAos+B5txzkvOOvR9iStoGT8T8dxvU9YIzwg97ORjSldai4FGHvU6aKk2fn8XrL+ycM
ELwqjq99y4Sg5+xZYM/OaACmFLTK8eyq1jAjMnNVP8PgqPk18JWRXLUEHV8sJI5f0cCht13Bu61L
HDkYuYNTX7Kg0+dtxvKKEEcJr/Po3IDmxhV0fntVa2Gx3U10VZhcpM18GZtrp7JuNoJbt3kvX9tx
E5KwFX/mDDMMseOMAczveAY46ZNpG+/W8k1SmCw+WF/CObRl6wV3cB/FtXG9DS0bfC7jHZ0nKgy7
SOV6v8ltsMZS9Oo0yd0iOtS0jz35k9cHRturWtunQkEJBI4NqP/NQJ2o2XDGIrg54WsDfEYyy1to
fC69PtVlGyzdvZo+RYbq05/42TUCyFnY7Inhl6s2kmKik/n0QGNSTvlCze5+PDIYLASPdyKQ8SBF
6SiG1tOJCng0TmVXZtBgapj3yfEke/B6HgoGf/k6KWd7TfZplDXNOV7d+zcPKGJPF/IF07lAtYRX
JOp9rYOMrt1nlsdr6VEbrGN2cfQndCdb1cZQzJc9fRpKsNvoIWGg9PeTvsaA1XYnUZ+Jioq1wvPm
/6dOAMG0c6odADJPE8IFBOFTtL0OABcfC5kZ9qz17EpWh6k3KpE+5D0EQwEMdnsGmlAralJhJAK6
J6z8ozUWNcmf0QShRQ8Iw95+xAxUn0fn4H2C3DAXqU3Z820XACSTsImEOC5oRHLe28pJ/DR0UCFB
JZ0gl1Q3U087aHE5BzFNMn+yaI0XIoP+PIcABlILpZOqoMFUgLdyKtvr/vULdOwBYVSWzFX+Dfam
px9fF4G1F9qQSDtCN3v2yOTUCsvqgTTo5K2jkB5gxF/SlL/E6NNg2Ln3iOA3KhwCqMMV/6eGhmW4
G8k5wO72Vl/6QkkUA/SWNsj+o8D1Xubh1PAWlbX+ro30NihR5PC33J9hgzJfy74IFHOByea9tlS5
I0DTEwyE7Onof4/oTS7H0zDdbT1Q8DUlZ1+pDaWRYA+YQ+gzgabfFOA4O1A8hDl710IGGMWjnsoD
FX1OniGPQ7F0jJb4g0oUwONsh4ToRg9NbrtVOnnaIHYIaDGJcoKraAd5UBp80enoqK30fUo8Lb53
8r3Kj0d11ePl1JTMv6SPA76CBHyTh2FpUSHZh2dBaj/tOqcYFPpL97ZJUMNlSCmSWE/gEQ294gBZ
2BXUaet2N/25c0K8N9Ksyi5A5ydngUn9c978jr/7Si3z82KRy/LGsbj+9huO5V6ZD0XlEkZemJYI
MiOy9rx6d0ySMZyWlhgbyv1lw4sfJ1I8tPXUv1PSfjyQDlUEEXUImBIkXfmoZRAv/88Ui3VXF6NR
3e00dypFr5b44nEDEjflprahdGCcU1p8H/VKlt3DZw15j+Jq3MmqNy9VuNg7GukgEfeVHauak5OA
Y3zUGTnUCxgAwAv+Ie4WtYU82fIWEXAZfRsnYaR6lTFNlShWc2NnhuckgqRCmhOOHAvzmcv+1VxS
bb8ItE32v4bpAj4y1fMRfbccrxyCIDp1/VkOa/V8n2ivQkxd0+m5HciQE7BLoE4o8DWj3dpIYpru
CbxK/5tsXKDNen+e4xjPmijhTwK7zpVpEOh3LnwD9QOGvLE2XJxlDMVrTn0WKJ3xHrP/txIZn0Z8
73v4bVhx0jSF3sW+1/CoSwRb6ZZCEa+i6WJ5TCxmFM0BH4LhGFNHbZkLZ7gc6FmrySiy51N+za6F
azwSB5peZAq98QeTwOkpQdKh3aUK/W42GdW96VFRdV7NPtSaP0I5Wv0a8hbYA61sOQvs+ue82QPJ
IDuHJxSDiVz+qPS5paUIdQUJjZ9PP0H7exLsQ0KzzHZn0lgMZZ4PmPmGAzffAr7FrjEVM88VG1pr
sawoSONGnS7R+6DPbLKh8Nqvwok63DWpzOnMGhc8DkGTahmvVAfjg5LCgpxarj51OMjbm/KXEWVC
LranpYUIuF+VSfMMPDsLLGSHVPI5bPVKmARnss/dja5GkD14ikxgJpZrs445QLU+tnupi8PlmsOO
xQxTSdtpRJhyoFVYUeOSQ4t4WXXGAOR4Phcp/ZXQFjcc5WpQzw5GBJz+qVdbWk8boicXq0CR8e5c
pWcQgnwTlMn9HYNswamLN+qOhME0SNoagYAU0BG0Q7X70qFEfjlLxV45ADMmyD+WqqTUD5zrXpKK
wsPFWsPv1xH1RSQQ0WVNOzhY856CxpgtsUDJTRqdCnQnG8D8gmkA0TmsMnKN0/KtMttoWsEbh//v
ltND2zdJ5eVdbs6nhwrirHXWQVdlYXMtfagEf4Z6v+lzagHWMHPCtxYqo/LlYhHOAqyxsOJpj487
/CqH+B2H1hxaYGt34a9P2eCThJpZ7YMkf0wJTduai19OYYxS+73F/bpRVBjg0QMZs0TQyv4kPUQC
QvXuSH1Y8yDzA1wGobcHC/t8Emiu59TCbT7SyDHmLGrJ5WLBoyYv+VIZRHbVoUpM79p0iLoxMBVV
KtKEiVfQsAuNYXS95gzIcvs+wCTLY+dJkFCg5ZNBxOTe18+4WmDAqZy+C+032CqX/idCwo0Ick0b
1MV5UcG5KaF3pa8g/kzT7Bh9wyNACyg0TmerB4CucAJPBO+YpZcvrKyE3GChgVe2/Uh2Rjr+00dC
/Yxi59var87YCtdMM7/1PtOCo4BtIyH1qO6g2S26FBXPQqorPBOOc69aoQSLTPGFPXExq4jD5edV
gVDX70QLuwCL0Ffv16VCgP0ER3WoR8sxYoIG9B1WSJc3DWMvTbFK2pXg+Vhy4wAqBtCY2YF9wK8w
2F/PLbT+M8WIcMJwUkqVyisBv+bOKKJQHM0Q5cwyhjaamoGOsaJuppIKzNbaQP0iMEurcQo3WCa/
+Vodr4nkLF4VY6gqMzgJmiWrX1e1tglNaWQtZ1kz+jo8dv05qHu4s2QvGry2OSFTkbDOgyngXSEx
TyLSw5KTho6h9/Po2FjPHIqUROT0Ocro18mL7wYzD/vJG96Sl0ot03lrcKV4+ywlMZh9a3GOXi0j
fOa+faWbZ6o5HhbYaMPvCkEiBMdS18eFuktxt2cXNrbDw0ciLrOml/4kiZxpg9u5+y2bEeFnR9Pf
TMT61GCXIMU3t3jAIGkkUVTVJ5xS5XuKETbQ9krD6tx1KRZdJ/rXNurElzMsQaDqVxkgHOR5z64m
nv/FP6Iyvu61OuTkxJtkWNiamhOB6UQAsciEMyJa8zBG+8EBapbbkNstk8+fNV+i6tYYvI33yEvZ
0vI0Xi3x9IQl2drP/x5ZMyV5kkXhK/E/wSONyYKtuEgAQBbgTG/WZNTMwI2hAjtLy/EGIB/qTnY7
geuW07u87+2NzKOhywgVjD/aobaxclnqJmqKqLwNYdgajKmWS215ScPEKNziMYV1iGePKENkeTgR
83YSyrfJ1X8alfJTbYONjSiTqZXE58osPPb+D0rZ7viz7IODFH2aJQcUVX9tOa8bksMBhCV2oSeH
siQODaytKPZi4JxO52NDF1YxOc4tlfWWibpG8cOcAJr3iJgYHdjkIimJzjM8ysndrwbwW9mYeIl7
5rV29H5sKKwDl/NpKM/ovAYE9olD8hlnQ8qLvCearOB6dtPsb5EhVi2w5/f08K9ovfE4qwLYUj8P
98MZZLCnOzNMaZrYeiwU/9Z004lhv/uXZGhGbzvvqXTOTa6anoThOD9qh8SuSNJuDUt7PgTnx42S
DeIBdJ4BKV6eKO4cWITun0ODRmW1UNwdXnAJ8VDZEt1yh/9pHGToe4P5eRo/0OVG0tXPZUHJi199
sccgN9H5Psgs63LE8dNZ80P1BFFXtVPOtIQ49jWGRdZ/RwbKsjib10pWgwFA/81+mGYju8H9QqNg
VeephkpDsscx12UuP1YdbLaVwhQkEXWlWxHNiHt5jc8cjI0234HEcg5BwQYkbPAW7VaRyBeuQxax
LKw9FSyouiodwoF4zAAsVxH/QHUd7/BESYPXhJykZvcLYkgGlNhzfrMVMgykFdbKvDnFj/Jc0yNG
Elg9OvPxFrXHmXC3KSh8/Njj+8Bys8J9UhO4kt7S07p7YtCnFKjAMx9kq3NSzejApVTWA5Qua1Y2
YwrE99w7Zfr3I6OCplefxb+V+muid9secvIjaqnwQCwreVgcYHwsfXRrlBOSQT672xyKR+EhLhNW
tmKg+YNWXPTaKWXUJ7DylIlqqLZOROmm4tjeiJrtKLlb7M5TqZ6nEG31ADdUp/zqJImKYRCVfsJP
pZHf8CDmamhEbSpiOyEm38Q4E6Ujd4jsRO3lN0IeoCbAnNXs1aoLkC341wL2imt3NnjF2e/c/UuA
m3MZKRi6+MqaBkK2kJWcxucwjGb7mqZcyXqP/RwJ6HH6QyafX2w5SCwf+zJUOZTd+tlgs0pfbsnT
Do/M54nkBtoy+Zt14q945zRrrjqxOyawNpxC3VPd7+eRcJtszx3DmBCLoHrZYx02976p+MqJqAtJ
1F1qe5vCZ7mYB88Id8JyNDpZOx45hkphbilORKjtjgsJHWYk13xpAr2cIPoeRqyJAyYTlo3hc/Ln
y5O/18ThC8vhdbZAbeXeP8sOWMPrjFObfp+ZjhzeLH3lEnopm6se/DfXLd+mRd2Nnoax0HV9uMoU
yCCYzxgmiVybgqjTLDoPNA8MpG+SVk0oL6KVIUBpc8O1uUqo913bDTopkeGn60S4A0IGuYdMVsFN
HglmcoHaSzj7anvlJ8/PuKIWTc8OHfUOgPhWwdcklGZyYLPQOC2S9YIJ8lYrDAraUI3Kkb5ColDc
pgvT/on9HgQLviRbF68+D1cN7WuGy+sBoC+2xT288tGNNJWQ8X2qXT4a6/mIclVGSf1lMZbIWBxB
iRIhtAXs3z+JugcWStRvGbbvAqQdN8qrHhLb7i2O4v/8g5Z24b4sNMsPRiHbDxNFqJW2Vj0ZrWWU
15luQ/wIMfpBs/vWru7C/LyXIeOIYrwrwPg0uBrDytbJhNB6G1W6sIredaKtWxDpjbSMGjKE1tnc
gSokP4Wi1ZYAyITOku1psTdHskAlNVmVEGrSUVibslo4BZhxt9E67VFULZrdWNUw9Efza/Lmu+r8
LKvscIJloAW6j8KJ66z8JzjdgJT6Cdk1pw8PDVsR0L00whUUiK6/h7IkcXJbX3vscYXE9ZbYRqvi
MZzNnzzX39a+8upf8WOLxep+Kof/9E7KRptUKrt3tS+qBrnfvgSm1B7Z2cpKFewCpDCRmlOaSLUt
9KSPIlF6CAcmD27jhMMBForLZ4Z2RbkPXAcqUX2/qy4FAsRs8k0ZMDwZP5ateUihWrTxO3CbNlXI
Yhp8GZSOpV9g3uPLKJI9FcpJKafATR6jlfZEQ+A6HPta20isyDqKqyZpIyDF7zk+jXszueG6qej9
5aPMR6GTas+bZYGlkoDn4tq1/pAvzqDf0GUnTCgXvXPLAylcp4jioRUEKp5w0t3ZK0iD5JJ9iZcW
q7irxViqpHmJ5+JTeGc1yp+JfP5YH4C3uGOQ447+Kwi1DtKw0fqpCnuLR1rGfxFcq45cNpmYSBhv
e48GXB+2Dfzd41lkVhnUQJ+BP36CGNhfYokfwKGNpplIWsZbKshlWGXjoTO1723TKar9n5fv3wBU
GcZiq9JUVRRHcTccjy/3vjI+5QFgjp0DZqNKW215arlYuNzyIG1HuX1bE0QhL/nacPsUnY47/mEJ
9As+o2XOIclh2BpycblJZ+iDR+c+dJfZtSiWX7EGKjPmuun1T9r+Reea9BGDH+dTI0tiPgyZGSJ3
g1jJlovJZuWPoJ8JeN/R41kaJkABMcuGSs5AussTXggYKElzNaMsqFmjV2xbdeylZXR7FwxMYeL+
WEHm/8ww5VqOQUTEgoddx6Su8Q37dQPUiO+C+nmZlJqANm4CcD0ZyT+tEOFp0jdn9ZPVgL7kR/g/
MHtRUIz8c85aFnDT/l/HsRhIjEpe9bxnU5aih6W2ItzEgwbXXmovTjmAutMXh1VXYhV69O2imbrN
u/ryviZvoGVwDDKmtLtBPOtQPP1K7w1/YQ1rhLLKpu8+MmOXv2lyl4D4v2M5Oo/ymFFTlHLkrMxK
KBPKPy8rUbGN4oF+IIgZYgDiv5NlAf6u8kYG4kADXdMJ5UmMi1cpCMtFoNSJJwLQQ2kuy5Xcx2bQ
mBnv8PGUFt47733/NCtmW7uzWgUQl4vP0CJ+vFh8m205HlcnTZc6/v77fUKm+tFZA2L6gxKU3jNg
cbFiPEL1J7NfnrzU5qZMk0Id9s1JX+5NJ/laacONDjP2VN/OJH54aY6JGTfXswGOwIJSZ+/2xgiC
2lB/rva+5DHh4ICEdP8IB9OYkwUWeYyG0WZuMkiPnxkIOvD4S4B2BvLfus4NKrtaLKOW6onbIlnO
BJb1YoUL82Xo7HyebT8CHryHyGsAx/ZCaKIm1SRPRThjKHmMDQO+va61jVgRs/Jj35N7EXFfxDFy
1st+bAozwCknR/UhU5Fyej1tLLVwkS8istxbPQhX+44E81Dp2ntKmzJONZrJa2TJc2M0P8wguJOG
efsyleq4BMZ23IMEDskeGI9FXxcqAefevM/60ZKR7DL1lW7wFczJ+Fuv6DMiwpvRt6MsM3P+sDcq
H5oBlQkoeA7Rn1mvV98WW6R8xTPP2vajTwMoVLtPp3M27iLFuG+Di8H+lkC1wH2F2zzXqkOO6VVZ
cuECn1ivKiWc8y6penPs1pz9xaNMQHKSg9LBySAjVe4YJZACC7JRK8UfO0e1wPUGO5jCYYeFU/hL
VheciXHlicoMUXfZbP4+yYke8MPzGLZgYovOXmCJ8EtrYAwgrzGAac3ki+4q7bGWTp+1e+eIFxIl
N36nK2/rssgww9JNp+w3yu0rwnejXYNyupjgN1uG+9pAzsHJcy3L3hWUgD36xXEh7zSOqpcTVzkK
vLfKty2C1DOOgptdRxZzzf0OCowFnai0T+r4/FPPDVFTYwaGR0JKi2ucybMduHAWAS3gJhxX5/Vc
iH2b3a0AUHJXuibA5sHE/YA/zjfBCeGiIS1l5TiSHxmu9Oc1dNvW2PiZ1zaTzWWlAwjLebwLyEdK
tKIs9hXrokEtjOqGCtmmESfmLKmcXxacZ17oauLud0gEWTpwT5TcWfboeq8Yi/LAeG04+QAb+eaB
AsV0xskPieZhZzY3SJ7u0gy7s6HmUx4ZeTTKdfWTg7i/4FZ3W5yTb8W2pqYoVqtH5DHrXh2NN4p0
zkF2iIBkr96dkpYvv/e5D3S5Emv8wCFBH8aJYGzWdqqwoNJd+ZRa5Df2+Zj2HVBMGelC8KKM34gB
32nGKlbuw86t7BET5e2JDtrgBymfNkSJnH3uMH4T1LRYj2ZD1oNcsqCu4VNIc+EoWlHkuXrVNBgw
BA3m503P7Kk9CMnmYsRM4VggTyMsnJ/DXERfwJLWnlNrx0Xjc2xyMVJk/DVm4AElqO0c81UsfGGw
ATWMkHiiGkhzz1ZC0tLbWF+WskXyxVG4dNituuZS+2zyqdY+xNdtUja0gOAsEFg1fBNeVXxSaNxI
Th2DI7gr202AMftUauCa6jmGvxN/J7SNQwgGd5toPMAoc+grsBvwidU9DWxNd7rIn6JqFtz34OAi
5mVJYqQJj7TnYwmUHTOIA+kuWaNxJJIb6dx0Ut4X0hqqwuLQS+cksxkNuzfp+9kGBEPXPG50Qxkl
0DCPz5yIbTByEGx1tSl+zFCji0yRyH0ahphC7spW7DbUVPQl8KvNaIa+XpdUqvUF5S5LiorBdJ88
Yj65Xe/2qecXTgT2E21ofccxHJwooYJJpM836uFYVOheyj273lhocLbK3bFXZT0zY7sCFvrsIfEl
kZbXUZRtq3+lH8tPghpw/DKucMU3WIyqj552RwauZ4tzbelixAwJEzSUza6VGZ8B6hecSLbxAY0r
I7I7SXcY25fv23UEip63sgMA+S8zTSxkk6AmUzD0HBGXc9FK2THUlRdu/GZuV/cMKEboaSO1nKJd
+WtfjVspZdnFejEjAX+dJYXir1b3bB/B0GWKTxfNGej+6uby5v6NUFus/9/NwwR671CaKfblA5qy
MxKDHMklFCzjkS4MkTs+kU92tNhpXSGI7vjJHAsyPPzU+fPgSgJUGMqkurvCblVozMiFuFcRQLXC
0HIEwH2+gKtqdbnOdNGnqbrqig6IpjvHTHdBF0urvHnxpxrBZ/uOycHiswv7007yTUg+8+IVRW0q
JuzUZLGPr2c6rTXWd+ENGIiexjPnwNeld9bpuKVELB1hTkQtJ5ULJWYStEkDgIH/8GensItum1ZH
7GsY41q9VyC4pLKtrdPTvQWU0AwhY2NxxbhEvdGwK2KkltjvfnTjjVHve1pd5lVj0xJd3RGMM1Ud
pkUDYdiZlFULZ/SLpXg1CH2Fy7dDSftIMyOIRkw0VoCCP8r/lIc5+cW3BH5irqJpBCMFh2iFUQlS
tNeqttcKDK/VITqMBFCwUZn174PvLQNYLM9oVma02tNa4EsBiKcrZ/u0jo/H7S+9i38yYN7q4Mon
XvlUkOvOcwUDb3aUotXxi1L6yp9h/NW3KSAyM7pvG+ncCofYyvPJzIwFHiWwjjdJZaGWASl8yC9Z
NPw6ZSmKavenknZ9vQgZqmR2oTMl/qGHHSWFXlWMKmIh6P5y3sV9+sZCLfxTqHLAP7ZU8nNC2jfg
z2NEEEsfLkhXvqo4ou+X0zu8jfnqMWSKBKimPS4wbd5qjbMnVETZHWx1d4aO7C8OxVRH1YUcpPcr
j+PxZcuGVC6nY8EAXKJhr2rB0WRk2DhdXH0y94wkfUNDxbVg8KlmuAQIIdvhgctm4+/Tta+W9++x
5eni2KHUuVvgsoGh9y1Xucopk5/eI/fDl2EgaLav66MNzwOAtRrYBN7qHT8t1tn2rNFP5g/84eaI
ZDF35Q2PvGpWN98qsPQX5WTsrwRw2Y4bpMC2VMF2sv8Qe0R8zSI5PSQ6GB9cUhOESh/K0eY/QbSC
UJ/LR27n2Z7yu8uQ8ZBzsjIbozQ2ma0JeQsv0vtLvMllgd3XmXnefqQE8yd7Y5taZktQZIY4BSZV
EIMu7fz+XZJQN8nIJJlt3lV1PL2PaWoNQJ0mfDB8LglYuP50dZO0B25Mu7iLJeZ9ogVYk/pkQxv7
Oy0sGe8nCtiYnY7M6hn0pL4iHqJ/ezL87JTXk8elZXd+NMioyVFYe3mp8EgsqzSDrujSrxqTTchs
nnT09Iw5aDPiVF65Qy4cHSrSzyQIiH5itvFHQeWUWRIjipxs5RQstjrz64G9m+3zaeApirDMAfGb
GzZHO2m02MaNq1gfgR/YAUbCpYVqfYnnvbn3pDTfntefW/i7/o4mPe+iRIslU7kJMTrXDEtsTfaJ
ya3yGU3VKvwa+xZgCftP0//uOH8LpZlkA2EKHATKm6ALi1CFzZCHIeOa/Bzyom/TOFsoa8PEkrr5
26PRPIqm02te4s2q4KWOqUoT4s4P0rGe2UbaKiJPoLbkuwCZioJRRZlZhbYEIXXceKLwRwV4LUuL
n3ZUeUanN+PBYCLQ/INn/23X2WojzPJtjnTkwW9YFinGTYCuvn+bF+hiavQ9akyituaiWvWO+LoY
dcPndjB58poAAyv1WojiLo4wfFFueFqKuWhQzH03035j32VgbHOsNn4BU1++k04quYDCpPS2HZy5
6lLMUhTM7sfFC5zVXU8kKqtdmXYcCM8Ye1AODMlb4sjflEcuFX6oS4C4b7L5v5oPFhVRFKR8Vpdl
ZngMWkAxWWSDgRVTq7+SVWskr95iInYFv1qxU8JmbKbVd0IBLVAq4cfebFk9n07re7DqHx6/7eey
YYP274gP8JVWoty5v0MZ8P+kj9yYzIbbXLoIrJrMS+xsCSPTr5KsPr0UW8y+e42VV4NP4QbtDAgZ
BFFMgvNIBYS+wVJGyq8cn/1rMYKD62jV/G8YpCER76Tm//xmRYMl2xRMXguo6pITfhnBRXAApEWB
4vWJo9pllcZY7VWngnnRM5t909wvyHakXHLx/+roP/lBNLwau+eh6hoHngu6l9f4u079/PATH+GY
2WRbAimbmEzgRn9nstgt4sNfZVlPYl6gXRxjlTQmQ9ZIqsa4Pb/QyvIthF4vsUsELfW7TpTkx6iU
ggdJ1ql+KFSn2IyUsjc2JWP1wyW5M5rDNYyZemKiqYOv9jbGUpYVaO2y48hm5MH6NbG+FQOHJWA1
ja9P9dF+GONRpm+EIFFoHncniD17K+Wo0K406HMdaTmzWrvVhD79eFD/rE5bN8dvwzTCq3nI7lHl
Fa9pPGpz6JLkMBj6zgs8V0GEtYMakGOXiOVRK5lf0+fs2gUg6uT+5SQ/sbW6J9EH/21WbsHSXnTs
7DegnQJH1rM3sCHah0Bug6CDwN1BfHLtd8o3ZHb2DGkD4ITtA7ilnlRB3Ak2SfJVKyFd+8RfW2tr
F2gulehrt04qT707MWAN5SeMA/u6f+r+DmlCZjf1svdHihIWszdLXBoZELysWHKszrdo81/oTWYG
Pj5z+y1nJJopMIQxY8lHQ8U2teWlH4m2aYy1vduj5o66MZ66QRrHVGsa/WyDjIg2kY4VaTDfQOkD
zlNQdwE3nFi2UF+atsiRLhk015BZI13qFP7lqJfXHh0U/4ch3SmZvHv1TfHqZeNJnbeI4ydH5ROF
FmTP8VKO43+Ndx/x3jWIC1dYfolbMCjpdSz9MDN9fGnjDMEWSmQVrX9dXlW23kBrK3we5/J3pD0V
WD6zVeXkedrQQympiU0UZbtaJAg7PrUUVNUREl2QMcNFW4aPI36d1IgHA2zEEeYlCi4kidU5zIfw
79k33rOSiPBU6NYBgSDisNxsmAwMpbfXpe/EItdTbP1G24YusLNl4j7fHQjkrrYv5MI0tL54UdxS
oPdj5SiHJQ301V5a5oHyHFouNtZ6OQxGoNp8ZrMenTyjZ6WCn8EQyqMrnvF+c7hs+RWJSXzGMpmC
MRMcWqu3/v/TwcQxEr+ky1s8YYP40dJkvonAiMnYLO1sXrpwzPVyRPJmqrmgjdxkSGCxogHugqlJ
1iqyiCQ64xbuvLZsMFZHaYT5KU64gHRRXFOjmFvwgk3vGEmK5XofmnfeoLHNRkQetLbcuE24ctDw
phdRXsFLDH9IyvkuY6BJdbFVAr3QrnTelM96VP0j/Xt0WRS5e/RR35Vb0rPsZPeCBke6xGaSkPx/
/aRiu0QNMee7Ee9QXteqeQUe91Qq1yhFrj00mijBkonAY/VGm9dXYDJ58mrTGM66XvdkHxLopax4
GEpjzujIs/uDI3pvKSnS8DAjFq9wYCTkacPMNZE2LCjoW3S3l774OoWgrnIJuIYGZ/m7U+1txtAS
eSISKbtp9lWp/YvxSIRLEhEY4GOmNvAu+oTsX3xxOIBK2Ir1iRsD2nT7ZR0jeKS6KQnGknkF+BiL
mEpGtnkRdeJGjJCntvxyeucGeD1/eLQ/jcAKTSNzfhzXbdVGjJPuh2o1OTI+LPiPvOi/cZS0T0nq
1V/rhICnzUX4cE0Gut+dHzAd4pN1cTPl5STfmGnF0XAUF63R5n8/Jtz/R+GtPUhA1NMXNoH4XbC9
6f7JGxCR0rWjMLAfDYXMxACyVr35qDXk35PVddeA5bCYO4sTmqiXc4xDkng/6k0zGciY0/TqcTgd
H/gJsVuU6c5Ip1qqExKlCdEJQXStNVYB8Ts107TcpxS9yf2Hsz91YNZtbfN1oI3qFxxwrzpoup1T
ks1S9AouaEE4Ijyv85KYSw6to9XQ+qCkJroKT0Br25HRcqoQ8KmQG7LGxVv+/MmuHb63u2G6W1Cf
BEheFMkhrfvQ6Ew6shRYpWHu4LM0HSPwBax1WKSzSW4yROIlqSmoYqasc5sGSgB5MpxvHnand389
jj57QUCKCb/VIxjD6Slt/NiAAliqXgulJVpaq+Z83cAmmDRueBNnjdFbGPxUTpvFer9Fkc81W+Q6
mup3Bk6aRbaE+a0KUOewXSz9BtWMdhBYNU7o2mqdtJMvTtvXtt2nXMOkRMps/gik0QvB9UAEuBh7
JjzTpgJgoQMP8BdK68H0xJtKAdVqHUZjxLmogQrjAR4+j4WTP7r1C6c/k45c73z5s0As0dSI93Jv
MINz2YbfNxCuC8QxeVUZRrufe9RiDD2j5A9m3D8Kqsbn+gk/kL06CIOizt+6bdFkcIsMxKR3ZKak
TJSETuAUiV0sejmbIXEUzfmriJxrCi87S+eGq4jqXmyU5zG1vr45CzJl7NXNMDUxO/iecZZKkPru
z2jzdq+0u87FVLwKhiLF0/clG2pczXOgoVf8r+VhNG5/RUKEwkgSh+bYQrZTIrCCgVwAyj8y1QM/
MnR6FIEe/hrn2O4ZlUMdx9js6oBfOv8475NsWsD0mHDGtgeCXHF+uv8FISdxuRT+hmAzyJVCvmMO
kliVu0cyrjcJbT9SXTa8eSy0JjKhR93eC3YM5iuYTG0EPILH/5Gjpkm70Sm5JAPbQd+X68FF7iFr
CEBAW77NYjOLs6UvNgbDM9LaZ6TDvahn/kYZYCKL3bAJXRoCEHfblWq0uVXSzGB7KF8Q+EPtDGw7
sh1FBB3ZTiE88eyc4G/QX6aVHdHYvlMLtRncjxOY6iGW826gDfP/koHJlKUkwz2Qh68L3PwVVNXv
xaxYYTOHeakNnnnUjgjhtF43mfRZ3gZRZYBKdd8oIPtW+7vQODTwF7fe7AJrBdohk8/OqDOJd1v6
SctCBwI2IjpTMDGUjn0TmjIbAB1J/9HLEEX1jbfFpMbU8yqyQFkoWA8hh6M5uOjoHNactV8gS2qw
6MGQFBRzkTBIydKtgndnnWBtCI0+2eeuArNJF3KcSfJvBLJ9mWA/HF02yV6cryj7riit7uKf/6Oi
qQjIJOlMEXZmH/x9cYq//t+YPJGNIQBPZ7azeLEbIS9GNgTx20ztoJMraNVr9oLVoz8tuIX0UOww
8BcwTvuVH/a35gxueTTzZXXzdOsfKH8nxzIPhcd6szih3I28ctq6Bni8jjOdicMy0iaxSi/0fA3d
+21p3LZujRKZ5GMhUTF6Q7sktZaF1Zfz73sbkBd9q2Dz8pMgN/DFeCraxqC1DeFPlK7CU7bhv9SC
OT2N8oH1OGz1XpEja+FgZUeds6gNgTCVO9mfJ6XjqnwDyDYa6ApOgWfQdfebzr1upUjpg8Js1kLy
n1M2yv5SDGN6CDILpNszAOLIitf09KhoJ/aURnVXMQEwNjWzj+eR6LzESoll1N0G6f4QF0Y1rlKL
mSPmbpfh09LclmwQ+nGnFBzWo+jpY0c27/NtBHtaVuyq613YIYa+2WVLK/lrCS4hOLcA+r8R6dhL
rPCkFChuaEp9JIQsShuzb3X7p5DiW+EA9sgkJ9H1VHT/fvHfgjJt3tD7+1SZp5r6wSWkGkd4JNj7
qUMwmMY9aZ7q0mx6EOtGJ0jh91V8Qazax8CYT7lNyj0I6aaD55o4O4GF2h8FaLidCZxHcrujfFOZ
0bgulTbusZHs5V/0EckJjQYJXx5KlvIfjVXPmFb6SfIaGI6JwDvqYvZ1TkyI0q3CxmI1714Cwbf0
kXYMqh6B/Y145jplhpbNSuiXmX2QbIkkczKJS2mhU09QBFZUBFZvoWyEX5XkAW3HTuaL0BeOevyi
/gGb8Gzj/BC/IKlIEdvYa00H8k0pOadGZ6Tnsml/cGo6xaTJWMd91V+10FcR/dnWcTQL86InwWzY
UJoaU+cWqUrDhPWfd09YS8bHgzlvYmR35nfvV/P6cjGeMjpDg+TI9ldaNXUoWJZAxXimcUGXN3vQ
GJU1ijOFLOCSuNUaAXSINe/+QlchDyEDvSkWV4CcT9gqY6SHVwocrSBw/qQRwlvs1o+JhWac6jFq
aC00QpC1qxI8JqPD0ajjX9aUt/8VyS8tKWj0Efv+qkVw1SgLypL7rXqdLK5eiPL1YwvS9XH5LSeS
Sbum3tejdzhFZpFg/zXGwMgNfhbHTbyazicFeHp07iYi0FYwfqNpueAMtIiVxgfLJPuOPUO2g4g9
cgDhX2h1a0RtJmW9k3MHDJyFWuLZzLkBHlZiJIGcEehW+kiHCUlnqh7ozfXeBYAvQdBSg/kC5iU9
vhXN8DJOI2TUPrfzdCHn9Pn4J95+CpBwvzFC9cYfF7Kfe0DkLKZNqn7Ba4dTv47xyefnarXfbiEW
JPJOABGc2IK1EsJ/vIISn3XkCCv8lpYCWY1qRyB+CAJNS01kR9kVgkPHk8LKVRJtwNLd4QvZDpnl
zq2ApqFVwmddLXNSG9QWc7kVCrWNcpet/ROUHGayjC4ECO/7yilGxGRxLhYrGXzfSDfabup/WKLH
YN9veiDbE+5+TyWKZA6Om9TxVuhJp0Ab9qY70WOvPIuGztx+spOtbPa8/h4MxbcN68lAfQgDfio/
0Dj/05P/UrlH6SbK6Oh7uu1uCtuIEU2KKvlmmMCkOsL+z2i2jTgfKlivXdup4l0hWyEFMBnkAS4m
bgKc2lhQoJZYAivfG1s82IxwprUMAwL06kaF71g03eGj4YKcLKslD4nGn+MZRXzfZtLy0BmLn1Hs
3UDbZPYxVZL2htRGVm8w7KbIby6oxFzN2SuUk9LL0bES5LIHyPRxOYCMMHLV1Fh/WFIPKGxI4WEO
Wn5SNG+BGM8h5LbBJncarHsRIv7XgiEIoKTOkghlsL1Y2xkdtDdUcWBbMZ5bSxMZAyPGk7gjT6f8
jyfAB1tMVEZGTyHdkVpjDppwV8u8FAHSnDOm02pocLpc+vGoYFOI6DoseE8mgTxYywV2IYgLlvm9
mJgxFc1qv9XnwIea9FFZUB0aJ4i5dFtoI6idfYEDHXy9jx9D0HJ1dnWRfNgS8fVi0Evim/30t4Ad
WelTHS7abxNuK6FjEIeXd6MWdds2ipF4jrUkysS3q7GLLmtaSpxiXV9iNgXSI7J1iPELL/C6T2Td
XX0TmKvzflHPzhDBWyOdzKIRVk8upLC20Nh8vIHmMRNtqKTgFGgApWJvX/SOoFzDCe9S//FnbSxB
n00Ae6vr1565b5O3AoUGFLjkFTOKzxcZp7lSDZrZO98v1WGqt1TzaJI9RatrleS9WKpBF+S7eNpi
xgh3T93OrIcielrZAdzJx0Pt+TVWdAY9dkZRwJUETxVEevFBvGdBOAzN2GyvJr0lQtVQxEGyPZZY
fy1D6ErwfYFDYJ19egacP7/3vKSuECa/SX07gzff4lC7coeVM8WIc7kT6WuPBVPB0Gvz0lOEnt0X
XrMHAn4BR+UfZ3tBdklaRc/xVVKdmU8xJPrbpx0yg0ktNIt4A8EjruTfmKbc9Jg+2KGTAncEqOJE
/+jn2Qv+MxzGsUB6FVUTkMM9n7wEcqtiCpKliOlz2RnIQa5/IZukxdLGxRWpmgiRWXy1rB7BV60d
cX28VahhQFEE7KbGM7Oz4zv88kDnNbKYemOkWDPqRsLWYvelwlbUy46jhcFPBtClYMSmzXy4nfbc
DLYVKgxQHvsTvVI+blIO/lplnZkhshNJwFg/OjBSWz7XPRfErUIYOQIMPwchSUT944OcfsgQ/Lms
GdCYxdpXsXQJlRfb+92iMhFUnF6dZJ3k/wZtJ8EICDanrIrrsKXuauWujMsDeXOY6POiy6PXzn3d
Qqq9NDNblyWg+UAc2BOBiZa2x20bdB3fGfod888AcoSS4757uffl7IFB1crkgkVL755KhtVEePtt
t+BM1gghUdcJxF8TLFyYKaWElancIsEN3M2jX3k3vvkogU45QafnJ2qU2m/HpoVkLO1QcgBNf/c6
Is2jT41XTSXo0RfEDbkfjxThNxxME0Zsbj+KFUsQUXwFQv/ZdqYtVzuY8GI6OIQVU4T3X3KeV4t0
vO7SX07EOvEN/7gEcQWixy9o0PH+ARE2+iAKQaBK6Z6rGws5GeQtOLQY3OgY1TD9FjrydsB4J3x2
QrNOz8yTSiC6QKWWZs4nFUZTFq4kEwXMN9p0Cam3QiNdbHaLBFy5SQoJqYRb4CkQQJVGj2xPjFrU
IrzIxAaYNbYtEgveyGNivJf8ngUMHABjpWkJgeryxdF5brOcbhpsSvJp7+X39/D6OzfrM0Dz3/Gt
AMpGCYXyUQxsKZlLzkfsbY+zbjRu0+f4CD2hwkcUuv5EBzQWez09wue4GDuyJpx38wmpFkpcFJer
0su3g/ys9FKDctD6FvW67R6dlrzLCkhXTAJc6ZUcsxpWTuLRNKbyyTs0DlIjrWjU8u/13qQmfDzi
psR/ZCqSfoz05hmcFqeH5ycGNrfz9jE3X1S6rLRVOCQIIgxl8/z0I7/vcp1p+CUYug+mKpA3XL7b
3PYuRHqfNOB3zq9+079j1XXwUfmizB5rNwT18BQGDfOJdwBsgZO1JB23vUhazhtnqnjvFUdg+W/C
NjoXIsIR+BDR8UcrmCCY7tuUF/Zx2jQ/M1fC8E0GYOVryiEmAK7cNsDyvZAI+zRJvMrUmjmzFcR6
QTUq9ROmfp+7h6HXcIK+U6ShvJKaTe+m/3RYqfzrU5CD4bxmsFvUCFHLADczNFwD+9W5s18R6AdQ
FQXW+fQhyYvzvDliP8Vm83ml83l8kaS31ctx8it5Y1tp1UPEgiSvxb+d1bMqo6pT114RgZZWJSsh
JQp4mQJcm2557pDe2dmlwJ9RD04RX2etwEye9zLnJG+YUXJb0glWHI6wIdPkN+nOBF4EnZHRtPg8
eR+fwZ8hZWlnm/knG63wfGiQEtAHNzIBvo3WILgMJAVw/bwxRUEsDru4odU+c2jiPkIASzWpdjbr
r1EM+771ccDNN+FnVYfI0u89MOt5xpp8bk2DtQs9YKyyPVD33epleidqAhQDS+h5TM7aua/b0vGI
2ElJGFs5Nx64EtAyP+IxTKPl0J3n0AmwYlQrfDqCCHv0fOwR/7ZlluxBi9wAz7zzxxRRanV8Bya7
iqZrpkzF0RwLbOWe/D2TBT5j+geczfkbluLo5KqG8kPtqeGqBWfdR5QpmJPQTpcmOkkpdepwYP1e
x89k23nFK89CUqzNEP+vnKdH0p63YGcWva0XagUi6EAXRjpLg9gEwVJJyWpu7o73VufNhWt9SmX0
aDE1FS8LvJtLaVRuC0poJIFL4we+U5C+3jk8fu7uKSOiDDPr2w0kkTUQi4eBDnaNMoI4hj6to9UP
NQn18+dMrFY13C7CJPBFeuwMNp6QMbe2apPtS5bPV6msANn7BRKWN3AZn0/2b8q1hleeRmp3zO6L
ISCJhjUTvCL6uNkS23poFJ9hAFFdurNMcF7j6aFy2QP21ExR1+mNuUbGk/qZqfXgXoZzHchdbg1/
gCRHSvMGQp4tyYjbm2hPikw9Vn+odfqVbbVm2k8saW/cE2SDZqErWkxWEX4XA9mN49o+kxegdJ8q
8FjvH7apr/c0ZnaqZi8Z0dhXrrbaYJGgG6+DL2qhJZl1YUBP12gEUJe38r2fox192MwRj15+RT/+
rHzh1X6wic0jQCdcgBGd3m0rTgKUBE50lc1VSW+tFCm4a4EUQLHnI1m6jRNDSzBMeKh1+iGp3lNe
px4mRpld5FAqcETdFkilC7/hLFjQTWUWaJAQwV05HoI8Ccu8RNwUJFzCtTJGYWK4XvqCvuTwmx5w
tC1pChJBylDIlhD1SC3O/ufmtLQtZUXyYYB52gpPV4fBCN8gipIsMDD0uw54+vQkucYR1q12mSTN
5WEGO/OTVuF2ptlrZUJPtviBfu7p/sISmd8LKtny+yTzSx2mj2S4KAL8zH6KqB7ZuIv/Wc6J8Jdg
IUAPbdyeEWEu32+mSOBPHklU/RsEK1U+e1qwc9dK5DW01IcOKf+0cePxzr4TrQ6KrAW7IRdVPCmS
ME7Wih6knCj+wr/hGtVnvTxGItBiAlJN9hRvJBfmyCUjthVKNhzNTbs5BAJVilkvEXm0hieYaOOe
k9K12G7TY6NqlgiDQDGctwjm6QwqreEAv/1j2N8+lkf5kqrz1KIgTiMeZedtISAGW5NsJsrPt2Z7
V9msuozFmeJlNTziGU3tDOOsCxBuVp87HfYOzhby5n2ZoGd5d2yX6Jj1osAPk/eU08vlYwt/E5Wb
iqGIcLOOzZrBTKsS0kJRv+0PbjbfKkr5ERsE7b5u2PkOxiTdRORBhtk9YjfO0D6Nj87hLcsOhK95
44z/bYGXTtt8CMJniCriS/w7ML66warlXbSLdnalXb5txGh9OL5TPPjGD10nTAOu0Dy+Qy4gRiL4
Y/PjKeTZuwg7rf57XEvC7k6uJktBCMZIG524J8kc/fNLlUUgysn6mbRfPeF9jsKLheHTzh7FfhEd
fVOGOgoMF3PUoGdNWsvOlNIRCcdIobIgQlA52PjeaN/iIBuZhm+kdaC6hL6SLnq+byPKQrHXiTrA
gnnOSIifCiWW0iljyWDm3UXW/vhdXA7IwDnPfcJInVJKneMatJzaKUAz99zLV/3pChRnnKdstuc4
Q0NrdWgOHBkSL99KdwEOkvQ3296ZNms5/tN8FWXdMQTCJmgY7jgNx5oNxC1OJQAIH7sWbwLoKdvp
Or2CipIvi/GYBqyk60V4LW5ToyHbnpRJdkKUmRJOmo8+Q0ZcCqmR92YeY4hIuybCKeWNARTY2Bli
5d4jRJ7zXbzzdZz4iIGMkBd2HPFaJltIjxp/H7VY9uk1dQECvliq+57ixz6g249XqmTFs0P2hw/h
H05Ri8ZB768ZSv/GLMrHWe8v1YxpkYlRz2P7yjq1lo7Xl4toTWdOlshuTuGiHORuyjHG0KYVd3RX
QM6O85UmoKx44W3jK/rMlhoWiHYwH97kIzg65jfoAvUOLG92zmMMPHKSc1hmzrgUustsb0LySK2x
Z2Tt5gjxsomQ7JKV4uOxm7R1oxmvnymg9jz8ajxbCrJI3YMICdG3ppUMtKtqMkLenY3pUIihSQ7o
Q98nmhYE82UZVxOioVqLl0qD6u/JAnAo7Wu4ydvz5BS3RS47hWCzVitRM8mnxQlIABm2wvr/XAvk
9halNe67LDslVdUsl3LHKOusbxF8hPBBDIsl9IZU6GlHTd6kz8IfodvXBLbTBqqvp91vPsmIVKBK
eiRTQHWm4KefwB5TqNN57TCd6QYtlMp9Nx/GS3xWBZME4xGkhiVCZpXGtKxMYl2cr6cmC2VIU4fO
12SIu24SzIsSRHnpQNKirK3q1ZjdwB+Gu6gZZwSr/rCcslmTNl3uOsT7PxGW6kRlhI/kuvuUGx4E
OScwGTw5qw73I2vbkc+dylPU3x9hVqp+MLJtrpcUEo4H6MokKM6qf2O8+GhOQxCFKIDbptzJVKsJ
9g/FWD4IcwyfPfzLV9i0fJVWFgvtuHU96svVZbMD9y4Q+yNV2kMIPps1sK8HfCp9LGCsk9dc9IWf
qix0Obb/NtqIN5Q46ScyngEs9CeFdhMYiEQmoN0ePD2E417nQbBpAxHvJALHIGPcP0UfHxuYnkJS
1FeDEP+UktWAnIeXToTvvfwQ06JnHPp2kZczL+/EbOT1U+wpO/ZGRttt4b1xA3DhqQOjHkd/yUNI
UtgQmZwroXPZm+f59YpzukH3FDknDAjKJ7MnvwXHRU6mMLjVrMlkgaG7c/LOXpNDz6c+9mefaJIa
7oxmfC3q9E6z1ZFA+FOE20JQkYVhWDP290JL9mmplMycffTXwaJrXOm/jrqUNGpH/8ePPlYGIEGE
Au29SM/O2uydczPLi/bHcCX8yF6E/UL/r65QNPKn0mf/HH80WLRVjfx39XR/wWU+SQ1y/FFyZjWt
RnMVdcXPX2jblkwgt0zb2t/uOJJvoF2ogLkXK1lCoacEyLoJBwqFs+nDb2c/bMprdMQN1YACxXJA
W0S7PTceJ+OHjHEKWM/C+ybYWULH/3gMAb4cQ399ij7JXLHmp4aUp3Q3Bg6zZ7BNW2jQgfVBP/tS
OTkrpBzw0Jf+dAhVAXihiwuJZ8Ys+6NyUN2KGNKx/A5jzrm/Gpodz/ucd9T4b5LfVksm+ltxFEPm
AjSwWeKROaF5lXb79Fqp6MgqPRGwsJNPmqdV9WhgCxCvnLialpYd+JM3q8ccoA2pj9xjV17ChPxr
7+zyPaX7zn8AeE014Uusl7AhCfVEfdOH4yZ3bH7VFLe1d6iToftplZl6cuLdbfPHY2y87LhHY6IK
kcw1rpR20wUn7j2quqR/RqH4EqYypfTaNCMElyRIOIVSZIIMrnGC3xp9+ZbhADOdTZ/o6J0lKmox
TfK4v7mvmTo4MW4I21LBxhiJYzZsBHtjkBIJlXb/BEqp+onb1Mp3cubBSELSdbcvTCSCKbl+G1Xd
bjxTnXWBv25ntw3i090mumSC5qVHy1qcCFvUJ6tEHXdyNQP7VKuJE8aiw3YFN7IOJn9PzT/wsO2Z
my0JB0z3TGCeN4qWcmD+KkeanAO7ZUBbNykt6Yq1xVi5EzhIfaEG1GIXdoB9u7OR+7OxzN2A9Xbp
0zxEH0EmSU+gwDpOz6zL4x5/8SmKSInmpz7Drpo1JX54BgcEubCgjS9VA46muHNXJFddWvEjh28l
Yc1n8SxLWSWNl4w+CtlSQvfhzy5jMpZ7QNJUbIrqOgCamwdCJnf77Y7ss+EYRi7CBF36UPmhrLT8
VRaH9sfRrDDhQ2vbNPRLmBguMyEDcxiHtaUiHj9Y8ycPYGp6RY5lEiUn6rMxN88b13W6cPP0bwWO
kStbfcJpE5EIfWj2OG7imh390RLzc3lUJOqaG5ox9USnGDvtYgin/JmQlQCJ3goqBBNXElLTaurj
QuNd3S4rsJjv897JCndxFn610TVGaQfHLVnVAU7Ea5vSZjXB9/LOd0pzk9DJ4D+7/x2KwfnO3/Ve
kIqwbndeiiVM4mO3jPlC2yA1dQ1fHYP/DKpnpWj12ML4l29h9f3NYanKf+XlugmqfDXf0dcOpd1d
9g5UcsLo2BzUaaHNkdGuJvfNhIhVZ7ZSBIVxFmeHvTOEeL8XXuhjFbc1VLFcT5Hz8dKfUuJuUWNP
dt2x55AYz4WeLbIUCbnaW2f7dKuWnBU85Cwjomj1YVc3t2ixSr087qIhpBc/T3xOZJCoIvkTBaYq
M9I97Qw/KHoYVPsOgqp4rgLbDCjo60aZCBJDFjMKUbEoOzcHEjrPtBBF1fm+NSAlUnTJR2cANHEP
Vg4Xwek0HGRImcgJ5duFRMmXdoQfN3PiB6D1wQjnZpAwznax2DPwxA4poTgC2X+4F++bWR0X8A9v
ez7BW5H4J34WAstIezZTrU5a5GqA8Vc+rTHIAmVmlVZUDe2yeLml8a3rKCB8Xc2MmKWNRIjMgs4O
jrvNX4c6tULQkUrKDuZ2YdrPZ9SIHgFfkNFfTebSVizIurgnuMEehUkl3OP47pVzeA8hPhttNmJw
ETzH21DlRFjDUBqPJiBe2nKu1+LqWBUM8x2b3pSCCwl2LJ0ImkTgV9xxt/eP70O1BViri+wX+vqg
XcfmJsHms2ioD7DW/kEqQxv6nwnSgCx4j6J9GZbxWia76mbYqrPWPjUxtnQQkeVuH8Q4u1wo4rYP
Tq/fL/p+lWRe+n6a+X8dIoUTNuwzPK3EuhT1XeqBip0PCYal+AUXVLdfhmstTScVv/2NwZrSrdEg
LQF7fqAHKueGjkj9bsZHCx3S6xs22c0bAmcfGCEY55Rl4qnKZrFqMDhHn1LMPFV3onnmYPTfgFQW
1mrqF2vduaYn68CMhse4zbvsPCcKngUVZ6/1ocUX542LgysVVcm66oa1WyUhtgFkov4xdYeHbRCs
072ox/bFiG+5yrk4mtJkuddsvjULYX6bJOFS3LLsSy8ggnO2aAFthVy/l4W3wM/anxsmYUdqQ7cP
Y4hLydpumh5tWEyOEm0frK0uvux7MRbaNtZLtuB0R3Qsp+dO5FHRygwMe7Ba7Kj5giHCRgEmB9nH
vvgrJqqpgSZN9hoqhVTVOtIqQfL3S1irz0L3Q4mzzbCLrn8QowTd26WSO4WzfOLirPEyuT27aVlM
IsgoHzKxHYJfMNR1x103ZsmpBWYUZk1p2j9TyYF5pyD+OWXTB/5Hs0HeXKS19YCjFKgxLBcOC034
szFjbGKIkAopA8166zFf7PC6tVL3PNfaZbBf0kprBtPR2aoCNJiid/8iw36M9vWq0tg5hgjyzq8N
ZVdS5SenxqNayxgaBJiMnWeOB4u1AvUodXhmtm1iUHPxP+ZKUZLqHkoVEXmCQcy6BqbIb2EIi3Cc
+Lmzmpf9bHrQFii26YVptP9y2BkMJ5GibkdJABgGCxqk0QQBvYfIo2prKRT/cLR7wCLIjej4d0U1
pfgptkzN/qy37LXQDSWQZKmFHH9Hdw7GvgvH4LQ7fkW5EJtcxMUo1R2va+6vt7WWuPB5fi0C1irG
OP8jIH9gvY7kWbqcQLkB1n6K7fAOfz3ZlGdKVpfqmYqrWgZjSfxkqAixiTA6pnY49DFI/bBtUA1L
UM70IAT0vBCOzgcguuyLXtZHzglaBFAR2qzwZILiLSnumW0V5P7C2Y9/x4EhR/dgG/Ozb1hyPeoT
+3/xWLbT1OCUWMXQ16jhis74G2Kmz4SPpfJKuOjDoiAkKiSYUB++eZcfyc9wljB5UL69a9EJUxbu
amTZsjD4zXuPc8wT+thfS5D6WPkVkYlLXowSn6fCm6hI5YUiPKl+7mMjCVg4OY9biNMsBf1vmFVv
NaLc633SjbuEukSdw93S7ARMu6WNvUn9UsW0urGM9qSsA+YUzz8rQWeKcZo9nbeBJTmaNm/KZYzl
h0/bJb5aPhG0NDZK3CGoC/wepNGfqO+N0fFIKPnSZc1nzspniSsET3BTn7yB2/jkHTYthLq4tZgP
0MT1tcOKZFhsfq3E5CzclujddTlUhdm53qDQW5ZSQKedYEGNIlw4n8VyRR/P0lnMzJkcOuC95drE
Jxob2AXLtXMogoYp4juM+MAkXnjGP3RkhlENJ4btq318dJuKei8tWf1Sc0Apz0U3h9LKcHE67tYA
tn9/uuSu8kOru0zQgBlKAeO6vVqYeswQWUKUd+3AYJLyyuemJCHtN0ahmzIgQnShY8reGxPdSPS3
uEXvJdFM380H4PmIPp2KJA5NWJluRxb0hBbqd4WMEQ0wMehha4nA+TwIbl6ICylQDsmGnIq4fq6k
DKuyB/TshpZ2ehQ11yh7eXxBfd2iF72CQCxTG6oNDs1H4uGdys1+bgv61ZyeJ7lLFdyQdw/uupG5
Vik3VL8Qhri5cJ5k8FLJXNmPzSVsy88Cci63qSWQcPksidyNiCWkRI6kEMtMgc/YhGIx2uzZJfHI
A/e1GoxCSy3bE11alXaouJk74uIkz+2GGA3mbTys8xm3QnDG7BpdhyOuYU0k6KdFHzQqazxKnMVy
aDLvSPEp891/8u9T6h63I5GsCvFVaor/DOJRXGcQaVN1RW9Njzsk3K4lS+jEcE9oj/eAs/1GfZI0
tQrEuUX5VO4GpnQtz2KOYqLRa4dhp1RENE+tGY6vSy2mUOHl81Ln/PQVC5tOZpUbnqrob+fFh64D
iCqazD/S1dvxKBJUPfS+sr19o/peVoBRN7v+t/V2mpB8cNPmrv4kqh0lZK38i0X59cnKTX/F7BkT
kybNaXX+Bz1bzeAORRsBsNnVl14/tjcONSJDRcAwcd8cIPQQW5aFxNiD9n5C2KA8zxe2E4PHdiuy
2jhF4JwBDiY1n3tOERHD3sW/G9BB0brtt2bLqInswHdtddL01npEPvT7ID+zMEaaHqE1gh7xx1HB
lUwKNaDnI+yYTsd7bUMDddN/R38Pbo/kanz3RC16pu7HsBrKraTFMthcxoyWKjfb+sQ2AXQXt0+f
v9bnr+BGk+Dj2ZZSdGgDlIbYnjfRlHxgNKfgsI9IRkxSILck3raHlx6dWQbnt7cm4QYk/pZLy1sv
IkBd6h7Ey7StDD1OQKvMZmgNDp8/w2E7ioGP2LKdboDhHS6ZNqwwxRiNVBhkcl+dnvCj63hUlIQG
Plw15UNWyuXVmPeJaJ84PSKjADuWkP9DbWVt/etjs3jG71s4SpYeOV7M8uLOi22YIq/bKRjxTqMk
SyJl7wxhDW9jMS39Kk9KhIlp8GWOrGy+tuTVHNtQvzL2dJnZ7n/PTISpoQmmEddkwsB8xyXXViMO
1GbrxWFna54c8DYy8GSqFSnc5hItxbKHSghS5rLIMH2YfH/LQ+9LNndGGxC27GeqKgojfSNxa2qq
yG+pDf1m/V348borgGWX9NIsdwVaNaU9OIrbRIOGfb9VxV+Hm8Zutsax9d1I/IqSO2gfm07TOZUX
k29sP4iJVQNgH5kfXfKR0TA7JIT0oAxqkpS5LRO8cJ+yFz5HuJwCY2cWfvqW5YUcwjFdIvMVVjXp
u2BO+ckgLlQkvlgaX+yxTRldTUFliHBpRCnFJQ6K6uezdf3y2N4TsfA69L91ay7hpqDtlkw/CiJa
/215j+0vx323GUkyLJzkLpQkeGnzNs8OLCPkUhHNEk0XA2EIaRAYYlGbc9rUbsUAlszz/yr7OGyP
HGsn6EgqdY6bdI83PgRJz1IamlFqFBHTRQcYJEImQzf0tLhu6KAhWUOyS+JP3xJVIy1RtPGAu1Ya
Ed2hgVQX498mk1FUV4fRFFcJo+xRvQsTdJQvp2qIykqj+NijkZef/tu7ZT3mPcHyjRYQpHiTl0Ad
k+0c5jhPmOIcyb9NSsVfsasbROGNZiKpTPl+6kwr+OBM+cRKFCnpyRSvLNwQ6Wdkq5FxJJXBE6AW
j7v3lSbMHGhZKYkVRltDIatXYC33tqDRFZCU36M6oQdwJcWyP5C23qtecLe18Y9g4MutGIWRPAO4
Bm4KR30yJLrV+K7eVuxxRJf+8lndI2wJAUyf+FmUXvxF/J2m1un9I5cgPT3McXGPO/bsZ7V4wf/I
h+X7XTydpZZeqhSYWOb+haBwKYXBLOnzb1bR3aB4tlUDzD+EDiXT0oR8IGe7TMhxIBA1hvYvas80
ghVZwYT+HWpxNAE6LH8aJ0yBas47+Y7w0X78TSa/gwhX5fJHLBFJVAL6AzhCDqBWq8+lWtNU3kMU
BW21o1w6ssM6OpYfD2P8D9qenouI0MEURLPvROCp1idiqsJ21E2lL94svaIdhMari9hT7RZcdW6I
6JSCDSSt73gWjm0UyeVhVW7iiMEPz/vXSy6p4Bd3BWPNAeNRF4Q/boY/rIVM+k6HLh3pcZB2yauM
d6fJlUq63WVLu4KNPnj5CXiWwHmeShjIwIuWP7BVO+c4AEy93bUJCovf1sUZDZKNPL4G9bScexL2
4jnpc1wZAhLyBIkADur8w1nItZRvkcvzZswj9DlIQrY2nnOr0mbs5sdl8T6ZyFaMYXAX9m8+NOwZ
01pc5vQ9dKYqCa4/40WyJxCu7VcgVmwgpvpN0uR81BuRgOMjjtdplxGyoHpGBBKc+nLK7F3pMQd3
biXDDhROjXbG0wMs3JiT1stZ4Ql9vPduHGi7WBJ0OU9EK31mVqEepw0SvgOyM3DLoVgV2GnDKMLJ
JHHjR3e7CO2pmpXLZcvm3b4lG0scu9OEei/wjSltj1/B/d12TpLnee4utV3fdr8T3zimWByTugLn
+kq/jkGCrZjoO0iSCs2xnItV3IwHf24anbaE94tD4bK+ckPueTXGB1wX8MKEro+pDQa2Emw1Geb4
KgxQXtixrW9ssHexCyGcZUw4wr2XX9LSgbPaK3Rp8ME843FN2XKi2M2HlK47assnffCCmy6rdotb
pwVvljUvs4gEixZ/JyePeKirlaa3eMP5s6mB5xrSvAo+l+5gghNGYKjzRCxzCvdTQ+1TTMHTB6yG
yI3q2FVgxeKRe0v0oQGL6YJD+hpwz+7pYRHpwb9bv8osnELpzxwrJmE7nx350+AUxH54TsQ2/sBA
UO+IyBaRZLV5sOKW0dC/Yb0KHEBjIerzxwZkLijxsc8pBqP7NS7idUNgt6XBx2N9nhL+gs+pj5lK
F3dY0sOQXngCE33EB9BCPdT57jm82bG+8hxhzKNQWJ2ORfYOhMInqjPhe9YCCg5HcQOWZaknNNBs
sRCr3eAqFahFhlRGIhpCHDxriY4sjh3RTiRt5QG+IUsLU1lydxdmBtkCO7WY+uWroDElXKvtSSmS
a5Zhq9RFcfvIPq8gMKrBbQhomtqzCSKXi3DRGby6Fhv30Phvv1Mnyn2n9jAe0l+Jeyk09tKs0p2L
rQpQ7uoUJUNL3T4o27BJyb1foXWZTPjk0TwvxySkpDlnHoUe12pwtS7V9u2VIpH15JEax8nV0267
LIpaVhw31ewv5ldRkXqskeJ3RufLmyaF6elMHfqgQOmMq44iq+jSdmuG7zUSM/BDnFoAK5/Uhhy3
TQqsOwHOaHL0nVYqTt1GQHmZFBDydiiOG2ZEeHAxiId6vszdwzsIu4sEkjr2InQorNZ/hJRAuXZ9
WPxSK3BItmZbr+9QAmX05Tt5S7mNxDDBNlM5EYKhxGepSL4OIfFitEKYlSReSw/bf/CyjjcAW68S
sXHDA2/h1RS4iLGqL+qQHiT22ZXHxnaWLpYDiXoKoasgDiLX8ctDyNQ4YBpvIrGxe7DCbqRPcQhs
AkrFb+N8F6En6ulfQYcw635iRhFBcXUYRKhhMbqeeivZki4232aUcmq+8v2xifsT+sKNhq9r6Aeu
YQxaHrFXIaExgmeDQMex53bp9fk0Wz5ND0QyRn3BN9Ff85tvVRnZBajJkEby0bjgxVowPZ3e1KPC
qvZFoQ9/SBYKda1cAwafq/3XJ0DEUIMRh0oB7kTSh4xYXslERRsIkWgyzXLizM8V870gy6OmCtJ5
jusKXOQcuQM1WFhccRMKaCVCEXX4VdwTxUmr5ZsY65jxQ29q+EsqRxmDXr1xtmG12pa7do6e2S7u
xs90v3rv2th0gGimfbtkd0pG1BSxlWKkthF4K5sKFguMOuyS+mgt7dzPx80pi6MvGdXJ0JzfUXQn
3anObOA82KXf4te4wZMuZQUUruT6TUWz0nymZrBIjEp8kJzpPNl/stbdqFFArIKb6IJoe7GVeDGK
yihmPWZvLzVulUjVLnx/kxVFqdS751sCrtsfxVyGSMmu2wnPvPT6o8h37CcA1Oacu10UDT6qFSPu
UHk6ZeJfi9irIaLEdMh3drAvKvpSOPpiBxblFhtiZFKqSfhKMIRNpr1WvyX5KKViYoyZcodVwuwP
4QUA29Ftrs6PxDuvZE3O09OSUiQfrUYzFo0K8lNBpa3NPwxMm6I06NXE4D6kTAMbqS0SvT6JJ5ps
yt++6LNSASz9IzsDzvmVWD1P4xG/y1J404MGy/NGe5ESDCae4Lh4TM1CQUFgLFBc0Wc4z8RlBVsW
gvY2BglGiYORcJZXr1brrEUon23E9uwf2aaluoZPiuilbuFwR2n7+n/Z+mK8e4tilhCILQVZj4nz
NYQTerMOdDcJKVRsjcPNEYnpAN0m1zGI9UJ995EBmDXpLmaNPX4dOcg21cZRA8TjeRruMp6R1kvU
yx/nxv7AD5s+uGwGoojJhoVT8cF2LzhWCGOc1U1ZPRpoXGT/j5ylyGzTrnA+XbTZcIm7qMuuEold
Zt7XDmmU9wQq15lDCmq65SK5TaA2TfbXBhVEiBHwJaHNaA9H8NtKhw9BNa3aRMW1VEPEBQOgUfVo
InjVkKqAgODx+cZROKDZLPKB6LBfsnoZQIYIRANr0767XjPf4/Y3c9XgTVKyfAxYtgTVKVX0EzQm
fpbkkrzT35r5uryixXa4vc1okiyG7Pc8MToFG90OuWaRI+Nbcq81GOpyaZagQI3Ho5z/oSY2zHnk
eEfaQpxoM53XNVDoGpwzgRlOTR5LT9GJF+HYp+1CrFcJuPr+eOKw1NJgjHHB4v9IRwZCZir3M2xe
O+sFBKA8YGUwF5hFSxY7Yg3xIkAeaseMzNlyKRW856NHx+o93wTg5ePgl788zY3pW3lL1e3B4i1L
xVBM9M4WGwMeHvkiw6QyxsGO5yBCadD5xBtXo/ZKJvdMtMi0a6rje+MLXyevXeVkEu5Px5GLlzC6
IW8HSLZt019LBGQVM7FigjL//4TW/01yCMTwMtBeHFBBR2ur9eA00OQmpFAbZ9WQzYviW0KpuEhE
08w+eWB7UDy0ciFnfScWYXiUOfv5D8kOEbi+gvosSRXbSs3rm2dJPb+jOQQCqC8PrDvuW65R7QBc
/u55t/vzaIJFzXi+IPoGRS36qTNYnlfvTs7qe1dHNlbZvm1aGmyOLZ082t7qNPcrUtFY7jr9j29g
56Y/L8OpBCmW4Kw3GjVpCFV1oSjstBmYHwp07eYmG8Fz6JkferrIJyZLs1vT47STYH2qBwilcgyp
HhW/Ox9qvoCEjtdvA5XLTp5UsIudoOQi1XlaUA9ahdPnwfZklWeIPcur5dj8olgtAKzY0ov5jgu9
p8dfarlPjeQeLz+m5grp3nAk1U+jqNmVfSO+tIf2ZTeRflMEh6VHgqMrXKdiK7I8Z6yvXvnv1IFW
uIL/HljCplhZvPReab2j76IgdIlE8oWISWWG5Dhx2KbMNS0bduqLh8cKNsIvItKvkWTaoghRTkR0
GAw09yMTmpD7Ug1wBXKhioDPPHt39EgFCo6cb4NukrI0ETIdwr9Y2H1Trzr/6Volz1D5qBv1OVJ1
8hzAVaH0g87GGEIQIzuKEYz6ZIIVwAXexuEKGRUezaJUa+0kvDu+NyQh4AbwzijAElX8od41NgsQ
vqGJezSMwz26uRLnmpQg+hYxnwY98oeH7HQQb7YtbVvYbG5CSW2Fac1Fp4wq+ItlD2F+7FzGIWpO
JCCl/sylpBS74GzP+PAgUIsT+0THILCEk+MbVEit8y7OFSQokCq7X3LKkcSkMPi5U2+1NKPfKQW6
p6min19rnMsGNwWLDHHZ6BOiAfnA0WKtEM+WsYjzQT71VIgYrs/XtRL6b6Y3OnC2Q0CDTIy+gxXA
YbA4cuM7BD6lgH8C40Lz23rwBV5lnYkVKLBdsIUwJuj1CfsQu1Eo8MTGUH8vwOVm4PWF6qONw8Ma
mCCzvT5nDarJCUZ3fTGHbBKPh/K00XiXB2XDitAiGjl/+xPWOX0r8MBMJaFrAI8cipKHnNCBtlKi
carjCpzlHdORsKRSceyYmcoq3xcMvI26u7ordCHBrYDLdqqffmU2pphvN0wh7b3QtBJ+sBFa3IJe
wsmliJ1ma2FpfHskr/Cv3ZK1Y6EsT6Zm+BHseWhtcXCSbfR4l8fY73I/8EnPU8iduVvbftYkhk/3
w8/Nq7EyExMEgWPV+b1+L2qB5WP6PvfTw3lg5lw8MSVUSWWcTSGgHMMFimht+h7J1+kuE8hwdNf7
DZVb0ipgU+26/bRtu+9BO9AXiRmcJHsRBrq4vDlyd29Dr1EA+HIReeay1arHtMsSaaJ7+V8n0RiC
K3VKSXmSFxWSSBC7qNNWJL2G4zC1TT/eue1X3VsgLcw3yh4cDCYS51fNIwUFQIPdfdLRQ0IR2jQJ
h97RjIA7KUFvTTU6vQUs0FofZOTeUeXwbJTl8BlR/jtb6yrYWvdISO7wPtdXVmu3FPLJJYcFLevN
whGtBEx/iRPH6eF3DFmCpmzJLJp3dsHOakFVt59o86ludaE56ZH/0DY3jO34ffGG5Om43YEa5fcD
kSR23VBfBX81CUu9dcvGH0kbbtcBzMDZnO8tOZgmGwfEwqeem4DTVS4U3u2m6PIZa06H8FPJQyUo
4GF0/s1Hwdr/fNadUKK8mOqX10DBFn27oo+6n/oZaK6HoKsC3+D///QVlIjj0iWF0b1qZZeE44Ok
wlmfrk7A3HIPFAeDnVibhxuZsgR6PclbWwFow/ub4MKGi1KVezcrc6zvijXnMoXHoBEJCQdrWBMW
RkELFCMtzYqKrjxVs0/mCFkq1aetsIPdbDR6e5l1r4QeWopTQnynI4wr+Ip43Q9x5JUKIKp625M4
p6yS3Y0mcvb9aV6jbrIuJT0COC8lUwY3QuzNPjiHe0NkAx+dPgCm5WpyVvLKNXyFvHMqDwEM3cOl
z/aW6YIRfJ7cZRGXLbza29pYKrOYCdhjJ+cuR4XWjb6skgXo6+rGfs8/CPEmhrhyUxSltLT8ehUY
mzh8BrDNUPnRU0JulZndPObG09YGRlk3F8wLI87DHQsSqymy/eCyYV4c5NEZCE8d3YakcgIAApCb
4yb45HlAuCaKnzz9VJ1r6hFwn9Ty3NqCiPebDfIdpymY3T8JqSV7wYqkou9WhYDGPyrqX4ibj7V0
SLyyN5iYZCjMrEi1/4BHORN8TeXfNfmgIlT3WPB3SnaNaslH/J3iqygXkZIGi+oENnADqGHPetY1
/U7VN4OPwvTfuAZkSrMlenLW8TyLFMkMYag/iZpxnmfVZylw+R0bfa7PGwDI/g7IVunAfoKNRGhz
adBGzoJvIc/BX+peLKn0QphJf0g3Ep5J0bK+KBoHdT3+tKg52HIAe3SOchbL9lnsQWRiA5B6cKTn
4X6eSjRpndfXhrhb8wBqW3dmZdjszYF3QIbG3D+LK3Vg4d8GMmPWYIXsi3P7MtwJw6BkkuYNuLFs
niWoxxOSA+IVCA1U6rj1TggBHYcImjB/h5EMbf6dYXglrl7C2yObfCS3qXZjRG4WI6eygSY93IVo
qGqBHoBjPa3XaladwU0T0B0dk6X/zogGdaA5PkVlcm1NCF7PlIim7qAzybgRDY3B9PS2HpijQdAg
Xw/IK/Vkb1Zv8i8AaJ+biex8WXlzf584jZ59TqhXwNzoPlRWXP5ZS2wz35PRzQzO7GSgt9u4fb8y
JPL1CMZX1suVsqT9vWTS2LbfJTh/QJ5M7pcH3JRh7R1XJHQvAUuYpA8ng9dj5q3FdQNyC07SSIgz
z5AW9ZaYWpnLMketS/gHcZK7Gd+EvnDwGTLX3mDB+RI7+BuL/g+6JQewk22mhl6lXePoSMx0nyPo
khjwMam/l49g+u6EGM6RX5lsGMRoRaekEQpXmxM8nyW7sozXimD5yJrXeDO/0gFu7KzhUfX+sfua
+kdqi6i+b2Y3SCpZA9umN5jgpEAHs8mqH3pbwqJUfMF4Cu3KW9AxFBhvddopaKFMICA4Wn13uPOs
9v98CdbCnuqc2GNLbNKjQXCHlJmCToLhO81OHv8GuDcohDHg3OsOyuNh3kpwy9FUXPAVF82o6XhN
MZ4KePVvK6V7nhhWz8k5+FiyRfT3oQX0zlftuo7X5AXWSgUKQubw+sllNd/cctkeBs7sYjbah2m3
rw23y+gd7LBxsuz7DyuIhcaDIvMWRmQngBtUrpnTSBhG4UkJRgBh2AFalwHm3YFXPj6VWBni2DdR
/NEKb1NaaYLRKkIWhhp2kMEUb1Im5yaRmsGiRslUN5Ea6pnWFcGBxcA1K0MIu4aVGPXmSROQaE0M
O3ddeD4mtu+2eUYo0BmxK6LTKW07P8R1tbQPzXMXZsRhSUyEEXkIdTz63O4fuKjVdB1LXymVduKQ
RDJFZSXv++skcILJe4Fi029Y7fSQ4qCsQ7Wl7ouevSPzGDjZrWWwXPBawZIqI3tTEzRCMEyeDi53
kGwAl0HWnAg9xPGchSBW3kRhjqaMPy7LM0SXPmt8nANDPwX8yYzT/HGcdwqOOeGPjFa9VX3Q0wJa
ZQWBUEYfK80b5w/PrxdC/1Hm6I4JPIzU9+He0yMx/DQm6z0ANbs2jupwq4YlV9rbMZYwnSvWLUDP
B6X3OksSilODmzhhWZqpYXfZ6AEV6UuGDVFiqRmkMSV7o7wSI3BdMqaDfaiXumUcKYmBoVJrbPCx
odLiw5/fsX6Bt/tEbyXKCqN5BM5CSdRAzt3PkCYS1tSkXV4taXiIBFy0ZNWjGFzxxB4auLX30mZT
GAElQJsonxFOOmWflo/bAzbroYDLxdBFwqtJBlIYEaIH8djIsDvs1mJeJkIds1srxSL9xRCJw0dP
mfaMPx2HMCNpMoRlTh0Tt+iFC8jqY7IknUiSZ3mTaZT+19S/MtbsjFwCm6fk9+bSmlXA65IWtkN8
/jhkN4sh9xAlZD80ePdF8CoWEQB5ZNEUMlvVhKYOMPLMBOlgxv8PFQWp0UhNhy6IANRI01NMzaAq
lXvJmlUluOAemyeFA5xcx/34hGY9vKG1gmBbXHKDgZ5ALHBSsbMeBe96YA28yTNJELMHf3v4f599
Pwii3pNO1fLoWDap/9PTGCURBUI976kpThEFxUg9JlBu2NdTGRYURAsp8NxRV+MeW8YlC4H0Heug
Czp+b735181rRNMyPIqJ9yjbLpxLJlE+IF+sLk0dqNZb/TSc8yJT0U+NtY1miHDJwU2YUFcpFQVh
e4hI3zVZ1idWQtj5HNUC82gVaOS/nUxZ3/li1YcXWxCYSN3zmkUoPX5Z6G7dWoQmOVjUIBFye7oM
v98ZjIA52evQLJtI0p4r3Ad9Va7yPJqqTgtFwjYU7ichDz1B4dWM55LGn8PhUgIGnFr9vXzkM1ce
rOgMkSXebgQwAT7SEQXUue5lWJwOiQfhcjHz4jxdTWB22qdigCrdtAdf8kIFy/iQ0ZeHdtWFvBew
c4o8wMbmPCY0FFSmAqLS+SZZ4ZUKjlLyfpW1QaUoYn7IWn23Z1MED6UPc2cL9G7Rv4nqlm6R3OIB
IM31cWt0DPebdSPehRigiN1ahC0JfZ5HPZXZTuTmdVaGhboNk5/6HDfqx+2AZO+pU9Yx0Qv3bx3F
KhX8r24Wou99NQh5H4mOdiBP/r3BcsQccv1wC02EA4iQvHjX71o1ngpD6NaZKCif4/MPIASrEaR8
RXlD7vmE1dd9Gafiaxf72FOWGDMVzSUBUQaoqDDVYTF6YRMi1UeUfKAPHAtzdxhDQJeS5WTXVcBY
f9cQ7fJY1vp8tzBkHhgUUMLHpl81VuTI6enIAtRMvnRw4aBBUe/CSQ+7v6xeob9Vi5+RZb6EvxPP
girxS1IbaYpgzdNF6jabHGq6ENgEp9VZpufzaUD7+MhXmkj3WNkZHsgyooGmwUgmo8Rw9D+BVFjM
O+LlwLBCqvvNZbxaFqDPYFkC1IQtN6oepeeKVXdogeh30x2QhkJUguKgSR58iO+aFWLmOS2gTpCf
vC0geGL5j46IGUn/dOs2Hvc4eyzPXc6OXHulvjmvFz7o7ctYpVLcJ2ySZAeTeJhlBEfBQZeawFfB
CoznV717wjas2JiBRV7Im+Fd4NVbiHvCwwXvRkO/AzN/uA11IL6vItXK6QtFpE0IlTezHlEdvWbZ
Ka2X9jeI5+ctIetS5zWRY+LdyMWdzIJIEsXGqebTCFNN8WKKc0PzCSllBvia+mIjXjiCPN5JqfSp
sZyyTBW836PAMGuKLqXnPStzKJocWmCrSSRvON7XiY6PNibMo/6I+IA0B9YgBCcAyjz00PNfgMZ6
x7vbC9rKPwD4G4cynYR5HtBfDjXCATDvydIUcp6r5OoS7yRCaV8Z6zEYmE1y6Zm0GLmNk9HTDKa8
QTtVJq6xyDa8+0f6ohkHq3v3C9X+DBlaMJuSHEnd1MLEI7SODieHYppSoEtZYpYPh7wDPd8WsbHR
HT1/NnYMdgwa1qklqESL75YaKgTlzGw+56asSbkUwwR1XKlOy2m120yUpbQUE10WrbbZfwjlsJl1
hwPYGSqrzpxDea4Vb9Qc7fMeXVkO6/U+96ZQLG5CP/OZI57tDJCbWNS3VmJhN3LGRUPC1gjoXsQN
7WW9WwJnwaZrjkd9BKmVp2cAvK20ZwBrV/S+J+Ibl8u7RhSo3fmTZ0vAsn4sCz1cqeyKVYb9GIm2
a7WIgBHO5zOC8h8v5BmhBDSjHpdXS0Lcj3ciMvABwNcHC1hWck5QKAeEL+e/N6g+8S2E7z96svcN
v9+bEWycNqNZzxvbz1yj+oEU1KhyFuhxA+1BxcHUKrCGFYxm2rK55wvPpEAFhxe71HBwXlNuWM9q
zvhIS93fObVP/HJci2bNGho0AVL3vaMRK7t4Q58662bFx6Fl99UbOVs9CnYs0bgELDlDvcmMIdPp
qgzkOFqYOTO7UmyJRLvfmnxyPEaasgLn2BYqAayCD0fkpBDzV7c3cp2skIrh0wq4tWmcY3gkdKjr
D9dMIuZYQ9RBaeJSNKzibbm0teQvtARKa6ABf0M7BpD4rZZyRkIULZTjo1Wimm66k5uwUseGghiL
L166pSjpjMz5/KXyTz3t9aOXw/kTzxl3Xr/51VZHjnwQk7ShdCZZH36lZwZrHLK2xqdVv7bby1c2
ScKkgeRjlozlhNAYVvH2kOtMiQVr/+MAeXhlien+/VAGI///8s5xLOH9qV/GfsRZ1y1UYa7xs2v8
6/elYYdKKzHl1tAc2JwuUDuqJaQoKvnekuPe8VotE3/fgCZL6iTJO39pXxEuLJR7q0UzptPk1+tT
SR25Qq3Tt9G5MhETDnE/mkYiO4gSJYNCSJTvVQGHVDsOuwxpdG5bLJRb0MwT3Gd6DZDB5FdlX+BI
PLbssM8kMiAOXLfrzvKnX0zV1V+Iqni2MTZMh4zHux0ChpC4Hwmmc/f8z5CciWBQHcAY+mqTPKGR
TQYAmOK5WruNllW7ctFiJNTT834O6D9wFBxqogp5eA/EqaiKNMMuRPOqxKozjSoEXsTaSbWSUULB
NXCGfS5xSJZH37q0s6OJ0WrGD9t3XAfrL/oug7dvWvhDNNajDAXQXLfS2quGPDwugoqyhLAZOcl2
CCEyPmC2XzTgl1JHvOyvJ2EpOY3qCiem7bLh49rd1jLAx3ElNpjJJremjmZkLnhDc36KOA86GUJ2
3UbwrMGaoPkyzkbwBqbrebywTot9j9Nzls1Zr7/9AvhFWpvm3RYH6w61BS4mDDJhYqTMAXIxrAPZ
PhWvJcBCiC5V/defpAuF+kS2sGrmj7dAWK4NSk7kdvA54pAdmr7GEDWs1YlwMBX7/N0FS0XxZNxF
9tjBOKgPm8auQQ/6LihWWoiM5H1h8Pqly4owxRFJ6h0J2UwSHFvt+AptoOTxH2eQUgUBE4Jew3Tv
b4I2Rmg2milQlMX0ittvZvJp0R59NAfq9LvpqPGjQta0CsP0cAnZyjWvG8OQGtw2nD1H6680cvmK
lFKCikr1h670T47J36V6N9aCRrax+1sVSOEmpo+/ncd19qSqrBZ80sFisSFjSExLkPyD42ZQGyG/
Z0riQAHbb/67W13M36qdxQz4Puy6UtisAc7mmNg372oLyU89SuSwEHVwknvTpbWWfl0WVmQ7LYC7
0sOUVWo+xXpKM0+7vu4wzNF/Svbz0uN6ygfJdTc2g5dCwPGYngniaqR2k7Awuy80X9AoHuE09//9
pFcuLQbLWeSTulGnR7CqOjWwoy3UInXy3MjX2Z9yEARGOYuobWEdJvBqX6huv9Eg5x/ex3Djhm9/
9ZkvT6ivl2vlxuhZq2EFQvfdziohSQCnaI85ef/GibXXAHPV7ax92p1wLM5Pof9y+oOzy3NLW1ba
t3O8tJWae307jeO9yAAjIIW7rtrRdJzM/nX3CiMGg8KGPR/LunNFunhiTYYgxCsCh9Kx8NVNFhIX
EDu3EJZULAUkdfhmjpuUyeDTw0QPNWYTuI8teCrPffKF+aXotLGozeQkuf6N5nFtEuh0cpQBruv/
rVQp5p+6mXRZGApytHEssvJlEvX+SUy9GE2hXCCa4Bp9ABqnF10UBLy82OXtuiVgHfRkyHxhrYHp
GHWNEXXSatuo3MYVyWo4ilhV6VJIDI9x62WAfEhSs00QW9Zg14za5n7ZV6lj5DCJPJAvgL1mFWW8
MBA6o86HoBUzj1NDY52wKVADE8hjMqT+Co9KP6T6LZdEG/Ay05gs/oojAT/356wmgrXt0d2vcOEk
2kUMe7oDjLTXxuon5Uvs2aXtyOjx7rhCng6KZM8G/+4EfRjhxUcVU3+aj6/et9yWW9miIGfw7CkF
C3QUVt52IFfdtJ/tvWT3Ng3AVgFxsV15GQxGPaNwH1Dq+AuwAqKkt98BB/nFLkgn5dFPs+VBfX3n
6EzYmMUeyBzxpu3zdpPjEVfksQzDdWH/T8RIeSJcHugNGQjfaTtcb/Z6QJkknOrF2QUAXwGbeZXB
4HgIbc5n8NOmaS4e1cCpjUHRwTE2ZXZI4YLdnOgQ0cSFhrtmL4RpQ9UYVz62KTaQrmqXl/gutq2q
5ysGI/Pr10L3rsPAv/TKP4diTYjInao06YCBl9zQujRZxeHFIIodRAPjuCh73Ku8X1pUkrS2H379
hdl6lisePS4iGPrR7X+ItAtBalcmxfzLBgRvV+U2PDGGVRndjQLK82pNDIp61ikSwms8yS6CDaq5
AJtpYmph0rFawkMQDi9dZJrsDko93HyiuJpht839ybmktrvb0VWTMkjfyTdpmtyKvQiA4Sy9/qNY
P/nBBo4KR2oCNpJY+xVX7eB/EzqsxqRfDFrKm+yjM6iMl90kXLYhIxb5CVewviAxXBlJNiPCzPUD
g8Fm8N8zSLLJBG5iXnElBkKfw6WSl1DoL88E/caAIEIcYB45hfkmMjBfOLSszOMBwMzmQGBUjI+v
IL0W3yDf7FNF+v8sr0Q+m/aMWAmG0zbIbfJCNj6midq2JNKIHxBUCTz0rGRdCNRlR9XBrM9D7K5r
V/UTNltuLtI/CnJyO4XobP8V41D+eMurwz5oojjhGglzAYrqGYjIHjU7ad0IwuL76qZIOwh+909h
4k7PR+2HW8xQi0/DKOp1mGJwwKlSfNWvGDIJ9YtwSQ2LzhCkie+7EqeJ+fuowTmIoB2lajKf2knU
gy7F2A7zM/+dhYJ+2xQjnLeBQJZWtZu9AxUIyZlK9btQYEKTihmJXw1pK3uL9yogvJ907Agloxpv
zyB5l3mm9FqFine8iFF2on+VALYMx8pHExqCToQaZXYcvLcvhQ3elpVLLoLl+trKNCAK55FS2gEd
G5xWtVMtAu++kzXs/HTs6OulRE/FLnTIdxTNUdSo3E5COr9psVkNisI4bE7paaaEQrGP3ZHrTD1v
PHyvulP2tqEorRdEfC/G4bNrrM5yJDNFtWPp1/CquI2NhW7Akn0yZN/e9Biq95UVnOyeeSMe4f+O
Fwy67OqkJyu5b7GvTRCxU8dYVjwWFyT/5jOsGVfChJJLaWupz8Z42kYE77nB4AOUQxX4O0bh0e7s
w/wGzaRs7aBs4EID0ynxPsW2d+Q2GErFHfK3CJbGhM6D9+MbRt3KgJIcLOe7YDpYPWMKGS4XvHj/
nmhGNYxMH6R3Ka4VxmtPllKgw6gUt6Wu6ld7rbm5niLANlBclvfeUrbc5G7S+5FQRY/9zcbhFwpF
zDpQ8/6OobvxrBOSATbrUUsVIflZxfI7W/LP/JgiSjuDNUOVApYB4SRB5P5oOSzn02ty/7cBWvwF
hdk/lN8rKZBbgD5U/RAjdQu+jGJ+OFdVSL+nnGSut7AdTU0d1c7rI6PBfhFYztpOak/0SIhVWhA9
gD3CpBmNEn4IPuzmjJI2t+dncnyI8GQO6/awkGvqnZbuu1MKqjb9EsCgCojbNA4wQLlj/jNMm84O
L750dpXtXGXUYv/OyiBo0OuE2Sy4y1ZcBEim3zLZUvXK3M0ERYDFkATspbe9GShuD0azCdp9Mswr
rWJ570AnEjXFJtdP98XCU+oxI7sLnR1wWm+572pE4EYzg66pZKa3iKBDxFATnM66RwuROJeSIrSA
1xy/D85+0uyWReiGrsUO9XT8bSebGQ/Nm6/sNSkgO/98OOTL77NtwQvcxB+qFIYLh5uMfwIa2/k+
y5Fx1Yirzecdf7NepXmUGYdXkOFW9xDWdv/bjWqpy+eb53FHclqRlq8mJF4yGLIayAFb7gSNMNE+
WEiZYpXosTc8vhSwIuJTg9rG5z43Rtl8yT7g/gnI9y8TKXr9a/Q4b/f0UgNiqWx0wsKrnGnQv8aU
ke3Tt4a9gR8AAumPLxHZSPXSz1KCKPcDnHAwIVBGQJejbFwoPl97jqVLJ/KomtRN7K0mZR0nZDfN
8BJg6HW/UboaUTCXdjiwewMU4VY02F5n24Kt0TFnARmlIrUTLkYDVDOaKy/yTzRkeboJycj3txAO
jgs+Vn/NUCHP+MGBZiUIbDEkvtmIXjs7JEJg09mRifN2e0Hk7ou4TAX+gwSldzXTfNuEtTnyqTh+
TzmDooH57XHvctqvde4P5FeVo4hvZ/+eLLmCFNQ2Cwt164hSsAgnu5ZUfNT9XYBXq6/6NwPNtEZ4
IXduvioihhWujcYSOJc+NUN9Meb2NEV/Oku0mtMSdhgPkCR7StSWijKXwGGMEZERqPPCUxVFjsqI
Bu+KlG37BV0/q0UaQ2dQRKqf9tPHBfNH02Klg6FfT00vXbL15cev4cyDALMQhLxScNyvQUE3032+
3CGA/wsY+CfX0vHFMxLAchA+L41iXYBo46l6o72bL3Dwkhp7xmRfzFBqByrqWDrfRnjDGrQ9MwHx
yC4aUi4dgQyM9ijALd5BdeeyYKC442jvibmQAsuXqRgjr0kWpAauxxCRbN8kAhVpWgugDf/U5YWL
g63ZtCN6eBJitDQJnTvCkfa7yAX5hD3nHfjdvWv71t3QpjWYfaL1sixFBbrfds1bOl+jQZxvqV/n
MZR9ORnlrg2TEjOjkiPT1tD1HMgAlEm0SM4LVnKPsH6INtOvt8pXyx0vadmMP7Wn71ANmsCmK5Gq
vPsve//pFiZak0VEZ4FNfYb4XOEFGE0NXsrcxvp1BdKU3O+5GHffEchqk0qEIHWkOCXkkEkbdbwA
zhLwOcpKLbdfM3BDlPbOB6jKjZLglaa3fDNksFf3Dy3lzMUds5qxxghJltOzEFnTspnqWHEbz1Uv
RzIfbz5s9qT6XaMAHn8udxttZU79pFTl9RRNSEWBNAvGBtgAGpE3tsFmHD/mvyQ1zLHmcPxkBIIl
wQPgmUa9sMl4mvrAPLxWGRirY9aPofMSFGmabBOlAH9FekGbRT27YBR4z+ablyEAEU6Aueqh+8ea
uN14EyPbPJXUi6ObZPRRLe+5N0TYwbw+KR73xVm1JerjFPz0fvaZ2o6OktqruTk9t5QhYJn2xM1z
s6HK2S/z+Z3zTp+g4mRJyi1clh/XbzIHYoN3PvDoFqW6fPMJqJMgy1CIp0MULh4Ykz4PzTAXzEeV
et4OJkgS2p/GfKueXamEZalzCESsoFb7LjzL9kmcDPlRgzKlbth+4q9wwQ6IHkoSKXNaIxp+DX1H
nJ/eE17l4966QEJlXRnd/A2NSoA8vZ1npSXKv6LQ4/hsedfOyax02LXnLiVJQhoeezZb/ZkoKOtV
009OAccfHY37q39NkpQZ22ssb+q9G6trWCVM4ghqwJNNvYAEHGTp8bq+hAYhd5JYQY5qHUpq8Dp8
8gzpYc/+6ADXuozqPCDIgBMXuEUQ5rcCHyjE0NGh4yH3t+CBB9a++ZyXowRmogxQbnChIFwvCWt6
RX93oPdVfQwny3ij8XY8+lxL8gH4dtea5kXLxTfsHXazUOQ8SC2L1yiHq8yNCC7h5DaDWLTHBweH
oYaysF7ciI5AjF7FbnbRreBj/VXEVezhmiriGZGHcj74OsMiRh/EfwVH2g4uKL3Ejtkf0jLkYIRN
ZsOgRHszpFm71nisBJ3ci0qNumhQ9pWEFZ8mKnDhvCGcCyR6esEobFcA5PTKTlZDAeypa2OC3SPC
0juNZ2S9N5OPytq50fv1bbHiZhldbfkrK+62d/ofs7tjYkQkrWRi5qCzaan6/eOKQ4ZTmIO6o9Z+
byM76fJvirwXR7dqtQUW+3uBMRKuG4KgqJ/3Uu/FtK/7uF0pamubLa+47cLPGptOcMbJkM0PGD68
rlS2jRlj6MO/ghQ8T0NqfAJXCuGfj9w5hTuLuLZC+gZ5QrUwXzm/6uGjOwX42OWnpui+1SHXKeQt
mwPdmaezzHyvNRD0JPgZL1WNdo528kaAUEjoOBtGhLy6mE8EjLakTA20szkQVPY2ZV3c8pw7uPnY
94QrjH5H8ZHQ/tD8NLmV9t/X0+GqcM5W+WggwE2BcDKmmiuScGxvY0WwLPxiMoijK5gVJBcheu7b
Bco/8tmFU+gxTe/yw4kJ3iLfHiOHo8Dr0+u8cDlq3hSIqVuYNAF4rXKALnVZ9GUTlzF+UDeUovj+
gTACWpFqJyRZjbkVdHWgW6ur2nA4AZT+S5OB3ZGVVl7kLR31GJ+8oS5XKcrJXzNhlxaIcJwDs5YA
r1JJVm7unC+Jl/vrlx3dK1oZdN79iKRyJUl6AbevD0E3+6f7shdlmNH3P9XMhuyuaaDLlKtX/Y63
fxs8bp8yNZksnm8JMtuqhzzsZJeXRvAeIvx10plD23KRfWZU9iCdpzI0NS+1YiCicvhdk3nhKjkF
zsn59SnV1iMgJsINlXfWKnQLmKDsHmn7zJisKMzMB92G5JVZjIFuw1pse+sYS681CWrnsI6Be3ZG
ybOmNDTtgBEe9y8jdshUSavve5L42cEOsOJ+xeTntu1gWD3mDdxbu+LbBc2ZVRfA4woVHFpk+NoV
6fqU5FiXlwcEZWMuQOIl2SRnoU4ylOvElYZoGDe0V9mL8P0KTF3f16wmP5ctNcRlqErJcjNfVXz2
9wypiL/Xu9rgza0XP+jQzi6jlNUhWy3qYJ8pSt/VYswNiB87WtkF/iLEy2Hmtv0QuBeIQw25+8y5
idIs9GH8IH3yKRSXDNdqkA/pNxNM4BSNvWMTYrZTzSUiyTHMF4EOUD41ukgXut7rZHcXDrXFVHfV
XIbqpypgS2ctf6pu5U5jyV7dUk0tG6JIAKps4WmnM4FLm7XO18fEjynUtK9Wtr0g3uotCZgBVENx
Kg1Z8mSud/EgfpWE4tWXwfOmOoBZJIVtu4+hL5sn9Vap67JtbZwyj+9/LcINv+hf0/B0yI/vZK2N
OrDBCZy1vvms/oY8ZNf96y4zZen3rZNTk7BtIiHLOu8Gk6V3u6PaZWQqgVQtL4PkPy2uscJN1fZB
2vKfKFqi8a7Rv0yCKRsFB+sd62CPHxLldbzxMf1PofdyeZSOS5lol4+4eI39SBfu/L5l4BP9QuN/
cQJJlL4TpDTlBZxXhHgKLEYLyjM3ue+4O9t8NF4udQgW1MuAUspxpoauJh2bMGKXIaG52ShdxcRU
ZWOYY6LAmXpwSbyPMn3PFSzN1rKDzuTkrgxrvD6MCmdPUtmqx8uJCxg3lNOCw0BViJ29j/EgGnoB
g/r4MHurQLh1Ekjpp8CHcpE6o1aYV1XBUp5d2aLcWgthEOIzbR4/EElthHe0GVmbUM3Eqo+51ujd
zBZPZjG0x1vzabaAxMvs54azwIJyW1Ypov7KCjm5YS7Ie4UdfkX+BMlXE2/2LhSIS/YfCtM84qSB
go4ifdhr2eabNa0Fx3jnL9hNyJsImoOLxFZQuLeHe7uy5HV+HLdctQLbr4MfGIy2ZEE3KXl4rs2f
ie6BxrOBn6goymc0n4jnjsr+q/bjTHTvestFMZRa9J12J0PNhMO4tUSECdrHpn1p9Z9ANz/ckMC5
qOr1gSp36hsTQxzavt8M1fGeHxjiHfouZhMo1oRswNbuBwWfiI5o8yCt3jVH23BEAprMZH74w+uM
ruOqeIqwIdqWHm1/yMD0bjG6eyZaINGzSoil/wv5V/adt7ZZDL3Ml7h124LYnUHnEIpPFXP81z0v
l4+SHmt4EFmQXYPhrpq2jp+fn/XRlx1IiGzy3sIIsmxJ1onoa8vklVZe2nMZgpmvrOOPbvCMfsrz
QPpT1TGCFg1Ym0M/feBVaoS4+73F2rjEFBBuKINtU+Gx0dFjtwTDe4yr/0/NYdM2Qwn9CMqOcXUN
UYN88AcGWXhSzWQbYbVDoT4CiImRzwoksAOWPPzOIwQ94pbkrEUDo71hSiq0vKIdeaUHvPsm4SC9
KjClZymJwcyNIiaIFPmNXQl8EuZNZ89Y7nAVYKAqshPCRlWeB0kzxlM/rJT+54Uqv7s73bdlyazj
BJteBuApxo1zb7OJPa4zl2cGSE6HctlssyxXKPP0rFmup27WkS5710r81NDXngtR/+6NFL8M99h7
My14tJ6TaWkX1aJFTFSZK8zLODMOggV9bHjE7MjpHiaaqOVwK39gOGLywz4d0O4nGDqi8mcrUIpx
yB3MIK+UkLFWNN5o1QbQxCUqUkNyCNzQFzg0BsZSoluW9rZyyRiMmRCkv94RMFPtJl6UF6ABnVvx
nUtgWFf7CsEzGTzjqwWBEnimV71riIvuQyZ4AqIsUjQwQPyYPFQh9UNcOEgYlhkjaNXYfTMehbFK
YpPbjl2BAsqc0bOOTu6LdiRWzHP5CIA9DRXIyVk16BLGBy6K25VIGVV5l3j2vmY4CDdmghOLHbR9
pOPVlARKkufjdc015gR/xPZBGkky8kCbrObHuMMV0/0g0LVSD0xztxrAtiIkkvsG+5+vdQDyh4ba
2/99aU+JfPtaj0gMvDDoAL+9SS4UvyqrLeqovwNK4j/0p8dpSsA4JTscWHe1PRK+4R0p043BD4mM
qf/3LMEE60eQOpDOQvssvePFRP6IPL4KeAcBfvPVxeZv3NyArMmJ7RL0u4WOL42a5Kq1mVcBc/Bx
uo2cgHV2MKn78mlf3tMxZcWNVGw8yeoC+nQDe3XUT1KzxMCTO4kKi+QxpHbFgmYTlY4Nd+jxmdQR
ntApLik27GPgi+QZFxvfl6SCJnwV/JkbS/nK6MSy3lbLrdsDSEjpzgcvw4tOM6ZRZZqwfmvSmWq1
u2/EnumZsExfo8xof4R2NhPH56MTEzHydUfGqxSx9TIrYOMEUymd4rSubSfnGS1nG+MXPcQXm0yM
Uq2hJXFVBf0f5nmZmGW4qc0kxLaA/PaElWvIc0aGcIDezME2G+enUqYj9a1GUErZ6WdG5OjuJ5xD
9cjrMZhUj+pn2YWU+toWsMK0idiCuJiurKhbBlcX7gsi3urR6RbSPigapRqMhqYALbBNipbm8rol
Lql6oL9JuNvMBWbNIvUPuPaUP0VUVPrKiRmMI7Ag2D9hL2yOGdK678FScvS8Z4NTPRKVloIXpBkQ
XL2jio+CkhU8DVn53rD+RLuQQFYOtyKjKpTkBrkKqb/fSeTAFvnJz0ExdaCEyhKoSEN0Hp7g2hc3
DZGnuRdnlZt1IUz/27IRm75bFNoywky6I/8VC8gQVD3iCgBKsLQiksXrGPw7Yq85R1zuQbi+ewkU
5VXjnul/YSjQpUk2NU79GVyepmS7adCjruKdyuA161IdprDYU0MN9tTeMs1vvAQUQtTMHOEzZKds
h5yybsKBgfqnWcrYSgP5G6kQaiSkLBGlzbVgo+eZl/fAWnWjxqk9UM+CKJP3zF56/ZoGtayWF1ll
iBYTXv42NVdfFs+K2REZ3rnVUPE+axxUBjSPi+B/1ETzZNeZSVDDuulpXGhsD0uGr8DSn9hHafm6
iUDpUNgiBbSwWxk3frNxbETk+vJWeaCNmQXeicgZCwER3Pr8npGfG/4s5UvXbpTgo42BP5F7GJ1X
FKPJS+hTUun083uw3dc5nvs+kqmXXifC4+ZsA75O9/nANMzZsrJvC7o6M081Ib67pFvmi2QxLYg4
YVXKmB8D0xlocR9AmzhAbRUuZQwohgoivvyleIOt6WlOfgZzkBFL4zagJyFDqeHePGMVadgPM/Lr
709QbdpK25rzyv4V2V0OjYqD1DIj+9uyU4N+K3qx2j5sCF5mG9+rO4fRxpqsPFcwa6k+M+Xu8rP+
W+Q5gB9iw05n4MF0hQaCQR2kbAay+12ypNi+A/l3GjkYn6GbvT1Bnj771lxDb81A6stYAllHCLUk
9xhlSqy7kDJGU1EWKi2JsZF9j7qBWCG+mgoum4X6/A1uSw1JgR6w+MkPBvhQCn1iVbYW7UQnhMh4
yzzrwa8Xi+iKbjJVfrXUkJUpYHGdbedJdqNvGYNRGec/Xh3BNPx6JbLc1W/+LFmMbUjuASlXGA5r
PrAkPkZHayl8Nv5JxHBWxrUmiqeKCE3rPRGnorg1Tkcw5ET8aUI1rOBbCTMPcfCpgEh2b90OcUBL
4oV760gccU/Srkrlkmy35Ggx84N8O6EtbqAAOMBfATl52kRxpgBeqzkKuOXCr2IZAtPRzMfgNLdP
qhEgEdfELOthA8GD8g6A9Fx4VzhcOeAHYIlHiox5W583wKERpIYZ6isvGFh0ttE1lwMP5JHjO0k7
0pO1SofpZqsrqi+OkQpp268/l5hhAWIfvSYF3DuFLmVsfL4a1wi/g1zw/qAtPZ0ux5kPvqF47XHs
Vj8UGB1r5fo0e6Cxq+1GfIlwXSdlHFXorGB8reOZ0rKCR/MNaNGwtzygKwJ1wbKnc3+YDIvBa37s
3qxJjf4Fm6rjIEZPw0WqvQIlygihPte5pkF6isoYqTxPCw3slQZg9GzPuQxH4nUrdtb6rgWr4GgA
U+bn/6g/fWH9A7yxyQcd4ACNYYId6hSgbTKsGLta1lGU64LHqd6ZILHBh6YLBliStFPq3T7CxLGR
lMfh4FIi8TdxSMWemReiDqMImv9S1SNh4iU0GhshYTNWr8xCTJn+6olKkXUNsFRp2AjfxzD8EZPG
ZMU4qrz96VEQ7ecSmS86Ws3BAuLop/34ipQvKL6o6zEM9UpM8QXP96Kbf86HzjPiqfM1bbw/NUTv
1UXBsvfdnSprqhOOblyf0ya9kPh7u+geKrFR6aI6S4o+LwM7uPSTQZCYltQBbDWKL5ghy6qO7EM0
GgqsZ7AcLUecCvihc/As4AXgvKXY5O1xytre1Q9M4ajDG72YOU4x1OFleHf555jmO0CSy4mlBXiR
/uorWTFdVFnIVnzejfPnc1jcMC9piYfRFEhE8QliBY3Kziw8jB4MeZ2pCAwb6zMsR75UCEHYorKc
J5sohJrzW62a89zUYfZlW+AffqXBLwwfiPCgDLJKiq9CU3i2sY7Pva54Xi+4t6dfUt/FaOpPqhFG
i2vxpoHt/u/IVxXVMVzIhhbQ/AfLwA/SFZfwiBjVUHkrmjD6IgOtn2vpsCNFuQQtYAhVjSTQo61X
hS+GNjeHKoR0WJslZIzbEcYyoExheUppt/G78Vp6HjWzUIktAdtzBXLi7iILxN3T5WUdG7nuNeae
Bzy/Q5TO8ujSZxWXgiIt5o+KRe0ig8xLQ7HXhwxdOr5PGQNukFkJX0OZiUqzsJQP4Pfnk6fiSKjD
rwiElCp6J0934juNRtjJU+IsIFT4XiRYnsSIezDhJ/sSvn4XkX2Yh6YsIOFXMIEIjuLyNsfpRSDD
NGBXRoo02ydE6VLgKxAVUM7Y1ulnmCIsrHA4RH0lCcCRajMvJxYUOAPt8P/NQk+gy0UkjVMXqKxt
OjONdopffle0oPkYatp7u4xrX17nRbqp3vAX0iTdpi2jvTGSHm3DqbucW2rxMGyYaSCM+RJBiM8y
b/XFeba6EBVwmhHvc5XCGH/L+g2lsbxY3euJrfrGGYFtmroVOyR0vLpfgjwD7YjnspzsHqnuxbxt
/sQCJgUp2Cch0YocKQ2yKKShWnON1k27Og7k8z7gtLL54uMNvY8+dVw5P1nJFC55RwfV7cofUlDB
QmQUE4QdYerXcgEHahyY2BwhXN9nd2Ow4J8Vf72exiL0UrGgl7nGi61uuvEKHreta+xAS3nxHW1e
7NiqG2ezwG6bFCgcNSbL6dgUb8Grdws2dBFDTJyIwdsGawz39O9l6rj6uarKA8HBFwDryMtAoWf8
bj+6j4i8qwp1+kO/oCU2PTuVe9VlRnsmBo4tSvIfxnqC5TwjdyXxq1KSsgPX8h1ygLbP9bGqhqjJ
dmORHgpTh3/t3w4lJGqaTosvoWTLQreMJCSsX2CjiafmV4zWoiI01iuRnwCY8k3m2ySdooaTVxqu
di1KXyrnLZZuNh/NTuNEWxf539+Vt7YRD2LAEd79f3pUwZYfRZLxI7FZU9mLTiYMPOiF6+iGUbwu
cKm5eDIwODOoF98bVDq6bAWlUiN33CAUZxobwSyn0UUxFm3NpGOPwKnFa5zDfHlZ6CEmTMkF2E97
+F1JTQiXaG8qfS8COxzap2hJLdaCmqwtq1iPcYa1e6tJVFeFApbyg/yuN5/9UW1l90qddZltgKnf
1/94vr+eMcatbCmAzsCsAUCBraK1zGYt+t4JBn6+56jZ/AKpjQ0rOb7vsUZFewNWVnx90pSbur6c
3PUVaXZ1/t2LhKBkrTL49oMYDjJ7Y560pMvAv3yagzX3GKAftlTeiQLC2+JTJlIy4N8OAlbSrSoN
oye7xeJSUNVuGarqxgCLQYSMAuUGT9BSbWDucb9yDprllW79GZiksAbe6YDQXjhhcf1nyRuILJaC
IfoKIH/XYn5BGL0/R/dnnuOPwIH5NeszazB/JeI7J07Te7PHSSaqaGD1F3g+Mgizziq8S4GxjGNx
h4Xl1lGfMmfcASCDMEAcWwx2dyvTEQtwDRR0SgEaalH+7l4pg6E4NkS+Qae5+9B3muTF65Xsm/a6
BQVRdOysMyOmBP09wE9yoS/5vc71oHuR1Q4gyt+PM7o2ITyuZxpnmb05pVzuovyOOK1/4tsa5XH7
iNmFxoSc+l1m+XP+mOfJxyi93mBWDQCVBsLtwxy0kO79oJ2gcqNqYFBLuQP7J2qRC9XrQDYGe6JC
H+kTC9KmAYaNjQioIbFFRHWyadhTuvqJ9VWJghPtyMkI3DjpTVZQn08NQxSPebGigT5WY7KoOybw
7h2lR7rU3C3W96o8nASx70IxB/jVx+sekrecI3ZVHvSArtm5EHbUsTOfftmrsGZGEKBwrdf/+Se7
4ybItGsvbVQ4v3tY85/6yf81l8mcNTqqnc8NMixqj67kc+2Wv4Ere24kPSFxs6BMlqG4VhXkKuj5
28ZDeKOerO6ZUn6jladXi6eaSCKrlWJ18mnxkgX19ZuC9jd1LR0NEaDP7oGONff/LxL/ZlxpUb87
kpSCm04UZUpFkUvJwL5AGB541CxWjwkz+Cxfl6YSEAqnRx1MpuwLYF7IeiXLJ/PAzr76VzFEsGkC
slJKGSRD7ox5E/ZEHVMuiN7ce9/ndzauBYl8QNQ1nM4FBA8tN+0ThQ/DfBnS9dT68f+DlLA+zxku
kRNQqNJ4SnwGuvIOa88HiCGpRcMtjXgRrOnVqUQi9t7wasIEN0pR/4c98rMDW3U9yP5wQ8R8RwXW
G7zBlPLuyVzdZmtZDN6RblRcssw7QUO6L7IhFiJEIQVjWkGnl+cmlon7gt6YIq0sUufxb3PtN6TL
s0ujDDjEEVLcMXMc8JhrRUuHTjE2dwzpO+iNCYy2A0a0yG2bgPrdBvR5Miz6EYyzTT4QoM0wU566
3o4JZFbCibatKnmE/Nv/e9fqzob1Il0Bdh7AKKlnT9fMHaEnQGuD+elOE11WRTHvyrvOSsfBmLdE
JWHiUh/xZXWrKI2Qg6jPH7KDhv09tck3ykfGX2NJCnGc0LvhZEfmPK9CFlKQ9uQf9kex+UpW94/2
XJTwD7e0kQYO/EpRr89Fx/aWg63mWlSQZXem8SwYdvaBriEJBroaxidM1OhaOaKtuy/fTqPlw3sl
OLAB+ASuExrMKhwZTswybD/9gTqw1kAR4jwWllHUWy0bIVKmvCNnVmLVPwCt4gLRa4W76lfT6XUX
mjfSJw+wkJc4WhPtdkQKWvH3eWi9uls9A1fIKvw8qPZ49zbY1LsKYnqc29sISLmfzD7Xty2Cu3So
Sf1u+sKm4yFBHQPJ16233FQR4+t10qHR0a338zD/zqZwW3ldH8JdBaRxdAsD5PiIe80uOVUn3/Vb
g+nNy1S1+fR3XyyZEWLvGwWhg9Iyd3Gnynq2EoY4tNYBd0leZynpWKSIwyb9UwimYWf00CqOaTCZ
RMVCgE/j6g9GEKOYgF65LzhPD3UnCg1ykyi8x+yZu39iSI81db9hay7H5P/Fuvg4ZuOkVc2IraQf
2hhfdm+gPpJ3oOwItUC9tcsYnlhbZqCAbVeSRahW4q++rMqVjO0Ulwn4nu2yCwGaU+yp40q3dZ0M
nxbpskHnar1agKl+HQrlZSRo5PeBkQVwL9r/X7IvR4aLf/5yAcrBGjIcURYiizlelD+4PO7eYsiP
7+PU5sJkBHKpwR1oPHP5jIii9AGnckXKG64huiQm82vPXep1oUuuVVSXgB6VVp25nF1YgsNh7z2H
IHNaYW8HxPaqFDud5jYzr/WqR/nGnrdKv/fG9FRar+bkauSu9Ptt/mC/eJc71WzJGtiS/Cd+n3Yu
AEqXdzfxAlY+EfPg2MDyOs/nEqxYOXGReAB3oiBYRswSvDI289/oa/lrQgyqEqoYWW1zpYgia+Xl
jQrA+Y7Zww3iy0VubBUJQ0sDKWDgSavGEdvwsrJUT11nYCsssEnK04Xf6V5Mw3K+T0LsVrCqgSOu
BicTWvcZZwGlEaWL12UtlrEl6u/T3w6PACAMeCDsmHP52tTtPMkLdxfejVqdKwDVHfr0//anrdT4
gW8Ozg4ax8XhqhKXEvIJkLgoCNGdBjhwdYW72r/GFUb+IciZXO9S/iaKnz4Q/cMB+4WXv5m7NyOR
Zu56a+zuhXs8hgF2g7dA7Q84vuZMVxjhUqbWpIGuN0K4VDrgl5JFnSi7wRIEc9tIo8m6r6wXTcNV
8bZWv/GXNGbl8VKptJbWL+09mIP24bln9VxFHFI/XPeqKv2gd0rI+HYLlkKWZ7tVx5j1aKrrx1if
tHGanMu4JK/ceVJVNC0ptLMIPE6Yt5AbdS6dEv9DmJJH4bCgBmfiRqHW4QDhF4swG9iD0NK7Knh/
XwJX8mHSF9EW2PhF/6kbLOD+/jsCbYA3CF6TzzHAiB4XyxdYDhG7S1nC0kMVgWxCbiLeTzYduowy
IPlWWwJCH4xDU3VR1Z6NyADAa1+tEbpSyqsUOdZ5xS7cRHaddeU3XyvvzDQZGiIEeWRFRTATMg30
3lwq+1rsrY7afMXXrVRtduC/0YWxEn+BHyDAxBvb4q3Krs9ZravnoChKa699YjEjo22jPOSaNlgq
eK3AfoGRzxH7/j+1zZ8CnF/14sIxIhJ0VwR4GejQrbszMW21oRiMGf7gvkH6ZsRUpK47mmdAx/8x
fxTjUtsL37Xbtfiq+XN2FeyLqfc/tuyww9GNkvIzMh1b7B1zq4pjTqhrRo9NorIyj5D1evghS6yx
14y05antvbYQsqE5vlpqtPio1l/5oeGWuzAKizmTwztkQJ2IXsGNQKHf30wLeXcybvjArgum/IHx
2qlIlzF7UNRujkodoxxwQY5UdhcsDuzqLNXsNCMURgY5HXA/SC2A/g8L0nd3Vb6L7cZoh8kUrLn+
bQIH9fz8rrTxJ2L/CygPpjEvBtJwYKPaE1IhhKzqK299OtiOs3be480pd8Qg7aWUl8lQKv7bjyKS
eE1y82ZZ8inrotIE18NFHbvsCiOXkHFks/Zr/gMygK0x1MQx0hs+cwjXUgTMH70YS7YYI/KnQAZn
/vPAdzS7uTTEV5+CTeWgjpLZQwD1SFkRTGu95t18jOmABQVHNXvCtfQK/PO46+7HiabIxVGqLXKF
76kAOY55BFsAFVtLJCSLJKUqYsdvAq14mVQX/r4qCR0DXAU1XEtS3eC1hxOpBAVSiWChcbJ68WRi
q/Ppg1RQi7THvl5viep0a+aGsL5lf6lPcZzCU/sK60FopmN50GVABcvPbnd1YPjZlVlIDe3Gx231
OrNYFK8IbQKS3MQQUzZ5N1j5ACX5oW9aKMrOxdIAqgFhmfP/yzEW6SPriovavK6A3WeVS7uchxsJ
b4BuU64Wm0vP5E9S/ZNSDMDh3u8+DM02+dDaydxCGoQAR7aSBz3GKx6H5XiMeqM2qePvrb5XpJdn
5JKUt/EV5zrvbswlbhX+RhU+3pO6VljqPRVpeUIzfbW2XuyxYeTrKH6pFRIHuBqGG9UOojsgQuWy
6kYyKKSCsrcs5uD5Y1Fge/Mr4tf5VLD1caxVYSfIiziDOL+kCfGABTB4PW0f3PMs4wAQU0Asyk/e
RUWFh4HXJqUxwIuE26NL7x0n0Qhsj6B0ffegO6iCkPJXSXeqTwUMxbQkdUcP0OdXMYrW7vTzcQ9c
gl+F6OFk7D4LCbWl1emT1YmoWqT3imhLMZLiMnrlfPDQ9qSeZSfD0Q6AtJLBAqNxrBJVtVlkLMsT
4fSIYMuZ6d2Uv7EZAru22OirKtGQyamIigymVz+1PCVuUp8K8pdnukHm4tI2XD4o19HDOWSRBEYu
GlMviVNZCfy9o4eEBx6Ffb4Lv/9j3YCWUDMxU8950VJqgeH8pIRZgSAJbsNpmc93vFOLhITnzjEW
VAUZSNJ2GT2QGEk24aTsS/IcjTRwKhfHF+iFtyd4tKxbqwyoqQnwgafoFIlhGwtE3k9c5ljyqUTd
i1C56/GWEvuYvYWoYwtS8MLNT1yxdX/bmalBVlqQETmXGQQR1e+q7GXZ8P4l+4dOttQLMUAUYihx
5u19GaGPscqlXy6TJAKWAkWBvW/CjMho0JsXQO07ogWyerT/AnMyO+gNWvICaaKIYfO1W3NZxhGn
4j5e1GISJDIzrnLZufv01wl4akf2rOnaJNnwyPqm9FQtMZo/85avx8IVRaNqT6tztrt7I2kBwWR2
Uey8Y54sA2pR9a1vvGOteAj6GV9nQQow6omqCfv9uPHF1PNgrUwfBVJYkqSluxvjjwJf+uVXYpix
ifB8DPiwRm9cSd5+8bpu3XZCH/MbwIOt9eZHSIZyLdDXf840VAPdaL8uytqJ7UTKiZPmpN1TFjrI
J9LvRdI7V+EnMgPOjqhF5xOrypyNp7CJilS46T0y70jqPb0Ny1m+rLWVFCIOpeNd2V7/x3bCmmnV
8KFz/XK2MQ9wtaWiuP1Cqms9Bp8GWPUugdbmRRVNmOwU9RQfDUAMeuetxAfKyxpJ5frcMf1R8XjC
Ib7UH/98bIqrD1BDIEzEK1K4tcJC0yayKysIqM+PuuCMiC/22JAdTrvFWD7JYwzK0RMNU5O4Mwvn
k0H4qnCtVxxV8zSoqoSWMJ+B9pL18eOAHHZWgcRmAqmqtdm27wSrogKV0BuNyLqZQ/L6ENgdX2Hf
6XdHoc79okioQacssPIX1OCGRP2Qb9A6AbvPT0CB3qnrdB7lFRjBbh/LupZydmKCaw3LX5zZ/7hE
x1sMNU+Q/jRUxbHYK5aYcq5zHNwt7hHhUx2Y6/kw3glmQvaR8ZMrjoNP6r0eSPVGx4eFIO2daUpz
M33LOFhhZtUjuPSbnVpb8qzcjsZrdH/ukWeR00OFz4pJz7ly9TR6yKZXPE2tkHAavQbGfuefvtgD
0hOkOEYZ1HvaE6irwtRhs3bIeu0Z/JzpAeNJ8UTkxVIQCUVbkR/wWGofvcWzjsosuJAB/83wTiUl
0CX7yaPHOAtimth89cPQn6A0hk4movPfu3kP3lxCKY51YLjzJu9Hr3Ce4PWQZDz8m5zmKceIR92M
466ZrQTf2GVM8gzH069e9sVZh7FBUJAOPkqp+fMJyU4LPZ3m9JvyTm2yYXNKEQX9mXoF7rDtFdoa
8O58OJET6a7dVTqcu1I2ngE+yBf7EVOrSqXupU+UagDAWN2DRSTnaCz7IJUWEPjIGINC09jCDfa6
sFXE37ZI/KFmtyFddkdlIrip/3uiWMq3ZvBM/tvmcothHP/F+mTbvjz7IrlLfIXpoqc03zQNLB8h
OsDA9zqaXli2MRu7b1rtjqfdP+j4RqJxIJmrKpi+lyNfHuUii4gk1L1TB6FLyv4+ODPyYfM/UMvw
5OLSCXqYEM6JBaDew9iKMgKC4uZey8WvyGpbZlwrQLeKDiv2BhcBPKxc4CWB5EWyS1yiDVVisYwh
f6ExRSKtQKUxXyH2bYDfE38Z58F5cwRzns2/oUAI2t9lQwaUE5jk5XGETmG4BYuxudUxNvnJpfFv
ij9T7MijCMJGyxW1A7iUFJKh+WdZkZ7UysqotYG9CW/LapWTAMgjy8AynTA4RVZXPkSim2LoukNL
bzuJLd3EoKr1nBA7Pxg6JpY8LuVUlGhZrmGLZnNK36HXA/tUoekLsfNqeJ62fX3OOQiJ6Zc62UtB
9RrBVFvOusvybMQivxhtW8FZr00IqDgbowW5x2/FcQWD0UjIRBEnQRM2UvJIsumF8MjxGcGFD1eB
1j1fiVrQIe3CTIhJqGcO3IS6+8gDWtT7F93iNXc+lKHqdvwhIGZDavqLbFfwczRuyk+R5W8ivHIG
dqBPWFyU5+TC29e3yuoqeRaWUw+S8dK0Dl0yusr40C0iZVZ9GOqSXvgp+JJjJmb7gfvlIx0mmY3N
m3lO1crmanTL1fUzES0w3hL+jDTP1nbtwybhohy2w1aAAsgFqaJaQyXggJXASM3LbzvVTQL/7ASi
eJDTwPKkOiy/WzEYEEFKKHYcanqx5gR30uQMI0+A105S2KLNHxykRNVujychQMDW6fDNbLl2dcsi
m7JUcl6bUoGl7j1jeS1eIJRWQaDZQwwh6ag9K9XG7Btf60zxawbtqhRbL09VBt/vNDprBWxhkOPo
ER0+QFCVDQcVtqJqRU/oFslGrYwzx+FihshVvwII0aYf9bobCYpHLBeAN2Ah6aXnP/61xd6HQm0/
538exCR0gRzcdotVpb6yLsmljjqWkrHro4K72gW3flD7FUpLix96vvilHu6bjXxGQ4Ac1uWdt1Vq
nmospB/IBuahq1vsIQTwF14zSb+0GWlhVKiCeyT+aOWO8CYy18u5OORa00vUk3Wb13CDjcUc20vu
gQXPGYNMiABJ9du0yN8H+4QY3jvExAw1AADl5c8qOtsCUHqihPyDXjZOWv+W6ouFbvUYvWceIs+V
/eMHmDC2RGLCazsUv4XCeRcFlYXpfhkoyqWZtu0CnjPakEcfhwF1rQEYRSouoQ1dlvPjCF6FT+NQ
ok+/QN4BAB/DBejZXC7VyNuxxPuhmb05F4VNtI/gk9+ecrX/ucZuTi5nJHZZTSib5rmfB4ZLQIY3
J5uZSQ9NhCBWjRccYZiRJvk5NvWtHrxCOW+ghBcuSStu6WWRLU7nOZYuYOBUGZddEb70MFHDsnu9
xTEDvX+oHtH779EyELHP5zD63LPh9xmFs+pwWXk12OS6+dAf3LttDO6D3wZeWSAO4I5h/YzpQxX9
VJdk+dGDjy9FL7xKWojXSNPP2iVLnoGyauaNHb0R/lC61/cXWQUTKdVWzDWuIjOKVwkf+cn+kQqQ
7f+qGzGxZYWcxnLS/guT7AltTnE7XOQit/MF1Vtb4iRpdNTy2vgQlzH921etdNaZUYEhAQm43Gej
PYFcwVCD7U0w4scIGDsYkmvxfJmLIZ7GUQpCGDVurLdCTn8JryDX2EqlFDfDXGC7Wyur8POUFBBl
vqRcit3hMBzqxjSWfCd0f+3QOsIMf29qdp6Buefpfs8aiVwwzNtbDJ91Pm6F9eY1Ifc9LiQmdxSb
ZoFNNSPzTVHgR48ac72MhdTAhQXnQmgDGVJqVTLpPou512onM+cz9jWbosHoBSPkf/PfRmu+Udth
lvAb2PeOxDNqfpqkH6/d6vK+IKCF/Xs7iJAopw0r3l4+EVF7T7k0IPOZF6JZjvmAipMZWEUDlsbZ
vmt10V6OAz1v48aCcxkkDcxLvebiJYqjigl9zHsSptKMYow3MRJRMyOaY3sJziHoXKp/WtfMrokb
0mGowrDpiCIelTQ0+EkR9tJ/WMLblY7EWyN+2V1p7K+fTcu+uGBIWNM2ZK/NemfA5Uz7VBuWHg8f
Om0i2YLLB6x1G1IFl4RK8JJSc1qppF4X54zASVx9lqWrokja/vCrrTc12lCI6eFFm23KrHQz7r/q
PveIRabebRjlaXprjtEgoKtq3XcZ9H70IwAwGaiuLn7rX2h9QMrdbuf6c990BC4BdS4CKRkS71kH
4GBNb626h5XmJER/wHIud/3k3XbOEzFGbCrI2BqNl+lvaSCEzSJTB4uaMzBaxnANEuJg+qRjWOeD
VOOs34Y8AweFVhrJheCTsfotupU5SDuhJ/Oa7Qt2OcWwFFEZT/0meORMEnK5M4wt81MnXUxb+9DY
rVb/fZgoIgj9fGHKq70D0O6lJGNKRvuQE3s89RmxuE8i6TsYZ4xcaxl4KZBtxngdwf/Pjm0Sjkkv
EXEpGfB0kaCdvh/2NC961f/ZkF0hoBBKMNhwwkvcyJbvbGfYwnTdRGSpST7U55ZWj+1QtI7l7ouB
5QUYw+UWQdpl+0Z7BcqToj2Jh3PGzRlNosZgDz/IuQfcz7b6lgEPvT8OH+Ur6NFiKuoaR03ni10D
4YIr+AKWCDGdLmn3RKzUa+Yx2LqZQJtqeLGuGaSA/hCuxpTvUBj8OK88mG94fQPjL8mBiLOxYlCv
uaDj3CWFcNBXCCKlayvJXmST0jgp+GwQb9sSyUnugjzdmmxn2DIjvmz+tNBRQ0sUIYBfvpm74aym
N81P2OYeZH+UQmso1sFmhBpGJi9a6AaYMNsVOKfEHNZZm2GYSRO+R2qDTH6KFlFdKr14Hwo49S8h
vf9oogVaNa2IWqlTNWrCaM6crNYNl57gGapHO7k4hGgTtVh6L1Ws+jH5j7kJG1BfIbLcXZlUgSzt
q+4Liqvazvwxn9HRR1+qIuPpwbYR5uSrV3H+qYzKscMOTk42I/uZpQdpEWV3ET8teSEBOZQQJNSg
Lt76z/zIiAjg/WfpR7XfTDvZMmFOpq9bFHZOtnYGSdgifyzb1IQHr9CSl+wQRJgisDbEaaUEh4L8
8YX/D7I3w8PyJQ9htChTdrwxRK0EDTukQYUQ94kqhBwbbcQNJDV4pw1JYE/cGo7q2E1OdWVZcuJ3
iIY/vrppzKvBME/6zE0XhaW+CCRezixqWx1YRxdf3fkSXKuBMRg9F1olLZvgmsieU8+zHgceZsju
RltKhiAe3nq4SPtrLBf27ush4rbmRHRhavLeRB9BWabeLMpmmNfAj2thDUxjCx+t7YyYXP4U+x9o
xUFRr6McppLDF/zDokixRSmWbnGPKxWL2EwrRhDH6ukXIcUPszHi/a8MAeFaVezDD9CGseSOT4dM
4YgdCYoqRpbLaGIIlWb+FoUmQJeFvdf2M/ZhUmDAdxwzm3VBaD/BjJGUeY09B+Z3Uw2NUvm/BFrN
9snq02/iKa2fkg3Nq+X+Qz87b3HRUJhmGBUeceemtt5rzA8TOWhY/OBDI95srRqFyXNg0akCtgUZ
APHc8pY7hWUkM63GJSBO2GDybOldxDCwBRIDwHk1l5vEMHEaYTxuTuDnrJsNpcYfR0I2meMPXCQm
90OJ8k5ssH7IFjc33ETLkvMJLKLo7eJu97cBl1iNUVHoxycfNiza1Tcqv1S1CTJChQZWlumOJvyA
IuaI73wk9n0HedU9E0d7AXjsy+S/KcymD5hIMY/NkGtKGrC1KY63HDoe5GxAIBfZTE1rUOyhhpjO
DWJYg0K/uIw/W4EffI1cOxKogPuo9qfvLJUeK7rSrLQr+IUL16Vv5dSE9GsoSwIi9cB3YCrLiw5m
dE5hnnxYdXxq+z/R3y4tZVQ/cQxnAJ2Dir2s00ZnssrKKYI6bymRaulT1AAx7v2fe6oMLq0kb0YF
iZskOP/18Jv95cNaEz1ReClm1cGIuj9c3YLXILKs+HWlFHiF/vHO/q4YHvtivy/S7GMpiydOP/Cr
enWijxUtVzpMLh56rjx0ysFst3SN6JSeITLgEoEhhaBqdoR2XYs8JUjwfZL7/UQnW6JusOOuOWyv
0DQ7o10WHPoO3quFyVJLf75TcOjJVrjLMUmo/ymjDf6xYPnZ5CGez2vW2zYP41mSknLItQgYghP9
iJCW0gHEegrXznBsVfaf3STzaHqFlxEAuQ/D6voMURsAGb9MGQ1/Bq+S/aYZUZZFIdbigbFctOQl
i4UcbrtkOgcNa3Zw/xs1QVSa4gBb+EK2vyHVWuV+bBiuJA7LtNpRFUBYB6JZu0NJEwhMXgpcBZn6
tYNAnqylm7bGlQPHaPsX5L5TK/UOHUdx1P22GTcOSAK5fdD7zIIfXiGZ+AYuRumyz3YjyUtJvHBx
BfyZR58YQKmn2GK/sxwVQ2ytMnLrtz7A5nrzRF9L+DFmtf45ldH62xpsobN0GBTVdZSHXyXYWpJH
DdiqodnhUSLMZhgSJmcDWslm53pH+m39TqocJQfukMj7YoS6ptNgcu3/YbEKII1bca/YL/tKePqo
6xdEspVkdV8wjxGKg9HK5SMRiWMrdF0Vm5Sh7NwMEykAbmKLmipv4g6VxJYzHNh4SKElg1dkE0Y4
0SqVvTr9KcLvtudRwLfYiaHot1ZM/VYclPcelqpN5JSXt/rv6/msjuGaTDxVNhh/GA7OAcD9or6R
bc8MTGNDt3PrE4SE+ndDA8Hvo17kgb8Lqg3Dq+Fo7oYZiJ/zwb2eM8WNkN+XcJpjvBjJ4w0QrRCB
fobP0O+1o3mllxbZml+mQr+MgBgnW8u0vNow770HPmVoZ2pJlYQDKfAgDM3HGZQ+xAwPRRHwRJ8B
uzy6NSioOeDLbkuRazHEmVX+hv65cFkEEif1UmXNzQVSvm+l6Jzs4RlsuQjBnbrJ+vSMoWYDS92b
zAWCfQ+C4z6IS2bPzNR5UaYhfwhH/Cwwf4y5kDZccaQ+bhK+1VjzKH3mQR6BqA9WPgZftNzB/bEZ
BvYoxBCOLeybbZ63oVplgPu0jHjnXKIF75ON/oai5cXv4vnU0hIBqXY854b/vnlz3DRNEMzZBsk5
3Nq2uM3gF4o2mmDj2CIE83coJiYszh1Ew5F6W1qAxMDsV2sfH9EA7Xaurlz9HTrLkOBXHZfZIgi+
HIFTGgALvGwFYEHQEKV68FssBhJhbiHaUOsYwe7uQ8WdKH7woMQWgAskkSuDgfivZFD93uvmXWi4
pcuY7y3xedSJHJrFoFG8vR3D/r05ReKqW9lDb0nZhHtn3nM1UQXBM7XeW7E75NY4LLOnX5kRwUv9
b5eksVkxyyXEiTxKfKPmqF44LJK+VX9cNQV6NdkJA1CMf6h/lAwWOy3VZkW76i7ufUuPt+v5KCsw
sTSM+AGVeKNAhKu07LYVdh/6+aLrE1zdSW1Zv2k6Tlwj7JfoPEj7IPqEybGT4xLKRdK/vUK61w+u
cNrlSe1NwZpMhoEi8U62zgLs5coMoZ4bCXl3qg6isjFGdqG/4UpjjPkjzt/Piw3kB08MgV3JebEL
za+LAvr50StEEqJ2Q0rmg0Wvoi+rLSy0JsP5ukI1N5WruLeIRV2RI2iOQSGwp0CyUXeOwpczoB2J
xzxokFpwU9vziEHPeBDnXOOYNgNJOdZj//EP6KyGGQ/jHsNavpU3fcqdekysMUk/Ec2ifzF0zrJ9
K3Rt0xr81BhXejgc1b1W9kpuPkas9eHEJ+cIpFRRhPfRxGx/WjJTD8ayWsQqiwwVuRZN/xdJd6UT
yMj0xeaVrBAe4d4vitRXsdpc4wtmdVBlk7VC3ax5D72ULxI4iOKIF7EpJ2s0ri4QJO+UKyRtQ6fa
j0z1IVZHPnakoJ/Y7u2uCzrjvFNunch4et3L0I90lOMYWOXtaDwJCIsyu7naBBcGmAxuYRtCYRP5
0Ym1ztLSVD4SjcU5qIOva4XheMLHtNzxh/vyiXDXnSEjN+FtgR1fyQdCtimowVGHS1XVim/5Jjvs
0BIzkrY7zX9CcSrJhfl909RGRpWC7ZPtApC6qJ0c8VHcfnTUDmR/vgfNAsJZ2YIRcWKB+YQdAV8o
yiAVwz+18aCm+/Fh3hucnLmStVY2wHJZAYD4PtogoTTkJ2guZWsaBUn2WMs2wxQdVQQ/WMA1AG2C
+3bx4aus4vUOi8iaSl4xlLbYfH2HqrY7CJsEJ8pOZYn6TeO/LDNiUST2WIYMG1wK5+b0TQ7X+KIS
lRQJA/Shz9Ox0N+/Yqmb6UCqGI/TfyLikFZptNE1xI6ZgojnK1ak/Fk8UUmSe/7VJDSAZHgRrVK5
G8K4drjTzKHNH5I6jSsz02hWL0pDNELy0hFBkIpD7WkYbBRME9onwsVyMqD+PKQ2GDwCBIehCslF
AViRVZkdH7g+wc9Fo1g5sx5tlTfzb/y7sqe3C3uYyfBOupp7sZ90ZoFuhykMDgKMX9pRNR8OIqI0
suLl5dLNmkG/mFAfXkeQHbhnkB6TwXIap445TkEGfMrvQPnOz2ZR65N+Qy9cqk9sMqOMO10G/FT/
o8BfriCcudqTVzuuZoBJJVU03myJ+XlLzosSIxWnzSjIE2Y9tBzeVi82LMDFUNlgRMgU159ToVSp
+sj084d9L0EXR74sxON91wrP1AW+8q8qFKIMfxwEJAo4tdxIjDlWkyFYwCGzNa9ExnC2ANYLIpCo
XuBImabAED64tG7Ng8F7YhMZKRLebnRausQKxw8Ggui1tp6RkiTQBWWzxD6bzItHCmYU4tdQkj55
F9pMtBFZlBULOEBp2I54h3NPF0RItFTeFRfAl3AnpddEvbejxy/v/Ot4fd6ckZktdxGQiQ8MuFlV
s5BTDfDGD+R5hFEwesTPfrROqpGGAzFsDpDCsxqYmWl+DAtBwf8wb8ZxCHx9yW9pCS+4vC+qmKSi
/fAe2cbvJrperVchwP8URiCAonqUWjNogfPwv8931mgGjaOZqguOBYtI8L/APQQ36VyNPbbv6NeH
Be1oJOeCkcoJzgDzPkKp4T+Rt+lmEtC7Z+dk1WnlYRCOmcSSDQZufuSWOQRFLydheY/f0CjjcHs1
edU0oHm797FbQjt/6IImWzK5ZhdzP3sL33UvuBaXvBA0/4BoWSTws9DCncmqJp/vLUgcO1ZEHj6t
XwAqqz9FbjfP9MUFFiR3Ttbo1T3muCo+9O7kXWxNKUuJhh27jMTwGfGTnYLEKMPSNVH5y0Y2z9Oz
30ausTbeL7Xd/IJYamDgMYRFP0LZD9J5gVP7csuvtboxEJ5l7F9vju7plILU1o/pFIA021lkrjHi
vQvMcoVWpTdayfxQei5PLLwtpirF/sMYdgCO3RdRuZCTfMZcxQAsmLdpcxJ5KyQ81D4VQvf1gbim
ofixn7sc3OiurFIeInqOm2FGcrqkEsfwBW0CCOnra/SfuS6P/YXkOpGZ44UFKNhyomYv6DZk07mh
pgLnKOvYP0eGb6p84XYDCBhBcTlm1Ekhl3ONCml3WCoQrF8PRTa9NWYlISZyOiyOEKpGPX+lAh0k
PPk+cFRlXeLejOunBG4Ya2uUbYpSo/ixcfsa8OTj5/CFEsniUehU5waCxJ/Zwnhoi9APFOleoyQ3
TxgwDPDwOX2L67I0JvDCluk5DUAhw+jZkqqIj9s2Wshhx67Pt5oXzOM2NCXyDhWk7h+r3szlMFVs
YJwjLxMmVnxQ2IP0gQyNRjfeCiLbJY6paVGz63vC1k8ot71ihwPn2c21YD929UjYHUC7rNgUNz2t
ixHTx7s0Zlm4PKTTHAm3z8EhYBFYjjKDK8dOUt8Xy6a+SMVy9w1oj6hgMNIxZG9JRIZo2T2SeDXH
m0GOBBunuNKHyNpYsKLM0e3JRh1SiTLvgy52XTqIdfT5SAwn9N6D8J2l2AiH+cxyjokkBzNyi1Lg
m7B/YWTX/qOW5Vo6l15Z7XiNbG3jc2PrmfFOkJPbX33VF+gT5tgQl5dHffXMfO2j23vnULzvaECn
uYalFQCoIAKI1ucaJGG1Mr6dpXPByNG5+UsFr7BLR/0XIeMrovH2ZscExK1BUoFl/Rt0SlNCK/TH
eBKEsDhQcCryg8OWgIduP+ARtwkGAC7HAswZT4m95Gfrlc4tuWNBBLHBLSw+lq9kfvBlzIzCM6hD
frrNZtn5GYgndrs0oXYEvcbqn6CAVVVLsgjzCVhS0skBYeO2i6HDSIiDWZ5hpKsmKNh2GrGGFwBb
wABf/bNt3aQHyOYKTom5Cs/aPlhce1T+8WSghybtnSkB34KAbFNpY4bv6f4orYd8yBihuO0B1RZV
jf5KIchetYmp/XK0gJqVq0a6ZuaB7k2jfQccmqxKs1aZEwPzRSxxd+Gjt8fXfabBlOV11yT+9YX7
06T9nAzI4VjGrSN7IxZY5c9ZW8GNR9dcuIXErCJDH0mBWozC2HgkH3EFnOhhAmohaGNXm6UKgJex
2zUAUD3fNCPZBrdJl+hQ4yAOIAoaPZXtlmoUh8aIwSq0DloehgWdfRj3PjN24aCMjmyHvN2Uw/8U
ohHHjWM1QDsq5DhPwLGKe8r3B5nJEjNOyUChUn6u18aDaOv6MOF0nxLAHvavzPOA/Gde3583rXSm
PxWLHui0g9ZAWckmyJt5cz8DF8WPUwMHWh+GVXIbSahZd9EvCnLzmJfCFSVYytFvv72FzMe9IYRK
9JtMJu/sBg1HAD37vF7ohPXVhNL7hH5GPwNw4seklic611WlXBcq9WacTAMkkcnhY/0bqT3LfqRs
ExyL7gDwlWQ1OnyTN0MyTTadKDn+AjyvI0ccPnZ4xL4IbBQx5zQ0VXnwnwSOoryoG8PK6mLfgELJ
2vGK5A6rrw3PTOE1O62LuFZATV2gLuaVVMjmPODRmdbmFcl29LbUyAXhzZiA+GdH4bLzqkF0J/Ye
LMWGDkJs7WglN4SjY/oWc/N8Wt2HzUjbrLLG8bv7JS7i1Uh8pXpRmMUnaoPs7zRCQ6tRNd8ZFQcT
SQ1S/zmwfV1PeLEbmozoZwwTcifMnKafv0XFkkSQV5xbEX8hmax5178/xxWZlsWgJ9+pBMngbmyw
H60q6R4ze3BiT3NY6ll+5EEKdO1D0FwItvYV2vOnzJkns0dJieBD30Ee96B9LovsAjnV6FE19C47
YiGRdtLgQObCWLRr0ipKChRJ4Ni4gTrojhL4CaTPjZoJ+BwNeYu4w6n+hY0XWJlN1EJNk46Q1lv2
gBzhjWU99Z7wc+gV2AzyRI4p/Q3ApNGtTnekB5sDlP6GPDvkS8n1NZoIUh6o+ItcZlq6tJEJ+7L1
sgNzHi2i+408ZxLMXY1Di8hpW/LWX48syYLP5aRIBUtJFT5pm/F6rT6jQBUKPPB8RWCP9bcsewmx
cdnMP6JJeFqdY+n23Eq9U8SYNK1mLhoc5SkntjL7ZHlheI2Gcq8alxKTz8hvBkTzq/xtXijuCtNa
JGEeFu/yOlnXw+khwc/j7PW9OLyKvJIl8r+C4fEUCv3KSmapsSEVclVwN36eM3d7Kr/w5mxOx3UL
eGByKSzXyixhYwc8YDffp2AgZjFDjKZoFXtHLJacJ4+57klqlatZc6jfHjAoYK4rf/AVN3JIdXMV
eT6eQ36wHWLidIP+LlVLt96dAcJJssFANZ2rhtwBTF1j6nwUGjmiCtsF3mhNPspskwvQVHPSsdpW
AbbVbmbNz/5blxBOEHPifSI44qYyz4K+OSnIumNeFzhmPwQ5Kicg0VzqiIQhTZgCsNllZQzOLoEq
Rd16ridxZO2ajr5r5fEI6WRwTYlpJXIVClrdlzMFh/2EA5L/jPRjiUmGtcdvTLxAXNfGNgwSPxbM
DziE7dgT12jtfxD3IZJLS6lLD2nVd9ThW+KUWolhhZj3EIXQlUioHVD/+XZ1jaEs3yQSoHaR+MWp
sAl6MIvL2X3UmuX7u3MzCqm8GdtZalzcn6ySmfZkpAi+f3NXHyX3OApXm6r1Eznhi+h6IK/Ju197
vazXn1DoeMTiI3Y58wmq8zgam7Kqv0q5ChzBWfxL2j8CacHzOVU2+oaTiwaxSGSPuPr3OHL7uG5U
zkEWC+VEy20GJrFkJwXTfwQN7l2ASWj9finUk0B+wRmBZWxoXDf9CcO4jgEIHY3u2OyTdzXMGMUD
Q+poX78KQK9+V/f8BG0ZQR1Muk5um3McFA599Tc5CSWHN1IEaaWsy9kzGnpt1m+WLLUZwfAU9/Sr
2L+FTrlPOEO2LRKVvjTIUtEnKqRgEmIfiT6uYn+V+2msMs33SSUyNw1UnaF7ONJBmAhe/ccNJ555
O6YHlvVo3OiEOrhg2QoKESEYAIf8QSAOLwefPceReG+6bN+Tifx1LVJyKL/4GeDB/EyYKQVXcazR
JJxN/ZvvAeGmJ5el1e0REo83h3PBeQAoZQ3qYRypG9kO1OmN7rRHBQ6Z7K7BMAcGAjKk3YE4KHPO
ZtLzTh6JYvO3cZ7REGZgJP+sYO2H8UhKrNERT+Jpyih6XqhXsT83hkr1HZxrX58ZGbCK+IHjUlmO
QQXjxLHD+jrtprTPUc2DOKOf6rvtz0uiFP5DOWc/R2v/IeMEBwOH9CFYUT0N98MxIXlaV7aIAeKU
+GOwTxcdyS+G9dAc63mWA+Q5BQEgiLP9GckDaBdGoPna2xLGhYKFDCULsdZgky5+9ZOsck2ZFFCI
ptcIF1B2M4tpwXLstoUjRUWqGOlg/rfXj8m19xiASTNO9GD6KVIRIMKYapx3zBrK6axJlZsBa1eo
MtzvyG+bssJh0c+KEQE2bSPuRW6lyzcoobQndUZbLLgJ8F1nDRiHjQ7FNv0MRMCxphC1ItoJ7U6I
tONY4kdKYyTV6AeuBGhMoEwFKnuwYAT9oyhNbih4zzg/ZcltZjDpeBs9NKYmDO0luLivjUT/18DY
/1aLYi4FtZRkmhhtqQONyBJ0oDma1eCCDm0GvgbNnnochtdIwkCcgiuoHcwIMu2OM050xHA+PCS9
Q+eMQFi+/QvyilEpbgR7fe3WR41Kp6l72lLGrAHNw+GerokLMjlYCgr1bNcjWsq+ySL3yxGl/Maa
7u5HHg6OPn4mYy81djLlWKH9mjXSjf/G8sD/CtdVvKyJmu5xeFZ1Ptnwd+fYcpqiDQlggymucSZF
blFssxTEl2jCFkrxXw9LI6gMSXhhmTaxJu3OhtnifL+0XHSkNaa7vxEvR8aD8FmJIGe3Rj9eOX9L
rRE002SSUl0qu761rlq2Oa0fu0L/Nuvi2hL2zLadkvDGElwskB7KMXTnwgOfY8u4jZuXcU09KIK/
QxUvVmh/mvFVEGgu7f7V3wj0HOuD5owAIhjlYF/oK3RCE9WYQ+LEwbjJ4DcHG+PqwxTT0Lg8hchQ
ypfwqay/SK75Ti89ZNjV6JLAz+lyetWEBJ7pPaoAb9gx5wwikIIxARZQskZeqW/w+VP61GH5bJoV
M/oHQSGYyRUvxOA5uNt5dhyXwWx7Ij7bsNPYLPq9CCQpCexwmB3Mrh847W4I6trporqk/MksIZW7
q0IDHciBekvZpH6Y9JoN07Ar5YXTVFCBi942gzvOKXp18kR+/co+aCHxSyIcOt/lW7SqfO53c8ox
QycvE+rYCDU4OGNbnLEC6KH5lYjj5l7Ie0KGTngwyKY7Xru1GfltYEqxxNdK5j1/68dunldwrz6L
l8ZRawh2JGEf40XTvMYlxMenF9/h+kfpbYGo0IRxBCCpbvCRHb0+IgiHR02eAjSKK/e6bNGVE0KE
WCnS4y9h1UX7c3pzbDJ3JvzejR06AIFrqCFstPq9pEM+wJfgSP1LC4mvth1BlMqhg3Yey8OGx7mn
0KovWNprIxsWzASqeIsPJxQNBoNrE3DAIdCNTAbojaaBSURfBPbsrE8auL2VQJrQQ6ViD9Egw/Wa
dc3p4KVRvLT3pg3VJ0whZIxEcyqX3OHW4jB6j+A9oDbO+XkXY2fCGobbOEo3hiK2TiVSoG61Zyxy
u2RrQxJrO7e0g9mxliydjlHJxLrTWIBUyorLeHUgUmyZxlBV8GT0eJB8i3x/Z8ROj4X05w9oTI82
NtBXTXnHmqKubnhcNzxnHScJGOHHFCIzomc3UZDVZYcOAVEHGDX+G7AVYsj7rgbvkVtvZgyX8JK0
k/ajeaXXgUDGWiNuRDwJvuzPpMKhKGgx5WJbXQr5pgfNlb4Cghy797GLxzDFqMjRkaIHz9fw//eM
45CZX1e5cu4RAimx/64T+MlQRm6zEfP2EYhjiGvzdAsdQNT/5f3u0o11jm7KViKANmuiLB25+NwX
+MPWAWeNCmVjfMZv0opUiQFGoF0/RScmAmO1N6ak8sT7rhB/49q+5SD6WX49mhtuTsosImka09Sr
yvm6yo9TyvbcImJv1fmBCN40JnVQUxGCXjgfVPvBO52Eej2PLNXldR3tSLoptDSLwWucJJTfQZq5
GE9FQYZuWMS40gTZxhiwzqo9OedI7A+sndgrgfA4tGgC/2wDPwTFAZqm2J0seK5htqa0Rf+yeiro
Ods1+aL76Z2rHoL8jp40wJWYlOvIZTJqm2vExV2W4G1hWmZRW/J4hAoUn5TiKhTk6Df7rmqsAqPe
2dg51XNJCWjEHOgU3+IRmTNcnYKyo1/6V+hfd+KrE7JUtfdf/tdrKxdCF8nPpaB3URO5a0CiMheC
1cx2npNzCzR9KU6ofqXAVtMG8NoXwIJV4C7adgZP2dHCNl/Eyhc/8f191REUt24EwtONIxvE9eZv
Mw725aOiHGNEDzu/3F+9tEsNyNx46tHoMsyiFhbxJVW82+BFxIidvrG8Y0UPzW6CeQVDxxORedPq
TZxtyrLgwXTy2GXqsY8u/b+NQAeEhJaaZ+l2GiL0Itg4fNNoERV8HvXRyVJrU6fFeCWkm8BzLX23
gPFvhTbG3T1GMYol/6c5DQHXyiazCOl1Sbe9sCqKOT8znWsDe679rZ9NOyu5d0YucLHoJ5VtB5wU
i8/508bdLpkKx2vZHiXTJx9/Xk+zfjknaz+pdr7GgEVMvL7Q20iUZlxI/Wpb+Z0P9gZycSpmDjxb
KAdb/xl3idM1R/cHIcJ5IxlXfk0Fvvcp5Cjn9kVXae8hsf29taWBPaTVRZBhjDOcxXtl8Bi5nXUd
OtSQKBuAhhmIxLmTbGDMZP3GpMXmzbTeBy6qE9V7lNRSS+zpIcnvfYwqK7DfWnN7y4DixHVYaTt1
OWSwN3ZcCEjbCIlPze3oIjFBhQ+FNOnMfBz0Aoz2KU2MhrT5YkwamJnLUNUpdt0G+wqjGX69/ELr
/Ui1oE8aUUOXScNLL3RxYQFzQuBsKetVM30T5o5qzcpO6MHvx7fKCRsuYvBxj3H/RQuAfPvhW1sJ
SpUOY+HrFjWFKdvs0l6D/b8flLzyxnFhm7hy28IxByLmcNLyiWpukfzTLfJ5uuFq73izNI9ZLJIn
hwFF/NXQsl9sMIpjXbi8BmbYHd7YvVpi+HAaQL94HT6UL+fL9e/psD3quf7ODVp62+ZKmTSH0B6O
hI322JEHOW6pJpCFJzLzTyvOBiAZ4ZOGjPylcKV1CsprVMXj40hpCUG6W5IXDqZ5dT+8vJ0AK3bb
6azp+N+Ozn2yTmHBO715DfFN9/d1vqnQsidY5QMxw/L13DJPr4tnOu7ZYp6GFyGw/XwGC00zDqXn
e+kryJwbF6WS3fhoYXxWftrVvsjn8XYIry6XuAoBuxQ9nEV6jg0lrthWO4g1aWSTrh4sIdWs4I1r
CRTzSgZ8WYiGTRvBv/8avyuFaKztGVQ1McrIz/02gPD5E8zOvU0+GSUZi+jkR5AgIb6etT9RXd9T
UAujMclfSboge+8R4bG62Uw2wJWdCX5u5gXXTYBDG/5jWgdhWsclPj9Q0neyqJ7iegwc0uu264k1
pHsV5eJ8eDHPiRn76cHV9/tCqzkADsmTQQ2VlHJwHHUkcXR2v+0DvuEcAjnU1h+7QNtJhWOQcz7b
DaPAWrvYvAowZoA+RGAzmqJWvqunQ2F38hhXgalCm7rf1hVEptZ9QTGlNRBXjmupGgH1blOGqA8e
PyNigY4mZ9cfPrjyVpREVoFyV7yNoQsLnfiB4TjSGDwKnyP22ZzdwfeuwWHpNKxlijPnEGJ/8BQx
ue68GaMGVZYMIdzsdj33rakpglvvAbfDOtraFRusJlR2ochedwugCguj7WO+4glbprUyWR1imktv
nRG+8PDZidvU7ZyimLtfQ53q8VJfprnWmxeMvmIkU7zwDPwLD5Sms2o1qkbtqp/rRY2j4BHalqxJ
y+Sz95EkgxQTr7GqOpBFJlA3FOvr+mQH/56S9dxbrscfvw8JLLO3GrjrQNjQTWPb5+hq/XMOIvPf
0/jeboKu/NrTm8qfapcXSSHN/+DMLTejP6/E9TA1+D4Xsv8s/bpGBIqN3T/rUSunj0dJQXBBI8OX
DwfjBnhBBr0CPtKGs8pyoaA3GtaBsjLiPdfOoS0jH+8pOoBryRyzgq6QxlUqRjlDXqsdoebPnJAz
6Dqo7dQkZ5y7JpI1ZpdgcrPKH9A6+EmKdtf+KOf8lKf61cQuxaFPR8Rr8G26claBK9QoLuKjDdPA
pJVhfPsJ6ssN3FbOQ3tir3rDHOD5sKh/XvRJ3uBesSv338gUhNV3My7EqkzRbkWfRnTVKaroOXo+
n/LF/sl9+02HHG95HwRjwYpmXlNT3g3axxjhADK/z1n4qS0tZx+tvgMulKC5RH0GJJykBRHnBOu+
+8hvUsOv3B/u7Z9fDljTGeDoJfTSkPORoINK3KqEXJEJYnpr5thl2G6EODxZ2v+1h1BoQRpD9aS6
M+R4O9n3gSkGL1OsGxoJtCMG2mMYqWH/YB3DyDgzEXhBlLoQHuqmtKM13QY6ya9s2edfKpwfXGdw
l7NLgOKsFEkbPqWsWFvRVfDD/7YgShX9QPUdgWkARr0XXHRPy3Z65LRsYWFCzYHPeLRc6DnGiNfo
CgF6eyy+bjh8TzQ8QlRj4IgLx84jKp+Y4jXYSnHsg4IDixQkRSrBS8+wkR/pME3mDamI+Tu/9CD9
YlPXXou8wHwR7JQv+GrwI/MPLl8292hsQkfi6SEoqFxKGBcTjxbCN1kYGvfBhs1Kwcaq4W4Y0q8U
UEkUQGL7w5zjVrXSYJxyRRdcJWyFXA8fX75vJwVm2TvFbMNZe19bCeOhrlpCpRazSg9JrrSvKpPd
qfuOWTQ1FeXi4BnYU/I3eYah2O7sPNTfHDaSSwQ9afof3aBiNadQW+zXeA8ludGet8sAxXLDwKME
t2kHw+QxNVWo6oxfmpuHhBjJ+BB8cotqg2vuYRSl3JtYN1OhbbzCNUm4MwKB/gkz1U769p5xurjY
Nyz5UfVqqiph3Z85U5LWlwCDFn6uebmh35isrJ1d0mQf4XpPXIqyaQaI6JQTEI/asf0+l/faZqnl
pj96ChgXSwZvEzGg/ZMSdLi+HpYVaC1jem5W8K1iZEG9xyd1FaMt7t+Xg0HmCYk/EsEDfvXnBNgG
huMJli1m6fgGlxrwaReD89Ank44029rRV2Om+w/y/8BQZzA/UxvNHA0I3DLsRpHegJsn1ShAismT
MpJUqweuLuCNbDEN34QvbrHiJkqmxpbZw+zT4NCvpKzdkIltGkUKzYpmBdLX8lm1Xvt58WHvuurS
G1buBJrWeeZ7IV0IVzqXyKRS+VTHm++u28aArVBpm0jVZbew4cOeS6FL6qCuEXbWfmWcI+/v/uix
K339Ao+wvs1mv2rSd6eg9ZmxpkQRjkE86BkoF8hdImEqtUsI5YYHlhwHZ32GP6HnK77n6JD8WIiZ
UnZHugwwhxftWv8JoIkMzBXtWfakDXfmHSN6AkKiuelW0bs3mz0RpZV175st5KzRsmFcbEAg9P4l
1jpho+FcuXEqCiENZ0jtXnPtwFpClCjfqJtZ1bLKaZrtmDH6RiqgQFvXkst2prdUeR6XlRibAQpA
ssz614CWf7xeb6PuGvFfillfXu+IFofbUOKsnKUJ5kzVL/5qJV2p7DnBUcnhvGwLw7CawLCk41A+
wEp9iZHqHvsmhRRH1buE5E3/0nOQCgRCExJCTZMdUsGiiwh3MtvuLqE0+fBaoDakl5+aCi/Yedli
aJWlkFVfBUa4h9xiOFpmTbQ/CUE9gh0Ht2+F+RJpAPlerlv7wMU6cGtqSe7bW5o34DI5Uwt8c+JY
XIbNPZgAsShxDhrNyeyMu4/i11nKR+3RnNz4PeqQddX+PB++kdfPC2K90PpnnY5aTqAcrrO6Ggmr
Ph1uFyzoaLSUFKPTDMuQ7yaQBhiC3+G6qZOpGRg1HpWSOMx8UOwwAH5qyDPNRHI/bS/M/rnFblUV
5gEUcT3HUDk6fYgQqNRzQmAYgnY7FZn9ohwswsZMKns7dN0H112z0tiUVGhBVyEg+IxCo+SMfCk6
XsZOC4Fahba3gjxGiXq7/ZTZlyJbn9bXdXX3Nghdx3qj3ef6DtyNKg3QAklPIvasnleNUsAaUR5Y
Me33hqWXEHi3Io0/q8ZAGAPeC+rPrbd+bGrbuwd5/fhdMRuIKMMbOq4CiGfYrzRMpHjac1tb2KfP
uhbsMzCftf7e4wGr4qJ/JWpLtKvCAAUsyLgT4nOLrSqS/TapRD/yTLljLlPySr/2GwRGSoJpI7H+
UesL+GOW4A1FgqZblEXnTIifTMXDuN24D/SmUdto2nl6dViwvLHX+MrLoCLcpotHcmJPV30Wfhx1
AGGicUbAmkIIRIRmyFFI6g+17ll75u07zk5RC7wmyx6ZAs+TsOo6i1E/IngfsplUT7mqqIxZZ9Yz
h4pDw2F5dfbiwsC9d1kuHFr+h0pcQ5cmBwdDfruxUurOAL7tvkuVJvouZCk7OmHuGl9Fjt5Wn7dM
3rOd9Xy51oeULNkGKF+rFfCnGsTMSA1XGaokiWEKPOnZvYHpeGtriiej0UFzUku4w5mkr8jPWD5L
T0df7i/udPbGrrSnPL4EzBLgAX1fiZRS56K0ucd4QTpo033xByEZN++FatZNGxoDvYtYPSbVLEAj
MLL1IbUMWNoiU5adlgGbXJOr5GCBjbkFR/dD/IQb7Lt4xp/M+CFu1zZ3QLDsx3CymuKwaiM4RsDr
RVsSMOyWYOYjsGfPiTzu84mxqALdsPg9+vQT/0T49afv9A3BxIbnYU/LCDi1Wk3fR/ED2XlCVTol
8sBmxHgnkpf0hAA4JyA1HJnFVAxNP+hILbZTXJWzIeZaHX3cQTW6E6Nw49/Bt21vj9mfHA3ThJ1o
Qvymo7jMG+w3ksHScYgyFSu257fLTXXhw/j4/tMNjODIu7WoJjfAyRviSEyUVhS6RVPzAsU/c68M
asnDvXctHzK/iRU7LzrUdTRfaFzNknDNWJSTja+mGc+ZNBvj4PMy5JvLE8AxOm6JIyNiergqtaYy
Zhz3hlDXiKhx/hp4SO8CIT/59BeQpNfBrU5JVP3ywXpMAL86Cn52ZHAuUhViUsAEFvqFvU6N5CmC
v/HoM1PYUqT2GsPT8ZuzsN1gVQbQkat4OA/CXE9+L42Vkl+yY35K2F5fO9fS/pSZrZhjNzSVGIjw
wRfFXvxYTsXj80axaBvlEihmIJD9jcyPJ2RSTR3omAEX1KrgrWf/XQNojQvbEod+du4YVAiW8x/m
XW/OHSKfpu5EOUQ3Ra+n+w6ITAxNDzhmAqkQ2SjCHzlj9b+avLA9AsnDRJK1f1oqwFDF44xLDNAQ
ljDjOqjck4spb0UFZRiM7/CeVdLgCc4AFF01n/dCbpYVDig9sJNDGKzC0lxG3kDmOqS+Jn6wgcKJ
k441h0L4aDF14US2KsS5zZmq/rWNDmC+qM6/N06O1YYbt9BZ8BC9BSekjR7ol6qTVgt8GbruESFp
QEkW3aTTfDR1uC4qH5KXfKvFbzylAsJAFQDqSQeSkDjFMDqkufZt85vSig+Z0HB1IQRG2ZPkJ5oY
Rh94h5Adl3iA52vTgYjpcb1ATS7ZrbW7i2g1BHndi7g/K3ylfz5F8I2ZPV3nv/4/qPYZl5d7NUWL
5SzUoG/r2QMQDBSuVOrNVVSzV+L437PsZqJ0Iu8YNLLXK8kshrCR0/uNYwBEJACI6TMJia3YLJ28
Y9+FDJq30otYJo4xh84uu1OznVSSXA1UDfC7PG7E8Ahf5eHPRZHlS/3oqlTPfyt1liDUHawI1Qgp
iDV2elzB/RRfNwaMnAZ7hvcfb0C2yKWLL/5me9ndfkPIUjrWjMt/CncG04XHROyBvGTZGuYpu4fF
GswAQje1+Nj1K8lb88UTmP7ajL4O6cjG269yLFmG4iGDMjKrQmZV6ERqgQi5wVw28hptMWwaeAOI
b6rCdspZXr7w5oyUvyUsHDPX01CqkqJVCDr/y3A5ZZtxueG2dDSx3o5cCLZH1iLgfO/B95Et9MvA
fTiz+6EmOUzbVpYvXrM06Fnq41wjgirIzqNS5IusvkYVXel3AszU9P85fcFA2By58AFrvZ2wouEI
rEA2Wg587AZEvMmr9jYkGhmxb0OFclXZrv4Tgo7b/x2ZKYAKHcLmAOabUiqjCypQA30kS7ElAjwu
rNEA7Rg1TI4KnFvtKVMs8ZVupXlr4+3oLJuLUMdJTVV3iorlGGkEpz2u9NvdqcmNm7O9Mv1tbw3q
BYoiEJmCQvPJ8mJmiJDHf8ywBI42nwT3TWj+IicpR5NHAxlOolodgoXYDjJh4I/dBMIjKIn4sDbL
FrhK3daLcYNrbf1WpYasXQY02oTW8VW4Wn/z2RF2Ce2NHQ76DdCNM0N/n6/zWV5XVCTL+7k+5zg2
zAdN+zmliHOQjiZPyIcbhRTQQDmANNi3fDQU63UMtHR3VTq7C2J6PdO+ynUUqA6d6cHz3NUBlr0+
xiXSBYUUtpzpVQyGUcuLrH6BSzyn8tJB7QArS0ax/9HbjqU2lZ77W80jG6CVFyxk9JjraRFsNZ8H
EYV+caAk6dQ6+ZtCPwUjBMBhfgHd5vzF8XwJfIkcdwPdTaiZCdgqYDTCeRDQxanti73qo4sJ3543
0YF0yg1TsYq+gSo8KO652UVtaJSt7aAKzWN+unmm4E6ZvyJj96x6LvECjP3v7IlaSyqMflfZO3rw
abeqOSc/BqPWjLZbgCZSnB4F3LXPM6LHLGc07rY4w1VHYQCDtLySPm/wYZ6OlNUwLplBoEPWpLTH
/LajOHS2LgRNm633JMvEM/5MJ4yTa9HaOTKyDZ/5qs+4yCbngbUG1FMr68zZS2Iv1QVXfAcNGOYT
7E/DCbiUjYd4Aqey6S9jqrvNGlv6nZys/62LtD/8uRXgzER25c3Jf3Sq18raBFn0KjK4MT2K0bf7
vweJcQ42L+feMdYcE0J1vIDk8ke/eFOSqvIl1FtlT0O9xUza6cCx8+pFSoX7b0QhIJ0NomSC4igx
uhsQP/g5/RckjA3ONBHFUmCwbmk7tferDQLgdCBdWOo1GB5SslbzYbAX285kol4oFw3TY0QHs0Tl
qA/sF0QCzuEo698/0ZUgoZdK6bixqeaS0/3RVR4ZM8a52Cp6dT6m2EhuPorrAnuACM1aiBZTkPI3
iOrbI66yqwYTAZ/j1cOXPHlIU8jSAo0P3E43nAvqDG78dqPA6N8g8JvSfeHx4vfiCTh5t9UijEi+
PBjR/+kSKzjDBCUQA7G8m3W+qvZc5aKMVmySi8H0jB/FQZcio1R8txOaYllERCAZlEXu0GkLL3yR
x+6sKv9dPcY89TWh3WW/E3TtLQauWjA2FFrU5grlC2pJvrDRSseCKilBHup9/L8fiEdTTACs89cn
T6mu1d5In12uEDVHfibyJut6EdDMd3JFcLd8QzF1+P8aGo4j6AnIliPmbVjsfK0cAdDxm0IEBfaN
5KD8Svm8zR/i22+1p4dl7URhExDwXnGE95MDtWM1E5BahyyB2GWdBdAlVP6uoUhLU4uCrWIg8VgR
Kxo6+dLh3E3PtKlbkx6RPgf1fQ0PCf1Q4y7w3XlPNI4/n+xtAl9x6Tn2YfOUYi1xI3UQzGJq7MBg
7I6nZtUQkKwrA1NGRGelAGczz+wKP/d2Hepay5VPyc7gssSuu3ilk2iStOqR40YNakd/2p3iD3jU
lQfTqMTW+GmVPsikFOJlwZuiPGkKCtB4l9FFQiAIF5HmeEP37YrNzVBmdjTepJwifsIiHG+r60Zq
IkgDkUXIz7kZNYs8N1KZamCbL/dj+xn6r4ScTpZMt+NLlfJiciDppxlnRUERMiKnxmgs7cpCKCkX
9cgbDQi9ERXvFgMYaVkm9NJJZbHLGCHIFLOyaJwxLlO8HvJxzF87ZWsF2mnq7UQxsS3Wc+MryV/a
zOlM0qPY1eHnbma9K/YP2nNuzwThz+Ot979WRgs7QyN6Iv5qsAfIdKXo7PVmHxKhwE9mFyNr2n2v
Ayd8lMAGNwydeHiaeoVki5TRD5lpMbOAEiNU/wgqxwyUyFC0is9a03yfi2SkvIeDHEa2rIaZnI0b
u+g4DS2Dq0L5oWsNKJ4U2qfoyOtaP66nRm0RmW4WVkOCDY9zXpzdAwFYWUtuam6SRfpcEGW5rind
TRevQaZuAfn/Cd5uk79p7bqY6J+gyw2qvqL4aVCTcBu4RdDhhtKiktAEAzOFTeGH6lb/PfUKGxqO
ChsqdNImIUC35dSslwMmmN6H42JORUEvb2FIHNu93e5SnSoeh77puAYEtmCOGQS0dUXweppNisSV
fQLR486Tzi4q0oCQcC5tWkepAfWwU2t8TwdVEeitcuj6oBYm4uUD59w3gFyLHL47QK5U2Mwauwbg
VTao934FedNOdZKjcLVmJ4fe4chHcwbQncFzLleIFsjN9LKbp8XKl15tPtf1I3hsTRwYQJvLFweR
MI98YYpT6jokuQM76utL9qKaJeOfSxMttMUNmUEKTsElOZgEE8b/LjMWBJVV0fJ57z4YEYdbmunr
8oROpLRSbENFYKhJ32tUJHN92OX/mdKBbMWfKWFisqhgJi0UcN971h//RH9wsLk/Ac7rmrjtvEaD
Ty6tQm4Sk6JJ0GhCrecf9JT7IUuApqX+2s6F53ktMdR/jchHPwlNNM68IB2Wrzl3YWgdYMSq1mQe
CuzTvZJaM0nGkiH5ojYCcdIKNu7tcOuz7hFx6rGcmIYbm2T/kUkyw4NcJaib0HSnN0TkGD9VU2UM
DGwAPoEEMV2hA+jygXg35n3anWoN5pYFlnX5hj7PIEQJfGGPS84SL+D1/7CkgO2J4gAXgAlFWxtz
/FUFYmNcTpmAxUtfUr5jENYPqqyS91rOLVrfAZ0pD2IHu8FGVe1l5p3bx/5V0Sb7IlqqYgBVWGY5
yMO3pvVro06wk7tT9m1t8mhZtraFFlLeldhvgGVLqPeLnwd3lSrEOJHpJaBhMRDeyUbyxbQlan3T
cQksH6lxUNdGPRcqYu30nY2C4nhyh6B5AHq5Con9pBgga69sNdCMZO/Ti5RQaDwl/vT2JqIvDOs+
g+4IzZ0OHz1Yn8ul06jFfep5xDDI2cimFxidyKW3yPkXBlQAtv5FPziruN2FitKYTtBNxoufMQv1
YqsnKwsscZ9EDuJAONCJcYDi0sgPA0N5TdCF/FSaKzxVRRIev/TVSdX2XRTmEEn+jZVRGHBpKqhs
xTIL4tQXYyIgIerOE6lu712/TJMEd4c4ehRwvnvY2eej7mOwkof1/89SVPw6K5ji8xPDHBuoG4Hl
sCs49nnefc9eMITJvTy9LPfUHzx/3uNXcqPU2ndfXpmWaVYA56dg8BM7lHEUJP+LOOQoMDWLqawX
v0/asWuGMFoM0sJnV4ogTDEj2sYqEvXD5IaU7yvz21bPS0o9v1BY96VY7oQvuu8m22LkFXJkb5PF
Q8KAvjqBPVwSrLBZS+8YKveyKta28jENDpdZBXR2Jj1iE48FcyGCctkDABEpJoajOvgTth3ssOAe
+Gtj8eJMTUbHNgvJASm+5S1AkXZOGeX3nou6qYxGfww6Gd+noeafg9Snl0CtfReTXNpOEavPAsLp
EztOYp45GQGIc9HO9O6iuhz2IAH/nwR4Gh5B3Fb9L2jKs1Z5gAqb2bHVzZyW11O+i9sPpGYbetx1
yzOJIElWCsWpVB2T0sT5r3drp/XMbr5xm9EPpq2FhHXlXzUaBMf6QRk4AgcrR/xp+WRRuRwkOzLj
hf+1z9rmPCkOFvc0+ZIupYDYN+uQjDVibw+1tjiSwEwFwpa0QTD9OA1w4pEeT4ddcncbPWkAz3vb
Vy6PAOQjXs8CsO0nsCbUgl/3MqpO4gra3KhsqB5bO80bw6gPw3+nMCStKrCi8g5CD0cQp+sxo86h
JM9YFXx4S7RO0jm2gTJX4eTpNrW2RhBTrKBP3Ljiqur+Mb1sksGgyEnBSQABEnTrrydGPNvh+SRQ
4Oq4zI/XnIETnaozzYSAa1vPaCE/ayprENL6uqAKgodaHOdqQMN9FfKmYtwIke75bkUet2kgDJFD
29eSKwTnr4sqQxXje5KnLS1/x0cLPaC5KDCjE83Lf6zToYgGfKj8BouDW0EqNC7/jJj+k85+aMTd
InyNHAm4f1UBQ2qhg/NPh6K9vLxcYvsYMbWgQLggBflbW803w6IhhcZ9rmfhPpnFEgTyLmfSUQcO
/1bPKenPaibZ7ny7QvTZ99NO83jvWs8qzPcdebVdZn9x9C/rh9KhlCjb5YqKSt2DrNXkgFTo+uQR
bUkBf/X7be2CAOVDcEaiVEnzn0QmtKXg5sO5HYfqG0gykhMeQEH3bqv/acBHDHv455c/9syQ+pBT
d380q7i9GR64xyvZmvui64Odcm0+msSJ8gUsDbBSBNj2UkOXWVycX7mNE/I0nYRT0px4sYgli9E1
ArT1ad4PNQnCgSbu3YWyACHibcAne7ef7gU65Bp9b08baboekl1cdHiw6/73Wy9Ke8z0YsJvpzWq
0dT5jAtAsHTrnfmTIYImxcwVa5UucuYTiogVF7hhcZGw1QK7LM/91GxGhtdb6lYN7ohyWLJEsTkC
qslIyI3mBTZMJSwBlnHeOO43j3AkHXVs9LmxKeh0tmzCsz/aziIfqf+gy0nRV/MXhqsqJFzIuHLl
6Eh+Mr3/H6ScP2aK0VxyVlmz6yUTXfr7KKW5G5bCaxwe33p9zstJPPUk/A2eBsVdBzW2qqOIHAtl
HpmThKX0JiBZx/qGO+zm+XllZ1iTWUKj7a+vVsL7oqkeSpPTWfGZjLVUzwyoKhR2edkKQCWvlBLq
MFlG/lAqh7Z9OIf8Pxs+cBwqLMKRxZiLZmv1WMlUXo8KU6BwNiT1pHehPQ8ny3pjd36EC+kASuYI
4qCzZ0FZD+d+p0hYxldKKyYat2ne/dSrcTmFTGueFB+UiwM/siD2c/QWxh8gjiDsxUCPiipKANhR
rEx9VeAwRXE80H0FCo3ia/m8qWFcR5202nYS7jisyYavdWPtVj3JRtloGkQXsVuO8QR9e7OEsDBC
ZyXe3RqcokbeKk53s9LdoosctSAKzoJi8xd/tgBx29FXeuoe2C5SFr7KVl/pbwM4c7ySnIwowLUP
4LVk/Y2IoBe18V4uw+B8wl7GWoKsCDU6dfPqlimv2CSWqPIp0BCGTmm2m54Pxkg9B/hxrQ8ME5Mw
OJrHnXETpbwLRl3QgtKvWbdQrIYSh6gas206+l+f0GDNva6p2dOYANdoTZ7kowIXrRjOFs+ziMTP
traUIrbPZlYCYztP20tLxEeG3hDtNxmqzBdrBAKAmc6sYMZpXmjWP0kPM4ySsbQid96uPoyBMfrK
Py/7lWVs9fC/ZWcjcc9aykXE+95xXVWewFRzFSusYUtJutRoNNJD0q9HXGdwWRkiEWrPC+9kosQn
4N0bs4gRP48OD2A+VDruf1HWxlI2j01dSoK55AbIWg+5uqdsPFoelLYaqJ4OcO5M9yjeV1fq2Fq4
Vti9aRq7mIuM+uMcpA6RQFxgdSLWmyFDbNc9rvX12RbX7apm6ASTKznEyIAJ8Lfns4QXD7SPOc92
sZ1JErqK43tbsPSmsed4kQbaVVmlqDr8GWcFCQHBxA6RKi1q10dT0DuNfiAx5vLO41S7hzJsJxf/
+LCjFIM6XixF8q1UyzzzxXzuyi82ogKYCUdtcjOMrX8xhbM772JPPEw0ZLQq92Fgebpt21RucoX3
R8hxOPYJiQ/bEjvtNSSoVqOzHHMjU5gWkE/q7ZkJqAdJj7Lo63Umh7ZogkCJ5dZtvrab/VVnbBTu
Y4blQ7uBVfXzVQngDR2wa6t8iBLFmFpzQ68XvkvIMEaNnQmYZFSPzxU//XdZuTktpSqGt024GMUA
W863ieqklpeMpWLTPvHXfpsymXYdV6fzJiq8DTxMkEk1WEzkQfZHl9KLMiHKJHnv3ynavGpHGHcd
0zqwDXUmhOD9A5zqAL7Umqk7cP3R6GWQ30k/hZjy/sszWwrfXfjsxjnnSF6uyhWRbm0FGk3VVvEr
dNoHetVg4Z8jL7WKaj43O5Yd+lp8C83mGhErRF8+pw2QN5P2nj3U2GiVPFq8CZCG5HxkNixpywpC
AQcSfrc0bXz8dHVSxQQFk1T90rLYj+vWZLeV+OsY2cFqMZ3nlgZpJfX1qpfOnqpeMkQv4tSoL89P
QDaz8adlcZAku9a230BWY41e7t4y24lOF3FK/xA+7Q344xRJVcw/XVK4dylydrbhbET635KNxg9a
awZLn6zOFDDTe0uWzutNVjejCDrKOZaEer03twFmVgX3Md6oLqATRrysR7M4kSqMPv4n1efPiXme
bIvY9QapKK0nH766m4L6TDh5INZ81eh7Wxtjpc3oQ3UXfsZJlVjuq8lTOVtLtKyUyIzEG2gJWPpT
BT8x6ltEAfmaYkl5dNjIdkwVKCTIG/zDQUqHirdc8nNdfmBlNEUDgfmnqRpNvYUejkmJckWmvlgX
Er1PBS5deyREEOqeXmsrP+S3WDXMN5DOYxYhyB3a9ZTe4+3mFTh2aqQ7sqEQgGH/sAra2iFDemG3
URO8ZC9dncf+7mVQHHhdoWqhC7aQ8C8XsOWnRoG3qpbRGObJkBOwsIx/jGRrtzM0UE0JW6bXv1ef
nxhPhSQwftt7OJK6rLjZMEFuJ9Wo+QLZGh/lqXttQ1Q6FkHOihay+dwf0xk72A7AtviMMJuuwkmp
Mql5dSKQRA9fH6Tt9qvjuvVTUyG8wenl1+WmadCZXaXCFPahjFKbaQ4YnTYi2ZrOTAIz0OThEsl8
GD4b5sbC1aWQmOJsJN0fb+3lx+9bI3F48nlsNsvPv1PDcAkpfXS7INkulix3fFArlnNNizC50qAK
Ff5YEpvUfdtCu+2JIfHfd6FNo9f6+X+23z2QgvyTcwhjoadN0yPgZNV/HN+WsQo8dSlGYTEqjsNi
kJuXvbN/vtyZLw/6Ghq9KBflhrBgtRzIgvNU/Jpj8UEiqHysi5jLYuRZFOH8yJxX7ell9WabFNfL
wN5q9pn9jAgFj5rxLeEr8e+rznAD6Q2aBQySSuRBcy+Y00cY+Hmh+1faPzoGwD5ikC7F5WMggs5N
/AosN+kyMIuMyZ+w6ODlJOayeQ1pphvQ/1y1/WJ4CZZHuEBM9jHXT2TthZ9/DfJKGQRHdaBYtn9N
rOiH9f39+65XQNHsPRu1Dq5qYxJoJ76ukimKIFPaWJelxFI6Op9pgagSXfM4tyD1XCczF0b+sJ7W
9dFH99X8C/i+BEq7VqOpyLvQaQZNKnRM/0TNrwlbW8DqNJ+nKNMUtMkHQ3fhp/lI6/jq+GwgQc5P
hhKmzceieXNeZbotR9v0g36q0XEyYGTKF90r2vy3Qp/cdEgE700Lx3fd++W6X7kMvQSDhOLsuXff
JsknkVIfn3z9aEeb3iNndZESZ3ZuBklk4WW11nV+so1qMm7hMu1U7AQcmGrQQ2q1W2jxU/5e/2O0
oMYT2ZtJ8/XKn+gVnzL0TvfP0TElaqPHl+GHMRdn3xcPP0Np2Diu3wfhVJSHXO/Am/08gF5ZssRq
/6lf6ISQdvL7Sz61O3MT4SibmQPe66uW8ibunV9Uj3lVcMtBGkwyrCMr/BfgfAp4HKyXifQX069d
6EnLn9i8W6qoN9UvSlOQhzWI4BbcHJpsrAjZH+9VdTcKdvuMzCCLdQ3zr3KPogH9/GdipeuLbg8J
YOah3pe1YFcKgYthL6fZxq4O5jQ/FWZ/uxWUz1No/mtFGzb4PY6WQXS2Y06e5R5m/YdDCJSB1R9R
TPDXh/z0nzT4K7i+Y4xE02R9N62PLEYWTm1BmVT5G1Sv94rOvmme0Y0AEr/557QqMeQpUwlNh0XP
FtoA/AkcC8f+nWZSIXsLDooanaZZ6MMMr4nZ3mxHMoRzgWNoofvHOG2+SdZ1OkkwKUKXuk1u+z/4
AgrDGrZifUEpsyqS/uMABaiSRTVq6+zOAgQoqnNsb+go5Ik8inzQE0UkWnJ+U3A5VyjLaPG9aSiv
W2gTF0AX0PrQPMKN45L4dHZERw5honw+ab3PRQVJ+0yDMjFT+QI2bsfpl3qm0yEfzNCpYQu7M81u
a9Ix2ArQipRUK/qFLW71JScHLrA3He2+Z/pxq5iv/MSZdP9sZH61FQX1Q07ytuanbbw4zNoat4Ag
D8ZUUJtyLlTY1OL8kZXvMRSJjvN9XSNTSTlglsGLpBB994pMPhN7foW//Eo7kkhf9wpxaG/Bwy+R
Gb2urqudE89O0CJAue5jkq2oAvAK1tbPl8QJ6MoleGa0R7fCJyiK5OCy37LvujoLa5pI+ognO8C2
AEq2OFf2yWN8LX2JrT0zbPHMJifksipRC7jqa55SmjvTtJWAjKXcsAIIfLbEQeV08lmlRHGT+/4w
8FQb3LeuiSOR0bQcbzNOsgErYiHk3d32whrfEJzz6ylPoQ2eTpV9Ar5a+5wgfL+NHyCO6cE6Mc/k
7jKAL1zGMfS3TF+oqxfSfTBBewxq59zcSbf1spyA8fN4BYR0QBl94hLL0UgSoRA4nIjj7Mmn4nW2
AwyRCg51yC+xOmFDp3HJbY512M7wU3PPb6kcJhs5QLzj5XSEuiBlE+Yg8VSgI+gP2t3LXLuBy4jN
Hh2oeipOgjqI3LhB3Q96eOdGo57uBWBa0ZaZn+IJj4jqzoG4OMJRyn+lTj8jzpRGikd/F9XntA4r
4xFgWvoTaOX71vZf6htDHNOEUZFi5fGeQ70uCWWRTaPsPkWoC2hsnyalTmiEIk6kXTOkE2sXQpZY
wCMnG+M19tAnqROoRMvx4Z37Ec8cXS05u8x3h24y7oWzaMacP+A9pnwRpQ+OxIihlaV1mkYRi/q7
ydMg0tekpRFhYIohCLSZlV93C//PZ4UmsDXGoF40qtbDjFsCASKk/kA5VzLqtdp3r83DdcXwMOar
BIckwQTvb0B7fZOW9TJs8nghOK0A01k3+vDB/fIr+oJN7dmFVuSIEGSBjvzRcOB/UyOxhbHFP7ML
Cv4/VfO+jsmi/sgoBvwQ+NkPH7WcbZmwzRvd0scLcgJOcBQvmzxSIIzarIvEggpxSrzo+LOrxAKt
g41dcuoIYso4Z+LTQ65yvRc7j3z8LOEUIQ6nG3Hjg/A7pNBIMVduuDCGuOkhsZFFHJltxRfTbsSa
DSyx0w0QjYfVhKl9HUTV2czhcx3LCLV7P6l2hUzZS3ZZcH9wtsQVR4URu0f1CgCJatIRP8YQNguC
B8QD0EKJPmSsLwxrzj+QTiG5f3nBzVy/l7ffG4hmLKrl7JN9F1AjcAQoit6SbZU3ZH3ZOzc6RdHN
H0gUzHzYXvNvU3FbFHhiVCxIvNar0yIvv9XwGX68+b4BKC8SqhVbHUpyxv77W6HO2b/bWzZPn8e/
tZpmPIz9cx4qnybxs5RGfjNai7veJcJXAujTm5eZNt+C16p3rk59EOP4KUEv9fNzzPO8kamKLNwB
1sL62cih+A5xFu/bhRsPsA60+bxwrrHY1sw/VQ7jIPUATWj3OTDUw898FJIbHr1G9HMfxDjF184Z
hadwu63/JbvAu56XMUW7T3jT5PghBHIlTUtejFjI4enkVH2RIYWfGxkc3cu7FgMMreFOT4/ooriH
OtmLZ/NLVW4mtTbZyJhspNxNZBOWmQ+7UJtjG3h3OeN8xt0t5zFfLVFsk/r4b7M+oNhWv4NsFJNy
OVc3dSd/B7bbHoHwVRcga2DFyftVoqK+Y/daphFj9ZyPBtVFwP3Q+rrWwauvBx4XeNk/IW4ytyH5
jLOjlZzGvvD0qGAYihNu0PnT4/3M2bHRmr8Zvd9jXGblca2aObXAWsi9OFdnJ1ms5ab9f9JRwCFw
1y9YrsA5n30bcs5F8bhHApfEvQOc54zL5DVWn74SWxSrizxR3ETuTR199O4cXLWwx1FQi8aXS5P0
nTrQGzwwPN3u97x7aLofffRfe7DD1BQDeDlwtem2rH3Fu9Xrt7oJ4/knPKpirHhrxfuEVRKPwAvB
PY+E/x/3pI1Vf+TDhP3VNe9brfqh2lVmHGRU+va5nZ9PjkasPveVKPDWw6S4dQpJXUDtxEDSlICR
+QOaDmf0KK5JLNpt1e/ucDMUz/vfGhHRxde980jrbq4HtEdrX4uk+c25CCD/NGMs50MGTxIhJRA8
WmUHkb3FKAeEC69dJ1U7/NBcx3KezaHesE86bHEqrUtohHeTjRU3fpDXFEY7knXHIRzyLbTuRQY8
F9ZbnAJGT8b1KtlATASXGbAOfxMilW/H+mxWq0ygvcUlRSp/siDEztmNqAInc43xNOiWH9iuGM5g
cnHi7IfLP109cF4o1GSh7GDu7jZVghCXfQdckL4MmKrYq8NTxqOvtJJgPpkqpxcKAbr4v6ZSktup
LfoJc+nGU++XXtuMU1PHKhL3Ugx6DHc2U65Xhkx7KZBSVC+L9ItZ30UP/P3GlWEzM6b2EKguleci
PRVXA4rVWTlV9LU1Bpl9dTXRE2ZQ5x8vVvhacmKUddsGWmZ35I4uZI+UT83K8JJduoN1CtFzEYw8
bjY3WD8NKZW4yhVtm2vp7lIvp42LPkLDN+fe7S7vCNwjhsmgXq+sAEOEMDKyfrPH9pUtnTeSRi5X
/TER9XzN+JhDzmYYrHB5Ehtj5JbluZ02dbwTgQjv0SnmfeGgaHZaqIwHqpf6NjY3XXz+ahUZJ5Lh
0PW2Vx3X/0NIsus4bEi4+ct2WA2Eq2FyyppP2oHb5fSSdQfYH8FQ7MfQmpwAyIn5yCFT648TUNg7
/fWZFoicyRM12FFzf2fHLQTP8J3oDiMJYEjxpPl4Z7EpM02N4yKcPD/cGz6lSZCCWGaLn0EfxjJE
tAUvL018cYRRWOyl5zEijasTkX54sjHstXTUQFLrSPgQG/JkbWY6gdX1THJmotQnO5t3jrX+3f+I
0F8pq3Q9xvafr+dDGfbsFAS6E40QyhyxLPukuFheLPGa0hplorj3rPbPQlMh8FbJfb2auc1PLTbK
CVmkhqGE2ypBTd5qYrf113ukmLYrKHxuTx6AJz7lvv+Tq6+7QqGA78LuwB+A/nu9dwjM0a4lGSrH
DMsQ9xS0FdFR/u0+gP3bvfF6q7VFV5fm042DAGPbvxwDyX7jkmcmFziBtbFRZbdlwlzuHu1ZnslG
peJ9sDj82p2zOF685byBeo/w7VIthh1p12pjFzyVojo8DFXWmsY52TOG/Le5auMHY9WHRuYvLSd+
/8XANdkJ8vuGUB5kjZx28kJCzOl4pjFHady8pKI4hCGi5ObRwOy8+8FWUlnJ0Ep22IKP+WHKyhkm
KgBcV5eFi2cgR/LNJ83IwxFXbvdsDYm7hjC1Ky8flVBxA49KYn21ZUmjLIsIaqRh68ZYWWpma6hf
mFY8PoZk3nnh5zUt/ugFWKNgm78wfHLzLsx9PKhVpJZmK3jxmtkCmlsodW0IEx6sR3c3si19aBFY
aCrxy6bkoh/iROWIYqsxYVtCKYwWwcfS77lddT5rMweYc3b/ibZXj6OSTn8skLGuxG1KvKM1SmJW
Q5Q7zbgWpJIcDQHLIQv2jZBwb1O8envKmSVqiNqJRf9M1OtvK8WAlLlMS81gJtoojT0Mc6ROC3cy
dEPs2doM8yCBHMm17eMrfUQY5tuCA1G/2P/f8PfzP2SLOp5JqAnka5rbWZ54La74XFvH3i6TOf+s
JgDl2+Pf3px7cAymYKPIhCZGMY/wsMowML0YTC5D49WFpdkgrOzlhIowSNMDzvJKOo1STQLu9ZfX
VwIXmFbB7R+zjLyFi7GS+ViOtzr7GXZEz/04v1Y7toeWTKzt0XWlbg+s0b3IwrwJZW6bSXi1j+Wa
4cQnsYdVS5ufXqxnpFBPK6XYpKnSfxdPKndLLZ3iijggDzm0wYj0ShXSBtDvnjmJTROeweAdAMcP
QrXI+0P/xieU1qc8Lk8EqrgdFT04qX0xx9QTVGBYhKcVneM1rqIR/DUJo7PC+E+kroeWnVu5nugJ
nb6T+gWJU3s5yeowDd6lBOEb6CAly53A/mZCrOu6CcNqavvUBb2JluOffIUrdO/gz/JmhnAx29ni
eOKHTxaoYW0OR6QqHBi6LT/rmNFOT6jbI0B9tTedb8s31uKipdTZLXUTaf4HC+WmMssQ65LVTt2d
Oq63JL+wTvc5tR6hhdGyV0oBuEYSfM88wuNhWXvtCWqSbInESTY17GN/3Gcyoqo8HCj9rdtSlChk
xVSxaUBfkg2TsCwJp7ourDCgoZYtpRw738Dw+kTkRP8oYfFgLMu9X1P/nrTtLQbWn8ZFSNDJ6f7u
JlESWASY5IMtI9d+nYKLIoFxQLEpNQ2bRtgFDrsqhwE20+cSWbQcRtzMdR1FSXGPpjaDlUVxXbZR
sAPTjYtu/2CX4QbE+qRxhJUzKdHG9u9ateEp6chTN//8LJ1X5Atx+Btex0XVS9fyZAcxXAQfRGUv
1E7BJDIcWdnWU94zeOuz2WTI3zrseorC3bjJmuZjUILUEyBicLcXa4OVKNBfHLqyQIPQYizoyDR2
SEfetKgj8VzYqnSFDzbiBtqlAb0HiMQq8V1RDYdoynLPmq2siPixU5avdUPmOuHCCqCjOTY0Sa+d
5Qj2pWw+lWYYmIFBhOHQ3BJHPw2LvBZSEt0qCD3+OEzUfhSSnn4YRbFdiujvC1NrnDqP7lF6OHM2
7a2SunAAcO8dHbv0lSxNGdzfLDDBU0V3t8LO27N1pyhpL1sDmersvlK1d/IPrmyto7tUJWIskxMK
lGTbpv79hO1T7WVV+3z47xMtXHjq21GmGLeTZOutsyR2tPfuh7DwhoxWENwsXCwrlBK0w19aHgEd
l2UbJ4ZG4RaKXEFgSoHHvQi1+egEcMTj4U+4UcpNfNuWp+xDhYX2G/p/NT4sdz44bc0Hgl6nz5Fl
VveA00lftTW59EVAnQ0vVKMZFBVaHHPWFzi5XZ20NeDMAKl0lmHlZtE27aqdVVnsQKVFo5A5iJ9r
gNLuyY7v5Nj4xt7/P4b4Tlh/fyWxz5QpldYFDL/yuTjpMpNESTdEFxD26hGQWyhtRtm1106fHQlZ
f990RQ9+T0l9wUSBGsoxZA2bFYjcFmoeX1zRZndMCJ0rcgz44ScyW1QRRpifTNzKslPScOV0NEqV
zNLP1V8S4v9dMHIORa5zZPHvT9q3Ova1VFYpIbWHhq7rim/JG9ic+7cDJrV89+kp4hhOxSXrld+j
XO6uuYH3WwnykgfDd3IxizsFrwwgjoPcR7LrCrLYjUEUXD0gT/EzQYPQrD1xHYoaYi0ff0lqQMzM
i3YdOhj6M0UjRk8EREyvqeZ43LpifOBzfgjEjCjHzmDQj1Pl8Cpp1s7sBtf1qJ6nJcy4lXuaFffY
NtIFSFUCnIxOfUaTosPn+doaXs9U6nixwjg/ucDQjAEPifvHTlktInrXCwJAB4bpBPduvXsxV8mS
D+DEmW7+eFcof9+1Q0ifzO0OTlo0i4cAE3TZcD+9/xVk3pN0MMNidYzSAbZuVGoMBDDVH1CTM/Va
90UH25hDs0M8zcuygwqFOzcx3fPF+bW5HN3X3bZ88zuJ1ClFHpGY67XQFleePHAjVYtX1Qs7+ZqN
39b79OAcADlFysNPB/eC9uIhtgnAR2M1DHOPJWjdeImzTMXtpEmU752q5dOrnFFA9hn/XFUwvGTI
WrvwbqxR37ADMeRRts241sfCJUGFHBlUEC658AMS0ym+tJTWW+Uh/quyWJYfnyOqLMRmj5ZKFcUJ
xTAIVxFbmzBCi/V98XJA5q7MbpkWnJIxv3aKj2+FQD0i0Bk6X3Cr06CPB5RmXOi7NoOyyOjrSol/
VNQpDA+K95AGVdcTy5ljozcn/W+AyvOBK1gqJRwRniPuUsalzZpzqqKndDciLqt9yfqmM2J9TbHh
HsoeJSO3osGuj4jUfU4z95DlzzZgiTgasfTFZAPO1UGeb4bUvKwnvX4aP41nu/RXshdW1bqOk9VQ
+zxw7jvE3m7mDfIzM50f/Iv48NHXSoBdVj8d0GST6svJynjkc3OxEL5kq0tiozQynU5hXSjlnrlM
82ogYCGmys0By54ND3BYLfZ01OTVBZq99Do2xyP0RLDP939pxh8I4A/DzPUyO0odAjB+zikpMq3L
A0bL2rp9ZHgzl8ye1J/Z4JlWT6sYFhdPGYl1AGqKCK5CTVFQbt2OwxYt1qCYBWkwkhpBPjAMQnI0
p4fY/r1VeIUmiBQsqJwkSEDfX53hsFUG50n1c1OahFj24wjV+wHUy0yFY0MYKdgisTMsZPhkSX0e
pZn+JumNahO1NhpxrkhgtUKO+NzxVvlLdzagVWEccCrY0mTp3FyiIuSxRrHY69+qUle1UAFbMdlg
ivtrKpw0LWUySeUgJsyT7KPJeXtxZhFUvxkFGixeKY5LaT74zQ6hljTjhBU3ye9fD6gMzwvDeIkp
vgcvg7m/rDQytGQajJtasfslwIfBJbdxPoffFVtfBHbaienNN6XKrJdrBaXih3PomTB/PzaGW/R0
9y4bDenpbY084+jgGriGrN9nk163rGYC5RzwQ2aaJitWpKcVcacD4DI7vlUB4unDlF/mG6b8LdeK
3sG+Uxhr1w8ugeVcT3U0KtOZlM+1Gf5vZjfEASD9m7sUbRvnu4c8loNNTgc1ayuKo++tV4k6dBLQ
h9OL/Abp6rqTzJ2YD4XSN92eZwnhld7sryCBTG0pZj5Cm/rSzo13SN1DzzWKW+zuwAkBey3xNx0h
IZ44gG0ouXBvxuyFKgrp+AzHUD63qJajGbRMLsjZlBnPuFG2y/FfIJJzYz6YFxyjXQ6Ndtxr34o4
2S7FVO5zCbBGEr69TNwikfmzWEpvDGjmdv56bC7o9UgfBjIcitCaLmccmqiuCKwIWFXGq+RzU0GH
86O1x3KbdtHfJNN6LoJlK91pXDETyZWSsc/wRdvMkLg2G0e951lsKCKkON88Mpi6UBIqLb3LMRQk
TLXSNNn+811qKrnE/7/INlW274eIQp6Kd8kiAh72QaU+ga48ce1LmMW7x9GEs0WT5YlKaZvfGULG
jwfF2GHkfr15GqhZVQ4JCD+4gPLlKBlxPI7KMKK3aXfvb501zWlvtl+WUlHtU+Ivk5PfdVn880nc
qCRCMlJ5eTaoEX76pexhZHFicaeIh/UY5QLkE83MZ1S3Mz8I2ghiMqUnaV4UE9O7LPPNubhLOZSv
h3aNn2U9SUcv/Ft997/1FLKrb3cw/4iPwspVyTupdEaBPDWx7Ltw2SxN7Xz63wqOVLp1BVxvH39L
ixHn/EtOHPZzEexpY86EMiizW8wIUVJdxAQeFxSWnwSyJRC+VUYku8Uj9gdkJLm7T/sOa1m3RxID
TUuOoWXKgCZjpgOQS0s7BLd0S7yriA34m1uiTVNxfx/XfeUiOrEGiRzNeC3OeQXf57Msf9vfxFUm
zKUQm5PBsdnkKgH0VLsU4Vf6uFQnCeM3uxpi4ZhRlHdq8ZYjQPbVlrAeZeZ8Z1A5WT8FrRcfQExq
qZUCS8qBghcsctGy0gKlQFUq1uRgTwfjlMhi+QkhP/SwRuOwxgKNM6dUapnSYLoeqBInwpf3cWVS
PVi0jfmSStUEeDUnI2rMGLUvMFItRc2l6Ib+W4C7lG++Thy0IOlItAiJZU90TgHTuYa8JB5ORlp6
cGEcVm//uanBWc+1OVmCaAEvdAQO303KJhfp5XFmoudmH5ShyRM4cEYUVAIbSXtI31RkiE8N7hdw
Y7lXS7U37cJxgl2tWumF67LbcYLPlkYPQZmJHA05iDu/PEiTUur9PeQAUdGJx70FcTE5PXfuDx+2
10ZjDOYGgGDkZhecV8JUmy+tCJNzwlHK6Ri9q82RP9B/Z5nS8e6MkjQH1Q9UqSEVnkz3e4/Aupxv
uiE7VtziKQVWG6W7nvoGtT8/oVkMnedNcV0lk5tZLKlIE5PAUbyjMxcDwUxvqt402n9JO5YQ+4z/
GSeK8wskZsur1RnoiWRQWw6/qkWgob1umkQ19oNfIn372HoHZuo5lnxoRJfx/kc5aTI61pHEMcPU
CoR5O2cZDY8YugOZJ68LDjQ1ZUKHdCCCUOuIvM3Tt+r2bTyx+lUSsdOZZQkSUelQz1I7bOBWtPEm
nycnJt/7jdoP4ZEAYYiB5P7TvWjSO6eca8jY+K4cXu23aQQ4WFiZH5pHJLmN7tvBAvXcD204pXa2
SXvkytbSXR8FjG2cYqQpSG+kQvyTccpMS2QYrvbEu+zNFm0uLdCg8C85DtoL8smDT6XM34u5ZzK2
Tji81DMM4E85Bea5hGlpRGIBP8foYmESsZuECUVzyNPL+rWyZpXl/1kT070AzinWBiF0FBcpQwx6
7D/eMAjw6b44mtgqdIVxPz+fHQ12McJEHnF5m5K1Mpce50yp+79Ur1nArrtU3HsQlb/S0ULK3Y3J
KMmO9NRbN1iZrMJ62u+IA4nbxB7RQ47kr9R8QOpu5jSA3fIIRTmOq12LSCrAcLA8vPCGEU310X+F
XAWEqP+uFKPUo8nP3Zuz/T4TaGIHR3ABra7nG0uEW6yEyZM3Fz8oWY/k/KNTcjyOrJtzE7TCyyoh
EUp5kYx1GqBCh9jYeML84QXkRHUCgX2dTKpj1zrbw/28PU9mlLM3mKfz8SNV/p9KIJbbaHKXl2QB
HgEs0oFxLunXeiumJK+nTDBi0eBeZ3VKglXw3BjNvn6FFqrAXwE/ByWV4ZS2+FcKtkRM1jpS9jcs
Lf4fYtb8jpM1HkgulvrVURLjSYLgPNGZknG/IA2OIo1FCnOj4bku6BeGtuqHKOA3pBJwyWwJvbVB
wceC+GzBUstYaXwGthNLgdmnWOxeT7l7Y/ijQbFHQBdmVwnfnx0w8N/TnkPFh9ZKo0Z1KvCpLw+f
zTP+vZ6zLgGmrJDJrK+kgevFBvAmxLNbvdR3LFkK89UXFSwxxi6XWmhtHZ0gUTi99h6vSLRiNdFK
TrkhgV/ExaVb78iTOfwKuz36YZZp0OJeaOdD64Abun2eBJc/KwR2RNf3WEp3GP7pXSGoAAQtZ3mQ
qQehkPTxwjk7r/b962iY4CoiQMloM7GugTbCsX4PIqGSwxGo3NDziru2T3c3HmoKqpngHWmNH33Q
Ilhhox937StuANpGy9VJg8eDEti0WbtVN5IvBFippFhptwMjZjxNrVMXV4OLNB0vPTOnOownhZQU
yPykn9sIQY5JC2J8jmEV2lBw9YxMPhj3VOrM45d3OKypvuLLWaLfJCJid+E6D8JldD6wnZCCpn3v
Wyy34kLd6I70g1lvruXB9ei6U1NXiiIvKEasHWJ7vCtQOcBL66d1jXad9sULPSQQNkmQQ7jnN3Yb
Jcbbpmmn0w0BGozTwm0QwFNJm8d8nuU8mODgirV8ewnIepCSxNZ8uNvkWr7sWbE9XPAEY09m4n2t
X/iO546mC1gqhRZXYASCd+u05TLbRxeCKWPxVXAcuvmzJFzBHMuMCSx7H/Dtv4tK/brZ/CTv7hfG
jRsZzlxPxLb4U6YUhzMyjMyA87FjLRGC0lkI9F1hvNxxB7W7/EUK1j9z6O4KzJ8Ns9tq4Mq0jft1
SxZY7dOgz7VGO9Gs22/1w0VBlb0b7i48a3yQnyMEIWZI2JabNAdQIMXdLbZgOGLCvJ88EH/+Urhz
Ia51mR8il+VonhJktmjlqQXhSFMLi+j18UcJu5OJz+rPTOrYZX5yqP/iqv+BvpS4p1cIi/7FGdCj
Jt3mkOgXtzSJGNVoLglvwlFCAX2IPnXuySOkSEpJfUy+uKFSmNf3EQFdwgJAvdAy8LjyTWGnwLzG
sJaGLEtpk7it3CT5WjwqzIS0VpPyhZVIYynOAy3F8z1t/hPwDBi5leXbc6I1qhQHKM2/msk0vacA
x6j+vgNBopZpno7vQmKnT6pQxhmUfbYiWeAEFwJL49LOe32Q9wSdF3ltarj+/kopr+M3yrTpXrjD
YhPhRMuQIfbpRTRRh93aAUXrHQAIQOhP+6+HOR2xNdfjKZ9ZLJdXpzwCC4uhCiatd5q2P/shDRuN
oS83LMrewgA8G8YYepifxXAdQcspDMgP2aek6gmlzILiAP6XLiEHBtco2ErqBPqg33/zM+Br2s+I
FMkzkxvslPVXwx3ySrwB6XbF/zNBJIKdaPUpR1cVd0uzl406hQ2PEsXtHEXAREmmsmehNx9MDCCn
5s4FWz8M5cLzzMegVjPSD6aqSijQ+uI6j14he7BXyqnVUNXNxT+tmmyw8q0R1VJkLNezapeAtMJy
1lZNeZPG233rm4XOjUtdtwas3uVip2+7cXn+SExoDZcbNSQht6s/u7DANtoxxRyXgtLtqmtbX2Uk
xjfwiorD+3ZdZpyUVvBRx8SuU4Zv/CcY2cp0UOuKEsba5feq2mn3Nv9Pan1aaRDTI+uDq5dL05QJ
zJGTwX9v9UurJIRSQskIN95P45w0kzkYSEOy+x5oK4tw3Kf6mJ9sTtTQayhfMSMlfftPo7A4Ld+R
cWBGQxVhlmbYD6RcW1uQTV5bhWOZWrDS3ClA5w83CLmH9qfvMlJGARnwtXh1T7glsOQ5MuB6GWeL
/Su24CYnck6/NSbX1ytXBv+A13zUN1Zs7wCmjuN1JFZM/nxKp5VUHUeLnHViDZlvVLF4KfSVBNhn
Mw/v5MpFw9RDCXrdC7wqJfouaFiPUK+KcWeuBFFSMBoB2Z8FHibhlkNa+OTuZK8tGs+veVyM8QLx
QxZzc5MT4oeeshUtwI2rwlUWYGDzJsvFl1YDP4qoQTDh0Pkd3VMJNE0UUlgyuSNFTBhAlb4BLN13
/s0bXzRINwBWXpHpPrz721d37owoMpSnjqm+dG7p/FSFOPx/BSwCWxHprqPPFt1QjfaaiDdJ2tu/
zxKK4B50XJyP3nS0UqrT3qbFmkewv+OdYzPi3gCK0ZxaADwKs9D3ilBIEBKw/oK3Cfpa/UhFFIE3
EK8kRNmO8aNQmXfCdIso0Ai2OHR21Z923svpWVj3m1OYezHN9i01VgnWp+gV5cpE/3b/YSkyFbyt
iMrUH52eNwBP2bUJ/26k2pbnKW1BaDtptcbUAym7DMJg0mhZ9aFayC8DBfeAH01r7DB/gfDpqU5U
c9WhHfoiYNRjHEC0HIHsyDEqpt43CbsIjsgNNMgBNLjjZ17ekR2r06ktEKSzrRE7ifhIz7qseRfN
ih3ciLj/tErs4Fiw4WT57IJDY1ugnwqmJJowaCd8KvzXC+3QyGhDNpnXzr9Ezx10L092mt8o0TeL
kCMSUSIoe1ZlhmhpPuUDlNzFDKyFNVyOOEccTUpqOPB2x+SbVM84gSFSyV6BDsMR2uubK+ArFCH1
z4yXpr97ZXRQTDQ0wI9d6dFhnLi2d3is2K+4Ck786i5w62HmU272pVC7sBx3hQjKfoOYTrE2yxui
t0DWDuQJlyjHoGC9McBucqls6iJwja3vZ3XxBPBknZapYN2OcjVMv9z4XZwSvw51wiXurbR7KY8e
NG+buf8W58gS6Wx/e8ooKjYA+2w0vmwbjjnqlwo+JHJQLqRAnpqXfz3g9WaVEdK5Oz8RQ2jxK8PE
e6RLHKt9wK7iJNxYKip5THzFdc+br7WbehWoFkRan1RU2IuFtFppODGwEBkMWu6vFFkE2ZMOqo6h
NCUuVaeLjBaQk3EG4mX6LfJH/7DeqTzaA7yDowTRUbMmQ+k7pBGKfhsDClgO8gkQ66V4QmAua5NV
P3WLkVE92kcIXkKa88PujSUziIZOD/A4V70CCScKVuiIqw371NYuQY6tAhL3kHndrKqqKjv5P6EY
Cb5a8XFlSPaO899iDv4I7ZfVmAF2wRTbaHMb/cDo/StqBw6d0VJf/ClfCLrcjdCnAR9U/rHXAiR0
BuFMzmRzvmljWDZd6oK3VJ3A1xZk3F+RGsnMmPc9ehmkpbwQiok3lR3jpHVVhne3sWF6GvpuN1G8
INI/yo4XBocQjZLhl4RYlyrMivQ9ZqAeyoPavZDLytmAZIZ417J/PtXTrk5tV0oOTGaStqC20irS
3/d/9DkP7hRglEDwBQjOMxig01ls0j0REDvWtCeZki2A76s1M9JupBR2Pg1noVtGefmrJPmBJXDY
df9XFtT2NHzWzeoxrZaRwBSkWIa0vjLr3NKckxjuBCqxndq2hFxUYv+WBlaZ0BLWnlbCCNfOmc9y
8E4g/BVRaTktc4zw2gRiYcMHMnJbWcGiyiJQb0MEBDgT2qdW6MYGWJbStkw+TNFXt1GtUydfm85o
I0Vw7Ge1IcFyw/+erRbcaiI+AC2W8eosB6UAuJAP0lfOHTPnlNvZ8TYKGn+XFfFB+XS/j9pcCZFQ
OpEDiU8iSJoqFC+SYlRlurFOAZPsCjgFdopJTPKQ0OJcC9GXfN3chDilsvz2BboN7oVBWejOhLib
leH5YAHlIF9mhapOdl1BFaReuWzz8AHN9PO8yRa7MBmKklacy0QBE6IF1EfGNOTPmFIuJn9YdspM
M6zCdoJh51FDid8yHLFiOWhlxFfff5s7pUtsMBfPMpFpC8uCmXDiWLOSShmqqAVmthOzWAiG3QMA
OR2OAuFC1GvC3/2WUbUoVG7wsr49bQOKSDM2iE0CPWLgQ+GUMthDP91JxRG+T1poz0xDYlLKb9BG
nPDCbzipctkUfY58x025VYgADKlT0GpTmn7FXtAYzlgfH18MFpEPkvvu6cRgS1gkuD0PorYnG8cI
YT3it90+kXP2p+O8AiQeavJNi++M5HOK523pjO1LtnuPVvrcm1O5/uhcL5IBP+IPdjAbZWvXieVx
naL6I4iztaFCerxkhLWMzXb0a0vY4acapaE09ATfJF8gUXbTawOE9yMLzJVvu0WfKafHKwHyVHmH
Jmwyl8YZDYhLAx5WVgwW21jKXMWqjuGZeEstDRHqQCgbWulIuBi6dn+hoXTpaxBJGoA9Ce1v9P+t
ThqB84PT40J/rd2MzcLGHP+zbV4sxJBrR0pt8A+Tin3Y0tLUO7RdO7Xls/Ev8REIrUivGx2tnDXZ
sC3DI0E50UsbhtiCKFC7AW6eRKT1koBFvKFwijWBrpy2v+vo/wX55J1Lp+yaZABfLhl+uBkM5ePR
FI5nzF8yVZLk7Eop/+jxTIPxLvG4zv6Tj3q8mcPiKx7+kNVkcxoggYINv4K2q1AK6dHzu38lzWNU
7V/xfXRcf1aPSI2Y8NZIvkObG0rrNCZtkpwkfmZGa9e9dAgIxoiEqqkpJIKaAPqmUVuf1JjMGSew
0FkWLNbWfKWNQlNTX/jgfmiKaDvxYrXXEcZhptrPnEqktMyT1MYBeN5FXfVQE9l/U1/gUGCeiq07
Ao5bSeTexOBO9u51PELyL898NeUlSzgKYkj1h0sQtZDegXl5NUO6PclmYtV1BiUTJiKc1vN7jrPF
SAkMMS4XHupwavf78jZ1gxChFj7PMjYupuxvp2V8jAve6G+eA8Tvii+r/oyPyGSaeAKNJHCqdL56
CwQK1kMXsuOLtnB1ivhjbvP/nYREKA6jg6jxI9zR+cpxqIAgmJNZHW30NA5T6+l5lKnAQ/OPgBV5
GLejifRa7W1HWcQSjT1jBpRlakuvttf8FfUj0W0ailDjE9mns84ID5rxnUdS6GtcmN4mnBoiVaep
KahpOjdjjHvCtqeAGRFxB0/Bmd7fxfYP3+x0FqHSOcEz2xUIWX/Z5ekNy8xJT63od+KoKluGziqE
qhQrT+XTm1m1Cy6NcNEazFGU1w1oM0futxK/HK6rmQPM+qfyQBY/NL6OS+v9HmtB0ZkcC2JauVuI
UxUnzts/FyqdyvWs43z7JkDMjxwBuIJWmdsgn2XFTLhwWgtFJbFX5yYfedWuJ5sVzUxVoxe/N8MV
rcLOGlXDpJcONTgtXAfVo8UKNCzqFbC6pCFXDoBVdj6RuWjOhFSH5TJ98wo54tsSv8BCXUwvjVIO
2PbtHpOs6n18xtENlEhXWy2nlZZMEAm9uJmSTQeAYn/JFzvcGqNBjDMrKpkTflvLUzlSexKOyXMg
jW+7D1CXVO5PlNTmFEgAvCs5UV9k10PorWPlH3AM66XG/QIFZTp9V4f9uWNi11sTG7QNQfLlwAuf
pWDxVPx45USRUeZB/t78RE+7ccHtwSI0Yixh9eZljwfm9MnyYzW5XE/TYx6k8M6bd8Kuof7ckEFl
EJJaX+OtGe+MPd68uTLuKvEsNBjdVF3q4cy6bVDGPuDCxBq9c4FLVyLGlODvDzaiLzpIDZ27J/yC
iwuoCJC/S/I5wqSlUTAwYCBAWvZ0y2ZKzI9C5zoBoBB5nI2KpvyoGDIV+NWkS9Dqi8bYDkZCAZNY
NWfrepJAGUVY8wyjw+AI/BcpndTz2FafEkjosqGnTET5lU71lhuMxCzZpeW2jl9oQ1QoM9nu/FYl
fvakyh5fUH1a4sExV2QPUToog8+B3F5AydBHuiOyU/Q/RdnSVegvtcOW2oCs09MfdjExaHSI/eAQ
lKYQDUI/Y7Vsus+kTZ0Mr0+2mykJnEoehUVKKze3JQ0EmA4KpbIquO3PxJAmQC3afjQruhw0M+Xs
qJb7flng/L23yq76hVlr5WyZ3sylf3RnMc7kT/zIFZUgEYyNW2C6ddG59kWvVKu8/DDx+sVEyv67
K9TFHhK+uwmPeRFYksD5d24KQX61M3uKV0mmurYhZYpYri8keQvS6Ps+73TPl4R5AvxWKmGhRyf9
c0e0uKpDBgmPaYn6EQaZKMNWhuEIe9h9WtznD22FjAcqrpCvX30yA6WV+kGZjJpZbLVwkmEoHgE9
v00wKW/rNg8uylHC8tCt+xIV4j09lE3ZdFxyo39mhk2BOzWmFi33aPpy/CbnpOMj8PVLUJhFcZX0
Bm7PAQvCsaEInE6r6J8PYC5kHX0jTGdo9D1vDGGgsz9zaUjp2WjI+iQ1szosXH0e7/L0fq66ewRP
WI6AZowFo550rB200UkRIfY8AFZCLOU9Y6RnBCV5awuU3fWe0rQ2Veyeo89zqVBd8heIeXS9+7Lz
RXwdeNdhwhfr2O65Kvy3YdpAEHUyt6hqPSvr8clVb47KaiI0NFoZLlZkyRqDi4ItxaNupDIkYkVf
hZXm9UJjZfZPQq+JSy0yx+6DUP3k4pVCXloM56YTjSbRHvT0vMLs2tQe1ABTdXjLO04ySrYv9sng
Ksb2Mabi9Z66t3TBUVCd16Zai7TP6Za949snzYRymfOSIp+75WBDhqwFZIC6ToQcr24gsNxcvH6g
oG/MA52spz7Bgd6QaGp9RzZtdUWAPuWO7UiEY51zFF5BNjfqSwT9bZmzWc6EK3YAxO3A/U/fMnWS
nXrA/td0mX8o49Hpd4o4aR6M8gtFKyFPyTvzj9teia2npyss/jShFQn3N+b0+gZNENC62fA+Wbdm
GAAimru3bjy5pP2pTYV/oSuWcb62wzltWRz9TIPco3gEYVIq41nYSq0YxoLaIl4WZLIUmfYDXL6P
K2k9aKYuy17CIxhkr4dOGeIjwMsUgrY1C0saSfu2mrc+YKIDDZ9noJsuc842IHDfv+5v1EVk42o4
HTJa3pvIvhZLw9GryuIX5H9W9+R/P/kM1gHzGPGOASXGvhMEDfZgmju13VpZNDUjiAzSuZZrRIyl
eFLELmKKvG+NHYU9lfF4QmVmzrNWE4R0iZ/C5CNYFWHcBfOsArmE4clVftBSRre/V8TO1pP9bFTm
B3xdIDXUT3FrzLNGbvPGmSbDZuUjj4lKjmmlDky+Kd37MDwugwcqyghxAN6w1GJfVsI8tR14Zhmc
rY4zKAoPPaGlh1oquPvmyRJKlFxpygd4MyEEG//nrhtMHciDjbgROagWF5Yc3GJn+/ODoa5jRb2K
OpuJnGjbA8nMdIyti71yqs090/aleLqCKZt4jV9jpccdfdwJLnqo4vSwmdVmtWdq8aa7B4rrxJON
Y55way0dTKz+BZgCq9iuuRQ2xb3XYn/ECS36OPL0OHYFdX7otiQIvoocbikBv1NXLfD8sSDHTPIY
0oJkuhdQRMDjQi+shDV2rABxc/xQ3c2VsXeP+i/A+bm33WYUY1VTj4TDDVCo/RSg6enZ3LGAck8s
VVjcPNQ36cQUhklh9MM6TZbX7TpQpLfT0BLN3FaH5FoUL9n/qGoNWtm47kFoRiBoPRweh29MXzHo
LcLEfSSvjzkvkSbEzYKa5Z6mH9Uy8ct3Rox+aBoOXlm0uXX9zKZpL9FZUjwwd/DYg/3TS3CTh9fN
xxK3AOTWdgjZQmJVz12nmmWaq+y1hOEp6WVP1Z8G9wx/8tJSuHSC6X2Yhc8ecckTxle7yI8koxNN
vRpuy90Tu6+GVERlWtnU9qkl2/SopyDc4mAR0kAiVJSKqjc9QXbvpd9skTz8g3T0IJnqFanyUS35
x37iqKFXTmlKuJUWhKlAsQ2E4kfLQzFiPd2SaaJBAHQpSznxrmiF3k2WTYXfcasW383vanfgtLJI
O4Dox+djv4xFLNzVTh6Xkdc5LVue3eJ8PCBEzHg6ZAm52ODuyh9efLT9bJrvReUa2XWQ9z/q4DIN
sSJkJqYw5NsY8pgVPeqZ1HBod1Syhe1kSciCscIOn50UMLATUXLGj3snE2dmaFf8mDjKz9GKonJl
oV3/h52fLY45e4tf5eerVdBGxLOKp/2A/UlVqfS2XEY1e6uLwHKU0YnEf9zPfKSzPWZM9JI9H/Ji
J7lVLr0Yk3EveKkUqy2rL+3HfNwvUWxXEe7t69Q7MeD9KcsTl5BZkKfSx9unfG4VyYKjWcHHEF9l
JKiMLqj3riJD2Wk01Gfjm69wXMtoKOdg8xP4hGvv9X0emOCaDfI4YhD+t9C+jaRRw026Ax6+UYcT
PXDKnbT60s9jCxKZQ30Xqdrc5NA+ODigu7+0akotNwsq5Zw1ihBwTqcvRd6IR9VCVrMI3LJpUUhu
dYhAIE+KrjgRznxUdxkMyCjsPUL39P2yrGgMYI8APs9sBmTJTLLAiL7pUWBBKUdRk5fhUlAcD3HR
RpRes4jKH4Cda2O+VSP5je9NpaEYbaunPRRvfeuoW8Wn0D4LpvPXYvPKeKa4Fbn3PFksWzw75WrF
bV8zhvMhAvEuKNY3cpPVif2sdCDt8xcSoCHzA5tvZMhaIkoHCoIJqjKgFrA2lpc5HvDxYbGL0YM2
9aewT8QozDSSn9KNiS+H35IvrlYfIV7H7cLIk+JFAFFMaXXCOzBUNH2sUglAggcAcczW6ZqpPLz0
BZoGMgA/CpPuQgeh8pLAvD3+OQYcCnZFQUbTYH5kl1CCBnprtonaV58vwZ2jMEySP8BU4tql5bo2
cs52u96l/PGespvgQdbSBE7QCvanRj9od5XWCyjWbgMYYMvVfqb3O2nWuKtHxIO1XzoIl9XmScbW
mz5aAFdXW4+sYVQU2sy1ZqiTJsR1nNqGJOIgUzEHj3xZkGvzxEahydm/o20cF+dPiYUBJz/ImbH6
4MghIZVL2PAiLJfM86FA5fyzxHIREZE3Kz0GTTj0Qa4ECkqCsHjtURJsomQN6IOJTSFeLSBoVigw
JmB3MhiqwMgZfuqFIgXc0ApKnhTMHd8DFOmyxl1YrZdG/dNTiGI4S/3SBag+FUQ2HB1G8FKD89no
wJBgCE+b+wqHXVx5RN8l7uVtuss8LYmJOI/SVpDdr4a/CepLCx4Z3bto8CTiqA4TqNXjsE6pGX4W
s7JrnaC3xirh56SUyAki2ZvNaZ3ETdUXF0/WTSaB4yKWz9HfK74i2KvZ0r4swob/cy048GBfFm+a
D41Q7w7HTdMTifbH94j/3LIkGVmI3A07jmILrVKoX/HMNgy6St9HLJkdup/gZQt82gwN2YkhFeK/
wFCXekGmWes5UpDeQLocVWxjtF0MQgMn5mnK8+rx7h1Rdxwp6WKto5k1Q5rS2yC9TxnQQ+g1Txi4
AW0CY1JIlmsP9gaIRvMY7+3W/07/FOAQApAG2vES5fTzjH/5jAadS5BYsUhd0tIZPtgeOtKe79Ra
q79mgIA1wrUB3+pS9JZLrFBgIgaA3svZ3wwI6UH++QWZL4QdXV29gsxebZkaZG8XPtL6YNDjd+Q0
ZPGqbl0IMM7l3TMQ5q+DniBy4Vl/bJ8xJ0jbrdm0er9plRctfw5n13D4TEQddmSW4RMKA+Nlqii/
wJgNhgGVc5TgUgAfc7/GJEQNci7jm2+Fz5VQSnAO1brTqrPDcg/48vQ2o+6WJBjhWnYBsQ4Pyqml
k+00GksdNKHt208MoLHlHkaCrCM5+75QV7tCTm1xP+LZL/d0nJIcWHujci26YLzucIpqFoWgdrun
gkPBSUWHXDJ4kiN2Y+JeFtbX4JOBEFnOFW/pyXtMK8IIiYZ3Ojv9oueYf6f1XbqgFnD76f7Dh5zg
ECyKHwzwXiuxsLWAFA6tESzgl6lzX8WJ0cXunVA6/vwKhcxvx448Z/Ge6hO6amM551xtJe8GULPL
socXJ2vKAUrL0eYzRXm2zb+HcMoQFUa86lrXISSLdyFO/ceaOXqpqRh3iw7w4nr+Rf0ciPKjuTd1
7F7ExHzp/7uB+42cZxxZjLYlXGz6YFAkO8XGvztKkdGzg261UCRJBDgm9RrVwGe1PzyX89ejyJrh
t+saH4EVdGAt1jv9WPIVK3JSRarMSuMdtSLcABSvxLcI/AQEsKrrdZfZDaDpaA4RcCBQC+ZXJBn0
50X6BA6xG9RftIvYNJaKOXLyGjZ69k5kwOZcF8oGyvM2jSSPIo4lF6//X+9S8jY8TpXKRgJ+oUKc
PrypKRvyrzo7lg6+bozsR5FCNabvngnZYMAtD8O7blq6nbu8wg1UaeCd/P+K/QcbKhJT8jHBnzJl
ti4Iru90LF2Xbk9wktqY7ciZSKN9XL6Pw0l0FSLtmqw8wrwVJfVVtUIAfv6lPKW8XxAwHQd4JbzC
z4OC4xx/jItiu9/OZ1wtQyYzDBxAA1mB3qX/SnXvEqQsMmVEYioAqk7gBkwxZgnZATix9qMlfn27
IXaf+BO9MgDBtQAQbKwhefoNCjg13xJgt4G+V7Mfq/Fl0U1+yT0pTHH0/Kn6Qq2HI4CQV1JhYwxm
Xyg8uymax/ni0xpNdw1XQEamrN0uNsRuMppFZTnGGsoEeCtYfn/9FavVzHTYUGir9GGH6LsCcRsh
4KnbBdQEvvqevgWLuIR7DyXremwxrp2aFP7kHLamN+FhbZVmE+5T3cCsHRSpRr9brcgwDEinnwUk
0aXcEpkY94xqxEb4vrqWJdLUndQ7MJPYLAHvkC/eB+aJ1pn5kHjEKcVSrXSXyrEd+ERcZCT1SD9J
mPQmdxdrcBkislDkP+Y81VAZfvK8Sg/clQA4K42loHwzWOaIP0zH9AC6VmBGhtjcmT7dBWHkskZi
VDp5K+vSLGx1QMAgZj5fMi8T3IJiaN1bpHZkclYEZJooK7tqtvqEROmZr7G2wUWhdoeRCbby7rKi
1XU2LiZYYHCkmcndd/eMmgEsli/RJEhYePOCONpzxhqOTujwdmIQA/femMhz7Q+kPs71GRTMJaWv
eAjZUsSTVz7dWqPjdhUAEHO6JWGle6jF02ziSqhKtkDirxxDixKrqXPPWnbHTas6JLp80jY81h+M
0jfU2alSMe5BBjavxUfBzX+HCOMSqJmupcxvoXOmk43Ph2y/1G4VLtMmHfPNH/Sm+UeFdQ5E4Zcl
q63tiPQ7UtHyb6rhhmuauRGDR3iX9qu11HzaVnGwnW9C3H8I3tF3gdDH8efqSaj/JdIKpwtl57fX
lXhOdQDFLi1ewxYGqNBsh4r9hh4iZ7Nzru/MZktq7cdeG+D12F8woU3R9g8FlX5SoSJ4HdOg7N4F
ahscKwSEx1gHxhFUbDCHMfWGVslZ/OOUmpZH4bveZ/k5Kp6dPMzCECrC7fdrOvqT3+XemK82LXyR
/RtfHOUwcSOtyjYHw1fH4G/irkzTJ1mVelfFFuDKYOrY0P0oOb7ieHIeALEpi1eOva+/2dYKpZgY
tEQYRdb+bIk7wLBu/vp0199F5q2pdEtDiG055I5/0Y9hiHDjDMysaf20zj4XYIWgvW0CCwBSUqa3
IHMDDT3dsyH4K19V6w4XmhKjM5DTb4Bo4gprQgcExQNdIwf+GwOgGhbO/VaV5KZtTKCHPkf8o2wd
oCg0FaSYO3qi7S+g2x7wqigCJaC+xWjnMTKD7LIPnFvVn/FdFZg1ito96GQVJ32MbUDPWWED/YyW
OwxrMMiWAyO27ci46mNTXEgI9xeESPStlB500d9H8n2yIP4VVvKfwA9r6ASms2uF8Ak6DkpgF6Qd
9q+H9d6T+b5DNCESBM4tnYxI1rgJHLvdoIXsQqqI9g+c7ZZ+TwP+ZOWsU+Z05lE2EE2YETOuXneo
rCCsiCK6eoh432/dbcDoo6kwOd8Ldi3zrJDThuvhySScoeSN1Q48WCTtnJzB7CVSuUOVTygsjBMo
x/kGvt/TSAMf82FEC0hzSxpXuFSHQkkvkkwqjnmdsQOSZaP0e8n+CxfH4QJYihe143PW/g4lv4hw
u6jvw/BPvZ2csc5L34/a5kfKM9fLifrMcneKVycxQtdQtV0ghax7JR0HxU4lnuvw82+RDXShaZch
8COccfztbJazgtsYnDjGyI/WKzI2H34mMhc0Pi9PTMyH1CfSmdhjJ2e8Isbrq4FbDgMx8O0XH1lB
D8pNyFUP5lAxaaWYIhHlCAqG+qt/ihJvCidpbZnLDr+pOxVWYsChdxLdF8ky7Vs+wJHrTKNgc1T1
A32IHe82xva0mEiMpQVU88hFP4gQSpMC53BL48o92VGOIZVGtB00TtM96tYbmM3ws0+8qBTazVNw
R3+o++nb2m0r8GgJrUj4beIVqX5tny95HVXxgRxrmtHruUvBZh8XKLznykjyI+GIsDE/QZ2jZpId
4WqsLoX0JiyOto80YsBJP/96Syw4wgCRMnWxZ4Yycil3USlDedFmPacQLkNnWXsQ3wqyJNq9qDJU
tzTCiKZEblRNwjSNdGm9DS1H8Uuvwb+OZlet3/MGIaFkpyJ+6NVRnFNkqxOMWXKGzppA5WiuSqgF
7FVgXUfAo11nJhnMUIdYJIpABKhme6qYg0ijy7z+og+kpHb35pM47QxGH5aD3TEQhlX0D1KZvjKp
hbh8JNq7evdWmf0ehZ58qSWozGLnAUZHr9ikmiHEmzfLUDVFxMHCRCDpuqf13guhdq0icHXFGtIr
i+TVqCKezwLxl8lZTFe8DSY8lKK0rAYrtSA/JbYm2g2rBA/mAVxyOBJmtFfjmHrqPuQoPZMLpWd0
4PCshpE0rNE/Kc7vbRjtwDhYxusUdZYl7ERBecZbZkkZPhCq66QpFnzyTe4UkMK4VHHcD1tAqr0L
TSsOiWH/7EJbKcU2dFHhtGNWX6ZkFeRN0DNwGWAFjPOLKQgwvKvx/96JKJDr6e5iT5tfNpXmdBPw
jWZG7WIxfY4feYjrQ5S5906mZ25hTdN6MUEjiX/9TSlfDCm2RBxqXDNSgpYaXbBIIjOIBg3matxV
4nxdUzlExkEL5v3lDv9R6QmaucRkh81bqswc1Afuyi70zmUn3HxCuXI6UCjhCnJx5VUY5W6/thH8
Il93TJ/5IXRhpAK8lsuBCv0yiEDm/A1Vw7/mNcqs43B6PEe3RE7ejbzyIKunlG8jM92k8Xhyis6q
NlsIa5vyd9Mg5AlKKaSVrAg8XH6S5Z4Nzb0MewIv0LascnF38U/Bu+Fc5+kBoHg1PrWK66P4rkVL
zuN6AKVZq+yKqyhNuFwLMVtUJTHEVDKQ5DcWwdxDLFAK9Xx/66kVlQOnn6A5yrDV9Do/mmSXBhPt
DWxoZAYNcAEmo1kqtX7SAKo0qT4etLOxEvvjHhJZfAJUuVB4jAA80SvAMmbUaLDhdG/2Hq+l96Zo
k1XOKfTUPpjk5LYWoXg60MLN8GXwT5QkKoHBtM0bRd2Cm3f/OnI5A+rogcvAXggOsM4ST0+KhUV2
Y+7qhJCGGRqRwmoPU6cQTtrtogezC0v4zazXCxqCPTbmmIHooGfaxeS5+46/SeiBWxREVLAwpGaw
3aUc7fe/12G2LkmSTN7/TSNNNP1CDZHHqO5DFd1OK585xOEAKg7/HvknhmEreyNuG1duhuvkP2DS
VC+/k7ZDp6lbkYsV3jH+4dvK2r3GWf+0Ldmv9xxhkUVedYXcXWc3b2MeHXKXyToSpIIZ6pieyYUv
zF5CZjMg0QASgErlubLRMnTplaVNSr6Ys2D+N1HzESzrsJcIF+4IS+eFLyWfkq7yoNL0SwzGxb4i
mauMsgje1iTzM9+8fGWqyOcYa1g/oQZZVkFJXrNCIaDrxT5fj+jz60gWwZi66vetdZ+H7IjRvHFz
Ae3uH2pZ9zXc+y83xUFU7nEgrn0kUV/Jtmf7YkKfF7k2BZLzb0tdwBIdW21SIeokrYth01vWNQXg
iWmo1HLZOQ+vPuckji1JpMaiBy0vdEpkY1SH9c2UuToy+wUD+2qB9py0Ul1cw9XeIov2gyihUsxr
tiYE3rAgihRQr+6Mkduh/zspYxbsKCcdK9mHxTWblui8ZvDCcRsiFjt1W/PjD/dcNjMNJY4fJKwa
XhVSCPR6aJCixBdju7KrN6n0fvdAVqHrRD0tAXAwQfHCUC5TaxzRg9z+cSRSt5pfTkW4fy/yZWdK
uF6fhYhwhOZh1U8H8/YIX+cnIn/YMKZLAu5VxIU/ta+VV6cQBxpzerPKfpZL6ncJtZxza9FrT4C7
N5ASNzUdsEdAAqKZlnqNh42n4rzmPx6eir0HyohFszWPqLExBniWOwBpBaS5QzFaenOx3TkvTXZb
elD5Js8c3E6zfEsb8+oaaaCX1x3MZgMs6qEvKx8M2fPSnBGhSpRQhZzUyUnmh9ANxXqBRymKX0kc
VGrS76pUn3Uw2XEW9c/CbHMu1AkHdtK/CSvyqkAa8svcAcF7m82flNl1Exgdd9VQvJub8bDUb6R3
6E5wB+sW0BohrekJPO7DnoBdQfx9PgSQo75Z58tYqj3YC9Ei15W4OuXTx/VSf1RzCTfRiGDhY6SU
gfNJH3ocAAHeV25Xqg6LuIddL1VLwUGffRw3PYODEdt9EYHw+5gMYgujp3DGlD/xY/cFxSkVY92U
Ugsnd4OJ0U9yQUFzapLh/5EMAQWt2pzBMCjIRLmltnPuaKDQRi4X4RplG/NSc02Ipf78xt+quO3H
2dnM9c/UZpqKRfkSVCd6e3a2cg1L2LcA6pz5pJKFenu408M0eQ5Y8hbAMaoNoEACBgeOJ86UGKly
Mx7bS/lx7M+Gqz6jf8+OJKch89SS7EDSEFM7kMsqBGakgs/+Ne0tQQZryHgxB9RwkyK23+PAUM9W
lMmUp2GzxI7DBn+lHvdnxTmuQy1v7GjkWXpvasnXTAZYxNiYzfZwe307WIu21RAsGPX0mpU7twZe
0x89C6dNm+gM1RiAZKNPRjTPKaKY+UHDLZCYFeKxk2Ov9oFmCLJeGqeLAEB83jIzwFjjtv/ODm+i
Vn/4TSMb+Q/7OFGaNFMmIZLGaD3LJrA3axkTGis/dOIu7t6UFUMJbqk+sQC1l17zwAQkE0+ptRxH
NHD2fx1w/PmiI+7twXXkhSEzk04iM6GsrF5zZ77TLxHJERk3xMp+gD5sghpLmPGR38O4+WmE62tT
awGrM7YiWMZYcT9Ee9cFL8q2lonFgwrrN9jtCJJnR+wh2smxMoTrzC5BiOrbcRVcbCclXaMy0Wwh
8kUwXVYedDzg03w81g01pKTHF7MzhypbMniNnP2+U1qxbsYE9Bg4XXJPGPKxFXU1iCOBT/XucnPZ
dc0YR/wmkIuLVu3SmrDqyzjpPCVDjkV67FI4kFz235yOI29Fg6uoDxYQblrrp/AwPC0zCrtm+5xN
Y+zZ5D+GMPBA1Zz3ZgEDpqUDLYQAEDkRc1otRBCsnH43bLsd8fEK2u7m/rTSOvy7ikPQDKnmnIX9
MXICEK7jMKKhzDihoq3NoYUdk09YtXCrXTsZE3Vq2R1xbQqjubA6eEItsXGB7wCXfndmM8K88lky
fdvnvuuhvhaZwk27FXbDIBMxY4z8N0skKj2r6Fce45/JNFbxvAI3fa6G4e0p94rOF+gvhP2JpqLf
+TntAQEO2lC2mJE/KZQAMFG7WWjD5pK6uWo8ixz4tNKSL+OLzSbcdiZ99/m50fVto0ghzp6yskyS
YZ8W7EYQORWM4sO50qjI1UtC46kQh+fbyDg2wxgNQDJS5bwCWSnRUiWfhFgXzklQ4QxjsYEUHfHg
iCd+AzwYgZts5vkfjJb9DMTUjSAMnkGXnOzidV7yxBRnfMfIv71YyVu+A/CS+QWnfdCYC1OMNcR6
6vcE10KrZp+T1GnMDo+6xFtJdvaQB7dSc0CDTxVLigG/+lcjkMJILvGEgyxnMZrUlDsqCg7E9q6k
qJHk3Mm3FXe6algsEvJU34O2+hq6HwioFxOvOP+cPGtMkR6L+u7N5NDcQkSWRp0BxOoTSMRBdtZO
1GdwwbzurFGU8QXWOXUL6WuHBUPb+PNiS1zbKlvGI/u3WXRFf+kF4VLgEqF73S9oNOqHn//sVoRN
rznzNE+wYWdxFpQAAJP2/DoEFx+qm32VpaKDBOXD4dpV/7Y4dZ17b2fhlXlWCGdTDBLwDaPTyOQw
QeLFxOPXfajsLPlstS0ITQNASVkDLQgzWqeqISivfr8tvhCjgIKL4o8voUTVm/MP5nM5kzlecvlo
o6+O99mnOhtijGYyX1ole1FWHRliv6yqF8T+Jssb0TwV0E5UeAmRwPJTxaJ7aCRp2T+DQrBSSLDc
kSLn7ZK+dKKsC4CIslA0iwdaSub8WMKSXnPqyZD+yWLCzJ4cLRd+IpxCCMJihdFSYCIEiE0frojN
HUTsNMV9QZTBg4WfnkKhED5PW26hl6hZt69wqOPrzQKOyvx33Sl9xzyi7kiBKY7p8pAAn75nTw3I
kt6pAZjmz4PRt5PlJnszd9VDWhFOdIqDrTFTbUko2STOGkeZXFkUTuttDUzp/TVMqMVSSbifZnUK
hEyq2krg4wTWE8m6voipwltJ8s6MbEg6JXew1ecW0quK7XDeqSqPhCjmw0qdPe0vzaKzRlKu28FQ
KsWlW8ZwlihRgUl4MRylvj4TncJyZ8WN/JlyKqbDFGMl9NoPP8ywCQ9zYXX2eOs51UMrCzPepWBO
CojLAy/h1OEilLpGRvnPhACz6XosaAJUuqOejW8rPKNNUbc1SdoyGGAAOeuE/3QzTbU8Xy87/PAZ
i08JJ2dKiB19URJiulINtZPS2Z4bK66xhixjggICr6ILe2ASLE8to9TLkb7qXrVPTm0P0HkC+aWt
RV3XehazqwTzc60a2CvUW5Fo67fHstatxBKHTeFmAuxlsO8cX3uwseE8Tv1LpGo0FmMZUGWdiUOF
7KMThumUUtaLfJlI6+R+yEYV9Cksut1qsDuS3Zh7pezOCnZZ21Wp7COOaXcfo1zOo0RS7IXhcGiz
syxPivwEoUsNvea7yKYRIVZ6FvV1KnQPbkDaa6cMvIVC2q8B6ZgDppU5X8hA0byKDF4xzZNTXViG
AMOoWJhXXycHN5Gz6dY1HdaJwQwU9cY24nvoouDQq1Zy9fbJ4NJh47vxyylWt2Nu8oD+Okh15Jfh
iBJlr4O41iTatOw+hua4y8uct+xSBjH5dEG49PW7BIbtrk8hlQY1eeN97QC+CMlbkVr/bMosBMMa
AG8q4A6ujI4gFUng5aPl3PeES7vPlPL4xb5seKp22/dAQiGJPJiVSPGvNmr/6tFy1hNOTcqG6YWI
R6gGhqFOgJHpzknAPfISgUO8R/dRqEJvaW8wBmC0yTEL7QgcEN4Ec8ZUHtDvwSkZBcYZundsdFvi
HsJADggUkgq4HaLJSioLu0DQ6aqWWWMS8aLueKUBZvZRH5bIavJb8CaifrD3Df0zVw0QRIi2Iwr9
wYQ6JXZKgNK6VRoD9kRm1Q08e0ovpNIVOU/ewBm5MhtKKBHpREOIr7y/zQs5cazjQbyDPo4yxkLc
AG9cet5BtbKgzMOiEipQgo+Y+qRpkWiwrhuCwQ7KvUNuQ1a8ZTMHdoZCU77Rpq5vWarJvmD+rGXB
HN8JujwipLEbSVJ/d+n6/n7ntLMyu4qTuFAILAJUeDI7YBWPrFDBbzApgTESUuVF0Tn8AARaUWuu
ZPDHYxSMesKU4oInH8dft9h6ugwoxM5lKEh4th/bgQLVcJr0sC+0zK5oBRQBnF6JSAGVLnSHM+7G
Pti5bmP9qRYpeVzib5J/LEJz7N5+3NNeCj1tsk+STFJ4ljvlO1RDjRdevCHgaPhCzEr7F4I2q+Hh
96SLObEIkku7d6dhg0tfBmCQP3HG/10cDfhiKkzj/y1x5bOhswfK1GVG+ckhyaaZ370rm5a0Rve6
E3aUivHPw3GXJ3f4FcuJQP4lP5tJVrqZT7KAxtN6S/L/b3RRskTmgLPRs9kiwbVpgWz5pquf/3OW
3u7GzUmFp0Q8qCOCrp9SGf7lDmpitFHIbLLocMovYT/oby0OzPFsjU3GChNyRcgeinlWF4n/Xl8X
auzrymWFGMnnWM10um42zY/mR0kxPBUAMNSrIW3DsSetJgwBuQotot92cG72bjDtsQnYxPiAx5n1
9DK8LLmTfCOlqdRPZLkcJnvpH4J3V3/mQTlNZejCz4vUM0HMtUBcidgihV0B7d8tX6f+KqlIfJKh
YzVX9JM/A6IYVcKP6XNKHPHh48PCtvT4dZA05wM7URzRZL1GnQMa3XoEkZCqsPGq7Ic2rpXfg7Kl
NQrQL8YUNR6XeXX3ztWWxGmiduuWwic6Ff8Gix+RZgt1GIAut0PfCcFFHk3V8vt4UdzWLmXPnQvq
1h4NbNS349Zk6YZEwSnAaYSM0ULXjPiJdSeiJyJTJGK+gP2nmFppDU18JMxcaTI6n707exTZGtJP
ar9WF1lZ+HGbwy77RdG050Ar9oqrK8VxEE1twl6pjMrat5MKg4fwn0JUiKxIerxcwMBzHjoL5t16
8OLmjSK8d732270PaoyC/oIFzeGtMkwMIc9G1LUw+e5UKjmKcOaO6/UZu3motNWGD/N0VAPMIjOw
cyLUsnjYewr/63qtHLx4+i1LCrCb+l6ln4JUXlg1w7EtuwlO+iIcMmefhYGijU1g62yNF5I6NwP8
VXeMcG//ILweGLs7RGMeGW8UyORw+RKSiiXEZCswBjH2d8XGeLNoQY2ln1yNftorWD+1VOcYFQSC
EzaITFDce0Wn8XLGaf/0wqIei8vzAMLH2jdvRP8U+y2d2VytsmuSPv5UujVTqhXwfPWjrPXHp43J
lueIBaOOUH22mS7Fe1Z30eESm6+uoq5vvNp4oZ0GmZD1M+n+h1A/7zIp90pQZaODnH3ozjlLTFAt
C2Mb/JbCHu79zSgcwUaGFfRbQrDXMQcLlJjmBjNMZrIBVJ649YL+dD0iSpILuuT6xvKVt8zb7pcA
v+R4KNZEPjj40CrGsTPJd4jQDoHN2QxvU7X27H9C8QxdgS4x3W6NryoVNJ/U/r96AuELKdPHzMI9
y1d/Z/8DR+eJg6nC21/ycDSfwRp0WCF8vDgcXmzRDDYP6SpNtapcyCF9Ld8QDAzlOS07fvP1wwaG
9uhoxYeZqbowk0/gc9jr07UBY/CwtsMiVlYg8VJPnvvs8hS+aCq2EHFuCRO38t4G8+cBZ/Tf8kIV
McYkW+8PiY6bKFdYqJC+vq5IfQBowRZqGoCVNHwZQ4xW3DgqH+e7am/dyXpkFV4MqPtJ0Olru4ov
UnTDGuQQMYdpbCidhqrpeIWvRjxfJUin5+xYsUAAigGzS+MijJbkzKm3HWmI/a9tR3NaXAnpDXKi
cc9/9Ko98aL+m7APtT9sfOMhKGigviVBNqJFggjtPrMrf8xy0iyZrnVpKolaMrBpkOhjHNw3NDs6
zeBJJc5r0gQvu7mid5aibk5CaUygkp0T7YVsA3iH+1S71fOsm3EnS1C+OqZ17qz/+aYtKmnW/jcO
qoB17W0rwbqOsP4jJ6eymdYJlJmSSsfDz1jQnxw6tJkvp7b7y07RshN8fimXsCcqzixhsUl1Z05v
guAnPwG0QKWim8NivOaoUMpCpKHFPLwt/+NtZg0VUWZZobN+BczTa1EurOzaKaX3gJsX5vOZPIaC
ZSLgqDQsLAgQZztFJ/DIUDp76tFyZlUmEqL11/44wSFf2CPDLCwQHAkg6Y0lo7LN+1dtG1xejwJb
ouO68+3dT08QV3Sw+7xg9Q9xH18Ko6/+JFbAjtk2pUDxrmX2/t0Y2VRpFgzltE7o6MveKqrhVciU
s7xBdpnsBghz6AXsxhnr8byXkvWgrs7KW6iowVf+CGQ+HsDoC5/pa3oPprmk5FCo35oTWoKUvUNM
RHNNS7v97HwFmtG719Hp+iRplcESIN4ayKOfxQ73AkU2lmS8zK9M/q1VUCGl5lKJGYXYBdJ2g9pH
wmmz6MM+jJJbwiJ/GCBP1DW6Np0SZwR3Reaj2C/fygd5fU+Y/zSDyxQMO2X59TsH3GCUsuDQUhqM
JU6h8rH7YLCe1Akf7HQvVop9R3cIroJ/kGwIlEFihkqQgi8/DqppgghhUTNsJa9ZMQdzfjHBt3tX
wRoIw92UKfgvEC+8v27CC8PcN3HSuclr6NVv7kwt8YSjjQDhCDog55vu6JvVP9vKeKams+5avflx
vc3Jlx60HQSW/7EaLZR16vfgHeFnYKxPfXPNccnttJVZYXyVX35Rfn8Yw+pjmmgacJaZ/FQgb8sO
JBVM5ccte3UdGOclAiD0v061FR25qFHUaZBMt2uyH9u6+jHZFAPjpT1hkxlTBYRWTj2Dw/PxVoCD
38oUEVabN1C5pFEfvRX3bn9QYeW8RYXn7po1ZAflI14icJJGGU5fxK4U5yQfNPHfG1bCpu6Onw1Z
MolY+GjgAiErimvdQy6zqjfcMh8TyRykqFyJl4XM0KF+QHMfll7VI4/Zk3qHtLzR6aNUgd+wGw2R
naCo7r2lVIdFO9uouzopQO9+0GzBwQb+L3rMZLzOxjHpqpx3Cs+//yKdoqbMikh/QY/23uVOCkz4
2Bfy2SoBe24EXG7EYKDIbI8PcHnL9+L1q08mm7Adf16k5G4Oxc+Elnv/ClDKR+FYsvvSP4woo0cj
n6fVkUXSG9hYyBU1aV6Ig82NdvrjlS3t0dVwWC4uDfGu32/LMK2YbTvKxyTDv44V0qdHx0V2qT7A
IaPPuWp2Zuwgf1veZsRUXQt39kFyhzUeV10u+LMI7mtleNBKUfnGQT3/Jgg7xpxbebSi+bcWPpTp
nTvWdZ9QY5Yvtk7UyHnJWi1NGkl18kxVXPmOi8ZtwU+s5Fl9e5oJfNu64fGW1Qp8NeztaWNvbX54
lqwwZWKX/nibfV2xaSTLIvqoeUZO+/GiKYbevjz5bXAA8cIF+CwnqaxlPyTI9Cns0OzYsa/PvjqJ
EfQff6EmHw2IYGtuU/BmBmY3irpfuQZGn0TJChsILb1fJf3CM7uzxYw98FrZsE9AO1wyoUIfOlwO
GLrTC5ppONXCCVCeem1BrKpNrXRQJ1oeWg9pemXU2VTf4k1g5YeoNQDdmZ27DlzkBOMsSF8Id6mX
RI1P4yFaT+TNdfOb/K/kFNMZgBauWfgSSf1EuzJG+PVZWUe4pwtSi8UbxiHLKS4m7u/WAbWY/P7D
r9h8anvRvfMlns66wh2Zr90y2jUTqehat8Ys0OEci23RPNoUU+1WJuQ463nsTppIitH5YkFHX2i7
oSnZq7mXW43Gp0KjgT2oDTVXMLfxIv3CK365/R8oZsKjR98Xo11WiZHt3KakH28NutlMweGXN5Px
lUUWjYf82iTYZSy8sbeGdmAIl0YH8zyzV7a+cYYLmoTyFb+sXESmBwxyXUusAcul8pq/dTjM3dph
YpzoE4W/7CisqYKCy/5Z/fOGnccZ0MiH1ZWQfivxDKkxFMzfQZuVWX8jnShcL5aAa3n60dlsJKND
0N68dIE2Q0TKYqT98SEdyutej5CwO2uThjO0LChm/SzhITRzfDHwpLCLbSngvQrjo4RRJMCzLIbz
AH2BuBz7oUCjqbUEnfLeyFF7mEEvOQTynXFbo3YOPKzE5RsD4jEFo6Y+osp1/qBYXnZIXFR7AqKK
kWZIjF2N4iV5anxLRsBgxdZEuBPstDjrR2zgvK0VS9ouKtZEqQE7/k0+8rTG7tg/r4QVkgj0Dmpc
0hBiyr9BKBilcBD6DLJNPiD32BcXZezg9xoduEUjnWRP61G/OJR9njWxywecK6tukKDLAravVLb0
kz5F/sg9JYXgwbxILUDKBQJhJ+iFW/oA2BINUjNi+6aBti1T7T4iza3dXPQry8qPfsE1DfdNtvno
HKcLVdFUj11csc1YqRIaaPjl/cRP6eyYqBQkqDlThT59jxdnXQ4qMUaUfg22UPLauyCxKxP1loB8
DH2r8CwMedQHM45aWxmzFfDDyydy02VMqbkb3yNgPsDH9mLu+e00RFbtHaNwczVhMVYCq2hBPCU0
QlFLIF68+JTvf+T8jy7aYm9drSkGeuRZX30ddlbcK9p4Ru1eTgWxfPunCr/uycyfBxQ/R0rpFNKR
WqFacZ2PmpDQUNz15+r5ceizkECw3csXqJkwJrc2gmk3aLq3lXnxi/8TBJItL1bU6zJUQBZVICrY
cESC38GdPcp9FRle7eO67kA7cyquWZwrWcoScfc7tbAXLDFZy2Mz5wJzfUJ4fOn0bDqWoBgOWPsq
VCCFqdqhLPGW3j2wgtc1g+YoCMFjI+DJm3uzNF9QbcgLhntsERsb2bRzkTBDKXFaazthj/md8fQ+
qWlyUiTbX2+29qBO9ekl4AqaHrw3R1m93ge7fduohoTxLbedHOlOH2tVfbzYbW3IMt7JguCUgn5K
PlYlB3lFPjYJho5byV5apohbH+XZgPrDIMq2xHkaMzEne2s6KuDXl6vMsw1luIuurR5yGAVrmXL/
Pidy3o0kX41MyuOzlgXSGMKokWrujXWIriLz9Qe/oy/+9HWtgoWpAGlSFb+kbo+gtOWC9tTEfyMo
x1nZOgBQapOTw/VNzqlitS8I3DbkOlH+5sDgrDZxmo0QuKmIdhMjuXFcG/HdUjakEenjcsHvUh2u
kvLXDLubhQTyKgxd8x99hpE13/B4AMr8MkGjh3YO5IwIAx0EVhAWl7uvRA95Wrj++TQXUBuFPSaz
Tjq9TTIgfMG3/P2caksa+y7CvQnwVZMSaObYZPX/fQMmHACFSXnO8TY9RnRBS6diljBQy++ZhzuK
/bqzJrMBS5iEf/71Oh5LDT+57UK3XI3iC3PsClJD7ACqmf/MFmG2GqD7yqnoQWIJoTC+jjMdm8zG
IwRibSGDkuAkSiBUxSqEejzIWQKMO2TP5mDri9hIXKO6BETfFaVa66GnLRqjX3ZdoBkomSlOil9Z
XE5YKsjHjLFEXR2IXDrZofdGbmXte5xAynwZW/Ca/Wp5c5hFNBnonblxQppP7WMQuQSsO1MWE3MN
VWXf7e4M1vFq9EWUScdQ6i3lS+1REpUjY03Y4FQLozXoRDmWn+S3PSGzTCv8dglH+c7K5L6Aethi
Lx9czQhPlY+Mpy2UsugpnbTxZm685sYJ+SA+MP8LerQUeeqAOrP0nesldCFYPuaUaF2/yo1R/3XJ
W/Qksb0tBRZQBJzKR5gzPk00AWPBkGICnDH/hH5oz/tjT61VDvEXQHMrt7MiMYHmypny8ST14d4x
kgk6zMq+S4ztPbwTtg/6wVySp0jrpFdmyDOUpb+EsOycAilbqWx++n+R3trt7jZE9Jkv6j9KJSbc
e6LAjo3EGL+Tx1Cp+oD7HUNsUeq7iAYm2wo5QZOQNwvmdDhUWmL2C1SHLGS0dQ2vSfjPiW09o4lD
cTVejeSfyxrakVwiIMvZgSoXttiEaZXKXXHyoHZYKdA9LgpRNjSRWX9PG3UBH9JpYrAQfITaoGCy
6imTLegFXvBW3VvU8uC3X+3RBpa2ev5nOGEWY8WCynyJ6DmvGwyRYTkaKhnThA3TKKv7RMYIHoAT
Pju+LHfk9VmSwbZs1xuTCTmlRZe9OHV3HocL+svT14OBTjPmiteMSjM5614+2I58yJdcydULaeK0
6s4/WtTPp5eOljinmanD45an0LWTSBPXFkIt3R/Vk4FwUODv62YpgytHogDaf8QfB4YmDLFqxu2W
igBHjVUyDJr9Om/7TWa2YCGMV+rtrZocnssm4jOv2Kk0gwlktey/Ngh9lG4OuxxBvBEH3MgDuaWH
RHI7DToN0PNy3sf/ceoyxfavXP5wGN0tKhbePd2e3r1tCHsp5Qss8VUZC8Y1p9BGiGxVCbEYXFNH
CtiNRXkNtxq5WbaKOi14OJBmqyTkufj5E2b9zZF9zYEEuRHlsFSoVkiKGD7ncZ2PMthKMwQaSUGm
uJo7Z+OgzwgiJyq+96bz73oyTPsI1XYIvMUV01UMuAl0KWVxaxnkv1B7OvWVtDJWQzWDoqTs7krN
nZuIZUSOjeJXTY74J69mbi3YGc8GT2AI36lVbHtWbdbba9VJQe2cFhvcRl9t3tlEb+wurIT0YOrP
++liKeyKg9T7FsJA8Q1k9V63O9c2mxN1vSRTQgAP9nGsx7vhuxetGZY+OGk0accedaI1wq27Hqlr
+FmU0mAIsHJs81+kU3NqL4IZIbo7U1MTyf4mm7ll1AMYgepcyloWaEN7B9NJKJfbpX0HmSOrxFcK
hP16EkLvdGPPk1mgk/EDM/q2Jw7P2mLy80UK78EpXiK4m3c0Bfoy8MlW4NyHMXF1quw5swuEF+ri
8aBZfRTfrZJx0fIXtiN6+vY4xKD3+UnWRYoSUsBL8xxgTn3s7kR2rEqjANH2Fy5SmGxDifrpqCys
LxySkdOY33PVafeTSXTPZ9T3I5dj+B1KgWcvHPwgxEWHgrLsWqxGfeB3rTWKoetEAHF26nQ51zQ/
e6mXt/sOm0RYEet3+IyBeTAoJqWoi0RjcH6GwcPjiizKqkGiOqkdanaWpLTIZw9GZulKr2eoTLZd
c8xXVOekB2OkxWkMMzLcbO97cCtU3inFU81u98hTes37JC1lOe/mItlb1zF62sHQO9OKdHSpZkEs
27GlKwIBpAywUNRUSd2MqXshXd2QHXFtRXKmcKEeFVeHksTedEnZQ43X64jyFdbVJCBt5kLSXMev
ugojkK4AiB/oNaiYQWA7clD1cXBcQFQOAaXDtj6yRCkvsKI/1bfKJysnbrSOhOVK1AW0QXanL/NK
NUW9Yt7WeWNEYp4BxNUMq7fgpGlzQN9sV3ea9GTEvPUOYr30cE2IN/DbPnQ2rGj1mvbnvrXzaFoY
zTmgckyrVS85dic/rWcz28dU99UksKtwquyYSnGYbB20eEkeeJqASmacbyqAbVLn/wglYR83781j
qp7EDyxFKUkcsnn3cgqgmtMOo4fMMkkLNc8ECs6ZqdQODniDIgxY6CHTMInwj/8MADIlZlYxWPi3
hv8n93uXsX8sfq9WpyQQHm8dZezSUQs563/R6t7/bSiefcOwFp2/+2hYdrnaYpWHQI5VZXkMVhF1
vLCqBKGBWTaQIOoLeH8POnxfiaPChMww3JRsT90jwu160ru7k3Ax9932jamLU423OA+j3UyxS/CO
ZcJEGQUkX2QW2z/nOVDxORaHAjVidQzxHcFBYfhVQzPDo8zmpcq6eNYNUs0k9J1EYICF8ZWZ7OmZ
m5AVeBxN2Ohw4a5bd9+WKDR66rKp2wOQkXSJWLiw/+W4bq5tWpoBatCtYLlBILfPfzOVYm+fRH2u
U9nXgv4xCEFYK8Kt+ACMrEQrUsJEtW543stThDfETO4tTnLvKJAIlu77QDdOaqtAmtKA/iRb+sdK
+PZ01qzVsgBAHRZ/Ci0hxPTHNlSz2CO7d8bPtiuTAGlqFKPxZIg2F9HiK7mBO9ZXVlEt9fA/GrE2
oL6zyqAbRO5h90lKMiSX7Tp1lFvGPLkcNyb1QyBXOiqxBq9fLpHUOol+RYoxROxA++lP5iL51/Bc
6PlRduwbdFAPiySBp+tUiNtyDAa4n3i0IEcc0UTKryIajYJaCA0YFLMU/ZYCt/GsvM6/W3jktFLa
pAHEsoZsM7cbfzGX/27eQHVNkQ6U3RqP9Hm4ewHWBLESyTz3DVfGk5rEpt6du6WjFQOXoOozaRMe
+o9fW3YguPT3LIeVJybgHUzyk4eaxNlrdsIzB7n3HnEVjYLOcTxRTgw35j0h2db+mp7FywEALbWu
Jh1DIQzQe3+WvvjieJ1+AdLLxqg47UtY/8E8AYPEsv9bJoO3A02jDMgZHeTtTVvyAcn5to4/X4MD
OVZIoMgbGTId1PIz5RE2nC7kIvpxzWOet9BiNIWIjYcH6veCeqJF/8zLy521sY/Ej1O62VUBXsjA
sZ6360UxFAKk1/UMk8LipQTHKuh0NuCPk5fDDhjKz61+sQrGiKL50pbXBOOk7NqnFxhaEHIplbUo
sA4rwMuOnXm6HkMz0TGbCVnnLC3xnf02bgQ4gBsGRnUNoBxfDixZN6dsDg3+IMfveLf2y2MNHe92
w3Aa3SOgNtCsmeuGDEulBQpiQ5Hd2Do37vCR0vZAvEXuzsMseWAGQvp0lFuE+pyI7lPyHVHqhIuF
O0Jcqyb8lXMvQxIo+NhHXyWtf7ZLqIP6Y6VKFdMBANEZqjJn10UlziQCK8SSv6/5/Ycri2t31SYZ
3+siBrE8GaIWr+WSndayahc5DMFN7JICpyQgnQ2QVMB7BwXG1YLtAyC67IhUOAj0omw7oQXa4rCo
6ZSDBEpEycFg4uCeLh/7FE4kQpgv/m76I1vxV/BEJy5WGo/6DU5syVJTrYJRwPJicPNM1F597dWM
9FFXh6AoME2QNgTTGx0539iPsdB6kEDQGUa+0hFdBWT7OmN4wBbyH2Ij0QnnJNB8oUEMTk4ZpYGf
NOCAZjH6otAAPzETNON2TWFjNySS4+gRfG8gI9dJHhxxFSVH3khKYj4gyZLkBDlNVXXAKbvchAUs
DtGnCT7nCezdUsXasFwF2UG6fqIU1LXzkSj/IV9XW4aHTA67HfuVXtvE6OrxkeNIiq/3cMPuHYee
P6dGueaVXpQAbov6EwxnYKHAYDHABq+59GwuOaWaW0+39hMt2MySSNsoHfnknh77UmCndTE50rSx
5rKjwpUHpesqG+pDd/dUYGuZ5yV3V338jFku7qAcpVQU5scPm2DKmLIpcRVjFB6rzpJ9Wkh80Jzt
gLW5j0hhrQ2tqVDXnJnthZ8P24wd5OiAj1StuYtNwaCHQvFNpd7onKQymhcyMTop0rhNlpPPWlKI
RLoF16NFxX3OtrD0MfRzqHnuzZFlmyOgUyRxn6v5yPFzCM9gMIyi8IWvbgVeNF8QpGGoxjkEPFzr
uMNq3J5x9h24+QoKgLrMQvWEP3g+TGAOZzlOQF6erbzNH1WQ2ln2Qkl3+q3ZK8mMBSkoOteqOeq+
Da49mmM0r2ys+UXSBEY7T830avkG7bPQ6sPatT+5sMMHplOiTistSzM99oY/9LIbWHm1MXjO+xsL
4b1gFahBgUf3KES9Cx33F1u/jrBBPdI4O6wymS9nh6Gcfke3nxIxWBl5cXDcbM7XZu09ohnnbV91
bKExy/o+kTZBZcIc/AISq0s9zQeTRMwidqqOdrYQyhhRv54xQAy3yEjMTzcL0uZ3/vjH2lX1UBGU
ti6T6mEdKHkgbNQVrCgdO7T2TJ9ASd82Z7pKxbqpJIQqPee5xtLFPfyOC16b9m4HaFi817aXMSQS
JhO6jmm2Y8NQOdzh9Y95t5UJ0otExJXDoqXqidBmBVgiB5Ufr6GLCNPuiYKlXqSYi5dplWVmAP8q
WQqVQuqVH5vqkDPIgX/I5QewB5kuLRS4PsB/zmjLjFz7O047BHwiTPmA5FtZB6Xe79mctVOtni1Z
zprOxi0W+TSU56a8GbE156OJcubXNI2oowWg0gDjMoyY5MtHigL1H+cAMdQZSwKgO49w/2zb95Ke
ou0A7x1+3od0Tzxv1HNvsmnRnD5H81Uk1aNvT4v01T96B9xJcyCJ4PtY+kR9GeI7AGJWz6Y5dOZA
7zWoce/C3s1aTUZpOyhdondMRUExK3mQ8HesAhE2Gmfa1k8I+JfPLNZRWTfm8dtgThhnE0m37cx3
9ODc9EXeFm8x0GkkUTL72hNfO3Rm5k4QrHebawvP2v9pU2h25ppXy+BQ6d61QYO28NTZXMJzgguB
9ngXWjZsNPixVxNYODCl3cecQeyUMCc07DCpP4woz3rIrEbbTz2phQkdE8evtvJL441zk4vDGkGI
4mv0sWfUB2ymDsZnI2q2YqLhBQqx8FNSobaYmRFn83MokqehbFXgJJpuDD6baNg/BsyThmSC9SUl
2gZZpIV1e7lc9B+KsRKlGvIn0SmOOq7GQhHOacnBq2Zk1KkxS89muFB7vO5E34Z2PH2ANXpjv24f
q4S2QpcCJhhVmIFy6ksbXt6r+ws5Yq1GwhTfMzeh6JoWnbN0bYhc4dr/e8EHYz9Izx7Jn+wJsqP6
bwZ1l0svrmKrk50a7gl/Pn/RUC1vHEQqmzaucfwl0Jz5Rmqo1QqhSVRIC1WFo/VZlw4INKSn6BZd
ClnYueXjMXrXW8nkkJzf+INr39QzcZhVa4q5X3eIzyYiF5gvuOzWNjbwLlFPJqC+BuzQH03p4IFI
JTRl1AemsEeT7bqHRUjJLP2VZlDvKr3nrSusGWjYe+CcUnYmFTfaPjYJFyXvx5HGDAQd6NLUtzPw
Izu2KOAscLvZKrqnp9qExq+z84O1SoK5C2kzZ8+9HrkW6gnJMBfBt7uE9Rpywab5nb46ptJckWyQ
ub5d+4ueEuCLPtU1yoTsV8N9teJVcBALihiVSRd1ssVhC2Ci3ghVJPneBCZGCIzTo1Xkc3KCFUDZ
lXkkbaJ8ctkI1mnmuigrHMCmKexQ3ppLLAqFZodC24EQGGhAwSbNtY7bzcQf89TAX1oCguy+Vl39
Cz/PGAc8ze3PLPobrLcjEOl5M9NSWBijL6u5WLOwYE1BG+dv9tdt5udSCu2LytW6cqjbXTDmQLU4
GBwxg2Bqa8I7RQXJRs77eyFjlqQ41sfwP77JyVcurVBH3mFpKZbwPXnaVUAiPUOkOMIhSfLZfUYN
BY8+2+OV6JZuy52MveZ0IoUJ0VaZ4ktlpWbmGu8MSt77sJ4mONtNohupno8MFj3M1q0f5UIM9kTi
FJz/2tspvr0ii57MAVGJBsKZwYAAXHnqPI3ViU1LnQePFVC+iYmXJOYCA2aMYgf1VLKEGi76t+jP
yLvu6CmR+fC9Qj7E8CbMbaUXPrRx9GfCgG0A5duQBfnRca/3s6rsYXCEoWdNM9irH0jXBuyvXTsn
8/VD+gL7eXKwr6xJ47LdiLcLEIX4RhRilaGdKkCkxls6DbsmQ0NTlL5ckcndxzZGxhildweRCFBt
VKbz/3dJkzI4wJOX7lb+TJhgVS1+41jcNlXwxAj5lJwuaRaDZq+NBIlr7q9JO9W7nMueL4d74m5t
P2ebz1RmwPE3uMvwIhWWhUjSwz/6Li+PMjFQ3/iqXHf57tBM0AE3m2Mf4cB94VbNcw9OyVj2C6wb
aoW5Q0VikqV654nXRUTMet8OoAhD6+Xjg8AjMITu464ELnRq80/hCj/HSaWjFjju/ng9AWv4aUZD
Kv/bxj1nLzepzYdwCENb1XUjdH2OursQaIxlgp6EYW4fLrU37lSvIO6mMDmexIwdMc3QJMXf5FvB
duzPsvZxPi5z9s9ePN4aMu/GsM+C94JDyXCMo1SV6eXLrDvo0nLfMbyII0R1sHAE8+W2QDnp3Edl
7PuNUoOyDAtkT/+7Kccjny5jf5pw6w/HyNiZPwNuWeZk6Kom5MmIpfWaSHW8bzVo+5rNV5/WtajK
i+sOjDvLkuzafCt+EIYKRo4kjTkyy6SjIYmXcDuqHXFV/z6b2HaAqEZKTql6xkBmJbPtJSi694uS
W6tEP6IOFX8l4c8PVzchCu/xjBCIOOL75d3A88ESMEub9PV2dURnOuoKyMyoxmRDC6n4iflpbrwJ
5WHJB4TkQrrRVvGprBY593lR8CRB4fUOCOL66Dc7aiM3pXUvy0Ha3LVvRh8BTNaZyH/U/drPuFta
Q4yRgNlHQmvMbnc1seL1kcWvXlTXx2jn9ThvX2YLqIJtcA+62AerwJC/FztvQCM4mK1LuB5VeaFR
ck8PhQ/l5HKhMlrg2ua1UpMbYHH77AMQRD+ozOlIUJcuqWyOSwOhDIXUWeMrdrwxuygloMu8bH4O
lzbTp8KDfxAQ44iv8aA4tllMfyizoOeQzq74YNRA20lOd4nTHflLMWLNy4Sars+ep2yTBjdv0mXd
wJpCI89GTc/4ROuoQUslfG5IgiBtu8W5+dqnVNy7x5QHb3tpSXNvRqOpVibPI0dPdOQwFuICHvnd
McgAL88uapCh883rGC8KC5G1rX3mWGq/9kU0z9wuAfxaL1DMl5+/b2fXPDmftJy8wFAAWxxT69R2
ofyF5qf9po+jBjEHTodxXhceJbIkmE4ars27B7LMXx2e7KVkKqG5wcseWdzg3rf+ReVffWLyH1wy
oBDfeSLzykTTu/RlPmLtX8EUSiMKQYpKcrfEU1IDG0RTyv3utGwTkfX2jZMNvBLTbus9CwZy8hgJ
ekzLP2V4c+NCVHZcRRJDSeoAfprJUCbH3b6VDdBy0XHjsKYLrSGE0dI7Nnfo00DC0GWf9GAhkjcc
FShmILc/S6ocZ49sH7xU/2ZYiRCV3AtSK4taEY/jq/M2o0rKl+8es5XqDm1WqkhwDM2YReXWYmqm
gl6aac0igXOsR4cKULyg3JiExazd+JSdYAwlsYLtHPHkbntN0cLb+eqyvdHTlu9xEQXNmcFiijot
7DqX7CRXJaaKMWlgTkmUGUHgmla/DSu5CBTqWADFg413tltB9107Btzy/XisZx8ty/oKW0IcQZaw
JzjU2/qeV4RSUUn/nQYuFrba64pbPkvYGpccOgRQkEeofh/mhNZ1ACjFJ2MhKIy7/ICrFturu7yk
icoNQWNafuuOU/CkbrKy8mMTIUlcSGdcWGlV5k3EiNKYedtIxOnK8kdYfDoaVz2NnwN5jpbiMYu7
u85K/MRkDYYOCYm6UJOUr19bnXYT4vBgL/on1MI3hH17X5JHqR25IisLp722JHLAd23l2Bg3P6GG
B07pMH3ElcA1aFjb/d+SVUZMbDmZPSDK3dvGT9jQAhyS/ZURcRnNqa/RZqspv2N3GoQeHt3nToTk
3psO4jGONgN1TVv6/qaIyTMrkBPFeKuViZIOO225P9CWHjZ820wUBevwfHKLFWnE2oYo2jIbOCc1
Qhrb48WdL6CNa6kzfxaTCoNSYSQT6cILr1omk/fAn6PBRau3VE2f3pkrdEfQdnB0Ylk4FAIiM9fp
Zy2I0NH+tMgMhyAXMyrHL4jF5NTWpjp6x40qSpNKnqoUX6j3YZlcEvUg8+THGD6a3ozNhXsco29p
7wwawIBb58vXhhJ/1VrnP4apOkS/HSNdCgeJumUqbjBRHz9mcrCFmH/oHa+ECQgPFxel1tmTCKGe
kXXjUTbVsv9iB7LYKT+/5uzqkxQQgcbunadZuUP0mpPlrSuC7Zt4B51uRl4izaffE1Uq26JGDpfT
WeGfsmTufPx+bmtdmefv1/iQJ/S0YC/1ZmNMicytBpAcXWhgtBvWrETqrk/f3IuGvTrhY6ZXFry1
WTPS2WCWbDxmi8WFXuTFMyWgj7ZbiConzLHfUECekRN1MBBcm2wUEGAyHuY5oXxBt/+YqqD+HvR4
6DLjYQjfIfscl+RPrpaKv+az0tF0sMtVmeQ9r/1CgRpXGrbD3VNi+YfRcXfh2jEyb8W826Xu91vU
xYPxZvg4CU+1XH/MGg0Hhft2wWCiiP3FLdliWqFzJZBg547J7w8ZvX8sPaOjA3sC3jYLEHE9ZWYG
IjzGiFmyBc4eDNhsZ1nshzQgzpDQOvJRt7XEJu+LKvZZ/g1MohOflKesH68QU8Z8aT4LBb1aCo/j
+J0cBO8I194E1LklICn90hUNOTJXx0nHxdcL4OsNCsB6ORxihh2RxDFocT/DFW5ZL13AGj+COQj9
ZyKSZpgQFAwkASaTIt+YRJpJJqJ6h5tCs1dhFkI+KJHLdaS7ACOBu+jbWb4EOj7rxCXNv2UvQtsk
NcCMe2Ej9/tVZzBdzNEcMyTX2AHmTHr0sd/4fmZCYUkBJp7Ikn80fDj2/EiV/PvXQXUV2C1r+dXN
++iUtnKct/bBK72LxmPho20J1At9fIJJLQZeR1TTu3TERg7Oe0E8I4sCPpg6Xgk4iGSHq7UhENym
9a6fG0vuoUTK/ApaTLv9vn9bdy++2rAXO4IGvyfm8HKBAc69OCPsH/6F29nl2Bd4xfMBLIcWm8cr
AEAqqNNWCKE3gz53kSsT9eNH061aWyL2dtikEnU8G7DFSczQR9QDHIIaSCPOtMO2nY0lCt806xI1
VbKE38JMekfFYfOZ2/9F45mBVW622yDvhXy0ATi1BfJyuZFBrzBPR/z0utByf8KkKK9EEUvZ2C0O
PPOUEDEPPoM2KBD4w1ff3NJjbwR+gMYdbz5fA9Noys/SxinAyn/CV15SlLd7SLi2dmScBKRCgxXw
TksxeMQFLr3YGhULbfiTA2x8XBzil8vGFeN32W6VlPsFYX8nEChlOs/jtqVVhfVqcPUGIbCUnyrD
8jUb8xDNNFcXlb+Nut4Y1FkkaaOyyHSbhzzy/Pp053w0MFDQplou3ahRGcw2/Yhkpp16Sm3ASRh5
e4jxnidym/QnTIuvBvtwWh7+EpKMpl1//irDjQnUYF62gdofKNsPi9ozVqhRi/RK5SaPHBf6v4cz
AvLNZE7W676d1DVrCxofOtbKXsyPm6mcS/Jmjh/UvZcB+iz46PLPSzYScj4xj9Rwlold/N0kZD5P
M5ND3+jIopJ+jckAgf/FBV69ckzMM9dXMZFaVlao/Alh11Hc3YPgKyrnoPfshRSyxH6Qh/Kz2kNm
gtVgJ9nXcQJjMJwSmtyxxUSSk7BFuh/LANQHL6921VtUmy+XYpW9ZU8T49nld0E21kpoU/+EB3vc
3B7pDEZeN3TCpEQGLNM/SdwCjBSMdZYeKinpjlcV+JZSmrDg0zmL9Zv3RdTccjkcr2hWKw5s9RwB
IfqGwzSBQXtGOPAZIUxyipazl2s8qXTU2TSSDoEWupN/PijkQHxPX8hoZZqrkwGsfHoSGRZEnMpJ
Yk3BPN7bHfDxris4P3vWmfntv4g7L1LyeMr+eLG9TnbCLbrNBl8sM553jraVMNdv1tnG8ykx8GUh
Ox0HW+Xz4XAgdCAUhEIMiS87OF0GaEamDz3xCQeUfrwuY50CNHXvIurdF+yT0A/9z5SEb6QWXWUh
1cq6F126Wz7d93B8ILp6z/VdmJ7/zMKJo8BzXr77a8KWMAFVL/Qi6Zx15e77wVGh837Y57qFdHEQ
N2+AKsroa7gk0iMcFH4cTeB4HTKkRA7NK/nZ+yYi2S7b0/eThEDunohYFUmsAHV6B90Bd8K2OGQs
uy15tfBzjK1rcwZC9KLThOKdIF7vZXIcpwieW70sD5K9clk5AMCMBpX6oqxQUgG916DncM5qvjIu
/9eruXFI1kSPZARjepscWEpswRAQfaQ4XxBOs2QIk3G81N4G30UGBVS+EpasLzK+QfsFyUXExNtK
1IHHyezlsWJKYLmatVzx+PKmE9ZR4rINSY6fTYjsPpMoFsy+7nID1FyV04lo/1NybYBwu0vlNeg9
RiVX6rVUf+MrkLbw4Q4ZOMazzOs7C7sVXDwCi3YKCGTmd+oX7+mkbVNnaFytg5cn2kokRuwubW1C
NGsi9ETUuLrZgiKHurAXf9cq+mkbmcbA/azlrmswpUMWv1kj3pQ0zJMewDKKrosm45aswQ3qSJJN
T/+IjbOXStwPZjGCcWhx96FWZ+SgfC9xNjEVPq/niXdP5Q5Nh4Er70eYlHw7j/h7R1FaKyjQEzx0
DhFiUjZyp4XomloeoWJdHP8l5O/IYep8oSN0ZWr0JsFulga3RXcjXI90eMEpJi5VPQoVTpT9sgt+
9W9aGSEkG4S2P2q4yMzj9eu81UG5iQkZ20NZQlVyDcMJRvi/x1SPDUnvHvYku+PiJGyT73f+1pni
ex0IKk3u9s1EXN6zdOAdho5n5nxh5gN+p4zpz8TQB6A1M1ZyFfU2YOv37J7PVU9pkD+6x/6tWwEj
uB/+tgG49LvdTM0Av4YWFJKU+rpW2yGizYGSQ4BKZM5GZdTYjMUu2OKbL9O0RLRO44IJilWTMfiV
aHBBtXt8+lTO5MeSNKJ5Oco9S9iK4wwIagE7xN+u/B6MT5nIj6kPB0im+d6t32yijAfes0mO01Ra
YAUPtbU5ofdyLfsGXcHTorilG6MUC9FVJKx12kWA50a5tUySyO0CwckI9Q1MM4G1s3FBIkge2H6I
XbcQwnwQ54Rn1Q0K8WnmrYzjjaHwwnSxbAN3QJsTQRpL5gpyFRz/V3r1l8UZ5W8LGXIxIMSt4T47
7gVd4tmUxrCh8QEhRtwVEpSgv9yfvfazcElT9dd32ZrSBoCRPQ+2xP+pUXLRpWgRxQHwBnPz4dMQ
b47BuTr0S/Z81LXia2H8t3OPRr1KKA4IAjnJAfg7/Cgj4pAYKq2l1pW8X2s3MjfV+wVF8ZG6Tjyx
ONvLGt1o2QI6Z0zKfd5eOppUsYCpfuAHU29FPZM2YSHJuTc4dZnTBnOd8tV+aSyGeagKfDVcX5Wb
9suhFikXeUHo5WnLL1/uwG/zdWtDXECrOP/Jpp6Z9cpwMVX14cudBgM+oz2BV+4LQiY/skruSDo1
f/1tTg9kkJVXUlPJtqliwsaICF/RzJq8FohTVTNQ7lBgHkfTjf6yCh3ToDJRVkode+xzBZ6pO3zH
GH0KbfLdBOR19dYh59vw1ch+xAsuWGXAY8x37UZ2hw5eM3bo1/gW5yq7Y1DtlLDkyRytULOaFj+w
TSzw65RF/RtxYIspQcrIf+E2cgyVJKrGh2gZUeUTGgbqyMH0lSp9g8XCt0V4L7X4TDQX2lkfss2U
ibJhvR35JBPhhB7N1FR2wDf67I2zY+SRPkSxhETKyg9HbluAmJtjxfzA1yfOAiBRvxOE04pOqjPA
b5kRaAYvoPIvor/mANLQ4bDfgkygnq327I4OHUGhbHAqK72cDiOZMLW0hzLKa3UZYYFL9mN58FiA
D6yXuZfUC87pdkbVmVOxThnFTBfl4Qxya3ETPb4o0gCyt3L3SN4HRLl7enrx2equ2OGNYlCi6MN6
wTlBhwBc1IlLpl+nSO876AGs9abfwISESSExRzk6PVCvGfNmmYvNWaqLt9A/JiEGDg+pNTfx162x
K89JJEoTREw0HdVQNj/pBeJKhAE2OuG/KO8Xqhnq2syEto5trbspnSgHX2Fo3ornNoiO3HdFgSrG
NXCZeMxDnsy9Zf/0TjScr8fPAAm2USvk/BYVWxjHJQZ0Hi91VuZbj6EoL/dURkMBNTBaK6k8uiKu
xpSaI210BzDj8H+ObCnTkHFa5885D64uLGJLEkooXt9OcZCgqdGsCNqtAuNOKytuWfDgno58U/1W
zmhkpm1B31HeVb7BDoHbdnJIY/ftKz0rSPJAJXWNKnBR//2vkoPA9HriPeto8i9OlNHsxZQYPS/B
zR62l1dYli6BEtmObaXtjTsRDtFT6pUv/XR69v5KOYu3dTUg2Zo+u/hHzkvGwh50bzY/OsJtfTNT
jUaAQ1B2JbDvBpzgWjEhpaNQavVhWBi+EPOs3QEnZficZhF5Cd/roSaC3Fv8DDKofkDKH7SZDEUE
mzuauPMS0+BzDHiP3fLj2WaT4kTaevbX3mwfUrn+Xx5jpQgPbyJJ7Lj/YNfMl0m112UhT0ZOVR9+
vae7uivLirlUIy/7PWPnVcgA8FJuae7/UJkJTxAA2HLdKJtwYXXehFEeIlXDXuOtdT/fgNwMoujL
L3Pz/iGTwVimCm8rDQY/8Ypq07RD+MwCQ6tEiUY/2ir39b5ZKR33OpuYiRrNGgJjGaaYlxnVDdpY
YyTXfCEqI04sbJA46kX0LOTgZ4niqXhXa0lsHPg/raMgJvfBFIkNCJVIiRMa+nVjMKlI7BnB8o6R
6Th1meVK1oirAWpYzE8SLPwgQsbNnSU4Qh6diRR7qIg+aT+NdmpEews39yUASd+riz18kfj0u21u
sAFKaHQ7I4rg/qyRboeJRriec3LKGrbfCLV5OUHB+6MYC4m9y5YWuwzXtinJ625+XEgSQU507o0u
N3VPJmqB1AQB2XThQUAkCmbHQ561+O9olMje4njQrMVUMPcumQmCiuP0KAmBScKMcYqay+/ZU8NF
B+768luL2WgHQe84G0d8Mr2zkym5pGMzs1NgTTcrCEZao6JdAQ7EBfNEq93IUxTipd7XBHVxqt7F
tJgk8emI0ViFuLphBGQTOnAUp73Y3Irt5eCsH5B9LJKIr5dLrmTfghtTpuFPWMM8lcPYxZJMYxSw
6ocA/ZBcMrey+e9bf+VHPJPAe3IO+aiJf9GMHRuW5M3CxBdvC3wHc/gam8x0fUtbwBVBrZAvLkep
j4IIMta4JSeJLwJyfodteOZ3BbdRvxoIbTfvtpu6NGLzIq1ukTb13IkozzE/q3qUbHpNFfTR72ng
omv4cBt98aF70FJ2vtdjAMgVgAUYYXzAyauAMLSPNzA7D4lEkGIeLRUmCaPwFgmvf0cxzqN7nxTc
wKKCMgIoyf/1VLfsKXYErj7pmYg92m1Tl861Qxd+X1HRoxuWCqNkMIKGvLhH+LRnnv0eyijrjaAC
ZXCl19VcRKuKGSvkTXC/eJWP5mhhYdUerrOpKRfS2fUEoiHDDXhRK1pamfR0GFbInJ/rpc6THsrt
g4iBuV+rTqBZYhGTTq9erdA1FGZ67TLbsWi14I7AnY8KzEq104UThNwcmGayjEz8IN9aXy3j+6XX
khe1QVbzlX/RvihH4fa0KwprdwSIrPkX3/b24c/vFU7gGGNN03rnWp885yEZzoLiVvw1mctQM90I
Pb2ytOdpZhRQ2taIxZi7dt0Jz39+//N3VkjhWhw7xBrCdcv/jrH7p8TFgJ5n6n4HZgz2gdIhmOiD
9Me1wiweBHLW+UCxMWyKfnXgVkqSGvp+fVjQpvlaQlBvHJQ2BRDoeDH48KgJr6i6nn6EdRxL9txK
i/gs2aA56WDpKjsqEd/TXn5Z7KUooLY8BgGVmJYKH6l0CoWYdlEtBpn5LAkLss+HOe6QPbvIRiJv
3XMu69QcGcrF+czbl2OMIC/oYQa1Y0cI87OZBBLmGtGeBVAkfksGn2uuOhS/+0HmqHdu4kyPDDvd
lg8xoCEl2Z2nvVAXfoR1z+ygbZPieaIMk4e05l88vRn+NgL9oCi5BTa6EOTu/yOoR1SScJUhQOTR
ZJfHbgUjRqg4FX6Fq+PWq0ohZqmkGSHRElb+jzdhQdXZGHHrSEOMXx1O7x5wdq/kQSpVoTzmkwts
5QVqjtDkeK4gb70Twd59NYHut5+8/lYoUw/vpKbc34bYirzorLrP28OI+tWPpf1T57k7NJd06g10
E+38tpNKBxrsGmEczasBJYQybHo79V9U9oHNz/Zo8JV3IMD6/BBHtnxueRwRfAXzSeLsBrOGak6l
/G496mYEdsJpeRxtxdW1LH8ElNKeljRZgb0V6U6cnwcu6ES2Z9oGT4LNCxdKPBbiTsqC4U93ct20
ugPxTjAQfo1HqWl17zR4bMTyO1bKr9bAdZ+MQ0yeMHGO2YrwheJLuSiKBxNaeQ+aofQOY+5WvDhw
o3Iokes8KYDbeYOyLEVx2R/Av735RsphM48yR1Vbe62pN91le5jUYMis4gTn0UmStEn6bYpyBL1g
LVKoRUZY9oi3XUdl2oUhDEr4DBszIyg5ZSXNmIEdIshwVTeI4JuTedCbD44lSTIwQ8Abcx1UvOTQ
I6s/cKucYYOZ8VQQ30MP2oWrsTyoa91TDktZ5ATJPxALN6+FWA7oBxvZUIjZqRmLxIIN6KE0dLqP
6oUOkuagXX+i9mc9JkyoobTDrpBCGtf/n0C/vSTuRHiQnN8hkNygLDF/Rvs3qXcNPkevgmv+lK31
XtqFKTmLS+hcVD/DgvjlNlY+0TYue59Fjx6ZDxSubnm8YHW8wpCC6SNBuNmzXtdz23q4SdVY8SG4
bnS0dDHCeHlO2ch/rPcpjReCOD+BgnUuMoXmgopIlBmrAL8GhiJcOTlDHcimw4KyrWemjlzEjx51
OaL6xoes80ekQIRiIPp2MIHtJivhcNz+MjX0/o3yWfHXEqQL2PeYVJ2YoTmJnxQ/HpPBjA2L2GUI
//oczNEzGbrceJB6AuauOPypnNB/cIAmqk9Lr1ime6kNHBYMzZwyN6rl2jqx/OiuBLpICUQOlFl5
xkWOHwgAhE9L8tf/YzqXypl9qoR19WCkHpuz1oPT9K6oAgpFwlQTI7ItXyJLzmG2UIShHs0Iwxy8
8z1RKTrsdL05jYlVQVZEfJLGllD6/7+UIUC5vyJ5OwWyz/2w2422jtCKKapM5AMFdHC3Bnw35iZ9
JNyetfIcwu6GyjUrL5bv++3HcAAipW9kaFzgOc+c/fzuPqx/laywflihOvV+CdvX7FDGxY9JAQZb
+c03HvEfK+EbsF54QN4e+lfcWTAiETSHBotaQsmBiHZ5alpuIRNCWnql3bX2zA3O/WRFLnThfuv0
P2BT+IF5t2hxp0332rY7tWwt6AHn9uw0Nl82KqzYhECI0SW26ajXQ3r0sk2js/Qwsr4m5PuvRE8B
mO3PHwn34sXBBZctf1qc7aiURsvsEz5glaH8wviEs0yc7YmuPxF41OmzoW2EMR5BvLkFdCfUS8kP
Mgp/xO0bNYRqegLFfUKg5vXD/TdZv60g6ElNNjoqW2IoIed2EeyA38qCujv+flt6HIoesF4K/Hvo
G9y50sbpxgpXS7OxY/jwAu5+5WtiVhjj23ohhiVzyzCylAq+sc8uX1D63GMyWiy0GKRXJueQYjee
ZhPDnGbRYZE4vctaJpBF4QzYdafuQBReNTNtg4QbZp6NDZMWQ67Hbl4xvjLMnb2isnYN97PHld3n
cLv7T4G3bd276yW2T3ZBw2DdpjD+vOY8VL6//i0fizvQIOuiz9wwuXhe6g5fK/87rlnzy9YDei5f
T3w0ORFIYrMrKKYjohri+Up6m5614SNADelxRxxyhXNpyYwMjCbtjbNkpNG11SMlLUoXOh7mTK4N
P5PON9fOajlycMm+ZAbT+cVarrHr031nPGE+AL1jnsuWF5It7IZmJKQne9TjtscMoHfHRWNa04Hs
skj1sCAn8ZoDs6n7usnfYkQcRUsZ7jG6RtKQCU95/FvIvUNgG52E8A664baFnyClE5Jhw3I0DIZG
eQF+yltnPKqA8B6rOkKWsdvBxpryi9ekQRNESL08FLaDwjx58DnMZKuzJ+Zhb3nVeP6CTP/rolEQ
6Fta+HoDC4QZAcqtlJm1NUE/7weZX0t3AZgvRLYkKjRW68dnExHrcNvxZy/F7CEBRBoenU5MmfwG
3/iZThLCk7f5W2XVaTCjsJ5prG7ggjI/vhSVmhlpwHvB/0NlOxQlX4vlMGWhJ346XXkHKUQI8O5w
RWXD9hoXUwQmZYmoFqv+cOTb2PQ558ZGg1HAG9ISqMj54y2aiShClMJn5xBunelRHA6/CzSoRT4A
Zk2LQt1oHP4KgwUJtVs/33mujLhFAV7h8K/LZ899f0pVNqz0+6PXBY/iMsF3xpKD5f19Zal8EuJ4
rhf860XdpzyKNZbWv5kVXlOeuV/W3dH1VAS0uQmVesOwN7sXs2FlMM6F5+gN0fB+5+lTv7/ZlAFA
43LWmjusF/d3JMGzkOY9WLovjJWbucII4xObyq7UQoD3a96JDP/xuCbv4Btk0FdPtjlCMglbXQnj
yvM5LhsJi+NQ3wiYHQjsWp8IFSqGxqvO9aJTldWBiwxTqy80JfoYLFAdnwcs6NDqMJIEOKnIBd3o
CG19sxx2uHBCEYKFxfVakmIdWLXzB2CNtljBnkv4GUoN7zL70AfrIXgKqxtr4hOk7pz59EtRwGOE
eY879nLFKpa/blwFhIUPtELpL6Xk8a+KbPCiAFc9Mhkw3vtp5Giw6pN9eVq/V0eDeESKtgOfxTe4
Rq4p/Dox1JXwDHowW9SepgGXGoSgz7CKoF5MUMkV5XsBcq3nUMdLOdpVWG1LnSlYGm/IKbZrStk0
0SwYNmBuv4/rsIl0p/FIuomfD72y11c+6azGmoPuytprP4OaYxa+PwF11V6GaYp7RKDrftkQh20p
vhAZasUpGPzrQkeuuwcHHcXhdhP42kSmly0tv1J5gzLqZ2sK/bhTuQdxWsyYbkGdomgGH6FEL0nV
9Abgl0Ufy9jaIPI98A5C7dYRUv1ljzD415DkOmxQd5iMjWevNktQs345LM/Phl8sGqOcERCs4A4r
+QZCYqxlLK1EzbtmWV0djwB42CWvQ1F3ye0gsAjhAK8C49Yprp5rQfsPOUdh3aHeyeVj7sKzfmZ1
YfBMLsLZT2yXohTh0SXb+DIW3tacI/0zQmVn+R9l2yK/6BrekH4l59AIdcVLip/PkM3pVU8Z0fxt
+w5L2eSlXuS37Y4C0LGhTr4TCoCfNMYH0MDpZAe5l8BE4oR202P/knG1bYmxpxo8LhgWKdlOgXLc
nxEgZaGNBuMYgsbykcXiEP88gJ4yxcSkrYCg7ApOLx51Wr7YLeHuQbt7jfg1RTHdqkceOL1QEUvm
i0KmITIzr6PIFeUGHIJ2qRBLBAidcQtOOUUpkDbYLcZpF5hTisCnRpnpL8fjoVviBsiarUe00B9j
uOv/qqp4LqGp6qOdqkbawE8+PKcsA/YpTsP0XYfoF6uQfrPgTrav111QLccUxlQiz6DNQ3XC5S3C
Xqe0FAJp+6B8aw8k+L0HbrBjWN0t90FUnqFjd3V+rO3r75B6hjRE6H1N7T9iADP6hcm/JFWfwgE5
lJK/IRVZN+oRzu1Ejr6n3T5Bh5Y0uRhuwuyfJ7E+DfU9ry3zHVed1E1/Tyqt7syCKzXwW+eTwhRG
a+kUM0/Cly7EUnaC8F870KEXuaJgu8iSxQEZ4m7VTRmjLIpLsdPy/0IJ2ZdHxm0zpWhbWYoDvlSN
47iLO5Pj0PLq8XRj/w7rtDiukvPyXoe/MyggOujrwim2in1xvwYV0oUd2RQ1E0bvCU8if5+JX3dI
5d1jA+cHZoVw6vI6TI0TYgohgF59uFbgjsV1+Ml4hcOtyoGInwgIw8qtSw+TK16rfkz+IJtTdYB9
qqRuvaGlpSH6leC90uDtwRNfKaXTr4gDY1oKqAliOGcgq1EtYsvxLRVcJaHv0+EuD/h8MdXCfv00
UWl8I0CPXEfJkrv7aIE4N6NZ98k2uy6cFYbZcHnRaoMu55Gd8FX0z6syi5OHZC5glvcjDCAqSqlZ
5C0m4fyO6G32KcCwJ5zcP9Cj+xNJYiGFgSQJ+dOfV9QRaIFSlfptpigeeKQYLL/2h6PQ6XZUzN7G
iAHVG0R89/LxiZskNz6F4Rz6po31GWOy7D6fUAVcf7R0vSCCzi9v3RUivyjo+Bb3RDE4H/94UJHW
b7J+taUAlblDSSj7VtENqs9ISuwYJAFS0Sf7fy5pg0gledvxwZgd/OW7ZGdwZkM9S6ZIlHXfbn3V
/IyKD8zaRxK23WF92hNmX1o+m3EC/dgSdbEwEpRv9pM1qx9gSQj0Q3zvcnN5CHq3eQo+hk8MPtZG
qrO2QLB7a4mLrIwdQiVCk+4dV55xW8aIb/8ts+PR7Ja+KXUarKF/9HMEkmEfCL1AND3lF/b+rslI
69CT8dN4FI/jllneWs2S02mtfgUXxUxasKw/cqSybm2YJAdYXh9kCz2hP07NYiIPk4LNvlQEsFmR
LM/srAy83JEvxmNZN5DPWSvU6aeyzzQyuJFjNl2EFr9ji6Wl/5mxq/GBNP8MvX9cYQLyt2Vb1D/M
A0vE9ocQk//khnHp61wYlB/QJ8KC4ZLXSvCwDdc3V0kHhB/FoTtU05jhLgT56bNbEv9NPrZY1S05
91MSUtzT/ZmJKabHM3CMAfAIOy24iz9Ce4INJcxN/PCogwq9Z5ZgbYBsAht9vrMzHiuOAw1yeeoU
kcZuNuudz4nMjwRtKB6vHdoq6H/tnUVAq8PkOh/DAqnNBTxh4o1rjvX/WJquynePwguDpMgR5KM6
mDc67wKgEIRF598UDoFCk+POYT3BnPOxyHW88pzoWRjhhJ7Lw0sZb7S/peVH4aDxwg8GAKhJOGEu
L4g8ekl5QFz4T0tEQWvEtz+1jIa5hM1hEgwasuB4MMvwsh4rBqJ3ZnorLS77pEL9pYr3Csj4qhs7
pjyxmOhVwYKD8p5wT8NST4KhwbOrEmCSRpc2WpPCWnq7rwR5cgkVcEediJH0SaEg9ryRwQ9HdLM7
3ZlZhdV/HdSpxVvy8sb/mWVZXs2MZkTN8vOj1vvSQ3Yq9SO9fVmiDPmX4xpzeJJrcps3GY+ALMKr
9HvqFVstliWSs/sE57u3HORFBSsTLPdIIuVCMVMg120d6SXZm3NpKu7d9ZkaE0fjN+bxnexqkmu2
2Md/iOh4aEOOC8n6kfJlSRayh01+Nu/ETFg6gLzdy0gcLHuWfxPkTUumRtUgVuBgit+PUUkrcxWE
P8e6HvxTHBBvWKJHfM/gSGfSgXR4ZLPVOoYALjVYgVzKkwcUn12ogH7p/TbcLUWMxAacvTnEmXEP
p3KCvthSORfYKhphTVAfRsHIVIeWtxY35lNLoh2gQm/4uNcN8QCqPADlhYX+LU9BAGd+TN9pzCaB
wlF7E92p1ujj7sqG2xQXQVkCGUwPgUesDAxDSB86mWuUmL5M0PHxY7CCdXUXhKNA2OnU88okwsfK
+w4IKoWIOGujXpG7Ru+OWrpL6q/92eeeOVRFR1+tEOmXvaOwhQtPnX5Sqik8Fg1pBD5bYQUYuKtO
PYFxaEs+AIPYtwdyampfZX5x2AX5GppCsqk3i9bpoaldrgwGzjQJpw/isqaIVg58V3AAvHOP+HEn
9zldgCqcDEChX8BBLbqhiUmMWA1yBo6dvttDon2qIvOEF0r5hIKQORCEo1MDPFCGJnDbCP9lDNZy
MYp0OKFNZeo4cqHb/PcCcBQ+FFNT7SxlaQ9+WwINWKXt4we8n79aEBdiDP0wwoTnSr9mX0qxnXmt
DVCqy1DlreEt6DGv8JMKaZasnW/8qG2fkR4eFnBUR3m8cK8bFx1HOuurEYluNgBAACrp/cTuPDOo
gN/glwtpRqdV9lsCD1Zy8ZgzCVWKg9J5TDu8JdpuQ/Njm+G9sGtVUsuTqfzKq6jg2Px9DoWU3tc/
blx54/8EPHV14cRbUq39e3T2B9GUJljQfrc298Ns+nM7Dx19H35vK8f6oMe8y5c95Pr5gWnFDQIC
AhdHX/tVcMgc7HVR/zk3H+f1xZ+RQEyce1aPb7IvoeNMGMWWdzuFFMDHx4qKiPEGxuewRHJm8Jmz
Gn/6P6zuCWIuS7f+3k04uzoUYU3ILtOINm5L/+HH8pRwFa3CmDyOrEtjfnMexZljac2m+TyadKj2
IHjnbzR7T3fAjNOhimAy2o4bScrytyGUL0KXMsGvxuMiqX3QJ4la8Jg0m3nVWpJWKUxlkZQW+u2J
78Z+szWiur3/67ll1Y1/3AfOHTzjzwpZhtZbS385V91iYl3gynrqB2mD1Vvq2t4NE3U64ebGDbuM
whcuXck2qamfZZ3a6Cy9/vpPLDqNhAMT5dJNoIlxaFBbLdpH0oUsrrv5Iak0JfthBrBXMCEnnE1Q
sY7y71bnM4dtxTkxle6w6bp5VlIIL/0iFk39DJvCK/6fxX99hv7cDhTm7BE28PW7TPMWJrUlwtqk
mw0JbNUVOn6SIfiGiY3LefPaKs2go9rnLx5+YEzGUC4wMdvsdDFotiGId2buO7PvrfHxNl8QPlJi
iWnoHbhtzN/No3rbMl+CO66voVmwXljNO5kHeWz1eIY2Af4EJFI8TFuiNE8wamRePXhPuyeQVi8o
mTBYBRIUR5lsrLOdYhgC05ZUcRrDP1X/TI3XxBBbfTAxm4ldj1QJlBX9R7cHeqShe2p2s1wDlPaK
A3WZISPENbRqKMCsK92YTxEygB+WNU35C2ymEIoUtTSgtgU+GA0MGL2hnLJ/FVCh5vOYUHFW55aX
YMu3rjOD/9aBCUuh58dMWHirPeKwJm4sgYbOj2mjlLsqurvIMddw69U+39WiFol5FJfJUgwY9t6r
Ldaxhbz0qxhCL1CjniZzvo7ADkCI783tnteeb0dqgdmmL7U4wLrTEg8sRqlKgufqR9NKD1QNbceg
opq+yMeG0WgAWin3LUIjSbTwDHjVzXK4PTaXhJPwFs2w+8/QsYAvBr/vsh2rgp8U7fXeKSxg82rH
585wmrSeIFO7hiJvmRmNb30Pb7HeDXnR17nSyga6QeS4QGs5P+H1tdvFrFoFFtYftpfK1M5DJaz3
OUx+Po0ZYiZss25HaQDiN9ZTlFF0nftLDyZ5F9lZs68FrnFQskEh9pZLSjnfUttiKw1bMpzieeWo
nXZCpr/23anYu8JEn6KU3WpyN4mTW2YINwc8ml27ot+ev739fWeYbmMRVAQk20xShDJvykk4NbnX
MFlf0Gz0l3r74nbyxfBy+k6WXIKO8eD3XVlMPNOzdsSAsZ3kvNaED/qtf2GIfNGlQsYEt0gQasiD
tWtYp12tFTG9J5MyUmeh7qvUIdBsG85r7bfKH4JIBCZzRc4S7cQIH7i/Z2QySau+g/CoaTWCWUpk
eVHexQFIQSjAuF9GlwkeOjm8PBSpuFi4ZVg/J70ZxRQQBGCsfJPN5nqzo3UFM/z5jy08Wm6iinig
Jqhiy+k6ACny+UmWA1EaqCl4TA4b8JT/71n8icoFEyTjkOcSmGFxM0y2JkOqSEUoForZ4zOA9Phh
Atj5mwiv5L+mX3dL84gebvxChtfWzpk6lY5gU4MjsevBv1+w9+y4DXgFvFJrKZdBKSI4sh61THSO
NrWV8hqIFDWJLJd4GaCeAGgrh8kLu8rKR1ydcp2d8zDumSB/XGn5XeA2jhffacccuKnTewXay8Dk
BJB+qsVArBHTzbWQSec+OEojyEBogGjeYJxVgl4ehcTBF6TnHBpj1nGmeqfzP0+Us6cIIBOfVYvm
1JqoefjJSbaM7PcLgDbJuB0vmkmYGBUtzsuy5DiAR3FP9fS/QcAsD0gSaTIvI6t3pqMBMWHjPk2a
D7MfN71stQ4k09awzGou7TyeTakdAVLdY8DrNj8RRzuT4ig4iGU60RhFT8T6Ahy1M7v5yEHGZJO2
xfLSpRIIXlO7JQpYqu6U/11e8C6g2ugjVF7lPw2VP4u7EjzIjd4mvUIkLVkPXsso4kSOgOlo6xZL
ga6P9UuopaytdB0eAIwCjYbeG1r1dtQgflPNiG55dU+WtJIh7FsaCPQAUi38aWF8de6QLw5LTAZN
PieWIcrV8iSX/qe1nQsSvQ/9z+MsC2F3yKS7Q13Rwj/JfRjikQi4/dCysdo4LwuLA17hBqkrCktH
+nVI8QmsJVNXnri9YlUy9sKah4RggcHTCbcwUEMZaqB5C8KjTVR7UqAyyNKsNSTVxIACdLjQB90D
mYBYNGQDtxQCIs+OO/msytfr0miAWEmWxJQ/d3iAFZyWvDCY10e5q76xin379POc9jE0KarPlYmz
IJb0X+c7mKTvGkBcbxyuwK8+xeA0JxnryVLH+nL//AIa5K6jOCUOe2cBFgcVUoMkrl9hRULK607h
JUyLezfniM6yeBHOXxD/0eaxFWMOdxzCHcivHi0OCXcmw11HQXbNDbFJxBsPsLNYOML/NMq4dxyf
llGQAZzl7WYHUIFxebOZ8GSzJqnvNWoEL/sl8x54+jA3ZMuEVfi/RjzQ6GvpYY5FfNyaIqWugoRM
BE9QYuEWUn6FZtHL3VKKYaQtY6pjiFjeEKoBbumH4tHdlA71sAfT2ylD1CbH9o8lCCwiD0/BNGTz
IfRpyo9614X5HHXiBjlZkj54ii+gyK3RLD3VdvWVin7/l6Ycuu+ROUTmssMH9B7E1rAvL0AewEGf
gvHKQBrmvd0mVtK0BFv++S/0EJnBAXFj0w7IGkVvqwU7eFcjade/9LOpDOwdrqVdBJw6aZX/Lkrz
E1hlZuVzv7MfvORYTxxaLrMico5eg8XYMuJz83CrWJxgZACXEGVjji4PThOEo69dYl8reEPOPFon
zlFCRubjMPskPuXZiobq87k1GjjM30B3v/QIKT4n8r8luJ4mHCVJts3nNugBZt2PLb4LluqVRSqX
LqHVWH31S1sJttuD2vFEoxA/dsMHLJBBjqHnq4LxCF1u+eQ8zLUAcTf1KjsSJ+LYSg54Hlci/WJu
X3aLmGdA3I5axfSqfJDSpgzmKOsH2KtXe11ZbuRopKJmPF5cloreqVoUBehQZE1Cu+AIdCLiIX8c
32BoxDlQ8pi+kTZFr5AG3u8GXcxjRdnLOGBQFRRAW2zge44bugFUfqljANTeVk85m1eAJQuE98bs
qjZEyvDkzNVCTMcXmUGXLUUvMadmmfe/GKXgYJCKz7EEELDDyWQKq/lJXayNIJSuekyg3j7s8+hZ
ViYwwB+8s6/aLUXgHg1TL3yn6bwZpeyOFKnWY/M9Pw+QaG238xzVa3UctqfSIJsefqDTlTmWNClu
fRPzpeQUNZKFy/P0tO0GFclgd92mNJzD+GtaOF13Egeq5Lh+9Xhh6VJRjxPC6Nk5pnF3AayAvHch
4mfvfz5h4bhYbkC2hauRnm6+An5bumeQoDSoqZxGKTTlE1qoM8upCtTn94OBT2PWbtRrb8XoGycm
iRjn9rnjzV7zWecoyUg51s9m3NEcIbXVvEh611bN7rtJAViwSrCDHCPprRzIcZPcHqiRuSwl+H0e
7MTJALQZHreb4sARxWqGuZS9LwA2QJmIT5OjFuXOPpBf6vUi4MZw0aKb2AqAdS8h9wfhN9caeP6C
1Nf1NI7CxBjsyUnByQDRLi+kxzm80CNePa0mdBOm8HlqHM7HHgqc0u51UOniaEk9Z9r8+34RIKxJ
jfHz5SjuDo19VcDcJwhtAjsTyBiFv7PrEOYx0fQQbS1yok/m+uIjUZrYRXSMdPIWM72oYzXg+gxW
P/lqp3Q0lDeIrghxvwsNIDGZWrItodEcwijL3k8wNhyeXmfPWqXn29QOQt/x4RsY2c1xQnDYKODm
uqfJIiE1lgSl3ICenmCOohdeJYk543SAtunUPMFFKJpJL1d7N4OmwqFBR8rIjetQfXTUrO729ppn
DmVnMxxcF2Sn1WEjD+u8vOgqRdY14ynu677r+ciHEepV2b6h4nj+ddAM1HotVB83u7jLbZJxuLqr
gLv7BL7vwE39rZOKexLnrh4skW0ZUa/6b3RxGnINfVBEcKfc9Z/hOqK8ZvyTuSdaFe4qUEDTAcUo
9AFliHCeB06IDfd9YBER3DUsY8yIhv4JQy73jynGraPhF5p8BjW1Dnc24nBjv382NZe7hKzz+ODL
+sizOXnQGaNtu9CNVTo1HnzgaE7ApH3+ADb9/yBn/y/NHihV9+D1mAXOuuZLzEnh1vV9djzyJaIx
gOrRkRCQKSPa+06QNkGOYQso58SWDX43gtut5WcW/9q1RUehtQUn6ndfVBLNKkxu9iKZ0tNJD83r
wVLIyVoLnOQGkTnaLEY4qHXi5l9L/yNzmGsOy9dnhQX1CMawKeMNoWp/syxuqq35Z79FdpKtoch9
lKENhJfxi/ajlQjHaMizWnQlQZjmfgbThs+Zx+Fv8eTWrgpgSRtHYrGa0BuGR1WkHyAHKmnyU3BZ
mOExxVJHQONR7inQP/LPsFr2M1z/kMVsQt2RBPhX5leG4FxlpqsLkOm57MUVf/rJE8L7f+4b449l
FEYfXJgdBKxY3kbor7aTEOeujjLv1Ji5t8mY9z4cI9IGU27qtyx0jxshYfiBKH8nc1b/ssIR289I
5QlYl7tquJ4GkAKRb8ios78Mks6QVw+1hHY2/QFpopqZiXsSoHdHTEbxwzFP9aDnny15obk/cmH2
/wV3n6IeLWmhlzqwdprMxsRsdV1zgVAMDbWE7km3bSykUCP1vk3LPBkIX1+TbSLDbrpK389wDcTg
rRSnPtEnVqWYRjTrehL81bqvcZr7mOhaT/VR/Ut656XzhtlenL7h+Bzl1zbBgtxE2ZY2yw9gLN3a
ZTnyeaUHG7ciWRntjvXGFUKegiw1aQO6oscqk4EQh+nKBcxazEyehAzieQ2WpmaSjNvmXG0lqpdN
ztYZdpxxJiZkG2hwuf/8ylXaHIIcY95sByl4oKZWp3VOf89Rt/GM+djRQ9VA8hSyfzyPxZcw7HZ9
p3/qlv2D2Sls+M67AO2R3jXA2UDprlfuJurYZqsXYeTbrgmR+L2cjfoss62mFfzQoobsvuak/WjB
Hoe4LRw1Q+yWmZFk+kY9cvC0ZDm3WvEAXrg45/6eKDu1vGwrdkuaB2wapOiHItuUjLlYML9EJ29d
pOTlqwLM9kEDDcWEFxRr1lmF2XhLVPbdZav7PQKynecNOaAUD4noiFu/0sxFlwBBnGN9UBOQXR88
52l9g0bVWYHlQhfb/xNbSi3zi/PW2EHBQO5Q68j0MbFlxqI1rDztvhk2qDskxjkUEb8tWwNyBedz
SVi5cqtO0xMiEtC491cwnkzg54BLpj3vTgAc8rsADB5EVS6MmZids/6WSlxgi7tUGAs0dbe0mtAN
NjCccUzIMRLDJSiEXQdrtiq2/okDtVOPdpYF4Z4VgTkS4MeFHgveqxNiv53PRvvDroEh2jXFntxw
UTuf5Kq1f/acPivGsGFqoZ0dgZEC8Q9+GA+Z0Hiv5orMpqs/8R3HHxwasIRL2EbsmHi2kmbay828
t+5/RG71KEqCIC+Qa7o7O25KwKSO1Zqw0kffIf7LGqOG3iWp2CF0ZmMEIxzV2J0qESZlKJYQB075
keswoMRrzExV2PvPjw2mSxofsL2Pi3KAHQ+XNFerEFgvQkLGLrmayvuoSU+vUCAyNHWiSPiU7Wnu
eSGQvtk7ZQYjDQXy9B78JefpJ/3vGhvEMKdKQpwOikGRd/mWltKax+tTtHLIYkulbBzii5+1bP36
LrGiVBRVSGg6TEiGMrXUSQCfmPm6E6m8+NS46BNxEGqYkfh3BJL00T4psgaLVs1LxRMJdB85YnNQ
fkegx0zgvDgkvvKdzfbx1Y3MW9rCGFo/+ljqVJGCF/T26LFcE9ZtkGHi4CZIGL0q4AMlw5fia4ky
P6Cwc5RF4OhN3c0vQWVC+NPbMAm9PV1mi4rs8R5fZYXQIFHWLoGS4zz5dMWKgaFk9YewVHPIcsYX
XNJOmNSyhql4ypFwF37eBmwwoDeDNIag11cDY/PFU8AMczpYWGo6ky/8tsZpoiZ2TLeeaqSkRDpU
g/v3a8+0Zis1qAXFVyxk4dp31heX7LDntKVV2yr5UcfWoGcXMWAxK5DA/L2SKdZ6lYIKFbOvJrTn
4WfknDR0MycCIbO+LPo3WuYlDhz46zoPCNi04KewFw9aCiFjqwGOYe2Idujy9iKKVLIjzA+djaA6
bdCSZJsyfJhDa9B6v/FgrN1Ki+DVRBg16Jl+kb8Xq8Zeb9CnZek5J56x1kOkP7S1Mx6FYLqC6o+M
DaR+I816OM2ShtWHtmG3y1VM2OMnj7hb9z5l8RwRnZah8mQPN7P41nJAiws+O4cSb517XOilsfr+
Y5cCuPspJUrwylJ5NezShUMqQeZFL6hdAaCArFciNPwHcQE35xWbfW/ZvwB2PTbGujz66dyajnx7
7do9qiNrjHOld3he4yz/2nHNxIle1u/Wv8oSX8j3YIr5CERLqW//at4iBYIJ91tuIGDfeRKR+xHP
ecO/8j5PHcFDkMEZKgk457tH4APim/BlFKqqNndkqpngExld+HiS91NtV+qMFjjjlMPxfNL3W0Kh
YqLMTVrQBVRL7YQkmBGEGR6MjgyyxElFXElXtx0YxE1PxoWMHS+nkkZImN+TpY4ZujATDt+zEYmP
YwQs6c2dTrxrlSopK/uoxjNTWyf/vnHHvWyHaBSgWodQnUDTDALEhWd6g6j/3B3XeMxt87vM7pRd
w5+JY5Q0DKDXQ/lPiAjUX9V6Kn5L3Ft/rmkhZClKO18RfRKCosUlfMB9tK1UBFPYrWxvG58IMC5Q
Nb1GJg2TJo6WU5jFt7cYz2mkAcynE4Yndh3PCCjszoEYuER1moUa3pny76QsJ+qR1/LRXAuKSxD6
UgiymD5gSGNnwi7EkepDLXboe/2amJGiRtwjaGrI+aIJsPfPRe+FxDWIMpzkUvYhMJz8QorJMbgx
zbCLw5+2EdxCL+UO8FUMWHQULaMt3Dt4rpbvtntNpQDpeyr0aTtjnb0ilBCjRGBV5L3oyHiRarFw
YZQEJ4eFbh48K6pvR5pL0/9LPIEieHWTTf4IgRm1n8Jr/vcDtYvXU6to8qg7N2bZXvsfsJX3oaNt
Z6i/WYHmho94OxmcMQ/820b4XcSy6je9l/jYM3mKs+AgbybE1oe18Oo+KCFoeJP9anSPjLeuOW6g
xRP07rMn81HF/eQwWMR1L/yQ1IQOuBH/iff7FNGBJ5a1Q8zFSouHWDGnmlfwr3S5s2DsaTcvlDSD
RPfZ9EedhsSB/spMkxTCdlhIdN+3nUaFYTz7yxSN599Pws1jyQOP9uia2BMYapbE/+5/VpiYXdB9
WVgj9WIYP8GEDNIKAEjQ2rJLYHO+3JdQ0yfXmzfHCBOKQy44ABWT1sH6ucQMaLEYhFhVdmQjcNHC
tYNhQFo4dlxi05Kz6i1BxXNeg5puCeoruyWyjN2bIb3U6oJyUaFNL52pzzkIdRV8Tw7XOfKsiM0a
/TKaXwEwDkdqW6y1lIRan+lnlMq6c+IjE3n44qQcB/1E3XPJVAkWw02BOiCVL70fP/gXANxs+4We
wLWmisn/sMrrNji6WcQo+49gdF2CvL0DUuztKkt6OQ2HtM7YbbxOFCHiS0SOp9HBF40E3sdz2f/M
zpyyECDM9n06gUqa2boeJ1rc+AJZMKzxL3Xy0Zg14OafEgvvQMRgRTW7oM9i4FpUgeaZPINcYJm6
0Nx5bsNUBJG54TWVc9A5f93n5u23LubwtMACO6DitEUGn0TdeQd9kb2r6NWQVUDYQ05I10cqhCPH
u1LSI6IABZVXos1r6dkRGPpb7SEpv+6yLQe4eSn2c+Q1RfMthZpKnnmIXArQ4Zl5PZxjnrizZfZM
DcSLNvuwUmLHQBvzBCp4K5uWhrpANE3R1eGRuiUGhTH2ZyU+J3DjtBh0gOuEm9yLT/rYh/pLjxuz
ZsXRdizAu4fkcaVS9Ou/pXHDCKp6/1OGcdINKxQVGpNa0JXc2x3c7DMIhixBlYF10pmm9a/u8hVi
TWMXawmRFb85fH8TeziTT8ArayMOV/uQZYww8sR//Q8vlRzhah+xu9yMoziY7A+jy/gEi3eJ9wY2
6rskfg2BPOmSf3iCZLPzzMGLUFlmaY8o5A+Dm4ffCrvAj+iLxNRgca1afO6en+uTG0d2aWxPu46S
WBYovHsp0HvHgxH+bdAzbpg1KjYiDZmkvkTzaYCODzKNPiitejEn0GQ7aRdqpuw2Q5g0tzfZ6SJW
wRRet6ojhAIwSBaGEp6Vo6flSaANvHSDsLwP+zz33clF+929BmQSm47hRVVfWxBlh5dMPAcGcysx
UsdXKsjN8aKHbQb24rYPKOfHo78fEBcuICJN+snJneynEHmrMJHc5JSM0GEKh4AWHFoxtWHcplgS
ptah+6p6Y8P6z++zvA7bnrBMudZlnOMGu399PO6dDoaY/QgNq9wiARbku23vAxyIXJDxKyyOhqyn
uUmljiN308ZSiUHdYDdAxYXZti+nsNWsv60cDeal/PirYzpj/GTAbKHdspkIgd44sX6oOeHGJK54
RFrov03jqEBggqsHMDE7Ep2bmnx9dtELFTunEKZNm7LCnffv4pM4H8sAbKMRKuXJ7CGUoql07A82
b/Pst096HMPDq+gJHeujl22+gSGBZ8A6XNXSAoub4qiVFpJJgqQjlN4axTGMSqqZWLyCpDsZWKfJ
jed89zLxkF/YbZwvfyLRJhEPtBi872H5TcKPOKDeToF2MijcqETcf+GQ8DqLqOOUX4iqDNj7GULI
9/mzwvjx/JqHs6inFKvpTCX8qx5G4qN2rIgN0S1s41sAaJQToiLlVOXizPLSFiEABacy1Ac3Ag4F
j8pMWLvTLgB/f7RE3zJ8d0EyEtciCjx5hl33sdDI4MhLQMtyBnXaaxCC/FHCo0iKgP6ImaQYsTg2
mn9KO/2TgZ6gvu5dMObXOt8nauvDfElFJOK3xOUErsD8Uex2MnWGUEdvDAhkTwRPPjfUr9j85w6C
MCcmxtxJs8oFSENzD9o9lzYrifX50LbcuF68zl4NvCEciFGcoc5n0yPU5xNA5pjYj31VexeUbtig
FHbC5JhggxaFmuyY3tagqAAA3WtkMtwGf8xJBLH60mHbQ29B5p1V71lldPbeBxr+rI10deM7f37D
eAoSnlTy+BrKJqtl//ODMzxesVjZmjA6c78wazBs7o/o1PxD5vn9H8hXUa7VW+Amas7Bmlv0rFvE
pO/hL2gYp2eaDUgDOXMIgyZbz93Yp+vfuKs6K6Ce4M/mLZgbdMWaUZd3t0toi6T3p8SukOKj5/6I
KW9iJzlxbkb+VLlXwPjz9ewGpTzLt7bwdjzWKof3pQ5Mi1p4zVBZQAS7crKkSoqBQXCJ4sdlljRQ
F43Rx4sPH9INfgKC3thLg7OO65D715F5y8o483PQvP7p5edSUDU23JPNZIUEUIEPg6iQTqi6VevM
znHOiU4f2gKbCDursocK8Z1rID44jLS/PHYMykRVrD4naFdWdMOcndboWzkmX4DcZCtGVwlSFFQi
zAoMyXsNCOieaeS0+ytNW3hpQZUvrE7ogXvqgW0mhU0DKnER08AUuNEaaohXPSTGl5nlMaQPVkOH
wEzWNR5+rvixOs1iCgeTq+dIX8pdBWDUNRg2oLEZXpiGB1dkt2C1I5lr6rC4xiXzXlFDwPkscFNV
klFtNp8sdJl2g966VaSDAyZbidUPhRdrmf0UGkGtW+VRSn62VJpUYhK4l7ZCPhk8NPpKUw9g9LGx
eYE+r+u+0rYBGuNIw6XfiCWlUcfnW9LTlC/OKIOap7KJTMJSwwQ0FeHTdV2KMyXcZk7JrsmmHVbT
3ZdV2ARhgrab8O9AMPeTZLvsDVz5Nb2O1V1nkO53WigB942tiJo1+ROeyHkZ04+fw/+f2RA+14Me
yg1ZksYDXxDyPgYaNLfUHWA88rY8Qvk6EMehGI/6aFw3FpmwxMB41qbyviYZcBiwQ1lA/nILFhnu
b3Vcb3gFlZ5/W41pZXuZVbHD24EWV93mW/P3v/77wQIfzHdFzyZC845dvRjyuBmMBCw834/Xy7N2
3ZkwybUgG3PP6RVyeyKKucBJXsZA0SCnz8UIOK4pJx9EMlvJiJZyneL7IUd7g1X/KpZFrhF96TB6
fuXIfTQH1jhh79alTEMNUQhYsAt2Wvlc6pUBt32KqRCysjCbJLekv6aWQAIRcDuO1nacGchNHgtB
xVQIKdjtGhXgtSk34lq1MH4r8rxqMl4rZtzTHS76LsayC9GuDnCW97F1g7QWhBELhT0lxm5tGD6Y
2Xj36QSX2fSb0iYeXVCPMtF5bRYCae0CbG012lZMfpFqYktfbp2bdkKO1p3XsIrVexJastuPwX1h
V5ijKaGywKn77pVRHVq3nyjnp8HP9hAOSSCUpC+C1oRFu8gBA6WIs01yzmO6YNXU8zZlC4d7sjxf
6YE7IOpPsPpzekcEsZhc8AoAHsSzSHsFtotmj2bx5x0zo5x3dxSpODhrLh3Z4mjux3LF7A9HP3Ka
U3arwPhYM4/jxmvVMQHHpiJFe0CAsrO915DUwPVyYqRrSD9VA3XyL51vdrzTMvxXno3rBf8BpXNn
jj0RRp6jhH8I/qOC0bqWsA/8Z3lGQuVJJtWjbK+O13EBHOtVa4NYN4qV0Z/sm2W9A7fX+vM4Pl6X
zc7Htcj0b8RZ80F4MCBJ947CCLV9eaphf4tCxATPpaz9tmNbxvJKSes/5696fPCL+l5QIuWBhgBi
D3WG5NenI3S+Aalt2ipr2Ho1glt0vYbXQFoISszupFh/az7+G4ul87E3l9G2cIecyJA7ILJbQZFg
ky4vEXRbGbmfYhbgL7G0WXGS/il9zNz9D5JLSY6Mq/UekgdN+qvtO8qV204puR3vRMkSr30bZTxB
bGlgbDml+Sw9ex7GUCLBycy5TuXFfB6PCYywmCVDlEpIpo2AsGur1lP30ofNNtRu1t38vsKfzeNg
UY9dd8oT5zufGtqzawY1+hSZASLL0v71zyKUeetuBtKFN0WXMYeSF/8waibhYlxvbr9/cjB21xHZ
ctUGPKOejCdn0oJPxmIidws7K2OuxA55DMxQyC76JYJ3xisJacZ09Eo1N3KHEH6YM/AMC41DZaUl
oJB+u+S5wQcID6dhzQJ14PuPQOFXHh8gOl3a0R4RS1N66eARxOBbP2Ao2mKl6agbH9GUbkWWTG0S
hXTZVajmgFJPd5vLT6PM+7kEV5w2puXBnq0oXIKTzLtpfzwYZvKCFBxekamNF+xn3+pri5M3gXz7
lEVtHHh5lbPlWWHYY7SMtUTIx213VG1xJYlYz/hd51qDESM3IP4xipdd/rxPCa4fL03IWjfGVpip
ojT4bnAikINc0CvtPEYHdzeqrwDgUSlVmQmF28vUhuMIZcOl+sLgKmtwBw16/OUKPhg0OaHprvC2
Im+z5GhwaSAv+ITFwhxxKmbgkSo2pt3UgUSg0H/woAiEfnjz3s8rj+OoUvb3iTXkQSgXwlreRFOb
bBXplh2QViNM1Zy+RC4wMDl2/kHcZgn/qpYVSCLIWZjV/6qFuSvXdR8icv0j+cN8tfSmnoYt11Sb
yhaDs+cazArPXRowhH/rNEBnz5JZu1cXFVMFmo1c3Ig+mJ4r2bmxcQu5Z3LE2JOc/Gs+tESqe9TR
9d3OrVfBGrwi29tRd60AEbFLQ0/7XCKJWxfudZ5Fq40x2PO4R2r6i9Lb4AQqHsyFdsMeCnRPhc7X
8nbd/0G4hVpZacdWG6nxsnwqGzA0RGNd4l9LuY/SW/Dohp69DvYSgY1rFZC7qzVys7oYKwvfM0mq
VbBpvSukva0699U5Yz1g4QUuTWekr7b3sd4Fj+RCKPbla0M1R89cUzpIR4n5uYfAeh0pB2msmfqo
e9hLZKSy34JAC1ReleojV/5ZXgGSwmZAUPu96MN/kmiFm8h3514FOryxYApHsls8XjPljf7EnYdL
2jajFLTx3HMD6TA+RgYn+V9m6sINtof4TFdmJK6yPFRIHU6Qw1x8KmW3+ug/c4+D4bWyPCNijXNo
bDy0MptJ8Pz2J4/RX6M10pxSr7lf3EXgv4TM9DPJD1Wn/oMYvqQwNtJ61QAaguzJ/sXUMV9Cc40P
B/rtm9Pbo6UmRxoUEJOBKaVla/FyTxQXMs8t81c9DEyKEPitOzrnVCD1W37aGdOfzBc2WNJ4c763
Qr/g/HiIPgLFy6f/MP7jlcBWY1Q0Q+3WT92aLkQ7IxixC/yHTbCl4WscKS+N58KdsVexbYaRMivy
J2yx3Nxu/CTnLmnzivy97bt/bF6fhvO8vS8xjjM27tbzJxG0GRCl01WGbtEjvDp0TVeabG6z0NTM
s6a/q6aEc+ihXiFFNtFJv6LoSU3MGYtTfZgqvIujyy585Ra25ZttIgsLWL+2NsUwZLqBH/Ex+ZnV
SJ2cXV8WWMqwBjXHxi3H/vNSqxG2UpBjoHgB6Z25rxg6uvyNIA4I2v0gHg7hAjBV2hB8KLZKELK2
7TRnj4t+0BcR0Ho9xlGvh2h/rAJg633obTC3564XlBjwa5DBTnN1QnYxWI6X5nUfoFMnsrKOtmTU
4Jht5RWJeYGBbCe51Nb2uGLWxXaQ/O3xFDboqd+XvBGrFGw5Y/ewrfeNSLpW3UU0n5W1TjRpA+th
y5zRQioKcuJQoqICKYnDvcnduMWw7mpRqF4FUgv+UWeujSb7EtDxFSFKwpDKUutlGncmQkkySugY
njXMBbjDpz7tof1blNxGZsa1247tDaXMcYW/I1e8Bl+tPSr9jD+tyoxzkXXZZKYZTTg8QuCesINs
Zaiyu42JxDywhh8cFVEd2f5VfTVa4nQ1jIgpxnbE2MaLnTSpZVe68eJLiXicjagNRcj8k2LfRKnK
GfDQrXWOpyj4ZyZHgVQVMdD5Er3mxImHEmkQayvTz3igOCWOSsCsh/qnTOaynwo9CCQv6M3lYsYw
nCFP7X/8sY8yMZrLTOD27DiPPfzSO959ZnwSfofvTiz/vToIwTiOt+lntk0tnzx3QZl3472+Qfif
QdijDCpJR36aM0Fqi83yG9MfAZiPhRlNoQvvAZTcPc9JIJVL0csZptL6Iei+FUBJI3VH2pnKMnEx
5IDwpStE5DZnmhYJYjJ+hRypcz3Db06ynTcQh48C1ymoY3FzpfI9/HVEW40jnVbUDBQsfvvb8tuY
CfQdQhKOdYxKy2BMNx/PtgLiwqWPB3rBilX3wrpN4ceJ5gV4AOYI8TLFzdVB73tqYau6wJmn+Je7
QRNmkTVjRPxhV78CLgx9hNLGijSX/egfgrUb5tCkXW6iZF0v6bk/Gl511+YCKcW1adwf2KWshdNz
wPeqpADz/VxPWtcYtwT90JDzCvCXoEoyrnxZisLr7iENttk5JO0mVrBnWdE+fTgoToQFPIMgufVe
H3NI+H/gLLQq0/JM/GiMf/PvJkoXPCk5OVTh8gJ3qr4bLnBPdxnwFJPZBNmu6TvKZFqF5JBXl+dq
g62DonbjAN7EJhmETpbQn8Gace8hiLqsQVjPzTcBVBldUX4znf1rP+r/MgMoG3KyLXPScBWHjUrY
LfOOrC/j2ZVehOFljqeb0pOB4HftsSqSxvtlhR68RFfpdFzUtAX470krK0CNqNMQk+wSP96mRqK2
er3gUqRqbNIjbYbKJD0LK7nviB59pud4/uTbUIwBsAol8OnSOswyiWY6lngMhL5IcpwEnS+udbBU
gkq0QppORM/9OAaGU+NnmqiqLvMd+OMnsscnmq3KPZIqtSZsFf8fEmZFaSMhyqebemgJmJ+WwcAH
EWB9cGMsy7WcHbJAufu/rE6Xi9fLUa3SB5sBWgEHCWwOW3hjMNmrvNJYXxZ697VpIQS0Ft+c6EE4
xnu1hpSr4v3pCgaL2Xo4PpIZFzICR5Rg7UuMFByP51sf/BDm1F3Bg2c1wI3oTc1erBvBX7c/FToa
loz7AhOCz2RE3FDuoKcdjirak+UFPnhUualNO/wIylBWL/Gdf+9wMLTFK7FkQckWo1z2nB0v2Oac
UAtZxzUcJs6ECJu+0wSjpeKrcOj8yKN2c87yWP5CWAEGYFGWA+eWInHbASUNMPISS6iTcFHBHaxv
8R0ZePxiCYl2qnq5U4x47zfzgc+ieriEyWkcfuzmFfuT/lByinlHJ+6qIXKqfsiGuJDJYpJ+VKts
uPJdKz+nmC+awJD2+ZLKd0sYb92tEFqflZYVtoBUboely8mNYAGXaBIVNGhCPs4oSgS7+Xk+6mF/
dsMTFy6+6VcUOBmB/M/mZb+vYqsSxWFByR/fHZFeARyJQOBXDW/sL5dOunX5IqhbVE5uPFYUAjnx
ww5pVvPnvz5NmUOnuBxJGvX3tpPtqeVwzDQPpg9uPJeaCborA50RMvmjdkeznix08tzlbmHinT4X
Djo0uz6QI9gSIbD3XHu5FZyTnvBrwRQKN2dqqt3l2WvNmdAMkhnYv5dbt1hzkZtsyDL2/f/XohzR
pI8Umx6B+vT3VTtcyS+UF3jqNJza9zdneUqrp0MLi4mIlvH+aEtiKuDl2wNgUm0x0wUr09Y1/Nke
hdtGsmOif/lAhFDI1FYHtvYYihWFelc/JmeVR+WI9U2MkkSTiufD1ats76ZyVMI5sRxGIioZmwhj
kiYF/qa8BxXDh71dP/BP+9vxin6kRBtPR0ThbWZFLAn/FI1PjHP9Ua0kmKNdHF3JaLfOKBP80CTf
vKfCHchH3qIQtURaPVo4V6nfVglNlckwzbL5A34oXEDVoLPiqYKH5QiO8qw6wKj4ggAxd3m3tyc5
lj3Up1hXKDx0Abq3UuiTRppwHKkJMKPIzqVkxOpztyyYvzEzlThcwXykoQ1ZHrfR0qxIxFEDdVFo
8yu0nJhgAPiPKlZvqCu2tXx2lohZl3BoukZwZuI6XkPzNs6yYkhy77LHCDq5QczljCpyed2d1wGG
76klXFORzxMGg+CxEzgjlWW1ecgFO8DosHV5zgk4GjUq8dLf1aB9XYopQTR9b3jwuRVdKP4VLAir
cmd3Rawn1z4L7R0i2f+f13dDwj6LAYiAin5FZR41KB7yiiP3n7NYHHlpiuDWrgr0NFeFFlahb1LG
XI1TnxgQNMHF3LTPFzL/DM1yGymJHzDPt/dXMRVVnGB04rDyunQ+XMdYJYhPMJXMTUCvmj2Cxd7e
BmG9eADA6w4v9NJ23uJUMNgi7lWZqFCucmPwnxeJwN0lKGEBHVbzW5y5Jw3iekpYL9SLAP4YLa0L
gGjROaas9PqpNju86g0f6zM5kw9bVNrcMKgKKh3cWBSp18nESbGQKSSyNiroWag2vxjp2C4J6cq7
e2ysiiiR7h+sRyg99G7F0wFcW85lZHwrC8jSxPPuwz5qygngv6KClsAVPYwUFq3aJmVJJHEZPejr
1fUyrXvt8gWBwhzyZshGWjy5oikwWZcSZ1g7jb72E0t4CpHqGsiVQ6QQ1+YJQpC507EzgowFx5VM
GefZyrgOvk4eZTnyaYRks+br+SiLki3wuFy6+oAvnzDovOQRkZ3PzQu0U04rAgeZ0F2DzlnoP1S3
nXG48OQVj/rABQYkv1HTZRW4X0zBjQRxEgn3SrvNBDauML7Y1l9HV4l9VQavG7Bk2+fFFtTY4rRK
TiOz2QENnc1r/HRk5U0SLt7LKiDklC0wyNGEIK/ehJEoXEW7zDdrK6baS86iViSiF4nSB2C/EfS6
bhqeMyta8ADzdlgfGlXENiAkbtjjBxQM5oEWw5+sK21IvMn2DThPs5t/SlLXML9+NGi+BfoaWpVM
NqXYWoL3XLAPHecM7sQNWAxqHEnsj8ItJZYuIDKFvTmKoeAT4QMyOmo5+OHcQUjEMhGOhrYn/Ytr
ufAhudt1EjAR5Y6aVT/kAfY4qTWZTuiRkqZOXDsrTs2gLszdqsLWJyDL+Oa4+BURRlJ/G0jHPFYC
4nwF4+eRb5f+qAX4XWcdMHr5tIYJaKnyJEP3nhkPW5blhDOuRxaYB2JeIp13FdxktyVVywykLOHv
W7FjwQWxxe9AD17WvR0Xc8XPW5Y2YsuPeAq+I5rGUAyz+dx7SfpjAJPmuEMiUwmRdUqs8UbLG5PT
W6R/z0ncOvv4zGc8VOU8eFD6pVOeUPFvrJln0ZpZqRryD1AzmhrNz6wLnSTwW0GR42d7E0ZoTo9s
ZoZTwnT5AD4s8o+b2xjb+8pxMrcCcgkVcqvb9FpFUrEJQgkqTjhWEC5AhMariVSYhk65f4sXU/+8
DQOseFYOrDwQdXtsCw2SK5HDeF5GP39EBw6LuhcVYuDmbB1kGTcO38xt4prFysLDHdT9pRs+Ltxi
Mn+IfdJhz/AOar8nl3kUW/w7oF3GHzlOOJfqGmZsGRU4USFVWpTdNSJ+yjz5l7pEnsln4GapCUlO
STZMlXtxYqO9wc8w4uAMgAuPuqKOvpX8+bUNNsb7uiyuKVQVA9oFWhv/gwlAfBTZYrr/nbYpu+y+
xlALzb8q/p8LSrORIlWo3p5ioCaeLilUw06neuvAAXtJM0wl6xT79R4lrnTlJJ3gtI1NDg0TSJtE
C0SnL7ix5YqnXDgy6fcgVqYUsJgUaw96v5/g0HlRtqAEfc9Ucza86Ngloh8QgrHlZvSXzPsBlst4
xoXcXkDvhu96PMZLhj5CArrZvAM5HgeW6wa+TL5WnsJOSjW5eJ3aabtkSCjHFx5kt/8IDUYVx1Fr
z5jkBs9pHkZRzojzxbv36lE/zTRfZZlyRaHdd1OiRMP817coe466vuplagg/4VXHbPio1SngTq/j
+hcCE5BUkPqQhcomc5lVXk1pjQzeun8TPqn/iFtocTOZvXy1cI8aR15nZu3boFXndO1tbzmHv3kr
VaxFO31ZLt4qmNn59IKXACxs2EYiS1+Od2jxwPrYkiFx+Kv+kcx+RkTgEP3BYU539zRvVmwSJonT
LZiopNytc+Z22R03WXLgrK2eKOhho9fVG1+Wxt42D4K68qOkInCW/njmKCNTwDwZWKZy2A/6qLSm
qoc4hHMv6mgNw8R6ibHiaYCTIXb62QO3wy0ZwZwvN8CYPjXHV5YNIzZBhidlPXu6/a+vKz/cp/yu
wS8iFHfNxZwkyvk+uoUA2G9Y4nd+R0K2ZjHlqVzl5X69oSPEe1WkeMcSjiZV2nz0lHni0h/fWY+Y
Sdf/OOP94YypP7+1pRP5fvuVssExNGKPUEyUUJWsVTFrS4brJM2mqlpJ0yewrMm52wX2UdH05Sn5
q0bqroISAYv8xstOCV5ffrxV/PXGYC6ikIb/2Jh6+EusSTog9Hm0O+A2cftVSDvW9oPr28C7K4B5
dxW1uYkWtp/I2hZET0WJBdUSXr/KsskYm5w0uHATsaBv/oQKKqfB+SzrBaVkoY4hfHYD7NeoCuud
kYugeplCH85WUOVIZneJV2EHlOaKvOjZgily8c74pBjQdbW9eiXcAIC3y3eFGKtfF4gZKihYKuPR
cA7Jqr2z0VNHqhQ647n63JJLeHtXPmoawa1XynNqtzNuGBOn6rgGqS2xOtk8Nj6CDpi4z7FTj6NT
sDCJKd0XLk/uSwtxY0bGlMhiaiB4WUPqbyZ+BHUWh3zueYffBe4rX3Mkq4iQt06CGC+AeIBqLAz5
kPrCRaiOuusPJArRkIprX5DkIp7VEQGgqQ3v7cbE9nNGCFjnXNP4EoAN0nCAcrbalE7KSN6OFXqd
oKpwrpqGrnIliIiLqLWhFI9wUycTkchaxT+cT6WsYL6/hD7IL6SqihP/rje9WvXMJsrTHJe6TUUT
TCgLS0CTg3SglO6qCPFPGGM+CKBqZFRLmdHjGimDmrVYtDEVBPDZ/bUlkh79N58+9KEum0TtHSZW
4lkD4B0NQvL4mZba8ykRe2c8JUPTdUZ76CG9iSfr8UEoxiX9uvI8l/fVpxCOITphRfTjKGZZmv4L
PsSQl/jfnt1C9txdU7LzHCkxIS4X+bZCw1WGE0km8ZWHfElGMFcsyPaXd5eJf6NYAFt6k8dimCXG
TsW9RYrX6vCt92OiYf8ejHPnC7SDy5Jross1Sk7gm+3ix8mfg3of3zOfHhZfkZN0gqltWnKYX16T
3iDnrQnhJo5ESIxJAHVJ8QGps38IUpmdOxyFjFEs1nRiH+YmBXbW4SNO/h/RQHDgvcuVgWbItovn
+KlGL4vtmsKoX42MaeLJ3+GPkodwNyYRzRZ0vU7dgDQLv8ENTq1XNpgwCa1TLcHkEhw30qBpQnDh
QRi8a8Kk3BOqyV3Ex1vPaaK0duIhCN5sZmLSviio+fZ1FNi5YJkJ/3NvLKJv8BrnRs0e5zGKE5wO
fCSWJnkNslMiUm/JujKV9hvrOmT6D8UAX9HKvHC43cO3NcJXjJO3CTf20e21hiN/ArOkHhHBdxVx
X3M9S2XMUOlZ3/oBK9OpewxL60oOXaDpooOXXivJeNh5WrJtQRedzApD89f3ewEPZrGMVfkMfavv
M0Acj3bJo1YpgeLFrgOVxR2mnj2MWZtAcQOK2RhX2PtFYXMPDJm1MR+P67HPw+TCN6yI1XvLCY4K
LTjqVjoWBgwg589AonqgGYpyQg+n+IMKasFQ0LHUXAdYi6pL5YX8s3BIokJwEQB4t2S7mBbDzq26
+RZi+Pnt1bvwJozhgQFpmxGfe9gYLsFsyRKUs2keUnKOYlrFrWQme67GoyHaKFcZzXp33g9nMGur
/50wUUQ856D+Qz9SJSxCgjN2FZ8D5EZPlslFL/d5/dcPJ29XMEyahWdKJZTt4ZZ3KV7ovz1sgu9z
fZY7n8MVqT8aP2CpkDCiSo9lSaJfftLkfefvkZUaQicruU9Qn3O+1ZOf3DhORu2QpBT3USXFlOZh
f2/C+/BZu2ZsZry8rH6Hc8Z2D3oTvXKR5r06Q42dX7lRZBxuKOKb0ovsh5v0cxYYqfEyTLGNag/M
r7ozDsZRg/K5DRvOlbZDOEpRvuFYBUpgZQ7lRJic3jWwAANeEqs2YgLqvNYG12SPLY7AwqN12IfY
8xuMnsRIIAwbK+JwFO0HdUBYxhHjk5M+VOL/+Sx90BqbaXYooaLBgfJhamaAEwedXluFT3QekCep
/KEcWk1BAPhIiGomQjig2ZSTBpWWRq3Eaa7CKzGaB4EeequSaQF+XT+6XEWDJ1tWVxIFVLoJMd6D
eYquPxcDtQftN0pxlD8EaR8U5rMj+e+HZxVOp6Kt0Mf2y7YlOTqmsZmSVhe0rYv3dtGn0VWrKLIn
ILRcOuiCNhsyW4alXJDmtzj+AGgNUgVYU8ni8caL5ICVDnEN6PW23lFUrynlCPsEyzGEYbzDKQRd
gnmGtVq4wQGluZ8DZI7pK+zurLOtHcrEW5mCmsAgiAj5iCgNlsbKMfFAESIrQzK9slyOwCXDmzjz
X2vUBcbH4kR376nMal0eQcHKyOykn1sgJl/t8HqcrCDrTlW0kZZm2UjuiSgKON4DsE5bdBsR2PlX
TMu+VGeQDEnsEytonHXZfgqOih+w3qlK6qbOH34CmoOXQxf09PoITptLa25LBpTEavTiys2o5M7C
MtNkx2gab6LRHlVzR8GuWQWXdIyBpmD0Qr2dwutKv7EG7EFnyepAbBSifyKFfb37L/88msecdgbi
7Tv8i+ztd9IPLivLx8hqAC+AP2QUb3L+ntz08XBN/V5e4JemKeLnKEyPNTkzIbcbtZdGRv8YIoAA
GjxPdtNoCvwB1RPLZkfYnyiLsYIlpmaRbQj5vJEYcK0ZejhBPaBnO8iU5xXFyIrS/7EC3yrnk0Jr
OXcJzXVlfbW21/Wr+glAjH47a/djT9o5RUwcoTLKzOx4YLAJWL0MBLe7UGIJ8M8ARXvSI8Ws4bqh
6TK4D7qP3syjaGGA/fJE73nUxs/i2CID2iznWr8WUkJSnBH++7EW7QGVFkFg/sZF8t3S1Bzlt3c3
TctPeTtSfnHdlVko9m7jgHSvzpU1Wr/HRHTbjY/TZPYTIMQ1jAMIrU2J/OaaBoY2kluzuNySLMPT
VunlqHkmwAMPrFFIapX/1GeOjbEX8YXmbWJevvycr02imzWTUCGdvGiOjOUbSs4l6G3tr90c/De3
nT1GCD+KqXQwwnuQKEcQ9JHBpVeKbFrSFjpDgJ2dAjFPOW8yTynd2rN1SbxW74+qdy7j43Khgl/C
XXpVJRg/UcunkeLFcihMD0tbZnOLxXFa4x7MYz17YyB7y+tOKcD6/B929p+ovbuHmFLqX6lbuIj2
zyek4XPCrCp+nb8Q33VS8IQxHCYmyeJJtHZhIwuS1qFMiJwdKaA/peFXswHrsKd7nfqB5KSZ+7IQ
HFkm5ytCq0qw6ltio97owW+lnZ5j1Jfb27e3IwIadflJri2Cm+wF/KkyC17gg3Z695kw/pN11LYO
YhvHZDtvVTitW+Lg7LOoOBneNQqfpXe+jfMomoMr0Up8Me5VBRSK1gj51Xe04fkMfPY4MR3wU9tT
bMEWrlGgJCu/vUdoLXt10r3r8SPKq2n65fzqWesWcJ/dLWno3SBjLtwnWu/hTKwT5lkkul7CClbQ
0kbmDtZLSpS8NWmy7L4akfXezSmQSd6GkYLjS1kkZhNVV2K2jxnLFtgUjvIQXO9eZjl7N3QWpiI4
Re0/lRZ1PDf1GKmOEz82zByZAef0O584VlwdfZhEQ59Q1GgWQPyMoZGanXX0ECVsHqaJBLgq5QdO
1rSlrOUnJT2N5FXA5AxZL3a41fXPkOdUH1RlPOWeaqW1LZ8QuvctDbInGu++BTm9ZyCEUITrS49W
0dFkWW3dZaPCI5uIE5F8Eg0IlntqNzTb0OfdrJid3WOBy4bcU8m6U8BJLATbRxAf9ne7a0z4afXY
Sb7ZOjO/Wf23yg1EUW7nLDdcvQxDMAyE8WwuzvVbZIhSR1RUB94pla6GlhokZHzNO17bnskxkUZV
v6ZCJc05/SsthVkgCrkYS8aXZRIuVJqcpBvX8qC8bGXD5B/5iEhhUttzdhc+usTqQkXfUFfUcl1n
83IpMFRhGUaAhquvTc1iWntPXc1sHPkCWUKxIwr+oCziW3Kp/AbYsaE09WJKLhxNBG0x1RgqKUvo
oPDVFP/xpCBBM33JMhDpXJ+lRfnn2gKfUrr2xjj2JP1rrayoQ0jcO8sueAUJnGXtQC03on6uQWJS
HbwZ1r3u7Tgqog9Oy18wgLp8ycBpLbskcIzZAtAXeVtKZoXFdhNw3wZw5W0MGXcn9BeEBaxIA/1w
8LXaI4tgSbrH2lXAq0mez0Ipqxzzrcw9kbdkkLaS7k2Y26KxBy1wzhkGBp0fDtjNQR+OwNCstrWw
8AwVFuKMgZAhgzkG7pASooX4eJPuY+fZJI/nlXFscJorPG/MK14tezhI8DO6RS7YxsWesQAJm8ku
9U2UxR2OPQdBY+pbdj4VSdWeFJWsk2XT/stwMuQU4Fciz5X0eNt2wmdNIR8roxJRF1BbNqAxBPv2
w/yz89xp89jW+KNeB0AwziwuQCmP2dY6uwXMPaWSHNd2RuUXChFm47ozsljAgz+G7PXxo4PyTXtf
YhcwxQwAhHUnLZoFKghcRMEVmPEtugfIYEMi7cigxoo764yHa0W/BoSCxRP4XGlzJR4HF11v/eQH
ZGPw1SplTbp/zkaNuA52cdPG3GDdHmXK5BrjxFSdsSkpAYyZ1RKlLG96AAnvVKehgSBTjNpZDceB
3oSZ+2YxawHTtrfcfFJJCmBmcy2zeccM0BHrMvvuTutf3Mnbdz6m93Y9IHnZHrS9eDw1ZebuPzzV
xkWiY/8ponb/PlUOS8jgd1IbpE+KsuVVxyveG4QFb756urjtoTUTsrg3lSKyh6frXoAJ0swqe1vl
C2zN40YkxsZbP3ZgTYdWshfXD+3YrItiSx2HEXP93S60schwjNJ0503ZzCWb52iA2E7f3QrkLbLW
xDlzoqARKIG42xcBLkC/UbMe9A43SlaemBohqEMzKvmv+fabnmuwm6S5FUrq6pIKokhJ95QYuvRV
T3d9t+IuaW6sW04RB/AfD1lezYlNpmIQrXIyPhXODyzOynE05XK/sqeBD9h0EQntaSQzqXglIeZo
NoZmwcD/8Kzic+J96KDBMgkxMJi+Ltq/hTvrh8dYiKDqLCgjeqFyHMZjFecu31MEJJ6SlqY7oiOW
AuRwOu1s4j5xQAs5cXTfzVXsXult3p+0pHA9/K9D2PglPV2/rOccL64nvE2rhYm8o/4zHvRauGAR
9GF8a60CW6sG8Z+VT5mNPQo9lByaf9r5FD0lNJwjUAQxbBh2V2n95DO18ECqhJD9UbTh/IIKi1YV
gPW0AENAtuEcJ/+h3f/oSQlwEv6fl6gaZ6ErcEnEOCyIpJ1ehY2iATnCabl7lAsE+sBef5HRH1mD
po7MovVebdixjlh2mEuOnEirLaLdFNmWXKoaqDye6S7gVqJ0sgjjAT33pKJiM/5+BVvNRTwgupJI
SlyuBbQwWiFd3/gT5hwtOjqyy5gmtTeVVFzSzDeIUuMglc9Yp943CSadmju6ZuIJkvA0jNugVkya
9eFCfAx01vdmi/N3t1IHDOA81o4hk9A5NosTIQpZB52GuCcM+ME5d1v2sDehBivybGbS2T7wzA9J
JgNji4tJbZpAUKIDSjRofX2b2RSYGMrT1EvF5ViS2ECKZQWAnl32HG/zQctxd0eUu4uJx/+87V26
Vwb7up2/t+6OtpI3GxT4OvsY1Sd1tE3W/3imTTqLf73oqxCqYljy/hXmesxosvRNoCWPeEOdCC9P
GmrXY/mjiY9voZMoVTkrZZ6L5jdz44M3QuCClwU8gQ8W5k6g1XFlEuGI1ocblGi5u4af6PXHLarO
9g/tLlzUHeNyehSyQgd07U576VCIaH/vvNxfWo0eg2hkoQEs8tEunP8ecgbwAtmGkTtsGMQQAxZu
gNSyfI5EFzkGaBtEuCK+CscRiY6Yfj33vwFGa35HpAj0pe18Q9f9i28KZhsq16gZxYwr9y8znlnq
Y944hS1WH/ONPCr1qhQM4a1gf2aryLBhfWX+Zl6LlLm2AOFvlDd5oWPyCMJeNrxK7vJvtrz7A4cU
W3sHcteq0aukD/u7FshI37L3aN01NPbv/whr7nP7bDo9KZN0FABj37hMsl5TIM+c2a+znq7RT2tV
ec7FlM2Yr38k0pQCryD5vCn1i/HqXQKh+BYfL/TUc2px0FpfynPNVxNZRKUquykZGtWwYmvwT84A
WWLCX17g0xvoO1qI5BqV71JyLU6Xc7LKDcxERlTDdrFxRF+O+6jUtiAp/KxjNE3kGg5FIcjMPjpN
d+fDDV/yJ6HwK0tU2CMVF1fAgqz6wF1l78TslgFW9R0FEwaupmmyMFF8VeHE0y/hIw3/gfvoaYeN
gCwZ1RPOkK4/PWFcZWr8BNWz+LnIKjGtK3wMbCOyUs86Xa2Xg9ZCkxOQpWk52N4wID2zLfrB9IJ7
jeavGv57TsEsbqunpqctwVYCibTkPeQkHTMqfJF07wGWMUY8CIzr2gMWDjxwNzcC+XD4t+o2MgKC
s/5b91Ty/+FDqiOwhqYhOeVOwInyuqhicqENjAjUEdPSHxNWUv6BrO8YHMA8OVCP03MdnHs+gaS9
WSZWQZds9h30PtFqXaELHy4lWGHHbNZGSEm3CLs6N1s9xa1YgeF346JNrBOHOVUwAQKO77zoP+Ml
UqVNlM6ogv0PGQEY30oLBPs5qgX/+jshr8CviLfaGKRjhOJ+t4IrHKUXsPghk1ax6kREeisfwfpq
6gDD+NuQXpUZCvUc5mVWAawcbcwlcBoD1zlCksPNezy7CuqvkewKMEcM2Q/vIeZ27SbqRWI9MfwB
q1o7AGx39EhjqISHCiLI8smRQ4E4W8/Th+asoPHaF1EtWu2X0FrBFvMdG4LYi4CQccPac0MzOR2J
nfed6UTTp884HdPRS0hxqyh3uim8/0ryP5JTfodf+Ps42YV4i8YT9nnUxDfR33ijUpYLxNnIlUTt
wZbkXUcMChgRG7MXbssNRkuL/za5EAdN61SngHQAQiOZweowAjTkJDR37NfCXPuRXiFmxWKKbhwC
vahtt2rP3v5SaLgGHjpoExJM9RJrhRyPfmQG10kshDYjEWC6ONvl8qOLdg+7sqv7axzES61ZoMfH
H3Nuh5Ir4uCqMrx6HX9npFx+ZQXW8oj1I5hdVY3aKQVJ7esJ5PLIrvAxopEGVAOWDnFzN9R+Hci0
NivoG8X40NeQw1/yyUKeGhOIsbl4t/cXwbh+ihFS+p66QEUyJ8pG4x+g5fdZXaGl3G0hEIZGBNLJ
UVW9QIn8VuUaujtb9yFJ8SilinuLmwQ8/RJdfYIEx/rpoLCvWUZx9nYDLNaLAqysOwXFiVJ3iXv4
c1m7IMEnAMf5SC047rxlPzfEVvkwqqe5hJyFf9kOePdn4cYvDkFpYqkQL+k1kis1J0s75tPCBcxv
BH3Fh0tWY8hw8QuGn7hyREbD0AwRFPhegWIIZalmkJbKhIJFgTUBz0JWjk4Dm6EUoe4ZEVbFBbQ6
ouYeSWfL/nu2mD1Oh1OqOuobkHiIUpEQuewjjmVLUIgOCf3ygiCtZa/kzz3g92RhtdPBXjKvgcrw
NOxPzPBMbRJqN7Iq0cleLFOlFHFIPM73W2Byxg3b7h2gggUX4+MWf/NPbtUSQHyYqMOzQY5WOxtR
zK1OxD5/Jaj5t9lBI0qegF1/Rqkb8oHK+6dAnc0Gu60mWehc+8zBG8gXFtcpvuCRCRzII6eICA85
JGLy81FY8lQSwVVvP2h+kdKlwZvJ4MlYEvF6lAdBdUj1mZcC/hxC9xjAIB0eu3n8POk+av98gDGi
8bhdeHspzS75hhCu3B8B29Jl8XXpKTgdD7+6sCP2jVCrLn8ZklD2aKdBMcsdus7pn3K5askZBASz
qZm/sqS8x5MqMlUv3oIPl3F7VldaA4MchCE4FcRPKygWYUdI1ooVafC0tmsbc6xgXGgX2QaeXzfQ
BGH9M7hl6D62vKQdeTCDarNqGlE69+nd7qeSq6oVXVEoJfwsTfl4+eUwJmltiH+Pbuudt9zpscee
9JKJVMFrs+SI9rNSZbCnmkfpGgFX4CMVr/o6WZsc6oSD1ndaJPLfhBKdQEcqzTkyheXGGeCMACw0
3sdwtfWIGoFkUvZ1HptfhDpPYnIfvMccqaaF1NOQGeEA97aKNqi6ifKg1+2GbWHRx7I9vz0LiK9c
HNFOs+Jmc2ypysR/duUcVWPegmJuvM5D4BKlefTG9w8u1gQNwQwNSrhh8cMYtQ7Re3MzxzCvvyMW
a48oXtBFRh662f4YYGhu243b7j8034W5raktONiIIIbOW0kgBiBgMcZyxSFihdz6HbzOlPOeO6X9
UeJDT3058VWQP8LlYIfj2/9IOgq+SQtV0fEmwivvX9h/NDG2qIlnFkuUqXlmwjxJ4GtPO8PWikzL
QLxt/9MlsXPysyamh0fJkZCJpEgJTUqZgU/qO5/jiK6eRTElA4tJpzpqQ524LSAYBUpzXylcuQx8
q0wiq0gmecax332pC0L4iT90TC+PMRGnhkcU2XdCetOFbhTYeMAPx4Ruezikc6kgGe6yF4Gscxng
3LId/LqxjsRaYSyaQCATYGKOGt4bzKNNr2mSoAF9RWFJBi1jUhlP2Ab9oTavDx9MltON6tf0rftW
8WcBPAQyNdiREhzNSck2RMQmX1pJootLS9mfp0MmVdYAufUcWuzhEs3K/x9/YjTeErJFLPx2YmaQ
QOuZ3rxom1WySVDE8jE0jEEKY2AOSlsjmdTN2x9NYP7EsMjzRTFwnQkWlY+AZDAuTcG0t4C7hcKN
bJDWVwCgyql0W1g0soeeEQattjCgPsGQhyBIbXO+ZoGG9agtENjrjmwnN85a+3nMazPI6+pLcGB8
lXSmYzjvQvxvGShkuHZi1qVVtaakDOMnVCoJhuL70COE44RM0UCrX/m9FWyNL0G+yhBZ4CARA3aE
wHxkod9qbfM4K2TCHCGIIbC+PoyAbhagAAHt3EcHWM3COLITUKEbZHazeHdZ/sl28v8VYoAf+HpW
IGReL4Y/fNAYIJZa+6dnYciOzj7aSK0iCYXxWuPGrlicsVsqWrCdzZKAPuow/CjiTugDtrcML2hZ
0kzMHtebikRezymGlOFhU6qn4VV1DpbLV1gfxTCQgNpefrWRd6EWO1EmrIydsqwfj7vbnCvLxKnj
kYkqGk8CTn63dlh2HRkb0oHBATDD6QoyXw2HIQllPUGYzVjg+G/jCkQXJVIMsvUbcKHK/XwMghoK
QIJMd1uRRcKi0qs5NW+3fyGgE50UDiW4aDJ4uwecfAkLKOdoqGNMEsmUEU2nv9We/IJUfHG/KoDc
tnm7e1Hyoug+LTqr9EMw71tS4kmdg5H0G8kyTNPBo/v1NK2cJGBcW/bLM+2LxmnhtKiHFA3onnlm
RDt61n7wMvL4cNT26U7iY2sFx+fjaCmSCrxfMf61bUx1D4Vqdpc0PEmsLTkA1+c0ioEHs1UFV8wx
MkLb40mdhOO0pUXrczHp0Fup/5AXTFj8mg2nvFa3OPwLO+P0JK2R5ZqWe1/kFzIELXc2ZrhE/3aM
TLA0o5ZM8Cc0gBK1jW2SsaDamQZadAPdgVAAud3cpqcIEr0R09qITUDeIhtn3CrFVSDk0e+Eczmk
J9DxKnDUolVKvCkrKWHITXiNZ5zADofNsq/sS5sqR4F6JBNVEwnBWekMQrB41Y2CMTAo2s21qWdv
QFJ7k5/oDxDOfvDJkN5IcHh31u9l+YvsYdh54PEDo/fhShW78Nw9mzgzJnkigPpza4Yr6SqRS9Fj
fyFdPLd28R+O5+lSxUyAj3/Y62Zidzml+qVudAsJzqCU0kW9cmbfXOA9AShx7O8D2m7CM3lEIUnE
5quJiRzJw0WYMnAabtpxwI7+7nHY3nImyCDegpeLxeeE/5aikXr0aUlCRcKamo33ussbauKHdyeI
nEv3QprSw1l88/VnWwcmaYSDciiy0DeyzUUcP15aDm8IdzZ0mj9UMTHHpzFRA5mC9gYLjU/bi6Ps
fpmVwuF21IEdDILWlWs6ccUSpTAzgRyN5+QtPJjcn2zXvyOREHW6SMawugEZZQzINhfh7QU9C36g
9Ok2bU2LibTwjp2tXtzxAXG65sZglw88H0Jr8VMduaSYzgMp40ZMbzIMt4c2go2O6xJIENctadFA
GLoDpZ81kJ5KGCFq47bCrOmK5NYxdhkkXf2TI/fyMlhy7c28h114T62ee0kgThoe23286jDTVGAv
HQkXHlATubzyK7LFvsUdS8j257UEg38+NvfjYrrDiyONO+7NzLsmRyrovAagIhMQ2MpZX1CoKqC+
8RCEOZMI/Ok9xS8MCx0CCE17eUwEygsIjO1dupwtGipaw8zWsU1pqaBXjSnhFBqgfnNpeCWXqb5Z
wcyTWIucqFMTTHGQyvHFJdo4snNX3ziQtUYutvznlsTZgJ+1FZyyblUnNlBLlISbD1Idt1cpDYf0
q82WdY2GRnQClbLXcWIvKqvaC+xx+E1J5X4+E1FUC/a/2YmsU74JDHCCqEsy6gb/oA/5iy8qqmJY
NfgDxmAEhIkvMkztQREacTFPVBssrcGAfS76tNy4MiagMfkbOEi+ausTNvW5OnIdy1nKfzkLaaOU
1vqnAnulM0w3pO8MPDxFv6k7fqvjS2zfyHIrlLQUSkWoSS7+smV6eOScBSJ//SPd8innvnyRsTx5
w4CdpzV+BjYShy6wfnl8CGwAJEn/Cl8beJXno4Sf0BNHEm64+hQCJ5euzviEopaJ4TTLSp72a6ZC
gcY12SHO9ziRFwbTgJWNg40y1iOgXAmOa4I17WJA/JQetnqic9E4DmdeH5XC7ih0qzpEk7yj+uDE
iPTRETCndHp6Kf1sePYlU9y95eg2WD8MRtGB25gaMvY+alT/qB0IDr1nf7dEjqq73Ij/M1bUbHT5
exnNnM2hOK9FBj91RzHs1TqGyUiMdo+5s9Usmglo5X2AAtjbTIbBBICxU+Y9k+FLtQIVEnl9PnOa
xJMMAfi+5cvElQ+/4trE9FXRexFi+R49Iy0PpgL/gAfCxp8S9+ai8q/snbFp1uSpHlnYCycykp+h
l3BA0s80ZG6P71KF3RyTThGrqG3ClDypbz0D5eO2DOwIQMWzZpyonn53eVgouZgNT6CUXPuEY6Dq
JWjGINRenEy53nfvdMl6E6ixsA13t+0uP1r9kzLANeRyIvYX0ifCLvFAh9CO5jsOcmQHfIlNs/g3
hPjOz9HbP5H6go/4PXPK8cpOwfvA6LMFhIfn8itPBc0rxIMxuQnsr1/LCRAE0HSFYlt1pAyFEYSl
yUq+5oSfQgJM+vjAy7Q/aTsm13U9tMu+Ekhb2HzR8e51OL4D6AHkXLOgKtvWtd8TAG4c/WLE3S81
XQvagl9ESJXBVV2HV8KB+Sl/3uHG9H14re1eKw2ypMYwfvrK/5si/5nMMrTYN566EXlidn352afR
yY4s7oZf8P1wzC54oNIVtk7plUB6nYXWl3uEmS3awLckF0K3lybD9DdZygNJT0dwR7gNH5gOc4lS
K5uhj391A+Zg723haPiRf9CFjuAjWjYCEmUX4wV0UwOyrakf1kqDFV9I0BqDeKO8bOM0bNpSnWTD
1pEZSnmKsK2gM67XE4XqBTP9kD8QNU99s9TBMGoo7R4q/cfi4iVuIKQZBUbNEBhujWLanKMWO/JY
VkItODN4c9BMNvs50qh0kJTdUVC/9EZ7fJbmwiehW0YF0Ier3gi/sQDyMf/XR/WeWW/E62nNCCPa
KcukENNbrGLurcZc/yRqLlqnS7/e/04OBfSTjQDw0/9GLd9H/cAI03dSKZwLRypBtf6FOQJnonj5
o7+iAiOsnTKRvxuW0QrNyl5g3/l5LmKzh+faE3RJbI23Ns+HlFx+bycRAvezRtVLlt/YT7vStJb7
3mGV1gTZGjDWsUUP/1sg7fPYdxAc3+A/EPq2hQvlpoivkDLSAeB7vMajkLRIcFRavGobuDnNGAYN
N4n12EDhmaUf2b0merR4c6jZji4ys2xblhcgbePoz/rTSIyUcujNssurUytFx9fquEkqiaINIZDZ
qJWJ2pVEM2C2+Uqy2nrPoRB/GxgKhEzNCBVicMu2HvzyQAJJN1DHNafsYYVo31jQVjeAQNCNVHAu
Gu0aO7YWsYiDWTeeCISJM+PXiFG0/GCsI51YI/efc9VVQzU/qBzP5XoerF2xOvYAGOrKuy88iOAQ
nv5eP1JRaOl1GKVvOHpJ86lOvqsKNLw6+5pzRBmn9btz4vLPpbzIuANLlALlf2vXLQmWYejaabsd
yuR5C5mLuoigj1eSGDh4TbUY2cyL2nAD3CqYYbGuZM6FTz3C6qn37DWBaNEeujOqy5WvLenx4l2a
2u52SKbeZ3R3vCMlmDYcSw6w96NTa3i+IQcUYyES0K8pz6xqgRNn2zazJ/Dvp1tbG5FBUzO1wpaw
dOpDvxAkPPROBgcbIUIzz0igIUf8C9yIIDDYdGsftUZwFD67KFNCppSkHudBObCFKmJhPavXVdwL
/YaG3eAMdX/OQIojmNbZ0Lhcp3dFywGOzd78IF8hPJ0eOdkDUFt8N47Yb2wFMv7PlWG3FjZzumBq
+p4tc8l4w/eEjPoLKweD0/YsCnUxMl+9SPCpjx9iQuv+L2AVhhZZFhd0bsBzAWZ7ExRpV9c31/GB
88vNMjhu4xabBohsDbGrQYg2eCm8Y3Q2RezSsnrpT1Womg/KwPsV3ZMQlwBHOrKQhFsw+Sz3dW0x
//HjcKddg9EUzkpdspoIAZpoGv1wBAs8dCG5koBdHgHdy9ginp5zThA8kIb4nYzhBsvnwDtILMdV
MqUXyWtbenZRXky6Kin6vX7i2rtay+2qHVUTOXKEz8taub+J9kKaPuuFfTrOhxoN1nsF0xeT/NsH
LE6bFALYEaaedAr4QMOqveEA013dgLbaCw819Ig7zagkbD2L8zNAcmiYl0xkxxAQ7uBHDY9DH4Vl
Wg6NT7e1fUaCBoaCC3jNaL/HczwzFSSiN8ms516YLjHy6sUOkif9Gt+nMaFP+YDARlYTRwntg5r8
DUTWxp+PM1He/NtbIYYDr3sUxQgd7RJCMc+vjTjA1zNdxLZEE8nJwlx4rf6bwMZdFZupxP0h+B1C
Oh9uDDo2z7J4+IgecvkL+LAa5VdU44AGrgcsfukfEFx9gurjppn9wE7kwT8LtOL5UrAnRUvlSCeM
2ZUyI2T72AngitrPG7Nv8kXrK+vQtf0XXlEb+41qpwJJRGFkQTIWzwoBPHjYomSJghKz2VrqG3JU
tR85ExpyJx3/S1zeq8T+KGTZWipzSVp3zqCp/Q5jE0YNs05Bn3Y/VgG0VGHEGe+yqEbYY55UQZQu
KuVyJMgZalMd4PjUjnHT4rDYcQaNYImykDJve3PHvHc60WT2W7lTXz5pzZ+lbdY2/zeWK1i0AuLt
+y/vPqp8+NgfEY1foAPOOhZD2a/dM2c3jzaoqQSOsk7LFUS9dgi+mkTt9xWNFkvumjX79zybHrlo
Nr1O1rxdR4rvLRm3Kc7Ko0+uNCN4JaIqLmolTSaxIgzdjUsdwwENbqYqnkQUNqcKUIRL/shDQeoT
HQzfOJ8ZEB3z3v+U+MeYYReqNOp/xq/XbYol/QHgbUd24dGmtH13IkG1wKGqVPB1zzvIc0L9/FsJ
YxIfCYLun7y5ZXL9U1j5WlnxaBA1bs35I0B9NJAypySXt55/erTI2BV4iSHXpwPdNGGxazGuIqU9
8R1SDvaA1xaePSGPtxqjgDGzcrXxBCOyQyaL4lo2CX7fO7U84RH6uJPXJNX8X5b7bHX2p4MGUh2l
vAaaz+wjeyX5B9d1B5NT0MblsIF1qF+J/36SX9ucEgH4gMnftGsbZbcbkjvo/nedU0ACpXLIYzLS
Fi4OA/rcE0kl9eF4E24b6v93AUDzKsjjbj7ab1oW+GAePY6p2zOdrN/4Dj2w4TXUDY/r3eanPedq
qt5dcwURkv1bT545WaUc7Bl0ZJVB+4Zmt2diDByl2y7+L3Gwirxw29jI/VKg3X2B5wNgEbbcjrzV
+2cgl6qW5zo1jM06QaWbg5G5d5uXx1wHBPbpoQS8n/TYCsPsptI0qkKLxsMIpa9UZWdCmp8HIVQB
xoGo0clGTjZPpUreQre1p6hTIuX0DwRtOfqdH3XMe5qdZCh0ZKo4WNQrrsx3fmO9YxHQqEQ5yyxH
CZjWBBuJ9LHYpU/3SiB9+NKPHivkufBBm2i1fLwg7uRHrwZ/e7X5dJqtnC/w5gGdW1GMw8JIb+Ka
lvcf52MGkVARNsHqYUyZV2LFkqpBZxzC019S0PRqdOzijYmLaue0KR8eG7kDGlXIKjcDWUJ1KD2m
C4lTFOdkEzwpobNrRMHEokVKXXJ1rkba6gA663jlgyQ1Hx62xOZt36R3XaNtV5/VEAt0ic4Vspi+
rk6c4KDSLXykuFZgOjI7R+62SIBQVavR97gUdBCh9HpL28eVzgTyNWY8mZ0kvps9jR+RwLyN+xAl
l6tBQGokFgU1GPxiEpwry563iHDO0RttsF1ZGt/gVciywgDHvjHIEH5WNIvTswkGSOHdTFf5/rZo
xswh2jlXzY87dKi8l2NgmBKMcySb1otS/8/hXXay/o/EidG5yExd8pQQ7UH8nIQKDaItSjzOkqVu
uC7H12PoGO68crEmnpPYr5Z++oTWz1Gdo3r2M+ZwW1WWsamc9X8gCd97oFGO5QNhdz93VTVxEd0V
KDIjBde4mtq61qMbAUznr9l9LzFFUISm8WJDw8sgASQeUzQqlD2M6XnXe+HmlEALnpfwv+NuoQHn
FVmwv1GgM0HpQnArYWzwEe7nPo7if6E1gscQ/wABBJmwL1YfP1QZDy52UZN5xVnk3DYgGYsoSplf
hT5RcIcmpxj4dk+uER7owd5kOgcKr8kanfC55VyDOHpsu1I30QzFnAw9DFx+zEWmfXwe/zWNX+Ts
n2UPUmVfvqu5gN0MZioGCk4PVb0g+TvaQrHkvlxIqAPVFuO65hXU0LnJQNqJBBqbe2FNyuXmWr1x
5xdL9mlrgZxcal4t4Gj2SITWOZpstRkRljSW1FgcPxGWq4lez1Yuh0WRELHn4ex8RdYUbNqRIAzl
EzCm3d6kRw6xzjd12JMWukYFY3yVdpv6W2eBc/mAxZf5yAMM5GY7wE2EUxy7vSt2VvLcwNEC6YH1
AzUBHBSLQYbs52Rfc9wzHIrHM8aJQGCW2s1dgFIuxNHya0GCAy/6P7jdnp71zhh3a0nVDZWFGlgB
w3nA3ZWbXOEpTHGsolMYxXwRqw6B4uqg7PnxmHcwgPAQ1MbZIIThImFrHSqgo1Un2AiBc53ATQXy
RA4GIT6ZbdC4xZq5wDln6st9VSGJIe2bykQkwpDRQPHEHlJnVsWlMm2BRsFcQmZh/QLhBe2cH6Uv
2hCG0ScJBkliD1ASP2K6ANo6TEuK6hOsc5EBVOnpniw80eC/D68SYwSNPAKJ3j7CKDS0dhpBfW2k
saQ/eHd7kUHObPXaL8nD0q7MHQ5nEwiV6j07Tge6VW9ph/p9awJoI0/kCpEcg03sHwPjJyV8x5SL
goAo52DKpolZiClAbG0KyT2HkrUPR1QmT2UquD52ZG2WfHRlRGcN7h0CeUPgdxXm3/hPa1fqlRvb
q619iSWG7kSCUZfu+rysAybXi0e79udK1pkfd0jamkR9oli9MplMKTAhAhnN1Bmqzxrd6SUsGQgL
olR2mPBiztZzZpuoQZatsRms69yB8ArjX+/i0GUNmdfRQx6Bncox7P5BGiV5c+Y7Zo6FakO7HNZD
H5AYUqe4qNnu3p3E5q5ZXEX/a0IBF/HaO+BChd4ID0K6yPYnn3Pos+nUDOgIMqeTneQFC7Ms8xz1
25uycMjAZ4JXZ3sDv+V+jM0TZMJykuutEV9jdRB01fa9ojMEx5xjf//QKyrcH5kOZAo/2bqeZoMv
64SJHtQYExRttOeFCIltFhn6/z6aTEbig0nIGJM44qp8L45AqEQ8SUIDLMnCh4e0vrheD3Ar54gx
bfCl2/lG97QoiOdJbS7RSNCu6vqhFQuHqH48iDusBHTRI7Qlz4qFORyDQn8mObbe1WUBn/oYNwbP
Ka8ACEdaQEEju4YQiEQpfaVOmyMF7yOXDljY4EZlx1TvkxMoFzUf30ysjFkJ7tCAyNA2WnzeAtfe
1/jHfp1pTg+W4y6eaHeFiP/gP3ESlbCxAPuoqa6ykNolF4eNA+Kxgue/KwhnklbIROzjXb3leBKJ
791Aw5MBME8bmnDFlZfRjLYwy2am1Nil6MJrHFwc7/eA4LWcaRtLInTGVcXYDifVN4FykkWu8Rb7
l9JLZMhGQ5pfdU0CwmYNBGPiHPXj1mHbRJjcDkBOIgXPfvtlZ1fhGOh6xIscJdzW90BDY7eqPwwg
mB/HOIRm7U5Wx++Lz5OvPB9Yg2i0u04SBZwxVHzyhgPycPURl/JiJWZeaQuFvmbIDNF097K3Do8h
fZ9ogD/ULhDkpOKKQnxzYqqXOj/Bk/V9Q7Em2fkKpXViZGAIWj8Hi64HrjR23HEFKyegdgXfvgKa
6evqF1+eOD74UEV7fZy5n0+Ud82c1jgOGPXQAwpZKeNBM3HkhZcWDSUZqWmm+XOs/vJFjJXb+vT7
5bHqnv4x935IXy2LyGnERKnytjAt3OR17nz9u8pI6Ugn2v1AxWepuXUFtEgxacijFS5MimBaKyzJ
iX+BnCgN11Wa6eJ6E+8gdBedUhJicsDayPPzpqWEeKoW15STr8McZ5dpNxPtyITK0yyDoMrF5Hvg
2UyUch5nmJyBWKWW1ybW1utgycuQ85zH2Fx26j2kHl9u7nTWG7cc7u2x9OnAPtKo2+kvRh0+wTKB
hF10AzuPOQO+a/CGx72UhlsQwBXRelXx5l1NUubXf3w4j36IKJ/2r3kqE1Xmyp44rFLSys4rs7c8
1jmrGiEu9iWCIF/1zUwf/Qw/5/qTyLUyZPclxtrenX3WmNq2AHwLizZDOSpEd+bF1T9gWb+7qfwa
+K+5uKR+Xiffs81pMdQxBEeI+e2TYbEK6OldCtIm388ZP141tKbE5jFX+06Bw89dTYUFV4l6ouPS
PUTpkjLoRi2yeQ1FeSvI359NjtSpNoSI3YukcnW7+ta8VvmyHVtWvfJXFP8ShQiBOQQO3CunWhJO
Zr5BtOHFX1X/AXhNYrLSSVr2MSXy0ApaNJ1khsFhXXm5QZHSLdaQWH0vAt8X5UYVF78EWAtTb0AN
r3Jt/PgW/ZxBQ2SBVgdliAhIqfK4xpa0y6uPCcY10JzyKrc9EQsn9bc3yKyFm+UyS3ohLqaatIU8
9lR+DyKBtCG2nDtb9ZoX79SzHclWWBjgo18Yf7ye5719kdO+nDLb3KZ9aY7rgqj2J9lxcCMxfrzo
GmllwXL/UZioYCR1nzKDffe06Lio2zSCDLYiCJiSdEOcS5q19LiZ4rsA2TNLkf4rStr8COiE9yQk
nDEAGxBIiJA3zxw5015DKyZAe4WrqZOfooi+lv2dT3Y2ENMYVjSDET0kJ/CtIrJlZdz8x3Ej94/v
9bSzkzWPxsQ8FIaqP4wF3k5uTmD905Pu/jXBNrGRNg/k9rZdbEq0CW12eor4tv4q3nySstZVYXum
KvdmO2UqkZxEANKT9D1L4WSVVWHu0CCZrNLa5cr0kgzDUBthlCHv7NGD9Ad76fzasFrTc6eMD6Rg
+ZXjJ7Zsmbx/febMMdnv0B/FFt4IoSe52mGNkuo9V6gITIfQuHpknkPTemrcO6yBnQ5ZsMPA184S
UhdlX/dJXXrwgbUM9e57RUVsXTZbVuefu7zvFTaMLzBTJTJja3F9XXZU5J+GwXoiX1w5hrqNYgiL
EJCCgjX5Vvi5Vmt+hGnPbMITWkw7QFyH5aF3qXibC7RqeyeL5lyXMF3SKjXyinNPsx813bevb6QS
I2U+Izj2XX/q06T3N5dSu6ctWEyB62NLBoiemLltCKNNKTil9BsNfT26Il4QDWh7AvxxfS+S94WB
2s3E5uqdFI0sfKwv7HjaM1QtzSue2Txfi1EZymHNkUSJt/g+geCtmzuY6barkCA9NyB1rxtpKcuM
ZZcpyBIbYNzTOdo9pKL/1wYyWoW+LSO/hiv22b7S6TRpNthjmSZVF/GhNA8w8cfr389Yened+03H
z8gu1hCsrKO/Tolg3W65YZcqEl3TdhHNFm16TQGQGtKTYvg7joKRGywI4Ro98B4qWGzn60PFjV3q
R+xhSTM3j9ZLBFDNQXLeh1ICkkxq5beq0KBAfDaT5xu/DO75PpFpuS5usRN5Mci2ywdz9ImsNM+D
TBh+2+1fo1tM1y6ibnl+jntYScQEAdqHhpVSllk3H2gtgx+8W2En9FxZWO+KW2qFk88v4LtmnXun
p8vf5ZbIraYil5qgfhgv6YQ+WOZ0M9y/Erev9GNql0QoVE0Kw+MVLw//1OPhBKUDKf5g7cRjo927
0MTNIWc1E4XDFifZ+OKQYTrmsnLsW70dItoP88Pdd0AAX1MxHH4bGv3fkiEOyAqnN7eJVGKD30ZF
5XJReCtrUBZ8DHvo8bjetyCzM6pRyWDeVSCOVaLIuhW4OdBYDnDfiLrBl40cuPYOI2vjx7xQkYNn
CxGdSh6f/BTF4bM9RaoDmm7WvBNL62W9Qchanz+hNkzLoKcnYhJiv4IYt4xoRX1cdkUEKpZH504v
r9BEwbemiveglkfXEWvwxgtO0CSbQ70OANcQ4QBcx/sphLao2rc7JYcfg/EqMjSGlBn0w8uaUWcj
6Ocp9xG1jPMSBwPeSBIb5Ryx7DFVUdg3wtebHsgwkbNDICOX0RLb6tDf7PjjbK2ox3sVdngFMTA7
xxRrH5kEarR4e9ez/vcw32ICYnfW1TBWXUhFX47R7jJn7s+TwNg6anHsQsBPBY5c8rkDhzACxbPC
CT/HBb/BaABtQC2aV/mSiI4WEU/mGl9A/XrWEraPecsxCLZcin1eMg4kFoSqRcZjI90GrFMsxtIZ
lgd5+RfkNNdOfYPPaumOnff3RP9RlQO1LVhkHMA0IgspkW1c6yreTVA/n9vBXLFleDOwXqRfmPj8
faBv27WnnIwiXZNJf90HGnjDck1N7sOg9KGjEWZPlgop7XaYrSuJWgXQ6zf6BY3NDxYycWkl/sFZ
q6sI5g5Ei0VjBJLWMS1cr4WhNrJQhZmGtrzXJDpVhmVkqfsURbDV2KiHf2kr+guNPfT5xHbmsE0e
aWnUM4hHqDfIM49x5H1VXH6+NW5VS0yB5iGC58bJuTQGX7UfYr0OlsM09/EW3h0BOAJd3ZUQqZ0b
EDdAsC4rn4bgvFRjn9QKh90Sx9c/H+lpLr/iKZXTQUt9A7YMs04t1UgyJ7RJtaEcUtMbK/OTNqAY
wNOF/Pyq0GSQOlAOYY9mJryQ3FKNYU1N0HNtb3xnEgNwmiPdhyBC88RHRl0eoSNu+WvheP7I1gf2
LZinikJulaU+WVbGZ6EC8YKUNhBX3nVIZT6AEAFQs5Rvqz/umNEUOuWck5wJTIsLie9Hnq3caHs4
K6QdxiN23HAMreT1CTFHyMVenl/HJdpDDORNKcKZW4daPj7ZKlbVsswS4d+Gn/w+8a5TT3H7Oufb
lENOS34exaJAc/csKhI4R5cTB/WDZYpAvmDTAZDe5qhIp7sOg2ce/zoM5co9May4OmsPPTk+eDcI
QhAmICC+I2yGHWpVd4zWFstYrrAByQT0cV46D8AAYLkY5bWpUNjo4zfJ58MPDhigIptsm/xMjx1E
hUuRdvOEDWArXnbjo7Ho2LxKyh4VoKsWe775W8XPaTgHeTb+mupI3l34VlkMgOsLrB6vyrRoXtK8
AaxJk+ehcGvCrsvBxkURq4z9KaoMY5Yhy4evi6/hC7YOxif1IOrfKSE3hxEMax0TtsumFwfvn0Dv
RZ+WXsWANfuOgc3+bdy7/1fmW7ci5bfZTGzVsPhkMgYmTzxawDJkAN34JhGntFSq9Yz16z/0Kor6
Q4zbH9EoWx+G+x48w/Zry9MgR9hcpmxJqT+/stUYF+n/hTqYfZzlsM9sp8kyIkES12Qs/gjIH3s5
UrHsxLQka4c6YTIQE8bgdESSTyCkqVqQhUKBc+DbzJdlDjHLOMvP+IbSvwBQiMwDnWNatiO+nOJ6
StbYMBm/15tclBKrFxYMsv/50wFN2sljPceIrrpO5QhOUSPIX1Vs0Pw/IFHzUaj7NkTTHbUJ0xBG
tjmrlxv7hjHXhFHv6oy3nY3T+W7C+PagExZlMo943xijb4ionohrkBOfDcOTFn2kRrnqZY+EuVlk
uT33JI5C8QV0CHobEBfO6YUxWw3ywpFe5RJattI+s1EY3sKH0F6H5L+Iq7fdGR3iHRVJ7yt9+9Ig
qVpzLj2u6qayhnoRVkTwUkov7IYuP2CRq883EvLNJWR5WMEEyRTWDkXDVKn6x1fDzsUyhBkNHa66
+Z9KPtGQkAS3gFUbLFckcx+/Ns2FYsQIGrPmMGpHX9X/nMzxfG5jadfnb4SVm5DHyhpenFVkELY9
C39dUV4ct8ZL+Tml8G+STfmUKSv6tJiXbZYG4zfL8gTRLNSdUCxakM9YsPGQQGBo55HO1v8kNFmN
2TrYDt8bEx6wUn+UsasEfef5qitqJypjFr6vmSwZwJV/RbeicOF1aCdQTRTzgC+YHJxNhsgGStsp
NWXhplTPVdsjHQ1PW9wJwe63BqnGrSvCZtLmTiyLd50BlfLiA7GQXcXSO+D7M7GQK8UXRGOlv9kn
H1KzlDBLoJHx2EmOOZFYrDG8KQ3NZuV7GCDHOeJOdwyuZuwXnN8HlYA99FYzXWzJf96/c/KIf3KN
v8nH1NrxdFAhCQ35eJjIKFetXxQ8ms5A3kaNDxTnucd6graJL77XLtEOS0E1K+lenu/3culCQdSy
SqTNt8/qL+1KN6Td7/fA6wAhdt4ADQ5NIXLQv7k33Sbm9JCr8h0AP1C7Rdgrc0/va+h9lYjVqG8H
Z7PbhvjVzQJpMSHbmOePPFr0qLKy0LPIMKwig5qguf5UDSPm0PpCezQiibt/lEaAH/PeYwhF0Cjo
9DHigOVq5aUU2S1NGV4OqjFt3cngnVZvXUeRPG9Wp4ksPsZo5F0m1SjmmqwZw79JkDbigNb+cFv6
VJdcPcvhw3FxKtBtNWg8VsGfFksI2fdSfmNBufD/iAzK/ru7bMX4X7yqTvUP2xVh3D7UqzH1dmZD
jOBdrrrs1SFSlvGXuEYWEISCPI3b9YLtww+y51ciAuD7AesxNZ+ymRmN7Z76g+pCdvXFQfEw4iK/
1d3XCv7vMOZrf6M+zGcVr+axNefQtIe/3UXj1X4nDAhgOgO2Hdyh7pQoPxRgF2LwLErHjNu9LGo9
OgxivZX8iXVbIv5y3Kg+ABZCgHkbpW6kV++IMICg/meOH7LWlioVY2kUHHKJm1FWfoHrl2mnNyRV
uS/d9Lfi2Gof3m3O9PGHA5ws3xd86mkziF0H8xlWPfCHbTX3gYqvoAkS17ejBC11sbHWu0Y8bJzP
pfvlxeAhVWF4CIsz60ippOp54CdSgNkk/3Ub0wh93YtiWO2xk9lvPogbANqUqUa15YTYsp0YZYCm
DoDL/lsqyOsmHRDMjBNld0Hs65yKEnJcNBKLpHeqXQVxpHyoXzzVP/z+e41IZnB/Uo5Sz1I9Wln/
24IZ4aVZSgpTucDUKcxDDyZpkpQEASJYrqaIeKHxa/I136KtPoV4U6Ei9OdThtdWDrZ9908aQFdl
2/wcm1AkJ38gXm0/ED0d3lxpjKd7adg5Bk2GgTCGY6ID3DpXms+BdRVM8tFRArrd32IRknD9xj4V
LSEKgrgKcOR50E7HzQ1u4L4a6/hjjZUKVEbUy+112e2qbYxURMyvIKPDZ9O8lhzynvlbO+bf3wwJ
T+K/q4PwWS3js1p2GxRPUB+iPXwmAKHkE4FQ2XphNrVr3kyjkNMYdQwaDsJ2oZiaLwzR/mMbgyuX
xgd9HsUJvzHCPChJYSNZFEe9n39VqELpGduLWOj157BiZstXzEzATevhAJ8q50J3/cqPXToIHhCa
pxi0QhPIVq+RB3KnTbUjAdtmInNmUjTREu9fZn6V+nwMNJfdIu2YqjSAitvDDCwxpXhXv/T5zokk
MvKWbPe7Ndf8siCUNJWdBj/1eJjPBoi4oKFCi+N2cxFa4jtflh23zWwwTM5f7GVKD4f1voCDQ2Wd
H+8MfZ+lSE0T5JMyTJeWia2cdgbn6xqVw3tQAt39NQG8WvMUQdt3PB/dRw8CPClXwkkj49utem1F
4M5YXGBohPTnBqZzK4Z224dMr0vfgIUClYR+W3W6lf5iD454EMdUe/XVXSEN632CyzcYogz5Wpz5
nJo7yXcISuUvuMvGeWpcfeyjU4gRBdLMsPbQl3tbUE0uxMGhEDa7IdVGgxZkboBbD3uiypEFimM/
QI8rJZtmP0WIkwoLt9gB1X2M4yTCvV0q3rTOkuORf2UvGRiSmUh2L+rQ0G3k4xcoHOeBrxuJyPSZ
mJMLpzQizjlOSy8Io3Rdual7+pi8YA37ilXFLu1uYx5/FgoFXCLZ/vWBh8yWPX4sFV93xv4S01Kv
BO5Cp4Ju+Mi4ADq4518zkfJlJBRvJvuFWccAQ1LsoFN0HyDHFB4iNNwhe2yYl3BBIasnu2/xmhlW
bLWBRL9ZiRbuFdreiauNQ0+qUPJHg80BVtEd6f4nRd5ZMEuJ6+Du+rfnpI8AyGN35jCTCdlnKRIp
oD7lEMVPTQU+PBYhkfCbFugCylUaXQG/Ete6ae05mmRb8m7VVcdTVQwVqY5AWPtySOR6BWt+VZu3
yh0SMWwdWZ6HdHOJMYupZ/H+044BzLsKfO+cM+k3CgFfsy2yCX23F+avGWudcByspHeUYxTZjHay
ym2s3WPnLzQTQQzFamkY83jdN9EAleRko6/4hDHHpzvyZlRYlKcwhVCTjV55Tk0zN5eXleB+kdnm
oW/Z0oJVxURVRlUaEEnxZ0ZxARb63deqEE0f1zlKizJ0gc//0PINnx0U5LYz+P5zgIUpItR0lJ9F
V08eONYiqYiPYEEFtXCVss+2qiJbFmn4Om/bTd4+cPwBeG9PldTqBjy3GcK04/twmiFy5JhDU0GI
llV9f+Y9t/v7jH+P+LG+NMz7Ev6BEUuI/BNHYcX23yU1BBxJOEPPrIb2kAT6oCXt678Q9L17EMW8
rjc8rDFeJ0Wpiky7zUwfoVKpIA3UGz16hOcYe6Bn7hbD8EnLYSnfwIp+cVD5utRfIi155CVkwMuK
kk0JzR05qSZF7w2QIRczLRF/LO3RD7lm39yQ2+R+WCFgZR8/1EEDF81YbZUs2thcKolEXTf1VZ/M
jEgOzK5NjSBnZK1Jmn6x2pNsYj4vlUAz9SVzDdrTHr38RPTm592faK7QVpOX14WjKZmRpr/6qqBp
Gq3Y2riS94oDg6Z9cKPDAFGyren+W/5NMR+FJBnWI7XqhH2h3yyrTq/JQXyU3vb4i11eGhfJ93+Y
NcMso7JNZVZYXoU8X//sWqxZDDkZ3FQ/a88noiaVbOKjKJTKz8Ig38caTGkIQuVh1zntZaqJMHHz
+CzJ/RujKgjm2lD2ww9zxc2jDXPUUxPGzDx+5c3U8avZJztADpGS/Yp1LGudn+JlY18bFzlkDxFF
j01b7pvyOGNlfzRj3mPvweQ+GSj2zfDLiRdDqfAJUGgQZOEv45XleuufXd6G5oCTItK582oYv03M
wKGmITLnlEmlIStbFOKUySYG4G5X4XGzPryFGmuhQW5Tr7/P5DxHdN2cT7qACCKTMquIL98F+pvD
ouvqE8vB+qHEhvg7mAV8yIsQVBPI2kxfgDKAgI8U1ebehJF6A8Q3TKOYvrJZhgSedh2zsvXN6IMH
bFnEA2KRr07maEcTJNsC7RGm+DPb8VVx2WziGbuMTRAZD8tmpAdA6DqTs6u7B6NZBuhiRI1aaKGt
qRDIFwM/JMJCXshb65cCo0M1uFsWns2073OCBf/mGzR6+1UbXVlQ4GWnbLFcCuJqDuQf8uNZiHE4
xlXilKjFk9+mJh8bNOFdAZpWDoz5YWLsHUkFPSqd2gKezzygQoFbCHPKsDEllXE8hH/r6qqz9aSN
gmCTj6VHMl/kruZm29jbYbPs/jDOHH2z0Fj94x0nInnCaLzkGqxodO7fPyqgp1WkbjDU14eUhiD3
YR+sVghN1BhOabqeCneSI/D/q9WlUMzDXuffKR3XivtBPfJ4YW3yc2ZQ0HYj5fqgQIhgE0CtnydN
BY6HFHQPBK6MljkzsyFFmTXYC6yrXloClcgsdZjm+PZ3nP3yO6YzzzSzRNjXP+L3Nisv51BeeLIB
6uKDcc6oHx145NcHDYP/A7pl47OTFoGzhqDXmr6IJ0qN0OasliDUPmoilUtNwTPWlNaxSuaN7u10
UbDPYVO83UwnsfG7ig41ucLmykiAd5la0oXLS605koVne4V8JnXJyTn8QRuDIyH174Rs6ZmYve62
ojXPQBDPv1JH8KDj/0oxWoTO0PpE+1HzXvGoHycgXwSNVNb6ez1yrtJ89WwQ3gf/iuSd1zcVsWXr
g601G4ijl2+SRSiM6hm/7/1C7DVNeWtkc8nE5JL7tpIjG+wRQLmmePOA+ZHKP0fpZMHR2i2Uh5O1
fKagFoCRk253q8d4Ga7OQsjK6F4jzt9VQuaC8JE1i2APuj6TmHrXSo+Lh0VNiGmeseFNhmgXwNBX
ZGHiNBOgaEDqTYznOV1X1oxCy1kERvVotb8jWHzR8Vkr1lJc7ejjJiYqzUQwfra+196bacmyKYNX
HWTjXQuI4a3CZ1S43rs56wVgiyF/4MA+xtMyzEi4N3o7lgAdAameyz7BOA+9GB6l4lFqJqUMcKTk
c0hpd1HAf4R8Rs8gXrRsEncez+OagYWdWgj6Oa+pYNxQeRMXleUP2ghTnYrMun7opFTXXn+sDAcK
TqJQi3pm+z3k9pgwCM7mLzumGQfi1sPIhXAssqhMFw8gGF20AZ67HH9FIkZLFrOFpuBqc/n7dzQD
40i7cyT19x8hXsgrY7AfVkVSws0I/do4MHIyUjpdpvH8HmXYN8tYPnEZ5x/dVn7K985+RGbztoKp
7vqiFT/cSG/ozUfDxjZ3nYo8qYcsj9kwz3nBnpyxxffOKFF4yuTMjxaxbu/jWIwYOaA+7F878bS2
UjEsO2bdTt6LNi7rePuzHO9Do3vkLKyqXhnBSmuc/W0S6NE41i+epGxjtwj2BELuE9XG6rPGY7Gb
D3aByYGzJcCTYS5MCtY/MjWCX5eXlquk6JmXs0bSOyij2dtyq4IM4lrnDpvUnbXhw1skV/Vz2wvd
HeEvhl2j902WKNqOrwgrevfcIWT2DjYXaspi9V4WCGDR+unTzmzCvPISryq+C48lYop9ev7EYW7c
a9msw/VPTYjEUd84I/4VpQzieFZK/rEvTEb40D8q1N6uTUp2nWGiLA5neHIOYgUADBBNfOD/MYBX
aDcl8HTolV/yQz60a80uFCqgbqgbaAfHcMyud/MEk+VNKVF5IbkadsNpLnjWIf5OMZUQSqBO9JyS
H1rmXBiVXx/sIgCnrYK+F11ChP6MkNiWoSVwsheFMZICm/0Zfp6jnZex/r+TVuxXvrIzOei1ruSX
znUUKK3b62oup0Fe8Fl3K9hwuyM0pwi6h/+agkyaXaP88cMRyY1WPgBBqckshhqUDZ7IB+gMU28S
EFictigvrf6KhJLFJhkgRVCCEDEfwJdMiit0WqBa+ZvzpKdINnXQzx4HnNspzwarbATpc/ZFegkh
GxE5d9HaWkkpAOgFYGOB+to2+iiK+8XclgjrRTpz+oeOJPSCA5tOaLg0JnWLmVhagEBkIn3HjKut
6yQ0ig3+p2xtQ8PRJmVLwwHGnyR12iXgt/k0VB5oeStZsBQSW+ob7xU8wGEyfPFTMNeAdrRRofvo
FvFEl+UWf9VkiSeQZTxqRG6wylKl89RRbHxf6xxTMY2f94qoUORe0U/ET+bnzYCvHPeDOZAT/QK/
GR64RnzK5bThV9JF81N7qAmtCRhiQod19/bs3oYOrKiSni6qd0BmPr8P+quOnRHS2uzf4Jy+AYMI
DlGjuZXIMPOY76ZSocC5nrBk8euIB0wN1tULL2Ox8SOYVqrs/UeGQ9SL6ckqYu53aYhFvjg291oh
pBv5e5GajzLTYI3t8iVWAAnGRXOAMfFYy398QorMY9J8ZRmtLSqK4YqPd0AF75w/xIXiucwCSfLv
F9rX4EWDrWwvfYkX0Ai38aaqKgOQbMyv562eo5uO3QAc1c0eCrCnBofAG+/uCSa5EGMNBOmM8N6F
Qs8TSYgZtkOp6L+KKBYo9hp00tPwSpTAy0CLZxKvbQ87CQXsxRbngatvfppQcZKF9eEtD5gmp20Q
0j8SuP0NIu33O8Yrpqr0ZjyrJbvAII6CCIwi625nmrysLNt4w3wqUtmD9CoqFoRwJAkf5p4wCh5C
ZxjFHKJx0bYfOicCLW6MEUna9d7Y6yqBC9PJ6i03lxtgGc3KoLdWbsOkhCmcbNhkqDIU23xmOP9/
ftNaizGrh1ZNvA3KF7seNlzXSKwyZD6SQ8eoOkoKD3qbzuJhpYPtVDcJCadfph6+Fs6w72GqfDqE
aWc9I1chyFARjiCjk03fJZ97GYrQB7uANZoYDXXYQgZeZ7nEXYeJ5gp0a3G+sIqA48IWE4/VuM7A
My7ixoij8qIuFaIaZyV58wKcKj/TkYcU/1UkmhkNCU7Skm/UlfMDKVGA+C4nOPdc5rSOFDDDKv2J
awF/OSQUKNoT5vfX7H/er5mMrq0GFhUSV8YDnuXFKe0dvAuSOxYUUvZmtUFJYm/AK4gUNOlJwnH8
ZdfImW3UC4rOl2H1vOp2s1roGpejNHLxISVBRbmccbxPzyqyuwF+pJ7tYVm9Yi06hJEKs6pqGpkw
lXkcVMEDz/tZiPNUbF0Nb9Z4YbnlvSq3pndJofS4CeWUvAXajJh+ZYLiB0BqGsBP17ObosQArqD9
RyD0lW3hZUnj/bcPIqJO3zpZC5VZ4Ei/NXfGIxrTQDbeb7uYSPuHsfwTWcCViteYgeytvAdOPcPU
bnnUcSWtfaJJRwJhndEbbV+5uIg5E6ShL9BA6qaAIwYJ/bYzdVWI4f6GJuDM3bjx2IuQqaVrIypZ
BJm15dH2rN0k5P7qCrUewpLUE6LrQOes+Q7EpS4G8C9k50gMGwnfMxvLQBN7P0NK+p7xA0syhJ5M
eiCpvQOg9Ay52ksm4H1+cV6iEzHIFm6Ocpls4Sa0LABNAa5U6fqjAV2ZHfwjnw/E1mozylHkm/G0
BG5dt9+RrPXlDXuUdbbz7gYZDaEQIroxSANyIl9tAZmmSmgEFxzJ62eicH+6xWO7Cdk1vsBhIhTR
T4CjLFYNWXkth34oxG1AVQM9z9cTnrd6TpYOq/ycsygVvvN0MTZQQnimQvTJRnPQT2RxTBQFy9Kh
unkmZ25ZOr9gnJNBx5oa32nG4DQ4U3vka2yGNZ7A1zomcFJS1aUyhoz6UasHmrongom165mkygHM
DEcHKa3fois7Rt8FKtPrE3wzdC3TRCsnnyIgpV08W3I8E2o2BA4pTojtbv3GalGZv+ag8ANNcDgS
AM4hBncX6feQXM2WZ0okAtU1nJK92zXLQB6aNUigMCMwIHiv3i4eE9r0sjp1Mtwkuc37QV0szZS9
ygGoCS7OFSczyRG3VmLJVVyJookX2d6DALfERNdX6gmn0iaq9dPJJvEuKrZsysdm0dgiRazbGC7u
iOEGbrAkEhUTdGq8pBWoxlwZiMMIi3q9Zv9FWYPbeAHh63RK+EGkl0kJtdfo6vmsLLnd2Tjstodx
VfMxVI6sYxIJ5m+Vw297knEYSMmG/gCnbCPRMRZQ2xUVmkET7TYsRF8Pc3NpnnDMXdCglFfy4cba
oXXCxjxJmKedbQ//VIECR8J2vj8FCKptqOgFqk84bWUt+/mLpaOfi+xKlwwIo89UpEvNMGNeKpe7
L1I1ACs1uGocN7MoTPNwtQ/bmKLvsr+yX6hKTxjy/iObt8I9oM4nhQQyLaw/aom6dMp5ouG+hoqj
8I4yNYMqSGNgXhLZtsaOBA5wzX6kco68TQBBsaSzp/o8B2SUPPM7M2PDRnGx41UtxjK/ncBk3mXU
Ak9/DiiFi33DCMQPhjVbijMD2LxFM+YmjHrcl29LhpR9z+aoubojO4K6+XorrmgNIfUMK2gzozOX
1IY7cFFYm+oZml6KlHX9OhRsSA215kFws4YsIBeb/+Eg9t9bgqaIp6Zcd2OjEYMEW0AtFJvuUD2S
12xjZfUF6i8YPzwWnL8ivW44zCDBraGgi2paQxbWJmG6xiaJ3U6PkiU6D1oBL4+bqWiTqDJEw2hw
ESuGhQJ4Tua1Rk5EbQWXMz4ghFvzFkqGzSaVjyowyMtfnYkACA5r1qoQwB+EJga1dcpr2vDUfy07
7UyyxKBSJXWc0Dnt9eWVuvPG+PXxtFGaQeE/VkFJWKFJ5KcE2il2tRA+33bSWJCEeKQiktRU8afF
SE3h24WaLV6WOE4btVwtUmIhm3OYmY36OwT3Iikrdh6R8MzH2g2sztfZBX6xqMQ210gjn0Zid7cl
KoXccTFYbmHh2pYd+LUP8wihm1fLR2BkLainYCu8rn0kvo8B9iKGHp82oXYIanjd660eLrU0AYWi
iKAap93kokx/QmsWofP49ktNZeV7a/Pg+4RdrqhgGgBQN0tXu4SyA6U9a6c3on4lmOFuophZVPYX
LrcvjWROeMM0cMXPDUwbxNHQjsVlPgOirkK8f4Iv+o+J659JHMTG2tI3tprcQD+ZOgFiJmYLKcMJ
2oLWgCKHjHBW4A3NtgXFU219fsvNw0awwIfaF60VM/UFEJ5pZ76p2emmpPIdKJyIo6Ua8cRhANiu
lgO41pTQNCO9mtYqTRKXIazJULhtkz6vG9tYeEpfWBi26Gx50qC70nkgOP14qO6DPJFLA3o6SHb4
/obNfpG+IAZVT3TlsvUZWoBQXG7lTUuqMMhNBsFzg1stzk52qXIiO13s4TLVTgTeZu4GhyGEDWTJ
MPWOlVSIThyZjK6MAT6UwTsuCWSO/iFLQHxjK3fpx+JQ2Ie5WrEW2iavgApfhCandP0TDCii8Bkj
1fJNMT8rzxr8sWhYX5gU2BUIA8/OskRco0YPaty8/ouUCnCXNtWGmjLp1h2u7Nz86Jv0Ac8JttJ2
U6ooLNSs11+74J+S7LNeApu164H89UhEpioitotDCLEFTmCjYXTiAc+6o04h9aujzrPDXgxoyDtG
9ErA0JPP48pjayrHX5UDDwAyNgeVlqVuLoIYXk0bOoNIUnLWVxWyEDTrkUlmGYiGcrDBYENXdHHK
tXqOYUdlrDxqVXjjBWfYSTYPFg4tzxvkmDRabHg6sRHAJoXwQPg9Y/qCtYnzLA6VJ3nDAkFYB+ec
M5il4PElBHG3TgzjtRc8rLmYUCnC4mbt/6rmVsWEC+PwANuia5J6D3Br8XUpSwceqpxjBv+BHo5j
MKb4RZQNODtyZmz7us29lvK0un2O6oxESwGSSg2snTFKTp/D4s79iYIZ0Nyd5g3JoeHj8Vm7MucA
xcL/hxMwb0gJZ3C/Fo7AE+G3C5xqY/7/ZzR+OefLE/Jzx9T9ke87Qzwg/mtoZoVnQ1wbUz9nLV7y
OpHp4UBkqLrgneuOWWoqZ5XsT0oOyTUI8QoQsQTB8VOrw7LOZPXS5Rjp0Mj9uSeXW84DwRf3Zqov
iRq/tQKyPusIgzI7gP6B9Xw8UWrXr5uqg/WNQuwWhzszXMXVDcuHSdpNySZPfmKZ1CI/iQbRiNYA
IJvYNu/FRQC2ACTM/KiEscPlY/I84A9en4wPcJc2+hh++FisJpL8Vkw0MuMlslvglVHUf5+9/UpR
kn+nftTdmE+4ArpC2BnLhZpFQa9T8D0f4x9jBQpe6QaB1BRNdlsXNOk/9FTp85rbLuvoQ7ubyQMx
YVNDbQElsict1UxsX9l1gvBujFpZgY240G42JJVfRwUZoaAYa0HH2crQz/xp9QmTL+csJLyX8vsj
IX0tZAz7LjezO8B0sqKoA8OE4j9AwZg1lpHegdj00wwB4VIb+Oz1qKBoqCavzXigbz39BUi2N/4g
l+b/hdFCjOOfwzLw8yB5sP0nDoHLnJFjONlBf4hQI1f6Qzi4r/0bcu7sFIyAXP+kzIJfSqY8K85n
VWd2D2PNYlrOtoECSrJ+Sdi4g73J2SAyH5uYlUCjVsUgeA6XfpJvLLTktLEX9LsgZkUAoJtVt3gC
Q/qksEEIUohUZnHad5yprf3ukaPOR7YS/SsWSLYB7LFmpnT0exkz2ErHiaiuYNS7K1I9oDLnjbp4
iEYeHne45Ngn13g9NOkHyo7x9jRIT0125hgIWNO2CwMJVEr0j7tQRSLQH5BFBjO0/c/9VxVaoxTK
K9CH9mYbxvtPPioDIuHhJ0oO4rl9TC6rmRcQv3F+u1y3baDg5piQ1ddU/e16lgJy1tM6tCLAnFHh
5TAl9Hg+X5/nXUEMMko6NIQBsy7GYAq0ZkRVOM8/NQk7YwzQvd46WWphApJor2v/7xenILzZuQ9A
GCOkQEXpY1i5d40ZK9KYlSEKfDFupnMxzBGHvkDn1tcKxtOL3wEy1hB0ms+4kSUUYb4ajQ0gC0xq
InXyCv5s6XLCxuXBguxO6Q1o82RAIt2BQa+WEklvGTjYVikw8NqdZkiwWuR+p/icdpiMgblKF4Dj
A3zjWVmYt4+UUivR63tiR0iv0cs8ZFCS7tf85jxs7Vl1ew1pOr5RdC0CqpSDK0LT6gc5qStV7uXm
TqywrlMx3X0LZCR/FZPyV77alIL32lcxr8eigjniREQB23An+d3P1SxMtwPTZZVU81EhMkld/WO4
tqq54P5ilfNsnkJqtiRwQ4VD78jIcgxEnnkjTT20D1S4o4Efgu8KvlZVmgVluyt4fmDCqHqIUwfZ
/Pld1iNUmNkuxoMCsohEVNbVsBIYv+oPIF7W8A6Pv1k0DYRnSf0OMjOEVmKeiO660JTq4FH6Owl0
uHfgwSkE9YfDxurl80cze6eYLsrFDlGSSXqJ+/FXOvja8Ji4avM9qhRrRZY40qb//2C17tunbOi4
o1QrQ8E8dY2Imf4RCNw6/mgbdmBryyiNZPEngN664j75TJOm6OWl2ONzZOUR+zORQbQ/XNDRj7W0
Hs1O5J6WCe0Ocjhx5JrQ1NgFj3bTgcqOlmvWfd2SomjmZphXG5zC7cW6yZH/m020d2FEJfB+gGEk
BbWek/tgE6+JRkG+Vi/+miY/Qj4pyWe7Z7u0bqH6ENPPHZk4r63smYfvsvfmbrknUx9PZMEmSbUy
Fyo9Kkerqv9XOTqJWf957ZvPOTDdiu9wtrY2ZjMrGrPmOg14MVjyhXDxUm3mOgTz6XIdqWNsMOl+
Eje+5r9uYZUNcMpwMgPYgHkVfajJ+EC+0y3jI6QfuKl4Mb4bXMmlcOprK6tGDF4rWz0J5bGj/Nzu
wvoKDQxSviQOe7UUvvT4+2z6eDuRlPVY9lX7R73Vk4AMdjw28GiURs3oMkAeSgXQ9EdB8dy3a9YX
7mpbjR/oMLEpPnky2u9doa5IfHdjs5fdtQbYobYc6g/iu+Kfk+xl15g5FTVR8DJIN//WqBWOild2
HVXapVnklbKbnYqmqpGB00P39N34Cn4Uzm7K3VgTL03icjuJBGn2qkwbF8XBr7gJ5Y2zxRhyke7L
OiyQT3bMpsScMKoSUxawdlcoy3aCIP2LhyAmzXeSTVNuSrA/0OuGMJDUWOvNtmC8WbX4LFN48F/+
QrBK4fBFcS97/T2VXxGTEJhjPaBw51Pct20UGVHyeFnM6kTJJJaTwsscheKR47qKkMXA+1Gnk1tc
zc0w59dpN3s+m1q9B1ESedqO3ehxCe50opTkPkKvrE3ifytJcfNhPqSMhjvsqCIrEij1UYYNmp0T
17jtUVIPItL3BZCNYathvxa9YzwIKiSstqxxiOdlNlT9usVd4NHxiwNYeMfnjgbsYNiBUQf6z74b
Gdnr2VxgYYiLUnt4zdnpWQ3yMkjJF9vdZgzC23oGRGlTfm4B3hhbYoUy3S08cdxg89kgMYG8wSo4
WlKC/TGnYpbKVmL52EzsPIa/hvSdsGMgbNGGGnSajFefRK73Up08ruGhR+73DDZTBrLiahdi3k5l
EoyNYdRfG0Stzu5j8CR2wVNl5z2YS9wYAjs6diFulc88CZx3uui7C2qyf+cBvYAktvmvolwRgu5J
/UNsmLCc7ixf4LDzr97+dhAJwK95md+eSexkQU55PmUOnfRAyaLyw2xt2gzDOA9NJNvahvbI1kAT
4Hss2QFkcOGb/3hiTYSk2NoP4H3dBJNHFZ3XvsHmxyZO2hMl7fwo4y8G7abiF7Ba3R0FMOGhDWZn
StuLj7YOYOlRcY+TFoemjgRA0udIHjMkkF2C5xRPaY4ycMDjuQsSOtQRC/6lNlK8rVfNfSLCMqQQ
4+3XoSi4hmNqbn2M/tmjGdewH8P5ivLwkL8UGU3t7lrGiNge0+G1eIfOmiWKVX2Cdt4iGdaYL1xx
kMNB5A2JW7VSNeWfr0nZJ9Wy+99+j1cHlK1ZwI+AtG/tJr4/TdOolXKWQfBkdIv9I/8rtu9lV9lX
DTm2nrNDc9NopaCshC/kc9J5Vj7yYWzRhyK/XUyXYmXqwVMs62XAzwJCyqKlKXoV7jUiWkB8TpB4
6342n9KyxFNiyoXTV3FjzkuGkOWmJEWgeLHyUUZRghW9vDhfniMuWlNWn2irWAINwkwOvnPkBUum
V9uibZpZcak5LmKqGSJ2arBjMG9omWkgsX+5XmXXPRgiO+SuaKc3A65bG3aXRFj0xIzR5N4Deb9I
B/UdXSYep1FBLGTfN6eReihQAWrcexIOJbVgSsI8f98wE1Qg8/LeXD++IVt7PRDqzLwq1hbRB/gK
Z5ms5fjunR+3gARqu1aIorbALcql8ZY8McIO6D9v7nyw79R6BborN/qnl9n6+PnbIYYXdWa7X+Tk
1xBFn8KG3FXdL1KeAXkIgWglo7IWo4S/80sEiScCkkvAHjURpFlnJ4PQcJSxjGqkbRC3W2si6CLt
vDTt/ucJqRgE09+EERNSylRjerPGb0glNDZi8NVip1iKrnAnB/fJOLQa6sjjEf7NuzCdct3G9YrO
VskUep8eCBZRmRltyBCIFm6SCXaLd8/tFIrN/RtkwcdGd/6CfySF4fpjmXSmg0olO0yIsuhRZVzy
tJVsIZcliY1Pm/O0WPoAY+V8R2yvsHhjH9ZPauOpM2UKdxWLg5vbj8LCPn5CodgoD3S44ZAat72Q
2vVNiNqEOZQxFfyLeMvVzQeRmHt+9CoiOCKIdq69t5Fc9aVXi2+fNynVhLopXD3D3CeYvO/NfkOA
YCGqu0jLgLAR2971dA9iImMNghJ/62UjDM0bYIxU3BNYTOFplj3csR2C+BvCQo/LCVXbhp4wELNF
n+IAKezPWe6idBpiAPRa408wr5YpuY6E/BOhWi1E4hj60bsyu2wTApk4iYPTqQUrw4evckob4ZrR
oaOkMWr2kahxa15sK+q/B355MSh7Y51ih4Ci5c/ocuSfk8BcQEBaukxkSuCch0ytX2PKvz6xwGvB
Kj88MWTwMr1EbNmxxroKg2AeWCy2GjMrMAF/7CVNVMvlmyrYuZ1HFPS6Ntl0StGqzQ3wkimAJg2I
ylVU0Rh7NXsBqvuHiiK1iCLRSougdFwgomyTkZ8Z4DeUCIOGs5W+FQXU5DlT+ROZEYsNvaZeQFIX
j29xbnJcdTSOvLhhoYzgtco9ZLSEj5c+KqFrxjWE+HHKtGlipAuaAezW/8zgjZhIrum5D4O4vqC9
QG79tB/Pmc/ahKJMolWcNet+1Kfpkq0GzPYE1D+TOw9Kn8Nb4xpxSiF3VjQlKntwCQDkecxO0ziw
UMRxkKowh4n0hc6IPrnbi3H/hiXaM2D+XKu1cg5fjbUbrEv4YLhNdL0Sw+gezjQi8Y5UYVAMYEMM
M8dek5pZv1FdbV9w3Tooq2SNoX1SMQr5KCYKD6K1wMBSbloiOhsTrN2UefuoGGvVIP+jYNL63GcE
/GeJJDL3VFvQhQF1jHPj3FMCUHIqg9JZR+sFlw38s7Ozw0QBsPsrAjpNS6vOSRDjdJTynr3VIzhC
qkhXmBhLiFjM8XH717wMEA22AvTN9edICJMmMJ0iUu25U5ZmA8O3bri5DLD4fqy3QMv9DnVs6Kgl
tY7l0B0BWJrvT6Z4uUenWAFyfrO6WCQlR/+5jsIKJOy9l/ABucEkjXK+kM9ajflgqx9Jha1S+9ed
7XS38WTiDV2oB2H1UO3aG83EJYjwf7ATJOZla8+ctj6zp0qvEHIRjyxdfWifMfamUIc3TOjq5EoD
3FFjRm/s0eXuEizpr/gh/OZH/fbxGMmdbI9ldh7FgWtEfQCCcEN5bAHURj6DHtDbhYHegabAwERM
HN1VaWO9rD8SWW6UBcpmDabMBYRoauSqV/xBYEF4CRlYqm0KtvSit3d2JlTJstFrysfosBkBkvYC
Qz0+F6p5i6FRWjaLdLEtQaeoBkWgA9Ent3fG7NgRVElPcw7dEAY9sTPDqlUmBOR5vb2CStwochKC
H5KxLzC90Jj+dAHECfulWLrbUMTP4wrwmgjoQzlkhc4wOoAQahkXr9OBRRmhtcDYeHDPHyw0OSBM
LTjdAwzbc4LW92ksIKtqTFKyqRtQgJ8naoH1fDjxbPQ7NW6/Mj11SBOP/3Txnh7y5bZY2g9unT6M
mRU6fqAhULLMhsOcIhbSbht6pe/BgilwsviVNPLyIx7IddwRCzes8jLgKR/ToXP+aT0FfniMkCZA
zeCg6ZuZWEgDXypjQ2UUX51wj35YGUM02/lCF4Gt1SO1lUvM7/colXr/wNkk1Ch50vGez+RMxyui
n81C+CP0JipkuWD2QCR+ZBCZVZevzgNFk4YEARaDqU3xp0aeiocPK2wj6BfjDP/jB60LkjbQjYLd
qKuzqjfh5MCp9kGg4Eg1Vpk7lGOEZV0zl8FQyAAAn0uCBNFKEdBfnvcT0HZ1qMZ8gUIuM6AkNqeh
8y+gy85S4VPi2HH/XVhUjkss/8KY6FgQjhKEdwjxV9L4iDW+9aTto1xB8DV/a437FdK+G7Bm6Hl1
QMRHtV96P9XbMGMXof5oTpvE3mbHKYSpb7UTUPBKWtXB1My105cXhat4U+f1MwhcJ2QtsRnpYsgw
bY+uIyN3Oua0o0SdrJUgqvYunWF5s3gtnAxC1DsdNKnn7aPSewvhISRY1dQx8Ry4ILUGUvvznyZZ
+tg6R3bKF77h841rJZRovGfqO3LzdRAcd1szT/aGN5JUS3jtySf3pgwbRaSGyNEOIf5D0sxh5baB
3lbnL34JJhGAu9D6LPvwVciCcWfTkwDmZ+dX8irI0cEdkTCjab8FtcEO/DsenW06D8GOja1LP0m7
5V4ElBGB9L+z5Bwo6DeFMY86YupyTRXnk+ISJTT0BuRayNdMzN1eQPpUBHgg/mHbp1k+ox4glhfZ
CTzGnvLhEgoUx15Y42r8UAmtkN+oipcIhKHjZZWX2IeTKWOCrwT0B6/DbGoKV8nXZQG+jN30n5fZ
Dz4YnhA8LFmwHQPoPW3nUu0nIdkQuVJoN3ogK42nkfdbQIfjeMw4XL/wm4nBjj+IfuhSXUfTM0ho
pnq9OwA+VHfFUL7TGJddFgp4hxvD/YPYyGybF2Z/bEiv4Tdesea8tIJIIQKbTKSe7DjRvSnOjKjx
pEZ+fVXKre+grBwW9WTzUpVFsXZpHLsQ6xxLhEgXru2WPHkQjuF8u3dz71VaEtyvW0HMCJi4qxQ7
MpDFutbI0kcsVfsIKXdAZFufv0G9ieJiPTwSJrdFUyf3aE8iik9bk3F670MKi4OyiJSzV5l/b9eL
Rw01UIhcJWbnXsSnYqhv1hTvufDmUkKJCDWYzbSuWH4XCStGz7q/42p0FPuHRk2EDBfKFCm4X24g
iJIX4YYdlgViijjbNIfs9+ZWS7/PhNSTZH3bTFu94wK/mno/6QLkJwK/TsJGqE0sMhCwZsMYCYIU
3QX7aqmy/dQ+ZHpIUs7bgM8yUZp/UH+cPLCbd8HiDRHGyvg9HcFWQJL9XMWL6SwgOHNYNirTLmxn
XgD8zgB4l8Qd1lcnfJsOlfYw8R2JWLK9U8Hf1UcNgnzWjqLTzkHsVWG4nB90noQRyCW8FAoD1QAS
hdeWqpFXUyD1B4Ji/4sKtzFhYJCH8NIydmk7dNiM6AkJvqXz6q6HGhtz9n36iNEAX8Uv6s5neEoa
dGOlOpyQayHYKRFuY58vhRHw7nhCt+LeYmvkRGM449xVFOxSH+mEvkUWPWMaQWb0o043w5EjHhhv
rTeLyPJeUP1d8BhFoPVKXKKXqX39z3nkKOMBcWYEthEn7ykXARjyXaWW8P7LghyOmyiqDjiilf8Y
dkkQYlq1UmgaFkDwejxyvraxOo7mTQw8EcGRPSt+dlBIaFjNhrMUQcb0OdmHkvg4Os84WO3jGgJo
qcY7PtseRBB4Bhg6at2s1l6ZAjhjHkLNBWDW/mvIhdj/d9ydmMzypVmtqLPtz3gmzMtTARQSsWI4
xTi7RTKjeMkhVUpgN2Fwxi7JtO8uGpJN6iB5wu+89x5lbF3uayp9Ob3mgAVdmnSrZ80glOCvfObm
gARSpuJPcxsyX4nAGEc7aWezV1ZYY99eA896e6QHj/Txr9rNLSlwcWdDQ/ZXINWreVYgz14hiI5G
WJlTDUM8pzzK2HyFQCxAxM7MGYL1dEKhKp6D/IeiCt8UeSrrIVogGQR+VrKgxSTcrENrXLivKNzW
1rv98BVslvpZJV0e6m3LEQWN5/l6Yj72Zg8mqNPuxmJCo/1rMKY2Q8pw8kFSYcvYJskbJpn3IxtL
LYduYFbG79dlwYa4hglOSOTHzaZ32/0wHz1t8dqeSs3qKMUziEA9eYnip/pIZ4xWeVLWfepReKa7
ryVHkHcdiavOaMWZ2GGhfO3DfZRiL/BC0bHq/ESt5PFv4K5SzNs2yxxE1zh9EJCGG6Vx4546jerh
9i69mX2SxWw6Lg5vIOHJfNLq5eI6KumhCuJINCl8y1he2PYGCecvcNutvxiIqzPW+xG/KjYsKphM
JnR/SRuNfMWFShKrQxtbKcEXJRsc6lJSIZ0OT/OTvGX1Uot45Kzd3X/zWI3IxbsC76GlHu0d3IZ2
cVvz06kNGS+6BPQ/13JhMlMiW36mj0z69NhlG0yJOnB5dR+HZ8lGpXd8bdD7vN5mIYdluatr1tXS
Dri3hyp8m9yHnhEjBE9fblXSEkl5/H7de2I734Z8uSqLKHNI3/EvgEppuORRh9lm24Mum4kv9FA8
xLkT1GpCI+iIdXqdxhwV2lp+JhGQDd6oQ8YMJXWll1gDJST/EWbbESrF1h0+GWvYOyBGb4pyIY0o
n9VeeKtgctH4mjs4EPT2eYlwh/OqdTVm/RZ6ENsnBHThsOKR2UpD9MGoQyR3zZsgwobSErUC2kZ3
f7Zg8L6OKfl+JiphTYeDv2IXsSJ6ndvQkdJBFQVeSrr4kA1uBV/EltXvkkpgfM6qIdC74RFe7X6d
fIclIrk+/skqCZLcBwhjV8kJ//3THLEs1lXRutlVy2N3D7F7q8vTfT+LblKKP6picQ+LT5znps/T
Nu7JEq+y0rq8WdusH0DKo6sfOQU1TREgYFdO13M3rdP5tZM33S4zfba2UpjHns5UrYieLuKyQmF0
IRJtbNMEVusIgBSv6FTIgZc31nlfod9hHQoeyerPRrhNSziHD2EAQw/q4uSbNZZn6VeOzGvjzG07
NKp3HOHh3MMcFsKAV2JF5YDFDdnt6MF2cKVi+m76TkTZakmQdChqptNMb/oox8fjLcTTQtlpU+el
IFSXrMDZFbuBtb9080P3IfhJ4exGHhQUMmg+oK1NQOEXmYQuMlp9XssC91bqqdOee5ysEXpiRzwD
2gb0QuJ7PUNsYjGm/bKrP7141LBr3eKlJwqoodYHPG1RZIeJ0i6TbQKn4fnVQ/GJ9l+slhzjmwlU
mDpkCoWCRgokMr7EgMDUSVCm/YDHhA0TtE6mJ/45VIyO3EL/pWPlFv4B62lDjWnGBEfYXYhsPRKD
Faen1ZV/dRfS3yMVFKi7JHnGW0pzlcskOZlAp/Xnxr/9RWObLkPpFSAP2nT3Uu2X/+xQsFlVV4iy
e7yKiW3bNg1dtXpMhxoirKmDOtVTIrK5DVf5SJ8i2hNvHSkjJVV2KfUZhUYn2x+BFwVJ2T9PsFDD
4NwcFFKCN80aN6ZGAcq8axevtWtAO3LMrh/k1VexCdO/MN5vUm8+ldt347DVyI2rmWag5ziEbuXk
9VLzbxYwtLAHCGtQsixV2qiHMnbBqp9vLK8Wmcb0qIO4aiKUYe81oUQcn4ZIRZXtwSvKdOVHSVTG
Xped39z0nB2voK/MRRAJg3h34i/t+8N0sP3aSKElqTuH8IR5NwnaIAevFf6jpAX+AkvS3kT8+NZh
YAjGciGp+fkiCiVdatehiU+R8yp26u9s9ph1d5Azy/jJqT4mdJMTFKOwLCXJXz6UHdZZD4o0mvkO
p0okeHe7DrPToNBO8HghINEtvSCqaPjOL3Ysr3wyrrF2niaZVuqF7MKmoyeHCKJmQ94LTj1E1KdV
U4JNOvPZ7sYG+hFQGqbZxUi1SVMy8WzWagVoheyEVyHJpq4BDmdUD5+oCQfdb+N2A3XBo2L4Dgv8
axiE3jSkBqdQlavuj2CDtMxulO0iaGCm8ONxusPjngiAnQldulpIwWoyHapHKJD2jMuqy+L6ER5i
cmnDtWoe/PPn7HLFG820UvJJHgMORCiRXUEhMqEgdd7N4eTzxHItjvLopXa9rzmVon+HaJN0P/4V
eoAANpCBCWwTCm1YuKg9vD1u1prT2v/UWC1vXx9w5oIDgWxNwBQfVpTqxjOJ9JTNxUBBUrpPwRue
XfxbNeRl0aFeBORMCGBGrsUMj3JK16Qr1TfT7Fzy7Ex8bx8IfONQ+NNDegf0yPsEN7gtH1Cc5azX
Xk+6AQPsaeDT8C+agZHII20Of+hHV1C6ZM51CIyNrJDHb04Tganv7PQ+CN9i7m2F2ykGmUJni7J5
te4+wUQD2lX5dgh/uk3eq3qMgwuknV5Fd+ssqmA3tVQ3fgBz316gBGVOEcnzrXTk7hmJmROiR0kK
lUazZ9c8xOBV7jxZwYEE0Iuc3RkIQgVwr2cM13ljk7Lf0/yY0vW4XdTG+NU6uB4BIKJnVkxITplS
FoOS3rd2/pTnT8PrQan1y23M6Udc05M6SPgGUS1lqgk3H1/rPVJAOCDL1buASFbgwNA2kYEwimzB
Mct+GBNa169b8pKqx5AbuUDZHFJ4p5QlMPs3Zsnc299N/suAFTznyE8EvYeo/1v/CyzhmoIoDFNd
JMPjLVo5ZkvNB5e38EV+1Dh0JCWBjZ++OgHPZR0gv4OyoJiZy3yhqmMj92xI1rsFgGMsrP+rh/+n
MkqCkEiICqjVcSbXUnolx98+cBjQgM6gu4UXbuBOo02KRcGHc62huHEvXcnvi3Jld0keBNwvdJP8
Ps7wyL5j/PyYiCQdoxKlFMhw23CwRl5eVs7vFCPVH04Tz9zrgi43myBv7AIFOKOeUpyoH44FVRAp
46QMeN2werCT146/Z5MTU+TvFMVhZBHsBYDH2QqHlsvv6Xx6BTHHvQp+A3XssITru6lHw6VZ+T/0
4H4xWnJpXhs3+mkIjq6FKUHYluulPAdRfqSULBsvsMq3kfjL+/45h3UpN1FyJFu0cLF7wYoVqRKO
qR0A44uIGqfxzFcC3vyYeaTEdWdN7p9xcrfbjAs+DttYTX2ZkAAXNdcMyJexkiry8BXW1V/Dk3yt
CKOFMPbl7idxgRKpaW1qE6tI1jcD4cbczvu4V+PCzztjtxcF+76+bSzNjsEfExkrzo13541lq9Yo
sZTa8++wo12aEGJ8PkMbGDcLkCN/udwmNbHSocAJXd2d69j8nmffv1dZJA6s7K5iv55OrJV4DHZ1
0jOdsbfpbEr7ddMGM1ZZT4IdGJ5GOaPagS9gniF1nYJ0h4EPc38uI3nlEDdGB9QnAS1e7veoYjUL
N0pPhk5URMUyKAyWXa9Bu2u1c8pvkyH1WJyqlbpSXFErF+ade/Jk4wT6QfjhaMBbivA5ytylpPvt
AYNg5rcwvWn/WR+15xeQKEFTdw3nTT6seQz47N59YkE5Ag7m/CdsOJpbg2nhCjrOEbbI6vxhEe1y
r2b27dRoBVjrM+kailTPLzfE4u2uhK4RZgLWoxq9m01n/PKj7fXNu5iYhfrziMjecz52sTMGKoex
ej/SMULcycqXs7LWVUGCe2HFD3pkUtzZI6PLbwguNCd+l6riJDHndyUbj/vJ/MhTtDfdLv006rwU
iYhFBO5UnXHEEQ1srZvRApXiAjPXiIAj7HJb7BVHCkJlPmcRWOr2MY4KXSEhYaP7GuyZd5u568MR
JxfDGD/ohISjp5JQ8sUlqRf49vTQ0Y4IvwyPrOS1zuyzHd1gTkpQ288FhmqYdTmruWSD/1q4Ept9
PkIhVXKv9FjLL9u21fd5z5SjtOwwDJevhv401s90mA49+/7cwAAmlp6ZBzGvclySxEJYtuoa54C3
mlBpRJN+hMKSd6GLqpcuqVzdMcbx2ELDWKEKGCrOtJ0GqA1ZWvr3ol84ugmIZlsLpEdb6Ks1l472
s4Hysh4U8V3JNvyoazelBzqBQbdnSxuKCbeG+2QihuFpFo9axnsR64fGa80UdfOKJgcMMpULwbc1
kVMRhrZ4+IOb1GP0+6bKKLhnYaoNK2Bj4umjWfNf7fjQqD+ekMBiQK6YcuZiWodpP7TMHz+1AwK+
MZsWX0lgGbuec015HKKyNi0qEjS7cNiRMJivaVtegN2w87XfxcdXSRFjN0YGb/K7BuMsPDQJiKR5
fmxf6BeDLgWm6GFQZKIZCG7O+sKGoudqmxYheIy3HdLMxbJJHv3xH4t2c0T6WK1cNS6K4i388tSd
6XL6nrshn/KWsXJSflDmlT11aXR+H/sXgwGFEKWvdB26gEpXoFMn3MMyOnJJs6zZglV+qUccWN8f
fXLhdhNriJwWSW1yOGFhtRMHRjqE0i53sNLrOxIF+yU9M69f7D5XcHuDuP80+bT10UxGWBkkj15J
EBVlk2JRyfFfJDRM0YpxC0Ff/H+zpKd5qchu23Y7Vkywj3kxU0gXa99xXBmLtmlH8n5Esx09IR3H
SPV9sZuUXrw1lmc4FJl3NkHwV+aXiD7xFBFwowKGQLeh8luidqGGewtgLKJoxQ1ZAuh7iJi5abkI
Gd7qcyCZ6n17n2TnEkEepArBEE7Th3VCOlJcOgLPVjedb1hLb2NgwnGlicUZh5OsYt0mxFNqcOI+
/vSa1rkzjvZ+pqy1jF1fPtJfL++mJd8iEyfj43pjdIjjCg9iyP/9ww/cGytlZ/AvHdkjh/c/V7my
ezCTm9OXOmmsUQBTgDnQKTmWc9jPTyYeiznr4MeIsT0i31VnMlQY+uL3+l+xN2kJR2ocLSE1P3ba
SlIWs+E/SOYpdnqWVGxQdrBBloSfwFkLDz8Uj60edTU8WadOlKJxVzeyiwgQPjwyjwQ9ZvgoyNo4
eDr5JwZE1Cb16xPcLH8HvxkoC+SDrNvlZfMaR0+POwY7EfSGAni7IsXYD9Zw8eb/phXhp4gb1BsB
RF7ZY1FXZ/odwMhWo74J/5LvIzMHxUQg0Rvr4XEktNpVtCfz11vZa3P89e1saEIey3d2szHASgLz
tFhp3slDc2VOwl+pOzirh4f6Wwj2wejhdgLGeXtmFYbpMpnwg7FbmuPz92RClg3SC5ck5rcMKVPb
0PepHMvP/YDeQvJOIzkhWgmVgqMBsKoidt4pCfZojRhjXhUG4hSXWcSsaAwn5G2Z9wgskKFOCTrh
HeThgibklEki+7gx4IoOGosLMzGaS8xyOkx86ZKPMeoPSYI4saWYR7u0BENdyV6OzifJu+HBuJjM
ZT0JlqDMM+YogCmstusVF27xyJKYSRLpZr8xj7EUQctBtvkxOKCtGnD4LTjb0qxICYYmwlx25etw
fEvDk3qWbg920wqwrVh5TzE4ZcQF/JNRdDXszjZ4HUViKIDgwUjahEKCxRu7drluumRmxBlaY3/q
EcSda5nUTTSzluMSfvAskMWq7kQaP4gigMy9DR76lT1Ejy/K/jcOoDeRoZ8g1pX0dDy5XKSzvKvW
QFzU7gk4SQnZWsN1sbZy8jZkp4EPmz6bVF2pQ4vatBipKgQGiJcYPRg7nolZpAEet0o5tOrT4YbT
7zUaN07SarCVT39d7sInpZjgA1uxZ9Q4tM1iyBslBDh7UXxPNhUrPPntLHVNy+bRO6K4typnSQiI
tBRyYvJ8dflzBxAfHgV3/C31cvQ1jFB2RkqcEuTjB/Ukyv74ZHI1NSsKVXekzxFE+iDNxFble7Xb
DFtcrD3449ybxf4Y0pg+UwPxuu9EhmhR3BMQlNviEgFle+uErm4sdQBktkO8iETJzYZKB1m4AATO
+EkwhpyWpXbLOOabU9CVNAhNG9q9YADYh1W1io9mW6ehhP78nwLZIwSrk2ZWz/96sYpdRSsKmxLE
f3bm5mopVSMbUukxt895VQ0draRTmP/b94CheA0pBMDeKGCFDLyNH1XigANQAZmyI18eztmuyzKY
qNe/ty3wvRQlbpn2O2DYRmqhhPyA8Zdr9bCHwDmDNEKh9uY5i9oSQbg0CGIPT0s37p5vOREQqE3p
lDWf48cXo3sAw/mG4RnETasrKyQZdQcOLsEH9EbSn0QneBWXPiNICiNWxa2ozvAm5LEFTLc3e+Vn
1vZwTZoveY/KJCCvIrexfhjeF7nmjM+l4nISo4jo2NSlUfMqrrjb+v/Kf0BkFxsligpIQaSeG8ry
cRgUI5AbHPzIuGTdXnjKFRVw7Wlz7lSOE+Bno5tQow7k1XIFXQM5xwDbuRaeXT6j/uMqSGmOTmSJ
sfUXEfhLdwh4znuwsbZ5VSFbopeT3tz+4F9gJfZtVMxPvZtRweHNK+fWkOVPaMAK3LWaVfvxO116
KY7pMKHi+/Xog94db6H1Gaf7Mw3mx+6ob5V5AaMdQu6LMm3TzepEVlhNvSBCbkEfT7kKOsXiR2GB
5GcCmK0Vd3LREgKiXEZ4GANKL/AVlo9MsTZqrCiorU6/sffkq0cx1c4s/g6HEz/EJHOkXHAxh2F7
Kr/+3p3mohOaV762lk0voEmUEOfE04v/sNdRc3GaO2kO0x05BLw5p1vsCncMoseRIjNuXwio4F31
gKlatLD2G3o2Odza1tiDXunuY0i+BVsbPwodZ9WPWUMk/4UKIcNUk2BkEiht5cz4OgBzT6p2a1Wd
dtwf8Pxz8H87BuHvpW83ZsEl3vyc4duruNlH/6Uw230pu9lumuXHlQBSLTyreKAHi6jbo7tc7C95
VFs32ILBWJTw9H28K043ZTrOeBNdfyzYgeUQl0R9CF8KgBdBSaEJV/DNMJn2QxzFuraZlowjIMMP
Yjlsf8PmasFGq9c6r1v/D3dtS++d4hXAGrmzPWrGu6xiGjMEL/WqALSrjFXCZVGrTe8qRfrKJJi4
tI0B0D9GYdgunppM68J88U9q1vFiIcyDUQRRst5ueSzNLM1DEpZr2J13IJ6qyI15FoDt5GmnOqVG
Ch9vnNcNUVkdEAI3QcfiEEhIe+PxlD3C9I/DNlubAWwdO5WuuJab4HCGaU7hegPJBZJuW828s3BC
PLyp1W9YUMrEj6KrCK8I5dGPeALurm0717JKVsqsqBSJBgNXBU5xRE8RC/sNetbrxgaDmTaW3YHA
po9aw/7kymT+FSm6DfN9HSFO6X5rVtjcg0cfWYe/pVi4usa5ETWSdoWNoKEg8OGdC8wHJ1K9ztVn
3d1uXdrPcgMejwlagMutNJ5IKiyeggGmTO7M9X96mi+WABLEK0c2QmQc7oyWmLx2047zlBJ44uFI
xzv5OH8XgbRF3xs/qYp138eI/fLCnBx03KHlk4lFPD6X5ZBmEyFOL9pbHqPhRA9QeYkN1ahVGoyD
HmtHlkptDmTXPH4IAFTYuv/XQuhbbualXhf/tA0NuxQLh2uxHh8JVZmD9S72c6ctGGH1sDiIhS9x
bDrHN29O/tZX6/wqMzN81nIF1OiQNS3u8D28Y0jkHr9xSfr1PFG7AHmFUjtScTJNmVjlA1sz6mER
Etn/HQD/Tu+U8kE1V7PStzFDAN39vfTFCDvkKxK0gwF0tqRK/kL6tq/30x+ng4BqX/xArrwvf7qv
yWKD17bWGE2eqtKqTR5aBgKLCnFsWG0T1M09RD49OQdeYsammXuOygH0Lkfh9JCbq1RqquI5ra5d
/tpORfH/XYs/+gJXhQOXWhRO/VZZ58wYTPUQpzdvOqiUyKJtMKyo2+aP9yrj5TXE8ASFqx0P34La
LRGV631x4RlwBtGlHA/yIL+YO4ur1d29Gf7oBqVkqnnUBi7hYdhGtzDyPJON1sOUQUH5Mo8uP4aq
HbN48KlQtUzkft+0yYrX/+oHEfLGsqrXLmy0XlHyWucWOdOaLK/oesEpksxOLaZnRmYuuvyRiKKu
oBO3MnlMPglPIqzenfK+ZjrnUSH1LW5xyV0qJuvyA7sfWrmWtCivY1XtPDdUYFqFCHrRQcpF4o8A
VlaWdRghZJlv3H0Orw/dc4HLw3qb+LD28klFNdCY5tAyFfXtL3zZhYhHzItB9kqAuuxwP3rD7Bdg
UmvIxK5xOEWzkdM5o0m/k7latkfvZSW+aGShF3hoU0og44e0G7ImgreTMDCXeRm4Xe8Nn7ahDbgB
lyrhcrcwxkocVjZhmp/vytFx2joLIcjBpubcdrGmxESMQnmBcNri2cqEVnjMLOUfatNwNWamdG09
IUMg+ICHrLq32LwwV6lwVdiNQAJMO0BLeDQmeNZjFanp/lVrSgwTCgFs58NV72B4dN8hVgiQTnov
E8obag2M9vWJeR8C6Ig08zdva0BeLVC5pW7rETTmwwavnnz8NMaH/Ul/TG6Gxcsqv2sOiM51XoRs
xO8Jd1sh+LL4BlpTGVehNgRAmmp3ilehSSBsSvs+RKsW5NXNkdSLfARkjmQdpnQObRvqbjxUZp4q
kqxwbC9bEE1mzmFZ/23A9rUG2vtsuUlN7pdgHOcn6QprkZICdnuqn89OAGzKzn+H6S407PAY6jHc
WeUVM8KoRaXSpJ19shmRzUyx9r0BQIyTBlGE3fRQzqIPR/Wh5O12nxSyxxQ1rbEQj3DzrthvsMrw
P9kvrwBeZtwV2msid09Fr0WAy5nn5bfQkALlqYrlG4aW9a3Xo4jQynAlTtoqKkuQLSujbFOgqI2k
QDFcHrMAhwuICKl7CoF8CxZ+1mSK/QDSxrtBpgP5Dr+bATVlav+YC9xqIPZ9G+q0Q87+1GwTvbJg
zHXntUXnZcfpG/RQzZvLCYhHBdCsgNEeX/7TWCQa1dN1OHy7hFX7LgDleY/ttYhSmGlfmF2/kZ93
i+mfeLN/h6sfayji13OOHc2+thCRmMuyA05h0rdUHq3CkYttMTWE9F4s+hSCNCu+Kp/qXB8TQ1Q0
ER4+psNqsApvCjpL3A27GGKyUNjdKYuPv/5pSZRir5rHT1HuVvtkusiDSlyJsdnvqInw1BgWTwuE
j2Bn7IBFPkWhkPBBHogRwl1OOUqyO7yAt87KEa5JkMY0gUNgeZPzUqeH1HECnWBW1w0XcVZRV2yv
g3TgN7ajVVbJPM/54NRGdozZCAhetksNHI/eQn2Y0Ny2jCPcM0fQOioO8dqGQTsIO7sCsxFgmDP7
SnrOiYykdbi+Nm3V7yTgO59mM3TJgpfntxUgIHhH9PrFmmslEe6ascyuBdPZKoPhKed9UL0S0PSc
oIYqYw2DCqqtGXAHiSvo9MLRJLr50sS/kcoIHZ9QglCjgHGRVRqfFpy41Mer+llsPn41rXdM+PMj
iB3vOxJc7asZ+5AW7WHa3eBgnO2tKYb4DGxJ23+5jPa8mdRs6LBX+h+Y/i0mVRW/fQ7xjvGNdpdq
QeaNoIvTXBj5DWWOiUlGnnqZZP6kcls66lineYSAvTYWEpgtbRFB9eqAqoqQqz8+DSHzLEJ1XiAT
z6kmN6kgangfR/KPxOjh7/jKtR+ikkWBZU9Hl3Kou33akK+ZOlvU2h4+J4cKjSnGxPwjI/XnoIFV
nh12bjUPaK/OQ6eRcQwKek5Q5dSohUy89FXEVWWODyDnsKW+6YBm38t6sa9BhbTyUpgQpPTPNxXx
EZtBjn+F7Vi/vRZayM6Jukf6P9X9sIN/dnLdz+12hrBV3Xt5Z2UXnu9/lAi3+ElNUV9HHa+kKrF7
nxApyTK2b4Ey6GE2tp9VgoOQTqoXuk2CsuRoHYCSXhO/CQcl1poNjlWVTDpos696UoYSj5W+2SYr
QEmMzknkWtsHSzkV1gSG1eSOENb5e65l6frDmfoPMGmODwJrgO9NqU3B2C3OVV/MQAWCjs4k97vz
vwQ908FrMhWXPs5quABNLb6wpJI77/AgzbPJOc3EM2iKg5Fixcs8G5iEDKw4t5igGh4hP6gkfoqo
TNmitDOEHqNh7zHi/jkUtKDIdmN8HgbmCvVC4eSaSqqPdrLECtomzSh4R00nF2ktP08oR6sX/7mx
fPq5e2wkcB+/b6ietQOweqPFEnYhpNK3S5Mi7PKDu9jXEpA/zFFUGCwfRK+fjmxHtxHeVlwkXUgn
nqUh0UiyRTGHZBidAVuodrLvJj4+qCHaoDZNB2Lyvc8ACGTsAJAuvYIVuKTl+3fvrLVcEfIHhBgg
9bZxmStHMa6cPItI7GPrh+OwDDZHaFkYPBNX97Bkkf8pkzEEIEbryLmeP5Hf+bbu/6gWE4K+s0xs
EMHnyCcjfGYYp30VSha1RkoFr6DjaSiwzb3TtZEHmSLjc2Qy2/lrUBhhRT+8H9y9TQs/KhKx3gq4
H7H/xpYR5lgpOLBnpAfS0U0Az5ryQ6StHO0i44D7e/2WeFrsCm3+GDqljJ1EJ1fyFNLwnV16ksYJ
FxJjuFaJtT0eYJeA+WrdMSNlaQSAyUSA1mOid12UR5a1iUPJQgbALeE0gfXyU1nOPBHTzX8igMfE
F7Z7PNxUjINI5kX4rTpYOlkXPJueBLAaKZ0ude1Fssikn8Ed/2xwAO6+9BkHB1Df7+ono6BN/usG
Swq5uAnBaKlQMWwA9AMMEKkEiBbJwS5DLDXA436nVygVEu6sjU8yrbd4eE1x8woub3xaZVcpieDe
FXndwVtIqt13UsZnKeqQ5oaa6qrUg72Wd0yJHVT87hc1VzIkILY98kZN5v7GhtRz97XDvfozkYgq
X9hDUmlVwy1Pz0Un/t1Z/FBMYmWXWTAqX2RcUrJLBB6rNSQ+B+iZffG0ex1zoUv5rJcFpc/WTfF3
4QSdxrB/F4X1Wy7UVrBckpHJLkDJgI+BA+bsxBRnbeE6iUnOphKhc7zHBOpjlHff/tg6nC+OSRvT
GLbNEA8rOj7OVe+XOunhAnzUdcbZGrsZbnPG3/YVnn6UbtRBzZ/ffEnyxDnI/Sg/h94vmASVcBkT
GiJZU0Ca/9J5krvgNrLlxErpZMT01sFKjigcPSj4TE9Tcag127inTFw+aMGqcpCLsFF/3TSavoSV
Rl4R7hdsSExhzRyky4T9fQrFHI1UHUFCIzwCNhs88wKvfxeH6uFNCxIrN7CvC6XB8Ng04Qw6XAph
blqso8ziLHR6tySSq92o4kOYB3fY5444pPFO/7PwxCRBTaaS+WJVwuDS+1aJo+FD1Uc0jYl5htNa
iBP0in+O1KmWyRzjwrUmqern6HS4nJ8yR7GETOuUuWbegENE31AMhYDScq/noJOHE0/5Ap0mtCME
YkW016kPO+sRlDsZJT8a+ltsSMcsHvcuHZbD9Fkw3T/tFWM+Uz0Ah4mv+CSDavvwf2qD9FuKU6dO
JNBMoRpLePWY/5ANj4COwvHW2X6NygF+bmEtr0iPg5xrPXa6TyOVqTeS/si0xdlmH/5Ik9EYJRAZ
+aecoOlK4mpDOWOBpNp5Bh7SPE1TsA575159ctVdulSajnE1PX/i6kLgx5/TWjL92zIxgqNLISPk
uD/61u00cGm+PMowqsPhhYm62Rxt5v5nBF9AEpqmT6QsR+BasVq8tQ4cUHhU0yDp0bLdLnekmQpy
jaFtEMhbq4r8BRlxqvGhD8A05SyO1CDPT2yDZquyOfN6CtYCE1Zjp7SmSqHIF4d72C29XbU+Ip42
aaSFSidh+Fr+4Q3jHfSQ7eFWDgCsx0aRHsbxJOzAX7ugatR/bXxas62GntdCNgnTncL7mbf0QEYs
PL5sIGisQSLYN7q5MxCBFgYvgS/yBoAMNikiq3dDl6uYVFhr8q6KAhH/7mmNDwIf4wk+pLd7WtQ+
KKlm3UPabrPmFhssJUA8ljmhwA11vIY/5W4I0YHkAb//2UYZYcJQ56KpIozonOR78Y6cEQkVVEM0
u5yKr3pCJBX3XTYaXdN3Qme33FzIPgoLfjwAbhjAMEv0UqyV3BC5DPT8MHbK/+wfJny5sxUC4ln0
muM8MZ4LWSlPXoDNkcHY+VF8PfyAD/M053T6xqkqqIpIPSXJXrT19Nj6yaAQm+BodApuZJpZnzer
dt2yM9jKIZjL+yqeEhX6FZTGL3GppYvIWfuehE61xAjP9BFa0RueedtuwqfGtMbfvJI9GxjacpxX
hTaLu1OGzGzVRy96m8RJ7xPA8a7mAtOKoGnnCY5hG8f5iXCgUxJjX3CmbSVXk35GcWnDiyhLsXsN
coPI9g51JBdq8v1bEP/sQUihFqUY0KTRHeOYZDp6ATpZXg5k3h9IQ6WtXrnJEAAWkuXUIyYAXrlb
n0n4Tu0jlS8X1v6BC4aTImUkWF0VCtmv9Rem1sTO+ofYlAdbefmxUfPguOarGrRfzK20eME63YRV
3Yv95ABBb9+SLbe8pxSm6NL0Yz9/ab/q+JeMeugl2hBt0ByX5fAZifms3MKMEULcvFlKsyhV3isH
oC3ofGqphFaeTO9Yfr/mTW11/Nh9dOvCQSn3YiX9dU++Ld5c0qk/NXrufjuunkix7Hffwp+sELx9
SGPLGV8JqDeVsr4w7HgYwBMHuzv9klIKd2yW2pEISmVJ+7saCzLTgIU1eWkTrXD+cXJ5dHfFGpqQ
CsAWIaI4CKRL1TPzAldC4yHVn9Y16TLiaJ/vs1/IQtdxmGUNMgCtZs1/g1w8nbfr9eonTNLwTGU1
iBl2gMRGgl2yaVLuF6cg0bJmYDCpfp/uCLvE+uV9rWAYEJE6PJSqvKws5BMpypHxPLNg+BpFvSI6
gN2X1GxsNRwtDAhtbXwOlKFcnVCXEm0o9z3PZk7nREEheMW3E8u8pO9KnAcRfwmD3gxlBA2KKEwV
N5TDFR+x4mESNG1QrLjZ5C62bu361m27CZCUoJPezOv7dZ2XlO15ZoOUrEhKYQGfX3Z5t9DGVfOs
g8zI4adopSshayiPbHedTIlns/At40YQaaDQuncHt2iFLGjMiM2cbT79w786poNHXXAikCxpdf1K
wZkhdcaAq7fLAR7pVODA7mDYaIGo6vaO5ABOW0NiVLHjn1Y63eQ5Gy9UqLRsMCcVgiejrt9GLn5t
Lt4C9y0l4QspJxyjs/h/ugVNMOIC1/oAlJrjlSQxa3H89D/oklEhW/nVdAFk/vsh7EOai+WyaL/8
aqylKTt1fx0mHoP8CtOn9TqlTlq74ZxQx3mY48GZc/FtBtXfoPIYSIZaeBghtMHvT4rX0fot7OIO
mzZGwUj7cANUyDre9H7HNFA/TCWs5nNGa0YwwW3vQwrhrZd8c6yEBM5fcpP9T7GGtnv4Bf4pE7sG
RyjUBg/hqRN8uFZCqnjFsnn9RfOhzjvZ2XE+CxoUalGtvUBRgvCR59Y/Lkxaeo02CNEnEM/o20IA
2QnB5zgUBYr6S+z+X5cima6KS7y0sHA+JCbliIfGJIvRO3gsTf/xqEE6nzsCwv/qLuOC72ZsFlC/
SUoMxVt24PCAgpjXPDvEeo8XdX+PlCYu41imDOWltUqP2kT8cu3P0AzxolhM8ah+VbsmaGsFcKL7
+BZ6LYGN2OkiphW0qWk5WxCc1RsrHvi+ZZ1y3Mt19GWgWOl6TYBhPmsiDq9vrcdDcS0QagrSJZVm
UWtxF8HfD6psFI4X9Ztx8N2CA79HE8GRa8u9nsDFEQ7z1As5EoOeRxbJwcM3PkWArS+lTolBaIuk
wVdi3g9pKaCH+ciJnO20slCH50roDHimKjAdcWQV/nXyyiUQPC1j+VVSYfR/Vje2Dp3Vr+jUgk4b
M6olkqhZR5vZYdM3dJSJ6qHzUSM757UYrQIzevA7FRmR8o0dtKxF5tOgAj1/DFsS5zTzoS+/EgI/
/q6Pz3NLbY7LOg6oFawiSfz8o3CoZ2o3P+PxunDN+2Fa8kn6tYTzQNW/Jmk2DSTp9fBFLWFpiThB
k5W0MorxmNtFQYLe+ZGWn1WhCHgy7Sa5HZ8c1qRQmCJp+ivNFS3ocVmBTCg86WRn0z/i0vSI5EAi
RXk4pSkwuxDwVCCNAmFSuPPxFJ4tE7WKQNn9VpmZU4uoEbjOU9rneJ+NcLhixB/Z3750ThMo1JRq
UlbjPKpOYnexyhR6mTOM+RACog2lQtQKtH00TjfgO9EDAuOzahgIpWCA6qoks5aCBEDYbTkkLB4w
98wqsB9e0NB94xdAJro4MQRzQ2VPLhsHTMRGsBlcZsN3VpLkUrGUrcQcqx8Qh896iXrHCbuplNUB
xVt+uk3yJFBHKQWdI/uQvEiDMQmP00qNO5cDhqsGCEIfUC0ftGGBWMwDqhcTIJss2JWvGhdEF7I2
ekwWPDnlJRk4U2JW4aVyeKcn0ZL1VWSpZha3kpvnbkO/S/53nR29bGLjgIJIVfl+b3iLgwJh8L36
+Su9uPpFaT9dbPxzKRxlBuQiKct7GZFKOut4IkeA5P4WM2S4KYUBfWqwnIPxJ0sW2eVHVFw5CRCH
Ni/PGHVqXhmVqrVJmbkZ6jYR2TN/P02u/A0EAVzZF1iVgsmbBNlzSLhLNciKrSl1c9W4GGwGw5lM
xMMVuC8j+zhbxiMopmeuGdHWLA1wa1gMUl4OPnywBGgUxk8ULpXNerxbPNBKgu8WL5Z6CVo8vSfU
cRttPkKOCCJCk9yTvBdg+KThr/DYV6B9Hlsl/nowvIanJoYJwltTBHlhQe/qWP1FHmrXfF9xMtkJ
aX4rQZUE5AmUZUutK+KCApOoeTBhgvXHoVQAoxLqnCcLQQI5BOAYG0qZ4IoHZCH6D+8MxziRTBqH
u1rU8MULV0QnYiYCHotFeRy7OkOhzOLjiP9skN7n+SYAh9FMqelX9uU9TFgaheO1XKxx2a5gYC+v
w5X0gUS16R/h63rMv8eXH+ry/G53ixjl6z2+vcNmNTSoqxVrnF74z9w78ETEKTcw889EsKqtCAsJ
XUGcRH1vciehb9p+TFLSqFjXZraUMWRzlytBHTakprSB2YeOY5kk2S6x8rMyg93dc7cpX7RU/yrg
naU10cx5Hayjv0b8ljnpyEtQ30qFd/ORwC8grUufVSsBqx/PINDwzO1N26GZqDU48Y28sl3BpszZ
BT/jjM6QL4ip9/jJfl8CuTmLx02Z/iQ3wha7n4hqUpkZ9XZQZ9ZFhCWu9qN0/hOXjuapmhNrd9bg
wPcoZputZRS9RCaXv+ZjXI3VpIpbTBPu17vnRWF+ASWrW+PCDGgVmky+Djaa8+AaBXn8NLITjHyB
ryM2N1qOtCrOzN/lQjhsx92gidWXXSv5NxC16VSVPnRMak2qkHAuy9Oe0ITIylYwddLEZ9zFHx2w
5T83CaAGWicog32xt96mEb60AK248IITutQWlRbFAqF5r5OMxJo891/Fg5mic4j8mATIHu5WlBUm
r94sdNzeOKHD8pTOdyxAQd2LzzmupDKwDjtFXEoq+DqiCc1vuaD0dKXqBXRLtRy7rN+T7jVrfMrC
SLr09/9FaGKyySI7/Y2giQLYOTD6JZJLJHY/d9aaw7oPbSRLt/Us71oBFdFVgjyvzSJoz8TDVGMj
l17c7CzZ4cJcPDHW01naIqZT1/duNNIXtwrI/wZHQ5l3SdGTSJBmk012jH/gxGZ67Kbu8JXfJ5jr
opiRxQY2E1fxkhrrELUuI9aPE5n4U/b+dFbcgOV/C8yjq+8t6vKHCLysBA1ZCg1y6Snt81Evkf1a
AY9GivpdXujagF4k9vkP9Xf4d/LeX2TRvSL92hRfV5va8U5lQvn4LHFabqCZIX3LTlOQn0/MmwkA
Uv6GyZ1Yi48QY3Y+HoZ+j7NnbmzuzqKldvvpSvN8yxZk7I0QmUIj+o/0XGxajcj6A+dzf+SvLGdQ
YXjrI3i23sdHapAquqJX5Y9vYL26HonwEQ2CWnYRsYNnwl2Qd1jaW9arNbnYLP3VDOjYneBvcZwO
VsK2ASQwbTway0qMxujwL8G+3FiqExM+JNLe7NZcFGWOEoWZ0WIDicdOkDmbW0mx4mfvR++krblX
yQ2meRLajl5s6qGHqGO37UDs1jMZGntRhZkYyVy4Lo+xdINQSR+1P+DIbzindXvwPHNOpOemomqa
5ESyrKJ0GHlioAmRb0rFVF1pgCFk0QooHQ4Q4NQ8M/YjM4ZPMdoRhHswcT2AvLcdDA4in7zXfgWQ
PeSC5VheOcLucPLJnza+7cKFrcSaul1NtvtrVsi4cx+GOE2Fm/BBx7wGkmw6MX/8wvKkrbl83Co4
Ry7jw2gRT+F5cTJ5wmry5jFf3PUXwJNzQ9e4smaI/0cvipLWLbd4bPkmq3tFyEJX9mL+1dsKPPJg
28yGdNmX8iKp4rQwhnZUckfwyD+M75fLwjiRjCiXIQX6DVfDbKyKRGFf150phBSgYAVQKo0wn1Ps
c4H3FKTOejxxXJQVz/dIJyveYvwkNdgDMMWKv8d2zLiZytNwBT+3s4YCFiha530LfcHnpojUkDRf
NkCbHLKOO1v18rCRQHYdiniBhzElaNZJaWRSPMRtRWsJcgdvtD297qiPvxl+lBYyQCBaXw1e6erS
8YIl3nbaLnE9Gmz0MZ4P7cpNsFQcMPTviBIZ+4LaubFEGs8vYQCNvVYW2kVwb1MopsDsSZfkFgSg
lyoVIke+/Ij969OrqwVgoob1ySQpp4ObI0gI0VVyvhIJm6JsLgcP82uL3ScTzo95VcZnPowHN5yt
0AlDuekYEKcuzJikyVOmnOfYsJSTjPj14fOgE7M4vkf7YLJTXb2EV5Y2o4ZVNMBQ7bJhn1KMucCi
j6AFswwlEk0fo15vYGGJDmiuIvWLTA/ppHcA7a1WwfecxQG0Qwv5cxAUYHOELbT+xi5RyyN1Uga4
dKVYhZmuqQGQ7ph5MVaYv7uu5kLQHumhIbf5rh+wTlFquC7Qch51pWCFMrlBmlwYbw1uJi3OTihB
y8RyWFHbhsL7FQU4xbsectNop/pw8qMuECu9kemDlyGK4/MUIofoL9yuhF9CMx5+NUw77v/wuNC5
4rlG5mM/OwTdc3YBtyfkXOKi9oJLv7tTJ9NIzJXw/vWI/xuR7UhObhuopwiZ/8rdWuYsaTv8ZlWV
jt8Yk2idWXSteh89oHocWHaqOYv9JItmqSYicIlQyJ18Wb5Ndr8YehB/p3QnMQrU9uIEnNH8ncN/
y6p2FoMM1hmr6VyLKTO57HSfCMYlDnrzeg65J1brQRJ+PG11skKFlJmZ6Gg/nFp4qYdIFjlOANxK
VyitQzu9QptCeArgEOJZYSv2LUx8sCOMxwhvladO1LiUlkz52T7bRvqYVNoTT9nLv/AcU0GnTDWZ
DjOwPrv7oNVQJ0xm+qlO/OjQE3uu0NuKW5CHg/iS8Aa9eLHgIbqtSHOy01PZm3n59mg8iPCXYrEW
KLmhJK5i8PIjaXVnzjT3al3ycb+D4mq+9q7HwCul/miHLl84I5ZmVmofYwkCBqxXivUp+wOF6U2K
wAZTjS2NxcXbWqAVzn+yxOnoRjFffaTOJp0qpTnt8UGsJRiZLEP/q+w4Na5NUKGm7pBCFw+f1eVl
pCDhWrRpTb9mHRjJUOtmntGJydaayO0SufBlAlCnUs6b8FdLIwgPqyq1Vq7/0jSYZcQWesSRIl+v
/4RWk+VKcyvilke093fyZJJ1lP6XiMfRLR/LwAxxUVTEqoZJFc2i+BIru7pBXFSIhzCD4CoCZLyu
/1qfVLZ5YEsex5jIDFce/IE5Kh/t1iWmuY+jZrXHNhqlgNv5qc5fETZgUhPs7du/DNovMQanwhza
C+io16KWfYTXJgzH4gzMGjAWkp/wZ9+CmCRgTyVYteS/8mYKs/772aft7Y+pgEzhJT/0Qk93iOQq
MLuEH5A+abjPjajlESma3wgDjA6WLeOL5Jhf8F9VXao20q8bzmtMWZSshAA33wsXG53Ci11XWHMw
w8qyJN3p1y2khnGFbS1X0gVzXf8EII/gwD2iu2prlpVXmp2a85ZTjZloH7h8UYRIRI41SignecxQ
vnA6Lx2BQ5LJbEQv5IcylZHKtF1pUyBE/jx4BU8MumZkhW8TekUzl5FNi+ikNWn2t76W0YbqcRS+
2jtsfoc7/rTjOc11zzKkY34sGZKSvUtGv77eix4DIRy8NflB05avqeq0/bSHg85Hwue8rXv1dJ71
qgWdwjKGbJAB2/vWr7STq2Y4lbT9jA9crnwaEQ7ReSb/cgr1r45vyxSfxl2snooTZdvN6KEKmRXm
+Xx5lXYTWhpqQLm0suoRDsZNVfPcK4kyqPoak7z4+vuGGuIsSr2CA5k9AITac128Vu66rfDLRRqB
YsHc7Bvmez8fBvVF+fv6Ub/vhcNk1VfqmD6wgBafDyqfGEw2AR1JdvK/QrW8oWERRSipn6Kp+HGH
D02Ji6quEdD/i+7a3/1fnI/QbyXYMxa3a4QvNKervs45YS81qFbJfx/DqjXJtGqirr/dbRrJJfEU
ZQsYBdoD36SocbiHij6WtOqPe3ZvIjGuW2m8pzYWyRk4O3pQ6RlnA1QTbChiXfpXRY+fj4ra8LdQ
aFIxd+SuMD2JP08oMWFwVmmv+bxDnxZFKPhEvGdtptfs1nPxZ0fCmkTfjLhV/J/nE7rqKoJUYJfK
qq9Ibqhw+Ar/S0UW7stw787Ti7FdvUC+Zzw4O1w+mLvmV1wiR2VpUj8vlp7dFWbq8sPNthcQxRjc
oNu+SgIGRfX1bfY2UDNFIAnBrR+ZgIILLt4iPvTgvR/w7dD7rxO9Wf8uZLjKaMfSyPGxWnt7amhk
6Vhf77T3z6hpMoaln1x3VZBrtwuQrNu9Z6kUaKZrF+zv63n+BDITzaYrmzr4rPFnMUMEQILfehhl
9cDgmaGYpHiN8A8BUJySQknO1GNb0dmtfgnvLahuaQ3wFEC1Al8bx21R/JR9ACn9Fu/Lh7Nt3Xup
4+qNCbNGo8q99mBKEjz7SnXoX95l2qfMNzwLNhdPHicIucswpQHAoNcL5ks5NhQ0rY/rYofonJdY
pJbvG3IexhudlRBtk04VZpRFjqLWfz0mXA9/xr7YzPG07ivHhypaOJh47mnXCxBGlR5TYTRXG1jK
6ByR2jCgJyVyBaDKkV3vhhViOxs0e3yHmg4JsZqG5jLO3zQg96GiUY/gOOoqfayMDmyGK1q6idGj
SQKaJ73QEm2qes8jtaZ71eYlBhyHO8xrKYF5Sg2N1QsHbQbAUdwhBvrmbC7nhaHdOJUFsZnINuxf
9X1yphr+Wx8OUCI904QPSX4e3NdBCRPam0iPd1w3455HrFf67S4WQL5dah7tqe/VYEwT+MvtGNRw
jIAybnq/xz8KJ/70+4GzVju2pS2CigFZGa+JgKc0Z4rG4Nwiy9i4NQnOfa/3jLVxLBz1Bh0/WvAF
SrOU8j/jD0+LoDB4+C4ODerFR2GjdIhaseUMkNzrxXTs7ySQTyeNLTJJ/WiepKO8R6hrnYaNRvSs
c4w7cdaU9zOodewUH/YRbaZgDDiTnQUsXdpJOtCtu5p/AO+x5CSDT/3ELNFW5jObWowW5dVYfLiq
LXXVMWQsNtSUxbI/k+rN4o3QvLDU/NaqixelXLw45SK80FAObXD1jccTVKH7mY4pMn1G3ic2FSil
a1bToJRooZB3R+jMcQpnIxv4ODIOrS6FOzkIBkJeC371XkP+Ho3fDLFbtpu3BEEJ3QOCzQa039ei
DmLQyKMv4PslrKcjfuGsXI5VZ8wxg51DnyuNPrQghY1bPxm/X/fJuwGOV/rWNRRF2zIeNt39IAk5
tlrG+l6Itu/pGpgZ50ZlsA2aoq7yC2vd3NSDeeoMXtzTreYi1f7H4GadSuNxdkdBYTSVDeucqlqZ
NLTSD6UJ7p8hD2hmPKeO5NlVsJQVRhJZpEbtd5rqPpLUBvFvFawtLv2nSx/Om38fbwnBuqlU0G+R
1fJibGhufZF/vZuMi8h29BHOQCTqgdTWF8Rzp6zBQKS869Zc2ZNHfMPuk4X0Kz2E7OtI1souHEFe
trYOzTBboNV/mkF6ERTuc169RfMb7D4stcqc9UJTJ5xKARFsVkfCpz2H/dl8GcWYUusQbZm0OlMU
JheM7HbBrWV6J/LAJ1PO5N6x6m+2bTE9XhY2VyRCnRRLsDWmnmRUesLVw1rCWXBjr9q7+HE4PEye
E+Eyr8Y5b0axTy1A1aqVmxUnpi1U7eQvI6dX4o8OrtBgl4X0dj9C86YPfjJFfz1LMaUsAB+X3cc4
WOj3mGhQlZ2Gs4oV+cuv2vlemsDmDU8cUDlLvSJeNc/FuuSpp4E9dMaQ/YPsDd7zqYaj9Bqr7Mcp
VAdvWUC9Kg/sE+m4HC2+ABbrxNleMB6d46AwViXmnnW++IJPS4siAVFkT2uXbxR6BWKeV3wyVBf3
CTotDzhPHtTONN5BLlcm4rQPvzYqLjIsOb8+jwYIIPyGG3Zrs9qZMLt+gaj34OnPkHEiQt7htWB0
nqxJ+26TP5BXS6kpj4GhdGqFclSgMtLsIosqhHDJhWf4wHEu9nWBoqWW2qw2+bMXn5xpw+LO9eM2
9jULXU5V92aYcuQafXj+SxAUuwLw2ZKWk42INaZFcpXaFMK0a4PX17uzGNSasRUHDRH7p0CWFxAd
4fj4eIV3YFrx7WJe9N8rx7KtehkaggjOiFCr1uiEG69DQHOy9uB7Nr3NjLc8BKgKEUrACwkYT5Z+
1Y+07CHdG18rHHswGcdU9tYn7R3kmR2D/EbZFTQLyRvojRaA6FJqWSEg+kjz+8CEJsczNxKWhxoL
peIqG08XcwgMB7wj+PKdYsVjCEchmaos1TaYQwbBOowjMssYDtxgMafkN9LGBIXY/PN9MjmmJFcE
K9+H6xnVnKj2yxYoYDWbbXIJtU1ugZ5DYjNb6vpHL9uzcqL4L/W7b+bfZ6NnQiDtQYHj+a7dy/cF
8inXoV5A47W958hfeYBCM05ytVUt0oDFyIL2X8S9dRihfJCG0tJZ2v0JEAfjSX/coQTR6/WwMgRo
YYZqli46O8laPitDKc49bN8OA5m28FekgVdsmBneYZJDAI4X7jGAQEpgqvWleGsKwcg2oevJh7nP
wx/2TWIek2a2iT5/3TI47TJzl6B9ZFvjoaHl+rlyTdDbHzUmI5uXxfLopDgMG1KjK+reYxsAT+OH
sOKyObkzWnu4eFB0t1WUB8oZLc/Yp5QEQbGtoV7reK7h6x1HFuV/q8l5PteA8VNVuJ8AzMiWYwii
5OZ1CicglDZLyOGQ4xuUFjXn/zbnEUCO0hCVhpemKVO7KD0jpIhS+IFBZa9rurORWqOWyVHAK6PJ
wJMbZW1punzfLP33N89JVGTM9P6vAyETXlSFZ8KrjKeTVQEFpqPyyG1VnpbRRXXFwMrN/zYc3gtn
EDF78bhYu/JevKDDmWOeIH4Sye04an2fScB1HwhjfRK0GvJiWdSLSviW5DkVEKI3IsAy8I8tFRJl
qx08dM2ighQ6Uw6AJrzWne680atzUYsUgrtWVBlhk4Rb0a3Xs8V24FrNkkhfbvQrBnoVL5opHTuS
xljfTQCx7cv6+2/PpIhTKUas1Z4+CoZbO8TgKwqVZ/2KsnbknconIpXHddmHCiM76ANcwFt1ia+F
R3PhVWj1iG1yV5V5XhfnkNdM8+LjaXR28c8wBPop9s5aCwKPCyugrQYST2erSHuPPPICf6ExIXX+
8BB46bo5qII2MXD/m0ComcCMyKSyMy3jYRR8OpJD6afx2vZBx4448JqB1fczGUKA7b0eIjzAZnVm
C1OrvdXzOAZLsVphvaF97pEY0SL8+eiry+WCRPCDwQtu2llD4ElrSr4QK5Jjxd354p1NzAqO8OCV
W/Anf6NGudTmizG0mgWelUP/7BK+ombqlI1oa65+K5u0UvSp0+76cjqIzzjmZGnxvv6NI3+GSO9Z
lzU8LD3Vdw4KpBNOvBHQ4X1WEZM9Wi5Kc5WJSbpHWga25oWaRT7dLaP0hmMhhaQOJ59ZSflC7vHk
Y4z5xujWRF0j45bm6kzVQlRuRRwbO++yr/oMWVQksRvbAQrUuHOzkjXzlZF7XDfFpgZVBu4s6yY4
tR0TkOo+60f62EZ44nvEKc0FtvIhpzRXES7aASR61CrJ7q1hRTtH9Ni71RK4Go+xgXEbmpNI01w9
pvTk9fy8J4z8JZMz06wt55qFIlAQB2sU0MevDZK1H0kzTgkn42dGYF9cKJFzpLS/PdMrjxY0kDlc
/oUBd0FyRJagYpWT9pGDaz9tqQT6BLnas05rRTcl6rZzq/TtlBSsg1E4wGXeQeFzf6ig+OquYLm6
T8AySHBL/1a+o6ZB9viqr0oI8WRxpZCFseC5JNMwEhmNURzbxkPKgxxls6q3iWI0HyUbeU8qaMFO
eyt3qs+aaX98t5p+BtiCQueRKqqOM5vPFpWlGaAccXuc3mHP9kfoOaTbdPcpltnUEgVfVhKHm7AU
BID6qN/ouJahQmZ4cAnc9f6XnKvcwW6vytYcSkvQB3R81YgkU4xse7WrqTJIT7vcEL+l29pZSmhR
0fHY0BE+JPbvl2Gw4BBWr3JCrMJEyZDcgIcLQmHIyJUcvzqNxctAgrphjGKZrka4+XPE/cbg9qrv
f4kU5BZVjhTldQWFzefjMp3BA1VVwI/reAITIa1wH+FppCnXu7MAXcjsUXwWyryEjrejn8c6PAAC
/P+HswjDNcXcO0Gh5zqVordYDLCACCej8dnxaVSB88L+38EbBuDIPW6CV2Luwc0ksERS+6HBOPiI
Lh7D2r28Qc8pf+oQuqGKnXCBNpN7/ROiX1dXTHi4N/h02o/ahtyzEnygwJ+9utij1F3WPm6COgZw
emS6N+pG66PDdHmLk8CPcK8/zJPmWIe8FWp9pl3wA4NivNb9QkZNrQkdCOp9zfB0kXMHBGe1K61d
r3Tu2p0LfbMeHG9c4mXh1CTaFiHr/jxZxgpf2nfP4mHSMi4bkltRQblYvMpGm9cy1Va7Nn9865W0
oWboL93K9Wm/ekf9ZWHEJkTsQV7t1TUTlPuwQST1k6XPkIvgeFanS+xGyKCBxTz7fYODGJvi6EUU
0XhEG5HA3svD4NbPNpEO4qgBYFkF69KHdBhFVT1sW8lCNqhTRCdhqxkzPYPO6hPX8ObZ0T1uAWR5
PELmDlFyMfRIiBAGtkVS4fO0x0aP5bBD0FKMNZpoO3Llmfe3aWunWBh1tcBHN/u/AKfD5y03NxJF
gU+i/M1iY4buZsf6nMGwrwKdUeQpZDHVN2bwK44OfyczAeYwh/sW6XTy1Dd2QWTnUNUmuOXL7hi5
CGS11gNYUmYGnb5rgBAhPjY9CzEth4lir2Me2kEQ8bx2FKKwBaiTF9luJxO1jIM3zzXV+LjHaHA8
yIuqhyQ8s7IS1xIN9pMPC82j+qZ7oWRVITM84ZjUPLGheLDQ94gOOljb2AOWSgpPvLJMwQiqKJo+
vtA5ifbRYJRYoPEl4Bw64wJAiad+YtGIz4zP0uwsuTMLxAwh2KISGqC+S9ogc2rw9tapFoWRUZ9Q
zJY5CQPoUb7SbjAgqwiEyUAq7sUfJQihqblsmE6rCirvkC12jQr9H5ohBOWZolWnkSZtUPdi3Rmx
Suvrs/QRY9k/CBMKKLn3fovshD8/lwDmcppQNy3pDEcL3v7Mn1iGstAQwr7sWjyoPs/x7rJEsRL/
llgOh/qCnLL2XQe/5yK0gyt5hJvXA7o17kXfp8ALZhOlJS4HTxTlgqhyA5Js6tCKHAivQWFBJR2l
icFAEt0Jrlngr7ePNe/mrIAhpJDBRu4X9lgW5GyleN5ACCpDINpr/G7Rijh5wNEANTPLDl6APEn9
89+Dr1UH9s0Nu6XEh0xs54DsrJNrRc3xfakO3asgZy9tlDZhyfwCSyqnrQr8lV4PpOl8V72l3HWj
sh0AESgkBFN1B9uo3X3+VZXZw2gVRaasODtgrubtpsPofZk8bOt1/R45V8DYuHRjZP6N/uZfqZ0W
XXysIB6kjkifer9iqdvk1MnBlGi+UQYQKgJrcQe+ryXnUim0xn47aKNgH3GvSmLryoZQ7ncM8Ocv
R+VbXRSQcoJy6+Ib5sKbI2OscfPm2HZe+4giSrvgVaSftMR+fQ6k11Kl3xf7B5f01qSnQ634/J6L
046r7VCHd7EuxenFO6IDY/mW3JvxxetKetUeUeI1d0xFyYCY4AfXoUkN7Mp5vM/AKU5Ytu5lHN28
859Fdbkxkp1C0zMptxBLln4a1CS1a/h9aRjVH+CXghtQZt3PJzdh/41danEjuP7ftXVhp/PZZ8Kw
mubgKdQG2Vhi6+i67UVYtRDYEJO1iosZ1sHEXpLTMzg6byGzn81el6nInbZTH8Xd+CZ6H8dQnohX
s8oM4RC9xlYBQesiOS5+fBgUPQlddJNhKJ+rH/nKNHaag4Ex3h5jSTSoY+flHXh6Xq6URkcMiWNn
nON8YgZ3OQ+1FxV2RdeH0retwEeWI2aWOh0ItzcNTamJm1dbwVepjUbKgFWtOE48rx34/m7SMhRh
SD/+wub22gYzLEkco7srerc/9+ySWpLYvM2SDoxoxhZzVOGMZ+0VzUMueIrpt9O0TGWWsAg5iHuZ
3PBtqDOADJ/Q3I5VpUcUeNbJHiibg+6g7b+jcM4pj1v8OU4czvNdfuhiNUNN3Cjy7YFhbm6FPnmJ
sFznYCVyr4qsaubi9uNNJwZho/7clwCI9qWBN08e8hitcqcP6xhRddcuBxOc2kvLaH6Z1nWAsbsB
APl6VX1XKfyKVRe6YtxqCLvYE2JRlzZDoF7ma7HeKptce6oH3h5hhFIZQ/rvybeVf6NIVCkYNB2g
AbhL1sRhPpw0bQS3ZpXtA3VcreDbNJ1anLYjcezMzpcyW5gURGey78NlQYDK2tSu48HlEvReHONG
XxWTbu7fozjgAaL+x0Ss8o+E3gcxUnfJpNGkF89vwbv9LXT4V0sfcxmMtn3ngndkTMe/5iNTvh+A
KEzJsDxTEsJHSRqPni+y/YynPrYfa/bQsKojt13To7dfYM4dBBvNXmbXgkBCKVcuMz9LTJLJouam
fwsi/SnClC8e97BD+9NolRuA8qALuX8H5c5Tk1+36N9jnoEUWcgMww8W270zzjNmIdmYmDqh0y+x
FeIbpCom7efiAsqIdhtSgir9lhOelxgzpCMq911cyu/GsjAkABQts4AudWrbvl32RP8blPKVWpX/
bp/bRqZFxcUXvqIuHQKJImGrwEuNqPzCPn765OyVb5sA4TRR8kG3TmF7nJJR+JqheGm89WLbwH+g
KBwImFv77r/GDRfgJ27JkfbFmS4woHMoEJZypuP7WT2ZV5pDEeQzMiIjfmN3pVve/rnj0bLxKHlV
n9xAyq+INbIAoO+PyzXucCJpWxiiYF9VHcCpxTqLJn/YEiAp/WgrwlyqTvoej5d9ILLCXf65LER6
yqUePO5z8rN2xTAhfZoe6/NpNz8tEcQnYzQF/EIlCyNpCZCoV0ikki1J3ERd5+JazxrnZYGMZhYB
WlpW2kzx++9daJ7K354BbVLqTZ3dyt049KTf2+k45QUt8WYTpZxOhNE4VZmV7CR1gAx2osiEjjoh
ADwoCC4z2VFu7yeq3HaMOXONKT2+5u3YcZ0nUFky3h+X4tKlkpOVfORvB+DortYocqVrK5asf19g
EyYdV6lpUfkzQXArkKwbMoX5X9ybQXYDQo31q4pkkX/u7US9J2EnnfXqEoSbkxiMQnWivGMq7at+
f16qjtx16iU+J2aIS7mAWMACZoX/eSE83UdEymOTfOQN8f06ljhpfjrsaXDFTY2eEQIDBftwaIkK
kpRrxBSKOuWhTgLq905nsS9GA+fRBvgo/kVeX18Ozf6mJ5qoJz1sRE46x4+4T3VR61PzGbm1syx1
/reRRK6PUUY7J4350OFDu+1YUYnCHa/SHfHtE4XxQ/SpSUFBvUapoVHmt5/6J1aVuI3+rL7nkA/S
xvUCODSz12abIhDsZj8AYmR0ETDqh0IZE6ACds+u/1A43duEh4Nej8T57XISYmszXcOqPEPsef+U
8zVqusUWnP6keU9OjRF8CW8Fzs82c500H722xZWfcwI2XVRlkiO9iymyZjaNLTWrkSAsHu7eyBam
R8254OYXu7k98h7q5rE1d+rowE6w7vzDE4j1X5Win4gUd4/9EUYPSst2CX5jVASQo9uN9D2L6+qF
7tfX29gMFiW/ZBTZdkUGAkWp4GcMe1GqAJ4cLcMKLgLn0NSee4T0laN6/lLPBznOFnvN4yvDl0gR
y9qFwe/hjyvic/uvhsZBylwXajZFfaqFEQidiL4pvVD2jGEQwST5cZa1zHbIzSRX5p/BFlPZVV6R
YESGX2JcG8ENqGBN7V5EYYveGiDUoPHw63Gtvt5O3DEgJPmnHUZggtDdj7odKjNfNi+4b9+ZHFAQ
HWfAfm81DHsKwA42bc1IALNKblyHQRPqxvst8N4o82/jJLPrrAVbzLRk7st4WrQymJx4HEu+p/uF
MSF6gzKMODXhX3jQ+UYOAf6wJLS6zUbpqUOHvfZ7qKSSahs++Gl4tMW9imaTv4oMiCykQ0AbWh26
d4qmlPuefVRLHb9gAUE4UYlsNyj/I7RS2bszohYD1OtOKA5I51uUZVIB2rVDcPQ4NuNwai9E+TT1
yYNb8Gqf66SMNLUMHv0OkdgMsD6yAJuYVv5ZirkQ6ghJvT8hncA6ANf++VSBxU4dakyGSiavx7h8
kd4R7IW2NqV/E3yhlqMOFG1iuyniDVdxAPrdd0ycJuM+dB2iAIyKh9Y1pKJc2Tov7oizliXzWWxG
QsSTJkkB/YyHe+zjPVn5udAdwyJdlfMPcW8/FExSgD9nw8otN2slbGV+pT0vZmdDLp0pIZ3+ryzD
QSSjRLUQUfo6whaTufPoZZ8Jabe8UePsLTskI1jsrAsiTy5pAhLYVKD+1LKXa6MBhhyNj8kw+isy
L7jFSaJBfqTZwvXos3FQ7zBUgI3E52MbShA1FGbbB9CW4qFfnbTIOinISeSPP9UUhawDGj9UOP3S
Vqd3xzIlO7+c/0jb0e8MWIcSvjvfc37OmQgpibGezhaWEzbSvzmzX1qeppDIyle0qx4XN1ZbkFIk
Vu2/1In2mBM9DhnixdDDq707CLSDqxe4ZNLow6bUQM7C7SA3XAroDifZ6RF+uAFO7V6sR8mAtagI
NLxBe2ClPxVhLpFhe9cEVxBg+Qrb0e5Lh5hrDJrIH2pquoB4PzFtZgpgn1r2EVAOy6kPf4ZMxfm1
lwr4h22U6gXh+3zx+2zNEpYpHHruf93ZJjNE8ZJKayY1tQbKMhH3FnYPzsNDE3P0tk/7oTeHluaC
haco75W4O0ktnWpiGjWIH+2yZkOlWKdKPNDoh+8a7zruUIgK1Pf5dYLvZfGsPsXcfpLVeA6BwIfu
rGNuy3uJeNqUL56dZRnrl33r56GvR1D3S5LLRZC//YG/1B2CmlsOATCtkdfOu4yqBNgrMpKbNnaF
Zp616xhQmeiDBJR+UrSjFZbsxQ6xS0YRh7n6kgr4zQ44yb/yiOZCGaLj1MoznuJ7womLOKxAK0mB
azIsQS2ZeqDd/gGmw1xGRfr83Nt+yqhMLyglLikpiXj7ykuBLuU1K703ufV0SvpxXfHMM3b7FflH
OB64OyKGPKJiTtCUwGQdF3NCya7ElezUR0c1MryXcmWXhBl21DwCipveaoB5HUJiewQxpdn3FDTQ
VV8rtXUtGZ8ZDypm9GprWwdPTxsD+xXHDi2ldxDhZ6RUJZeHvm8uOsuPc0nij/RDr4bM2ogBYj15
IYjV+vTP5dA+/89VvwFXtGQOKcXc02SOu+cgkW6UYBhInZdGGpPSLXZeGu+c78xlE4omJTUSIpnw
IWvXqXfTwXUSQ0uuUYNZbKRKF/TVrstF2mUxDLzg8VY8fXkESncPPg55Z1XocnQsnp5xkXoAoFdH
St3ER5aOrYHyP1h84SGt2HvwmOmaiNApNYVKfSHyy9pcCR9KQ6Fs+Ga1AAilLWQMQTbW/VSloQRF
NgPubXYsvgmJKuXH6ahhYd6pjdyjWjcpNf+wLB8zbWDqmlvxSVpYw0gMvYkQR0MDDBDybLRunn91
c/KCy4l4GSxB7hmd/8Q7ZeL9iHSmOkHwC0L4PiRk2OosTC8eywt1DR7dzx9Q4YL/tDP1axX8YQk/
AkYpARc+X9vkDGAYSyjgflP727FyZ1fuF6a8bN6T49+9+ap8Tc2tKuIiTiouB+AP40EW4H7L1884
hDR/OiBbEIH0RUJIPFv5Ah2br3QbipP817knzrIuc1ZjOfKgVVx5oLGritmNZeARohGSYXVNBKQl
+SgYQjUFN9fnw7/DJPLIrp/tDFTYM4Lc9KeikXjOVX2r+EuoL/O06YPRbQjrB5rKHJeriqr7UBdj
3gx6Cg/obzxULukoNLktkXPpXvrp5u+24KdCKQRa2mRLNmZUaD7I0tEkWLiCkZ89uca6d3ihv57r
oyaZTBSPuWmL3QcOD0TsP0qSILGfjh20zTiNEyp+UoNJv1dlc6gxIkWKvswhOBIHiPXKSDZ+WSua
oKNb5EDYqZ/kZdToHk/jejm+mMyanyNga1mKJnOIExXv2/2/6HQEWQnqUzADr91E3SUGZy9DNIfk
hc7lsC66LLqeialu07UDBxgIwv5IlQnOUtNX7TpX1sq2DtiJj9sPw1vp+s/U5daAe9TE+Pa6kRX2
SJ+Mqi2xrB2c4dwYPliM4lXuJwIzekLnDR6Ffn5aRTJvZbm+20jU7wftAQDNmz0JrG+fwBD+tklX
UxP0KD1HzUxOZeKGQl9Dgb/ZS/PnYN8LKdiOgvySRibHv2EI+JcUxds4aScjDQvMYNvA0jMesqZC
4jT00Ri5z75W72L5l/6mLdNKcLhyPLd/E1UkOud78lYVjlhqyhVRLgccWeRVYXv1oK38I8D+BSc/
CKUDVdwPcqngWpD4QfNqgLtrNRlyAmwmg7vK5HHlEqHWTft96IsGuTMhHRq630lWHC58EV6SSa3q
6fBK6IKTmY+HUNy0Bn9797ye4WlkMMzLuIGPHBnhQtebfUu5ebv+ggUoUzG0iSOTKhaksbEoHtoc
6OuLlonhmn3hA2qyKtSxorLYl8F5jZzX5q8Dmd6c+F6rdmtY+1fqBQm4ukYv5EsHILbBcbUJdjKU
4wWrB8OauFFBCfcauT5KMONadqHgMei9+1kMertYP2x2lUu+xyuJCECjgsGTbf6R8lCVPgn1DK53
2Utl8278bkp2x+nBZiYEp6S8O7ZzOP/9ixApWzT43WCS3QQ8FKBLvOPESAucAFQLcp5skivh5Np5
+pX+00thSO8oF1VsQ0KOIu+2lQ9PIc4gwOITaeEt/wAFT3Th248QT69pf7gCngfjFYlJAiheyMqo
HjZcmrjzxsIIMWhLmaNQk/MNVFFfTLDKFS1h939k/HEoA0DdK7sofKrM9VZBWs27lG+i8UVn/L5u
kGboTNez753lF3TfNAqY66bM5aa0v7HdyFXv7bkjg4vtBfM86O5vzMByZ9KLsAAMAsIO0QmwTmbl
S2k+oyBkGS2VB/Q3rn23L1nLoib3ualkWf56JjyuN7b2IM0YFX8sdHRi4RJYbCP/VGSUW0//tDKm
YkQ89BQidn7de/8V5gVtr/VM70JbEnVJF9QxhIhJRkrtJKg8x8TMxlHc0jBhtnD99oZML1wN07Zd
hKx7ua1EFEHP9nqIssctYEcVdw9IP7y/2cT2QIYqizIFsex2PcubvetnmjJYklmpwC3VxCTDrMob
SBOfpn9g5McUlHO/Y9GKwpR38aZNPgNenINj+6QarVY2QqvgBih3OahCgiK2rsZ4dVzZhxgOnL4v
sxGqtDGEwkFUK5B/xwl0Q7cgSFplQLNxbS2ChdQnvpG5/n4xcNaU2oqvCHZnrbhDUmzYRAObGq7a
zALhdjpR1kFugLHFNP6BccIeom3YxM+vdMh/WYf2gxDy/1bYttwK0QCvZwX5cKV9k7SZL793TPOh
feEKummpHbLmRNUp2K+y7sw9c7rLHIH9ByOHvQeJRkJkTEG7zeUNo3wYMjQrMzFuOeWSHlbt7iyX
Tq27bGSGNEZXDHPArX18b+/txZTgJCumnhpuThB8QuKaFKe7PG6lagINMRiN/qk3f48x0JQt1TlB
+OIb9lCmpRlGHfoD9EjqX5WZVlHOftgdRU+GX57XNUmP1AXVAjseftfDRb1wz0D9dMqncDDAp46V
K8og0DSsxORa04aKqO9k0A6OtyzgmaT1hKJxIbXLbaTx/6ZScDGTaRfuhjBoczPIj2P1f6FX7QAa
FtLiYoIGQmRSVynQa85uV8Q4aN9EgNKzeUUA1o+vXoHHdX/joNIt3fsBJjPqUSwVuvewY42ybXTs
gjszPR5oA9ccMPzEvkW9mIYnstYLOcUpPlQDKCEMaQ8/rqc7bgu/EoBOl8SrtEKibFBP0X7fwStZ
BuSc+OJE8cvtO4bc1Zt/QOuzVReLSoQVW0W7d516EE8VRjucKNW16qaIrrqHrIc9BW98atFUdhsg
X16wXIEHJpVKTFhDE5Dd1o+HAq88MAbAF8ciVo7PZIen/TDNTzkGvfij/IqpMLkuVIwwHL3udF4q
Yr+QisW6LR/zuNlL1pscuk5PxeimuvYYw1ypBLrnJqUZEKaYJzyWvnlb+B7gAIx8owUp3QVIxL43
Pjb+yBhfUROVRL4ROFCG9HBefFJStLnuIOUZ/w32ZxhzmcTyXwVnfHdgICyG62yOzEYxgKggH5nv
A9HRDWoUXckOUEgmjFaqd4RxYvIgEy+9HhpYgUMJRa98tzBLR4Qm1iyCIQgGbqtHogNWgpIgKrbA
6Zrrq+zFX5WsrxUTOQkF8F5k8px2QbPktgn0BoLe8gm4/j6CwB4Uz+/psPeze/jcYMay96qFrYkG
8Tb3lq0aXXlhdvrsgVnhy7PKiVFOg1zDsizEa2H97jD/rBsX+1IA1I5PAY5br+Q3MPRq3j7z4hed
feOVugf0mKKlnrtc49wR0z46I8w/uoDunUwuEAzES1pVoUYFYlTtH58NEvhFtP4ck1KPDhWXmVg+
3Xk81bYtMQuy9xGMwqa5Xl1MVhn8W5wTSlsFho09rPZ/IpR9QV2bHF/7n6HKR6Q/6ABuQ4vk4r+E
3ICPv4oxhqnHf0V03ADFXLn/z7e2ql19yc1T5a4E37xPv8rhLH6LZ0iDSb9gugyMo8ZuUbMR76ww
EEJ+wtXhcvJPhRRK65IhQdepqdDiZdT84uXZSPYxG2kvaT4FjF1rwOV2peHDzxqJnN1tozSnBVuT
4FUT223m+K/MSPrcdocB9oQcg1Kcf8CeCLhiQQbcuSrCdG1R5nvewqKRSqu03ppdsMM/CY5sX3Wp
9+IeBk/edJ7bj1jasRokKhypV6dqDHmcQjfsLVcXNmYIRu96856bqkkWAmFKhV0mBOZRAjjppoCI
9F0ug4PSi3ODF2pqY3Fi+U5fKXp28OENHzwo3Ml4zftXsDnwVe3mkYU+dmC6m67EdoVRHOWtLUGP
AjTraGiYAaMGVeTzr+hWrmFg2J67YGCBH+wDaogHXQVcDBkw7UXKNDbtBeUdQGQhhrNQPgPn3IiR
cMknZ2Kd3cxOa5miNNv0toW1XoGEh+ppb70F5664r5DGRmyS6TnRYMclBM7pzY1w/Xq3GTXXb1an
4tODy5/XjM446T6lm3TIdPtM/zNhqkBkOOqWJKlp0tnSmv1jnKM95/s/q9ynEsbA0ln7trTBn8b4
xbJCWrUI5qtQmF/6dSZBP2n0dIMFjF20OCmhtKJ9ZQIUwx1FqqCs/ICfN6x+mJkra6wEPKhLgK4W
POSPwoRdC2g+9khLe40fSSAxm3gQZ+tvvmfIoNX9Et3XLGDyI/nLuEVdRAiVmIoo8Qe4W9fWk03T
8rfBpgfJzH+jFvJy71oUt3mKMm/stpRBun0NJd5fP3Y2TIZ8CHNN28wL6mHfHLItmMsl7AF+4Q6w
s0A3gqDLSKs39dbXPP2cT4sc4ZT5yuVWdiZmQ8+IAKxvjRiwGm4q2VwWi+gi6rmC0mqDpaJ0/ZQj
R43DuuGcO232CliNM9xRe91njbvdbiz9USnznCFD1yAPwn6t3Kofg4fWgfZ3jVgUvaK3CwlDvOdp
y9IdYfBbL1Y6n1MAn/PKGoPSUSP/ASUKyJY0e6l0fJm24AdKANVQgC/CrMIwuypSI5sicxD6Zr7k
+9PK3FsNf/ffl6uYl45t2Tu7ACZgtpK2xEJ/eZUbaEjjFOHzgXmcG2z4vG9oYs4JD/X4xt6vh/QG
aG/ewA0aCpyyPW0DPijS0PizKgZjXB3XQYxp8vtwXmwusikDHdOUFQE1fXDvWoIqTaXarm3gBbgC
CLPXZAH9rE+ngda8NEMASg377O+VTavNFHfTzA0KjqDYdlXAzPjKUAmkoTpihiYlCxkMCIlivGnU
3wfxRJFkFaJuNaDII2EKc/i4bArZHBNy5yBFm1FYk7AS7p/xNjRAZQZvrdEC/l7O3/JhOj8RAvdg
fLGnQLDtTsR2wl3MV12ZVrVQu1/6VHXcb1EOeSaQoh4fBPoNaUlcG73LGtZXyrVabvXyobouYwzg
hxrYb/zxLl6U0f+keSabnuPqs5CSQYfVeIQdisqcj5eHriJwnrYQrg5XLLtuB/30zZ96vXxi8PVs
I2Y9KgyreEUVpodcwLiY8uGW27iZOsJz9wT3fvNWC2tZ7FxH+cbakYZUBXrU2rxATVXCVKB+MakG
YxUUYS5qcVWwvL4Fc2VJzakAE7TkpuT6xbJkTWZYHeUpZK0wjnxLL98YFKIa0pCQGDVyjuKirDhZ
QDDfXpSasUA3Oc9WNjBVCM9SkmGTjLrtP6m3uKVwUG/JInf3riHbyTs+RbZyzyNyKOvK4cqb4Wr4
dQ6IheBMpQc3SA/DBGjilj9LackhUdYSuBsQS+8ZO/gaxdX+EIxtb+5QP86p/WeyWGEpBlOjGdr+
ycIRsnbkLecU+LdBhvVNz/GYvkSHWCavG+xyD9ePoFRUJnpGhg4Yf9TFmDYE6sUsZOcRivdioEUp
LLkqOHpyRFYfW6k/5T50Hyu2/jgv58a2Q1o0KrjFDFBPs0XVG01nWa3X2MV/eY2BcDO6m/ZJVaD0
IwCNE7GA2MY0CVh0RUHW9i0vD7+QJiToXD2pekatrdNUB9bL8l0yOjYfMQickxhql6u/1iW6D8o4
GpksWcEYBi09NCuZP1nwq2PC+RboXNOOs0j3hVvHVboAc74BXlhK4ArzVqPcrS2fbrFO4T2S8wrD
3NFW7A1WRmg71Np3irCakb7Bu1biKBghPZQ1+8+NVtSPMcNqqtbze/1frnSqVO7Z8zbWZCDs5qgv
1V/Sg3PaOf3t2FWBorb0XOwWaXHmCTzmtIJ2N9SL2HtmIPt8iKfiCaYPrXrJ2N9JXgquJc4lNA3Z
Vi6vrETP9ZRz3nOC0oqbXINGWiHUzxwFfWRTZA0UrE0EG+WOlXfdO/Hk6U+hFwqg/G1HbPt+k748
APBk1JCtVWmf2iyroG35HOKjGAg8YWIXFQ2yhtO3UR34yTNt+m3eFb9+5j/TEBwA7LWC2LB4dc9e
1kfHjQyOb6gug4SFuMl8JABts2/iLk3bAWkZj33O1Zzu64CiBh6i3mJ9cQarDr1ngLHEzYpgrpHW
eifD9J/YMUuk4SESEtbVXaxfNhgoeBpIJ1a9Gk9hqmlt38d3ABebEU178y9EvT6Uoey9ikBm9L7i
ZK3ns1E7J4EYssgDRJKp53tSRoSBtxf4l0OTH2lwX2BxWHl4s5azdPAoYUfGFn/ST4oXeFCZuUEV
BQoFYHfEby0hoLO0C6U9RKzlIkDc1YgZ6xK6XumRSG3cXaIwY9bJXOAjqv18LCWDTZwa0BAoBjHk
xDHW2Fr+emxyOf8AZ1qVcphCkA3olCmDIG9+z3iH6Xmn0PtdGnnpTv6OjvKDtLVfDgMFHkvnmd2S
PE4scbMv/dyuMG/rUfyGV5mWE+QkVbWMk0jFHSaz64oMj1xN/TmGOXERTVY8A6U04LsgZBbk90GS
3fOPW9GnpRvas3xuwSA5l3/wRKGsrufg1wSDQWtFX+yR3yB867SWszAJ++DJZIDpHv/SPL49+3Po
YhULl9ggVONdv1i2VFr+XfRFgXkLydb8j0y/QLe0RB3L/n3bS85cmcVhBWx6YdwKalWfHFHLOxqA
2VpIcyxa9MZKj4SPYo7g5srbnmc0AeogCSNZsLVfLFo//ivT66PlyVxTZF6VCRjxflyRXPYuSiKs
aZk1j1q769kDB6/NUo7lpU3Ib1igWs58KeA79xg+9bZRl3h6XTpHDvWvDSjBRnQ2mdhG74CQXDN/
D3Afnu279nEG4gufP+VOWU7ieWIOfss3BS4tgqz+7XLVOtOVQa5ZG0fqkl/P5p3HpaYyyL4oqZet
AslSayNWMaW6JfHrck+m7iMyKOqIzX+4/l6Oh0X4lPF+CxHp/Wm3kRD9zCXuScJdZsZUt5RZshGC
2UM4zAiiTlP3H9mnezq2+0WYbJV+lNO6i7U+Fpy3tk5Z5fDMjzVg/24h7F/6VsO++DHiNd/FAmlU
1uZjg8aGY8HydYSMzDVGRWiaZWuxBnpaWFNqEjv/1ETO3CJunlLPzzCTQNypGpH5ngOnwWUgAr4j
bPdNfm+xJj81Mk3WuJFqywg9UZWD5JNLtEkvEErRIY+/nt9oMwzMCt0KCFCm4mkpzdvu+HTnPR2l
2UjHCNjxZ0Gd1ekABVT69dZegCO+Lzle8w1O5A1MPKItwyR1AcDr6LWAx4YDJ398KhHleuPWmEC5
STHC2gTl6mlR7O9SLskuiNy8ULh5i+cXq6HdnlkGBnlkDIMyI7fezBYPABEp98KV7aK9NJl7FqbY
YmI+hGFg0QfMFTaCmeyQ4RJIvjjem2Fj2OYubCOmHFA+pt7mr0tES0EPt2X1NufvRqFs8A045NxO
3KCHqXfolxHa52OXbft8BIyZNWMVDOXkDWqZiudXHABAWKnmGhX64iVi0NhEvAkesksUiR3H1kXQ
Qu36E5bxKpMobvJ0t5tiayVrfN00KZX/+I/112PAW9Z4IKezmFJvNR0yec15TfiqiPaoDcZubtm2
+yUGpZUZkK4JrlrYhVqXISvEW7EbQBfz0EIsXmmmtTZLoyjUd3IilpaJkLcREnzcRSUkGDy27Yzb
62/PiO8Ev+8kWRqgR2hTlTYc9PBJtsSqS+MbFFNNVTonkuuCsq8xf4D05QzM+CN8zylQXm8ILkwW
Ib8D+N1BldVKrb+a2LkErmo84kbfnQp3J3fNNzwzW+QnJqFGliqG7D6PiBm6+GR+Nn0dNN6cTEyl
AIWA9ryO1yDzeqc6kHAXtynZDL2TVafBnLlMZpgtrmQ3jmO70lrQVwSYTc7AQKaNSR1vnz83uFnB
AZ+LR6ssC+Eixfyv3bYGtwyI3Zf39YJwlqrRleo51PL/QMgU+xlJf7r6NWH0rOlY6CPySaRAVahr
cX4UuhJ6ZgLicGa/Ai7CktZ+kt/dA32fVgogDo4VduNiHrXLvyV4IPYQm4OSgmPwkI7uehYgccPV
7BIxSPJHqtm8FCcFwfZm25GdJFSlugNv3jGauG15IHtZCy5HgzeYuJg/vKVzFtrf1c+x9DygTp/K
aU4kbq2II5m2JOrx27XBTMuKX3RRffvCgeqKkpY7s7iuGrMEsSvbrmf+vNHSx1CG0jdyzN+YXI11
HpbynrEt6hCM7HMfHWjuzu+0acCIBZ+VyE1HksGGowD8+tmnaSpfJDI4lDEZZJw8XlPPUu0eSjYV
WjkmUbYyeZaRMDkMXAQoAIxuCOZFRz9FzIbmzxBntqrA9oSNX32J/oK5Elrqd5CHZDny0FyUosOt
H4sQAfIQzbAyWSe45n/NxNdnA5lO0D3Yt9eyl/fGafJMJMwKooIOY1H2E5piwJmFa/6loJCaTRw1
OgPYSaK3X1fMt23/LYKmLqwdPa8rL4qWlLNqTbcRlpwcKxKETyGlKiiuyPBM9k3Y26pJWU2vh8p8
ehl5ITlJCQcjGDXphMFKGQ+k7sInJ/116a9kg5qwhpM9gmXVNyBXfiip258tT72rWDqOCQykJn+A
KzXKFEbxz5Gc60KWuCGBUw8ORA82eY92AMYDWhN7BH1AJ22TvNrkSlNKXFQ7j+RtpqtbCIPuor2v
CmPFk9/fGUocn8ce0V4AgmC5Uh2Lh/cqai1/eR1Jw/AmVbVvpBRQ0x9Ge/V/4NiqLv/hg1k99TdG
544ewyadeZkTnjqxDfCBrqrtkxhdATy9LJz2kqgORrb6iI+LZyBQmzSlGN8LLAtHsX4E6RshnJz8
aoDqjLScvyEiyHZ+ibKql4s5mY9f0QxD6HThcFrOyIYsjgGEOuYXZ98aus3XItLMawSYeOXsIxkb
mAfkRdmxwo+Dgbqf6UY0NovW/G6tcYK5rj3cLtB6EoiMbvtgvFyuQhE8WO+/oUu9QMOq9VLdR53p
fLB1w7JKQgBQ52NyGNeEw3jqlIE0RqvEzqsnuw7cPRMsyjTY6nNmE2Q6+a3Q0mhxxepZkeG5NKh+
CvXodukSVi08Krwo8NgmXXJFtR2iqtCBuu23L7kqTlKZWKFoN7oi7JwBMGrw8+o+a3BgR+xAIy/G
EPKoVsIUVNuX2k1gjP3I/KL7TRNGvy441vaequGDlcCv8Nc9h2QzNQI95c5BeD/ixqwWc/RE9dEQ
pSLkd/D2OHwGQi0RcgrvoeKDIQeG/ClMsQ5Ji6w/ZaI30lADsiULZIyUqq/1LQBjYnB6bGr7NGGe
gekWIi+PBiBM4UI72AxOeHdgZuaLnyR+fbAwIP2H25OQi5WwtkTzOdEzoy4+WWVgDQ+//Rum3Mdn
7otRWHScONHlDxMN4CT+B7ekaW/N9Q1t4lO7K0DsuJSbb3uX3tzr73L/AMbtZ+xnbeL4ekpNVdUw
H/daxhQis9M/4zZlPj0CR3aNpSceXOm6LrLKzMxHBQ6hea7PzOMrEhF3cUBJkuDKYwKWGRKrK4vs
TYBYPsHFL1ECz8sp4PSDDrRnFkPlr5cOGj4T7qhp4W9xhb8Uf8IgoLAcvKEwjTwAABKbukFcU8EX
YE6K9thFxVg+/8en+sJ4VbHMjhQjoFChOsxkCCfyPlOoPWqLV8H5XvfDEtx/GccFSRZPuqN58Oph
9YYbBA6Tp46dBW17/MgEuFf5lI4+XTqWaXUlk3YxnOFvpe47ttBi0t7mVeFaVKzD3TtxSfPsqd1Z
KSWrZxuIMTTVtZgOIihtMZ3dtIjZda9Pvs9G7ehXKPDPU6DvupGdjCa/WPOSo2qc611VhWmOuXLv
hDncq9zcwPh0Cx2lnLIvYfTirKJNI4s23hOpRYSykZBJKSmcf5z2P6C2GP2dNoNkMgZgp/Es+bP9
pqpJii2hyGOrdQOPSmUbj48T5tXCqtNSh7oePRytTkzP+AiZcDkE94tUsM9bbTyBxD5GSPcV97Op
N/uFtm6z6zPoA1CdwBlShsrCW9e2sj3+aqPsN6X7ra44lhq+GNkOmX4yRxBmlJb2DBM8mfAlfWhL
gkcxMvtRQb3T502NR7/7zdJAiI2lQgNIoXkqclU0HinVv3ODKdKv973C9ahW0JAoHV+f0g9yDmf1
/QyoN2f1cDXDVCjWN5xfjPsVQhvaSjjprOvwUyc6TlameyPTeR+Wyc/KheH04d5zeQ98muhPzXH8
fDrSAgU4SPsuIhkaqsBz3vRP69XhkqCmlWZJuXEDDTESzz2pYfindJL/B/iUnlIGdejmMWMQx5zB
YzsCv6pLkr17JjxvRxpmudvJUVgPgN/+9TAtErsC47lHW5jyzrRbjpzUH3KAXwttW6ICbNzUfINs
OT8oT0DzXyAl3JnDAESY7WH7zVB/WahYNK5cJQNUVFxv02pzUzIVwrUgkSb6sZiTwxHt2SuUL2tS
tob1NAvBxuAsS00r8REp0GVg2moBtl3Y5eU8wSpUhNgxB/tCjR/uF9sVtA00G73ZspYr1pL4BYP0
sjouB/JVVocKxHkycsnfxnE5FvziUG3LTBg2VaMPrFwTxfJRqMKp/TBBM+aga0SR+fyf/m2RM3y8
DqG5+bCxZCJMNLeoqu/Np3XdvbJSYDdfGiLrwyhurb0mQxBNbJ3lzocWvDGRJ1Gy9F2V9qjo4JCm
fMqEn4xvmDO60p9MHCiXiat0kUWVxW4k+QISobEaDtSmjJB2XpN7JEJVN0qkZBk4ntwxVNmn0tSQ
z8cTtQB3EnLfmaZ1k5sSTp3OQ7oAOCn+sg6fo5zwISyqVKfvxWRHRMgC3b5JIaNnHkNLzaMO9Umw
d8rEzxYb4ICCRWF2JVljmsT7z651m1wu6Ilx28mY8ZjfCJYXxSFmZHUSd8sdOr0BMtNnzDQ0mas1
XVwRtA7cdep3xfvoQrUYOJMfCVGkSyslsDrDiyZeD/t6ZrT8BPqEHM2+I60Ndim1HWDrhQ1JaXer
B6pCEMCaTdxeZskcHf19LlorqX+Kke15TxSSijjFRD3jSquTCqPQ/Z2WUBootucLz0gEUCYBw0Zz
lyQpl2Lyfc1bUCIOXAIXwWDLGZ8ulnSe+L50OtdI+j3KJFOSP49pvKugwsRy0fSnbmWEwU8zxDnj
+xbm0ejxMtqIsgF+X1ZXpEd44cr4qP1MVBa9wElvDRbDx2bnoFNvo0c0CuuscizOmSO3qiN41PO3
f2pUs9jpJcZI4y3EDXvcSlyixlpcx14XFEE3DGK6iS8DZCLI3yl2i4SLnw9uX2tuFwAPpNYQcuh7
q86R/uuCkgeL0GipfABEKDvd90Ql8W7Zrb+i3lkLtCiGpSqd81WMF7von6kqdCzuFZ3pUSAkuE/3
3EvE25EcACkIgEaHkgHosGt93KltjnH9AtiOE9hZl4G/o/dE5hpCTFProNpyz1XmOb4oykoy9GWK
C5OCB4AHtMgmj0VaOWUfaByYFEtEwv3osGr1l9O3r3bZ+r1y9lp+HXES3osWlHhI6k/Fpena5b0O
l3pnXYj9jazYDv06fuZVjqHXE8fCVt3W4NFWdihXCTrCrZ8GoH3wCoSHGgrUSKRjTJS5kXRIbiD7
EIKkWhBQ05kThWcS1w91jBuTXN9uyPgLiolJmBxoPiyEjk6H4hu+dCPO3QBaA2W9zKycpDQ6fskq
WOHEzYWsw9efjRg0LLczvJfFjlGywIT8eyUWxaqFBNTpqYRBToF+424No+f+k0eTouJxHw4sheAk
Ux+bnjJqp76C+o4MmAIQtiz0ZYgvjKT5YVhTOYwet/UM+X2F1ls4IYrly/V7fPzSKX6W4hkvI7gq
DPnEf4k0K0loMRSorbkys1FliqwDPMlGcsBBsPs9sFbQqew/OEFtZ/vgXrGZ1amqTyf7L+zeswrh
9+oUspcfjVw9aZ91/ioXGgRzkQz0tqyXhK8iYDmbK/bnZM/M//0U7+EQmOWRr84j2j9KGa/JKp4d
FESoZM44J+8xYDRBNF8jHnph+cDsbSPxFeYwNNe7kzpTtAD/Z0eMsNHohR4VeUO7ZyTxvYKM1RLX
pYCjfSoxUr4LkGn3MHOg50A9AslIT7IFhkphw4OBcNkppLOmUGSfKlTdY5czhMa7ZmckJm+FnPtR
zSae4U4hTbjExtNK3fnoj55dYCGWbjfjhPno/CVMnoCbQ5WPzjdw+CENirg3azBepPa6kpWRBs2K
c+pfo2XPp0NZ/Lx5ykYV8xgtnrbHOmBh5ZqLMX8oBEZe697I2QzEB7CE9ygB3oARqRLjlE9o/wJI
U9tdfVGmqYibxzI81XHnU1F/HgYypx/WpaS/3b/xPYjT1U66Q/FUD6eC/QuhH37MQoe7fLLgfmuE
fVmj3YqIrLAVt2GyzPiz3Cdrkj1m/hDtygLj8cUeU6NBf0eAeKIt0JgwnNLfr+2aqtIp5lDJsb36
Yv6EufcIEqjqM1d1zT4Ji7TE8BvEkfPwj6nnE67Fv0x1Ufu0pAtrc/ZxBALr5abxTPQ8aObe0tv8
cVZtk4LvMtvtomE+fc/Qkoa5SMkXiUK54mXGJGXDaooXDYzARXcIk5YQPfe+qn+J5UVuMcy1z4f6
8D+MUOuec6BTzKYAXSqIKmDc5yDp1FKSmfq6z1ElaQR+y+0DZ3YaOzLicgX3mFLQnyRm6ZpLbbvd
fBl5jfYXpYX6QI/GggG/HyfHtSEskiGd2kXxvbztkaDFC8BqxjpOnI2V1ArqZr/rbYvAN87fI6HC
m1OKfLQLMJ/rmGzRL7KgPwbToE1R1mN5SPFQkBc+OROWWNxdoax4Sq8AllPaCvqCDkgBbFVzrMd6
Jk57rilWOZ1wMQG1o0R19nXIr8x3YQ/0RPxpbjkcxD9/rk59ZSJ6GorkzbhUbGUpPx5G/PZ0dl7u
nhd0/Pp1doHGVbAIiSQgjhzzTZqLFsXXNDeOKzwNxFKzZWpHdviZxoUCQF2be3gakHfrWs5oM+3M
/0w3XqfTlE0/SnvD1TwIyUO022KblmWZM5lsx3+GAwBySxvg39/bB8qrSusZrzopjEriTp5McZyh
in1o04aaEyE1/7weNuunV3UVHtGPeN5xCBN7SunFZW2tIVEuMg6XoSwQmWmNdnuqfoAhXTgXmkyu
GlaMn3zptH1ziAX7ogQp+fnMdlPT32uLKwWt8swzqGnKowRAzXqMEXpdmvmZIqU8ZGQG0XasZ2L5
G7VvEQRbmCNmqKndpGQGRk9vvwtuyaUX4d6RNr38ymWtEj7JLB58KooxeBDb8Q4XCgYd5IMBM3hl
9Prd1QoXmRoVLgjngl4Tlrr6UDrjzmeD+hkkH/cJOfKX7GAXDgKJ7FH5G0X/5dLRY6bc66KK/a/+
dvEHhsYKQrqaHlidQtA1yKECqWq7Q2DDcTOSUUbZTMNN59G9M1iZu6ypbUWTO4ARkUnjmyvsIH63
x0H0c3X2wbRiA7hG1pRMvDTBxJnJGM6kEgfkybdhqwiAhd/nv2NN2yijKS0DUoXrCEyhSmn/jEOG
9ntDjSzuf/O6YIMFNfEDzWcuMXO9tjEqxIOQ11jSJThQXvwLSHo1RfSeEg8gHYj12Q85SLFQQVLl
nCGVUzYvY/FNt/BxyyeokGpCd4BYvngvZ5BipCka7rURw9jNValeWuo9e3Y4Tarcee5nOTz7Z7N5
PuMl2FzjI08XUkTJoAxkzgHqV4iVhNT7UG43iIHah+YLO+9NrJYCR7bTEDc0CTEWWMeFgy9V38vv
qFyQGx+Rq6qFEWmteLnuZUThgYZLGBm50nKSkjeDt82WxUTjr/N7lgWfXoN84hNBGILmkpGw9zax
y1C5AyZeucsavOMJ1lnmPVLY9V1J1kJwIJ/4mafiwWH73mVrf3Q+5E7ap/07LViRdW67kq0MrTBS
iecaMth1lsJX9rcmCqGOKfcQrTW+PUnp1nrYF+DjaH8YL8x2ix2yvHk5xcfdx3vmKXYXSgAgz8Fu
2Klpeq/UO/F80jJkEOE9d7oKn+F3t7Vslcq+cWxQardE+Q0f12EgjvdM2Bw0GRh4UFY0eGXWaJIS
t85q7mBcoQkNgVmozSwcMBcTWSgND3aJaHrv8jVCyahCPRYrdbPTSqO1fYVjTeaO8bBkh4Uamk6B
cU6pysUOAeLBy5qSxvj3OtPAVgDR6mhOs58jVg1uFv9Geduzhu8kib1rQlps+edpFcrQcswBreSV
HK8wVxklgd4cR5IqkjoJH906TcplCJYELI9jRdTpcDvDthoHZC031b2KsIUYsAbLGui/mxKGvPEj
Pye/FLQWkS9Lek2yUkI+9uyE2+qpU3gRXGD2F90j2gOMQ2LRAiUKHOb/go/S1Y7vH3qGgInx0xN2
I38tYutMge6150GYRmKOXh1N4Gh0ifZybid4PXiZ8jxkMjS2tGFfxjxgAY5G6wTueQT1MoQMxaUw
lFLyGOGaHhSrk+7BW7Z0uFVUcmHGmlhc3QYX6BUtvS8haQA92az71/vn/aeiK7+s7V4zo+Vb5mNV
1o/UkAvUYAmfAjMs/X/y+UH0xVTWytZnM2fsyms4vRWZXJwxeA9nki7VenD+nHMawdG+i3IYX5mO
8H/1d4MSHtUsxpYiVhyJBocxa4YIbx4utrLrpzzeun+91jv3p/7xMDJzRbebjDoI/AI3I9Yy3W1u
4PWQHv2+SLlrUtPTVsvk4bMr1LXzwrIgz/uPwkLI6vQznTHJ79QUPpjFyNYderRJ0ZqzGNlmBSRT
ijp6K7yD1wXJvOPxpk9VXT8nJfLpMAEcc7dkr5ssqaqKSMg3aN1WDJlpiler1Q3nuy/Cx0ApmEBB
TTA3O9OcEwr00GdK0+L91klfRr8X+RfCGnEzKKrHiO3OsCaPmz8lhxVMA1REFqIVRHa0UaTfl9BB
o+to1uCu484PikwirfOUu6Oj8yF8E7K0U+YR1NgiplUIlEIdkI46ecgu84Iz7YxBnH7Llb6iyeYi
IlTha51cKsZkZngxYmLlQIJcsb2M4oNSRIIw24gw3vAOegu8RGxNvwKwbNwXp8LqlYvGiHfurJbY
G86VYYR3eeabRPp7+7UvVl6kkYFvJyC/3YzAu+ZE5R9/vZwTPp8Lsof4aBH6eY1MFzichGnm1AEl
EODBGzRFbZtvOdqhEsfGL8/VnoZcoi0Hy/AlqkLaps6+RG+JvLAvIg6OOxukBxQMzCj1sYGW3D7L
IlQHzkj2Na6F22oBUL6XmCGW5os2IUr8pf0uDXuGTN7UTSuZ5Sldh07XY4pb9Vd+zVE7mlia9+L2
9ykNV8g54wSTUIbXV9OUMlaOiw2wf23AeoyrXRefqflzJMR0L/763rVxWkraakOQ47tF7Tmn0dHd
lj7AFMMmuReBDYaoFk8ut08BULkrHP2GSd5Zs/UIzgflxbVQnXjEtG9ixboNhatExEn3uN1eOaB9
+eausY0D0OC7Aa28nA+Qzgi7pznmO5QV7c5uMnF5iUlUVCqoTBPxvaXwWLvJuvJbGdFbWlh0aQl7
bAB1Bz8DWWGK3t2mRnRFBEQnfzZeStGPrIPvHx9WY6PE29SM6DdIUix6YcAiGNJaG0lu1h28rga8
ym0Z7/8sizzxEJx0NzrW5Cmnz2KD6qKzlqVilQ6cPxp/am0ssF+0s7bAI16cX6JgFNIbtkazKYQn
tEnXq2c1i3Rg+MFkD1RrPes8ADZZ0RbIxqQQJ7ThHeBYzs/ImVJ5ZZ7txMQmgKoYzIh4swkZpbOP
tuW8Nz87p47sulmjvViOrxM6kBxNXCVL0YTDz8Nd/9qEngzNgwrEHL9zf+krVpKYkL+qoYbKU9WV
DDRZaLQEd+8qx3ghkwxJvTG373OnDnEwRXBsAbbLFR1WjYb7JpEJ31nOvfPPC0wT8x6BT9L3xZ9u
23EnKpAJrXFWklx5aDK8L0hEABKNu00QC3/jgX1WDE8S4+pteT1LvGg4Ixa4tA7v7GVrZUAKODYS
f1USfvHCf5pOuEemVmlMFNbSjdNZ8szWtIWD5490GA33zdr7yOtsLTPLDMJI6qHHof1sXr3bXvT+
kOSDqiRJkPnl53NeTecIZMbr6vwtXhmVkuu/JCC3fr2WhYWLvCLm/Bm62Ubchitq/Tz1ivQCzzJ5
/CkA5Y5iwSlIXNzjV3XGauqvj25vlMjHarVQ1pMWxUC/pkkTvGKRlRvagqYWmgHmgOOvAkBnQW4M
1pg7DmKBCXiWdnLxMjoBBVQ1r1Riemzu7cCXWv2sHFl5zzPIz0Aqt99IBEXWuXT57z6EJk+iTNBt
a0aVoIP9ORxrzDu0NqjgiJEWghTgyYqM+IZgy+SUxSZDNSEFekVET37pF6ZF0OJNknDTX86TLXFO
fDKJp1NClmsx9dcHhYcPrKrzJtakUXOt20XmB/6+IiQgA26uIEC6kE8zb6KFwvdK8Vgud7tsZMic
YEIQJVUDR1Y5axxaF8t36uam+NQi7Q8Pk0NZ+U7VKg+LlAH7z72sW9qKHTrbpUZ1zJ2ZplhZmP+A
9suPS4hPxLIQQcdve1J7y9AODKTpZTSHv6+Ka1eC+Xih/mSnLciIIQRRvD9XpjBfiD3+TNyfeSPy
gxn5k/+BpkkuHx7fl9gasaLkLfgSPWtccW/ZGHfzgBi22aNZjTJLoaW2fGikUNCuMH68d4MwhchP
c9twes+nr8N2pngl2URL/L5xOCepELWMNcsrzoFEz7f/onEeX3TIZI/DtWs2+K+9yk2eSOcuDFK+
xft1lBeokd0fofjs/nLPjQK0TYpM1JeMjureWj8Vs46PAGfneTY/ZDi5UAx0yfWq0ONsipK7+Znu
GShxuVl8K1W9IQXAse0HISMk1WOUdGGX+sk0ZpeYIsvTfZE06Xy270QnxZr8WSdoI+mxQyHz5/4H
KaVt541/xeO7y6QkT2ihzyxG1yYf5Wc0NbFsWu7MhGpXpuodHxVkwVu5h3769MrXjSYj0WjKzEg2
d9/jOWDzBELB/njOdStDc3vFTyzBQLAnPpL1NrunUvvkGH97D2PhXpNdrLqzgEEk60Lmqj3dpfNt
DKFJih7YfsVRWM16CKeAQ5Vcn/Mt2pDSvRGKSAOGW6mXee+7OE5iP5ZiFi00o0v2tdVwZTdWEiii
PWLnNBRMhRgC8CGF/ZItIu8AOJiCXD8tTTqIMQFC45XPZWLeaYaoCKF5cKJl6QZdak6S7EONpIKw
y1QJAcTYbmjPmFTrxYJhm6dg6Xc5wua5i4gaiIOLjpihDryZiiroGwuWxd6VcR7TBi9i7Z9pPUhc
HKuHomwHzFXJgfUiXS4nSSyCHPZAzHPJ99Vct6XQiXYUkSfWAjLaa1hfhAjZNtVPPxrIpl721Gob
e4OQ7T4CceNczLpjeV0jLZxZwJNKOKJE7IdA9ruf91YZREseAtUgHSQ52irX6471cigIftd3OCoc
L6yveUBWFowgED/ZsiJo5xAf77LX3Dd151wYjMyRgE5SE84MWsoHp5a8faSYOmYVI76PwltOvpq1
VmYmhhvXT0sDtjt4iVMnRubpX4xWMoCgtTYCF/EzqWn1rxBgVkH5JJ/8LjEFCioeCJGzbyGBEk08
QSEwAbo0M7A6zy8AzHfhYMJlLVorPadyGr4qhaeJVwiTUSwGnD3Ekzr0U788jIv6fsbK2MOqJTKi
fXThdn5LN18LmiY1z7H4+QRtrZApkMlQQSkJpCrIybx8jpvHy3ypNSv3izDZk9wG9bEclsJ9CpUb
L3aIchs7JBHCkEB6xHLOQq/fFp/ZsiNWaw1cDgCtebasUjUvhEGm06JyrSr+FT0T7lmTfQIacyAn
ROT/0bgw2j8fOB3NSn7iAoo5UtAhNEIteitSP87Xrvd4IZK07v1DxqbvyNNT/+QHhrHuzTKHsSA4
Nc4xwkyQgu02NsrHNpquqGwPGItUXsXrvvwLe25MvqBYUypMVv3d/SRTTRKlMg3v/6H7PQDccp84
8U6mOytvgsKifRGIgy6IM2bNqfhCDjChOpVT8ZvWZ/r5hDLLTGaSQ3CeU8pbzq5trD7o2aaLdd1G
6Y8LW2hpncYiAmF+UNGJxHz8U4ry6S5dMQ2OcEDZpB5DtJhteKDMfqhWy3+YF8D/sznW3HU9AArO
iKfH98ihgiiZRe56X7nezZhxqc5vldsCwF29bItcQwfQ63QOQhcLTH/eQh4bvuzJbu/FENzZmGWD
1slLeb/fxcSA86qPTOsJ6+KwiAEpdgv0gBuwl9gh8mAenI79ZAQnHYYjj6oZO3eLUtpYghvxepCe
yMAo9fBEyKTFPKT4RY+DTtzr1esrOy/QzeBOsxSjRdzZe2ufudarVuoI1ADFYEFKPE7+CKVaC/C/
DXP/QzExWFbKB+h5/Xai2vGwo1ZKLN3iHze90Gt7dNLZQJOSqYC/wbUa0pWehEkHmBPE2KyDDM/U
447NBR5pZlJJCPYREcrXVqOlP0Fm33JCJzb/MDZcS8+mTmEt6KOWYGDvGr5iYiRJ/OJQPEaX2UNm
BZrVgJmg4jMHftPM0WLV97UyIIanTqu9+0YccUOhc9r0UIMJ5SSPY2KvxA+EpYi7O8juzfEbkMSm
DPcRggFjsfdrmcD7atgEeH37Co+SCz1q5uRacnNigEk/af7gBX3KeD2cMTDVGxXWeqXyvOsyAm8n
TtxvLeo8O0La1YweqaoEFyhlHfTu/70GGrU5QRAhD7UnRgIvjWNSEIW2+dDZ9Vn+oQh9j6ztfTdF
kd/kFU8Tc8rHtM39jgCbKO8qrEwI6aa1VgXyts1gS4vQ2MATXGarRAY/FEgz8hw7T+DcJCIutIjm
D26kS0MzWZXiYY/W9pnOoWWCaMOdH+iiivq1w3VD62/O3SNb1RIWyiFTKFHSR3bam2hggnkSmMSa
VjxooZ1zqF/q9U80keqboCyhc9wGI/357FvK76PZgtuQkhmaTR8ncO/YEszpSrRObDoHKJldwpRS
daIEqILJft7IsdamO+YD0ikghNQYBHo/JotIIQ4WYJ7nX1kffdVx6l4Z9vG78/LYaHX0bwDWhUlU
LaTdmQq6+W+poZjWG8LVfqIy6/dQmpuOT4Vn9wb2saAEPugKfS2TKkVsuU68IVNzg//Xj+D+L96X
B/Ny7G/71yWtxh3QJUodvV75Ri5KNZfL3qxzst6hiWwaiGQ62xep03pdIZTuGaj7C0VGsoI+4sNW
E+ieLXlg5+UmlVVm7lBzSkMfml46AKuvqArlv41rE4oDznvvJmzgh5WKMHFioSaykd5MgAu4nr0o
ZZWC9w0FLE/1NNtY/Ef4XrRZZQOgskTteNCxfp3sjqt7X8tHNv4BB1oHx/2rNjxiZdgaF/G3qKYp
x/zPwEjpPYhgpdNoWjSjuFLiX8UrIPESvkCeV4D6NsIDAitsXGnb3yu90BqoPi4aSHip4O/9P+nf
YReGEluHwrkMfvIOCxh0OaIbVOT6u6BHiNuo7i26BIfedHER4m7lg+xZ8ebM8Boo+z815D0OulD7
d2dGHuK3otCNWtPlEJJo8br2+IqpglmZ8TG/S31SCuc9AcVMpVPHk6mZt/QulqVswWVSRHk+qCTT
B31QjXkS71WWPqNfoGWAaULv0F+W5SWwDqprvCTjIs5iCKTftxLB7B/dxlsS54mAhUJDiUYExRHM
Rf6yw3oEP0k6F1nnaE9G7ULcBJ2nBj6+8niT4qXXIbU8pI6kR5WIvydeC7nfY2f/VY2yJ/GI78Hd
8PzKUZOlu+97GmtohabH+mLWDE4CN/rFSTil6liUYYeismkApUPM+we1hDRBrYnvtBvz4Rxu9SvE
WzoD1Laj4k974hjZgaH78CnIxqZQVxNqz8URlTbzb0Ws+vHUNAnxhjbYGNvGfDmv0wsBz7AveIzA
fLsEbzsIsjCk029m/5DK0S1qh8ckzM2qySuFBrsP977S0EUu9ZpNh1YC5j8xpFWHYDjY2AvcXthQ
QTgkIh/4uZKLSsRrqVVAyfbLW9BVd7YSsTMd5eEZkpi2nLGddZJoJKeRudAvg+uDAhiBRx4Ve82C
mD1Wnl7zmaReXYhs26m+1v/1+/WlJHpdKlAAk9n/eFwFmyBo8CBg3BB4GVcTdn9Ryzpmdj5V2drk
AFuB4Y/2KGpEsZenOw4Z8Ecx1YyNmeCxlFUjWorIYtthTMsc/GAsj0T7FhWAsgqS9gpCpRavAmAg
eUcXxNWzXZPAC/KYz/WFp+WHeu8YGm0IdFE1dNkFcpY3EvNL471xN5AwKnEn8KnbD8tDdpyxdU61
dNBPFdsv/g1lpDMSzJO3fdDrLRp0wkTvKEv0gs7f2G6i8UvqTWrD4qQPtur7sRhMSBd2GyQMT2Bp
Zhxc1tNce26MXWROn35/i94/ECd6fRfqOMALiyoiBWv4rA5dbQpKwrraf54/J6FO0liColn7lI9b
cqlDZAnxsuKsaGApvI5U1Vkmx2yAMjYAxV0ixE3g6acILMDWw3A30OWWOEK+xk4o2s6O804hcHqx
Htkv45PrTrcKSZVvqAsamEf8XMFveO+8rry4Tm5x3GlDiv8JtZgLQcbgGXuFOai8Fe3vaw0MrWBl
xXK3NeC1ijMF/1DzrKw4aUL0IOaYdqMr3ldQxJy9OQQMVIXBS/lItz4Bk24CjF67rQhLUwyPelhq
cfoWHEMuaSO/mi9RZoWnnhEX9JYjQ7mA4vAG43CAHfft7O+3VFKpLR6FIPAaezRr7bTAv2qI6pwO
H5PCasaKIPzfKyac5jFiWtOdkljWuNy5WlWeO1IDqHv/pWS36AIE85OC4wsdKi+ZOdwk44+uxudm
qC5N1Fwd81g48qqbNw9O1GreDe7u8mbVss8C4UJqlenDX1EZBUEwnSgc0X6AfVsh2ki7mzlli7z6
TgqD2htWPHEOv4kSBnqSZAEEKZeQ/u4KDow7RB1juVLtwmYoUK4dd9soqvLZIXj66dAEbDSctfry
45bp8Tz3e8Q2MgIK8nGqgJRQBBbXW0c+irG/oIooXDudfp/JAVidy5xpjQj6E1Ft+bLUyYURa89n
Qx1mlFugJ+bZpXK0RY9prIVcJazw/bvG6YWK1m+VOn3Jbf1E8x4weBeoN2cwB0yJOea5FZvXhlMA
ejK5KHHm0Yq0AouDnmBg2RnsphWIUWBhyGDqcssTpDkA7pIYpN6IcK6uhnM3DTHwqYhGjMfLOZ7A
YX9DUiCMjCS93p9QR0qcn0BZ6ECifsH9latQwKtBI1ZdUdgEJBy6sYEnhCiPQlPLRW/X0ftfye/S
kVm4wDhUvbrvpJJ/tM/TbL0NFI7auUG7ca8I8y60cU8Rc0Je3u23KZpreXTJDYNg3WNOUWDhvnbS
ptSJ/CUfBHglSTlJacqEYWaxAb3zCIr41PkbhzDOLJ5ivzW+wwZb0f4B8U3aoyKxkeVNJHDGwvzb
O3WrgwZlpqcLlKTSDi2asG2S/+X13s4goh+MrfCXJp7XmXOoHCBAeOWYQgbOq3ImYizpBoiUeU2x
3oknNs0KQAWRZ9POyQvhwi9Vp0ryUUPMcyT8/mmzgj8WmBfeXiaWb9f5WCsObWp7XInnGd5OYq1H
0vEeRLaDe6+h5Z1vdCa0LuTyzlIUxuvlQ/UXIF4WjREwoBFCuEHp9h6I62lWoXroZwNBfivE76lS
o94oGYUKdE3/K7RreZ+Nu9o+aUw+Jy2Mo8smMT3GIQRCuVCnElxDuBDIO92rCidLam/JsEUZ2Vn/
mjPO9K6nMRDqIsvtl0JF7G3/a5kTM3suVS3tJFYY+EIVMLnkcUK9zeH3R+Q/bdcAjKvLbdhQNPcb
sqC0Xo7QZtHLcEE1sulBTMsz5eNBdbdFx3edCE2TZaXJ/MTeIF6ujtPQi9SezH0D6vlzY+9mOHiL
l7d21Uw/sZfh9F4ibSfHG/Z4kNr0UlddfzEvgiokXsdNYSUJVQ80SAbn84nFrROsK6TvwTYr5X1l
tNAmoqfZGlRu5Eonsu4zK4iLiG73pHREDEELkozA2xxn0Ne9eda0UFk+Tb85/A+jTYwdWiZUfhmZ
3AseGlPMDl0pqi08hl0+W9mwg6y03VQyISm1M1p+tBs9hwgt9XDCAkGolEZYphw0IkkF4w7zrBQr
h/kX8OAJGXoOYDk1CQ9s9oUgJTX5dTYm67YMLIInIBpCrWB58xY0iqI4uu+oDxv5jN2anPZx3u+V
tQj/NlGo4g9OQKXCBeyRGOmWzpgmSEqB/KRIsocIjepYG0Vr3Aklfc4G4swbKH2R8cgP0GnUM6ZW
SZa0PGu2BOH/4YDlJu/xM+sED9Kj9sPAGy+Jpx2FGi6gUah6Yznaf0ZKKuYeI8Ns+ygc7aDfS+/Z
eHAWSedgwFGuMFURr2ddBi+nSYCEOI/69+Q+681HrTgLsAstToX4DKS4EhKzZnMFYsXyhhZbYO8W
n2miUWvwSWKOLQEib99RwJ0Km99kbOTQNskN55840d/I6Z2Bqpa34Wzs+ZjhgKEKeGR/a3mNuGmc
qjAnzF7sgp/OaNbhSwotmYAW9MrRJkwq7QElqv/Gk51KZCHAhEd/w9uQw+UusUHqTjxMd3dfPkV7
xhq68Mw420lt//3RgolMjTzeuTrx06eRYjIhvZlSWAn5jqiYFYYpWWGNXyGehByavAWhDStLP02O
e7IoT+iGEjlHKfaHClIfJyx3P4X9JMqjKWI/op2KQuCfP6VpGr4pywnvN6xQX0B7QLX/sqbCmArC
8rAkX2YeeXjoW09FPJmPOfkOPgc3bLgv1O16peiV5dSWIAEN0x03RTZCEf0qgNzfzgbC6wLANRDs
1+6qPBPmXi+t6UclEOvu4IipmrqwvgVA+hNzElzQhi63amEAJmGx5G0zMsyafcu7TNXM9YUejt7I
59wSNE/tZqlziM67UlgcYNxUHK/WKsMsJjMcqmzO14vkg8y3r5is8P74wfuZGxiGM5d0lXF4Dpl+
DqXuXG6t4Qsy03i4pGIi9zG0eDeSUQl9P+DAmJjUkM7FZmQk72ws1MsMRXCojqD4Hnj7gWA3hoZu
HPId1jL699r3ZGECUK+467Hr10jHK7jSPAuqo3n9yZMoTk6VZWFEdPFWhPQ0VZd1iRodLwwXykIr
WculN/SdOQf93VWzgLkYN4E6sTqC+TfP0xlNx+qKJogP7YNinDJLOY7tz1lvMZuNmScwrCB1HZJZ
P4OFxdxgY2hcN0lvJGX3JgiCMXwRXLtAOV7kEK3EKi9T1xvKTVmrlPckrNt/a/Yn+MaOoJeSQl6V
1NVlNVA012AvKO4XL86wi7AZoW8s1yxvy3yxiz7P+mLnyOefNCn2zrY7mpKHc6MN+V9XJ6sKhJfc
5PLQ5E1czL2POzOkWzwiwLIp3YiYIlk/J4VZEXXu1fbeamzz16kvaXQfSEa6EcEhQBJm1mD/lOCq
WNqRTgONKkKtH1vpiVRO1AKGnjWNS1ImhrzcNSmqltT7Y2Ho4YpAbDhb7SMaOwodbRdP5h1M6dJf
X6wB0DAmu+MQrhWw4rI5XThoQRn3/bgTg5mEqvACjY2dtB8iGANUP07NOL/N74k58XInaHYTkPSa
fROBO+ycDdZEK0TvPOKkRnfoH0pTnbaXtnVhKJYLFshsXhT3/423m00bBgdEvFAGID40U1inI0DT
89r1NZdXsjJYCLyq4iEk6JVXYk+fKYh/UCCyoYeIS81eIOh2d3/AKFmwWfgET8tLHqk+Qr+EsmcK
QX11ve0Ydd5yy/j4XCRcTt4GK0cxwO+c8r2DkdRhs3xGFKt5hHcoWaoNGOAtU9MOp7hp1Bkkm/Co
OB1PH1GMoHUtX18bKLDJ9wzpPz/iXGGjqDhhQ0vBZQj91I4hDKLfMvTDqSBkqAnZPICE7XPjg5lM
U3gzCmhC+1R14HoFr8uGeezvIJzQYrTnLuuA29fVwwGXsfvNJVr6J9ToTP0R2VYWG2PxJWjRrJhF
LgKt1Rtb4Mmsfwv68biTbCwrioSo4WUxwabnprw9S2rxT99pInajiaZ99A+mfgFPSbrPnnZIF70t
2vUkfrTBkOEboQJkiFFomvP8qHTbSveWPStIrRLc9dsH25pUeD87AcrpcUG8hByTRDEmvqV42/FZ
wLkzKz87881uW+LoRwWcmJChwC0XWY+vl45BqBLcfh0rnMFzTU2INEb6Y9Gu0xp4LAHTqTCCFWph
SoKprO57XY9cxSXt26v0JO9aJKhwE9E+//FgvVNxNCih5tiB3CqA64S/mgojTetHJ+/ZNOmQAvQA
K1Cbtso+amQOxD0AtvyuPfC6Z3N2ME2c7FYYaX1HHRZ/kbMcR44CQtoeVJ/hHEWp7FAtev18X50i
W86DQrXxccAXCSwXBRzlyPV2HluAPs+w/QfZAyOH2ABM5G9LPOfTHXGeUJArMPTGduF4bsrpcCf9
fs5uxFb3RYLFPxCl3Dr8mv3WR+4+FA8DJlr8v2z53oI/mCDvFhxWVWnL8DKYiTAwH4rBdle1QumV
IgcChPFtb+4VhNX+BwzKhlAXgnfxlXV6LRZ99h0GkKEagL3HLSRNSfJMp5kNBfJLvHBxUHlTTEyT
JYsoEkYZNcfEBJwO30tfBZi42rf1ASUSS1yXg0GtNCOFUaJ7yh/KRKkV3b95t31KDJYLkzzA6x9p
QrGFV1VYu/kgy35mjg0KsBjjV9SIcjf4b/ZFjCXfdewDvUbJNbVTPelfCg07WkuA7N6DC31hACF1
CS0vdRSMf3g+8I6TajcRZADklmnqd2NyQvoK9AExZfRhqeLdlrX4KdJYkr1BGS7SYMd7NJTVCj0h
dUFzkIwldSNXkZ0qBmZ45ZFaTCx4P0rqjvJoO3kQdbHe/S9JV0ITp7ZTOC5cBl5kZHsI0mR6YKNY
USt1L0bekuQW4Zz5LIEITIrzOf7V5NapI9nwUp+m3BgAnYP9/AateMaZDhfUrXdBycz+nebYKfnb
y3zm08F3MZnlyqplrzp6Yw/EV367GrWu9S+/RQax4Xe1ZJEUgcnqmLWE4+HNurr0P9xngVISsjFt
RskD+jjDlDKvQCIBgAeDxw8EyPt278dSK9YmIvtJH0bQz8i3Cn2ht4IcFw/lIhdHQqZgy7+z5eKV
y+quA0Ngwp4SkJ7zVk7mE/mhhGItLVPORUeyAI4DgvFmYgnkkI+mEI7cAiNzw53pPChPrtE6C2RS
t0ebo0scnjszLxvkA1v0Mwezs+2t8uZTQUFkBRU6OGCbr3jph+UebvpmBy0pyEZXvVqe5vbA8U9x
uJZVzfX0umcTwOUXXstQTPMcQ1b95Ha3ov1jQOOb8NFk6Y2kwbiD6oB8ZFoUc9hnVTvHGerxTXaZ
ieT3S9gDgy0K2rvcy3pMJdddj8f7YK0rN6la5JkjsuRdHsauzrazXQTFVdxG14WJGipy6ZLR21sz
QALKJKfuJdKnem68Qo9/XRNC287XcYvqsJUcbfw8Nl8fOzOr98+CcMypHq12cDj2stW9m3KcFyyt
p1OI995THBMWXyhRU8/VkJ96AS3ypfp5FYluhh09ucQFqctod/RR9D/2CNOn66GdT9AivLEGXtja
koET03WTWouxOWtAjSMkehAHYKtg8gM+CoS7irROoncogZ1Wc2+MPW1/8UXQ4+FmYtHfOumepQtY
O/PEH41qjs8pIl2dNmkpqMZtofBHtWHE6nJVOYOqgZkQV9wvQX6Y5tR1ClqD0FIz4xJcmOS3TtAX
JfNj9p1Wq93PAGlfn3zd/64IbfTb5rsM+awznyZ0FWjh780HG/00D8SnY57JvohA2elb9/IiksKC
an7pBBo99k5G1+DIGyIiSdkYOd+5Odod+6EbqlBLaRl3C0TYeiqLmxTNapwZV54DGAkTOVdjeB6y
y0RQW6pm1hDRf29E70igjHkVPttYX7WEoI8/OiYNnyC0ak2Ti1sYEr7tCmnneNuJKuKe45FlMqPa
FsoIUEWvPuEYyNppEiXti11qdHIQ2QK+0GAzMVGqY4afFyMiAVbAvgI/c38QDgSmZ1VECp3a34fq
koZbVjdw3j83OlzA2z9PZhsYYKHnuRxJIKIA6S4+lYmkQbP/20NQ+8D74eklau8KWuRTeDT2mVs1
4/VCi5JJ+I4LGkaOhtCLEwHAFqErEX8q0oFEJwI3061BWhZgp564FyB/8pP+HY37aoHbbhoJxHKo
WU72IVentBvz5ee5OD/hSZH9tjC439fRto/U638OjI3hDBkkgm80vmvdjhaSNZagCibNzQzgY3r5
cob0HF1hvam/IQQEjDGc8gfCyhXTnEwyuVmRLl1YfqtzeIGTqwPCf0ojuJNqNTJdrsFTfo4Kt6lG
szyGpU0MDLufMCeDkBSSCu3ozSlXqKWcG0qbiEHnFDWXllMr5qRdzdkKUfU85e7QigNakfpy5aFM
2faEU1aQfHvOyW375REjfta2cD/iYpDJDDP9uj40nGS7vq+KB2Qy6ADZCn3JoFWQLBpL+zmhjDDP
qOaYIbCTWHzAv9hVcBV0UXVTxfq+qIETc3eFE5dmZF+soxlky4iD3wAQExAqfJAGcdDKT82o0qIF
FG7kncpujURI8QOKt3FhgYhfMDNZzYtNwUtdoZV4TDikSlUxx7n7ScQVn3ze+pYoAmfGC2wABzMf
V5spEhhHMhk+rafAFVrhnV9KE8Gl8VMgekKpdgPCPy8p74OaeLaQcimXFxbNTiOyrNm9uuvUqdd9
xhEtQXGOaAUcdgmKlPrLbvmWsqmBdYDV5426p47nfINOBUeofpF16TsYgmzdkY38b3KYtDH3io2a
tsA1v7O9N9qzuZvvK1wIRxKiL6NXCv09zJK9hUv0cCZbBwfE/iCjTPqi2IT/h3L7zh0mW8KZidxy
mdDb9naHesLxE7e0kZaKl8SNuorp1R7hgzmKg9UsNqGl5hXiG/mOcUjaqGFukwyF621oQjYPaiqq
loNPVjDq2El84YWY6/24egwa2x1mG1HlsiTrJlRo7MKO8NpfJ7CsqOWsV4ugIArWycI6bJVARKDG
e2UuOuZnAOMq4lHbShAoLe5X67PfkAM0JbRZpK/fMiluFxuYRE2g0bojh0oMuNBpxES5PDninwe0
m3l1r4ZJzzImePCo3wfQDfKyLGuMHuA26M2bdVCn0ZVdMayGt1WXEjzTsO0IXzl8GQjzsWF3A5IP
HTg4TY8uf3t+kuvl5pfFAf+sk7yNMOVgvyN3/BZ2oE199/4qR0wJwxHzp7Qkjl72AWZ4+s4pBpef
UIpUx66vfq0A3peQpR8QxzLy5Z5lkSR3IT0IAxyKKNai5k5XrhdVmDidjj5R+jyI0rEiLm1F1D7H
7lmY9ZJqyRir2u5Ykc9CqyJPe4y8LFZee4MZ/8JIjiE6du7vfap/WzmVBa6kY9vHxIso7OTfg0Kr
dcw5lsNji37pkjh5mUvWVVMbOghADV+AGdMN6XJU5w2UIigohISXwSJMdJw4v/3258SY3IEiotg3
1qJe8hfJ19Yaqu8wOAVzMmhfYd94j+ZVi8Nwvv5H5PKXyB0RqMpwGWSzJyjixYZV3O4hADB/kECs
6WUH2cjORnKKbJmjBSJdka5CWNlPBgH9/N+HFRTCVxNqZTrjgv0MAbdazi5b+JT7kJK7/8LzEEhu
91vvHIPfqV2aRt1qnz24/128NbdPr41EikgaYDREgU7hW8SEHcp1nkBHLgcUIsRC5lmHcmHR9gVy
W5183d8fVKUYP2ofxAya7PmmOO1VLc/AsPfDuCFynb+46RP0seem2w4QaWqf3gGS29vxap2Crus7
d/AcUM4zl32NOB3mKvSQwmQ/0/V8k8yDTChetwbYajxlxQVWr7aJhstlodKjKJVzL4Y9oA9VwToK
IAmDsfe5rtLuWazLmQ0YQSBLSHXCTIrBtmnOk6JRhgObcKxHlZOv2BOfbvTsKna1Oo/HfjEqVuOx
z2c0UhDdL/4W/U18+ZckYztg853Z6uxaX1a0JMaRr8Lj4Vdw7BXy7rpIKxWbhS4vd0oKws1jmDuf
phiU719DBPGBjmVNYY6bOM9VwLV5jE07ECKRP0LLPSkh5DdXju/I/8pGYHfW34LyWw7HVXpSkOkB
dkTwiYVZY5KQPJIda2GmbMqbgSYCn2aDIFNaBAAUkKALBUoyzGj+JCkVV7ow/i94cp0Mz/sGdc2s
Do7laspSna/jrfnYD3vnRGRcAROmibzYahAvDSoumLZHQNqyG76GFsS0YIQ2CM+YbLN9HIwCNNpp
Lgv6Di+XU+JgmDudYfS4q3rF/e/WYIEJ5NPtLA/H6DiMfZNwEsdd1bKT70XVG9laCtLQ3dNnTrUb
GsMY6pr8+noRNMbkXUE87/c1MXeHqzC7dSsr5ldLAUefdxXo8+HcwCLspbQqE/GRsQwL0StA+BgY
WUGZff4jXXa7s/AXeXbastxLB1zBjKqUw5nPt+YSBMYK8qXOEMOtqeJMPa/iszvi0xwck8f55VU8
LolSdGU9IHO7dOgvquruLTyiCCExgMjLPempWfYIDNPS76MglrQ+S4OLOJmTTTo+ynq5MahfUhdk
PPHWnkhPoHmQdI/2s6QNPRUHxD8GMqXctq3xrNTfJPjOuf3t7CuI+0W5FHBlwHkOJuUUzCbul5p5
r2XOnMwxDkHPEBvUbRhLdKU8FQvqRMI8YsB/GnAPGz9zux9HZsmt8YTmf1R9BsWKletVRn2+CSMr
mqkCH1/B6tY67ZyX+d3DUb7JJtF5JIEKkeiduUDl/dJzTBZtawLxX5RgikzmgwRkQr98BBA03mko
/lKVNaFjehZ7aOQmG9DGxj1oEUVWQiuMbY3D4CMEyLEAY0PJdX8TPFahn1QgsMEDBz49+ZPaqVco
Q8CyvYjZrc9IZMdJ/nEG1sP/m+x73s1Uuf4LO9y2ZgbMjE/trUNALTgTp/A8l+oOFULzGl8/ukwa
sNkLM5dEvXNtzrqzcnl9YcS7TudK3eHKKiD/h5CyvUyLAmCWtsgGEu3JOUhNx/qfqMzZRx82KZ8z
tBGwm2k9kWc1LSkPioZesxiSE0ywO9+oGmd3nsvV0XkLP1dABM1AhnTnkVDcM7/p+MMBjSsBUH54
UtAysiMuYIq7dcXt+8htKGnP7wNre52SY6YvQ3aLH56efDAZqqnpJ/MZ2VxR4sZ6297purSNRa/u
YTWTzZPZKUs/cJhsPsFe1nS/hIjNvIAxyBLWNKNwUOs/E4jdAqkpkDtv7vn8HDlOcTTYhuVPbbzL
+l49gOZDS9Kv1FFJtr3hPbVQkmoe1IOLOGdrmWtaVPx1CJf/yBaJ4EqOiYX3iwqAnG70HWZkxICs
ep7842Jp8U0ZsRMORM4Yf0h0lxzO7grOwyPn4ToLlOWnieP7VQYlt0e0kUGfj0Ywkqd9UG8AMoX1
XMK8FQVOWPjN8/LX6f0N4LUV06KSzVsY/BmdytE8OKYtpD7KcnQvE/Q0CYmew/aEZUMmXkNyFkqp
CYjVCrh7UNA/U0VTbHXaIiCATYntLn12VLPeshKUF59b+tkecyy9v3MC92IJRLdCfsA5PRP4M924
Imip+vPXj0KdGvIF5dnrdcWjV0Ml5bx9U3fdgiXoFQq6yjwbtsyOVY/SWLSWO5+3RqH3Y696pYS0
i+XMaXAr7EXCyice8jAVtqQqTg5BRHyttwo9rbLCKmlPNcPGOkZuGbuhC1N/Ier2xlLgqgyk5PwI
3nq/FlpT2hniM49VyCBAyA/YsM+wDLoOI5Bl2WnZcyX9hjuASEhnehu4m7cS47uNJIqtpreuFV+Z
F2GYA56+NTkfw505QUXbTgCqKevH5FKoQm7sqWPYrDDaERA1aI3GegyLR7QCzc+ICDigUxgzylr4
T2KkIXskZfxyy55kyOqhDdmWUMmTz+H6Q8NskwyDrY7WqUKYelp7eKK92yxcTS/WkiYUcpPGRe6f
tCyXD1CnaM7gqOT2LLsGeGIMiSej/H+bzMBw618mBbQBdaX2W4haXCJig/z6AypyKPKmOR7klzBq
tFUt/pHYGMGeBI7b1W0QJyFqPlpBCdQzVbFNNn2/0eMrRqKPREpV6lNdYJZ2itiKG0tQ4KhJ6avT
dZcYyZg81TgbHst3nATi9ddzIlZpivU0h4YR+lHWs9CHWmwxi+XjgKdubjhrt6dp+w3FfwkAf/d6
5ttlOAo2wmzbYIrXxBYEBPolXcibVrlqNcoTBcqy9Aem1zFjGuvnvghnvvxc/LROt8A+5KpD67wR
sZPjHEVAQFIn6MwjipdRlyRLD6hQafgH6VnXm5q3vk0ak/3jf82Rht4nQgJIiP4qPtnqe62WaQzR
KO7CsARk7tqBliFvfHVASHx+NFa/gJ/13iJsyzX+NnAS95Z824nH4djK/rm6lKrReGwhm3A91ouq
HHVokCahnU0SmU/4f+4PMMmlaTMikEAYLTycqvo1ZAm8KxgkB67KpnDEsNlCX2p14wt1N9CutHVS
ifQzEPEEUWY/A+q2TD+jZsGZURyZAfWqdI7Mo2E/2Ke3Y23TYL1rrAeYipnWzWVTezGqXkVQOskS
ZNKYJh50+Dhpjer1Z6wWSZ7iYL0CQXLaI6KNM/1nBNgt+Fsqhkj/IRzalCRkuDjNl7O+5L5OEuau
iOAnsqZO33Nu+YL6BlleAbBXnDl3YK+DFzo7J5sKcJCDQeHnqbRKXtaXr2NBSifFbe2YrGjNHyEy
6XfXtfw+y1pr6ASgdpx4uTjh27iLGDIHkBtL+ne71CQW5/OHXwNWj/DTpj/ciwBcxIhB0rNOGLOC
4A+CcNzcfDQFbYKwvKMXSatpjtCBpywtCG5iW+WK13zwfqqamRtTcE4eYZGU7Po7/mUaXczEfWK3
qeUEYEq802C2KHSYQUqQBeOLq5fDJfrALaueLaWLBR19iUyghFEguXnX4ouNdO8c6d7h53w7Mrg4
QOvW4D8QBIeWaJlZd6ksAlSrw7fsdCiQopRCDaruLbZoK0zz4vSyWDzapEeSg2WJssp3XQWbKs92
zaESHSsDMBbnH3oWBCUBtJsBHPUNGizDyVPRnu1iNy2Sh++DPStdPFn5/IKsyC8CcpCvMqbsXIzV
xejN8lxsjE95woZw0tPbWi/M4jZ52zDgi8NhGHmuJlttaz5+K0U7o7yf40DdfCHnoSXGQnTVKAWi
LuDmpSPtKWDd9vrW6CyXGDZh4I1yE5hxhZwgudMkHHOqveWXYhMnBUpB5aY9rrlNOU1IrUI9Kr6Y
gsgaLFxEgtrptRQj7ySgLGDSfB565ejha8ocMfsDOBL2UIpTAM0WXL+VtgG3ou0w12B9IcwCbbGa
hGyJYpZIGFd2/VPovu/QyqrURnuwwf0xVy65oSiVYnBi7NnGXlFEFiitDDU+dHCplYSZd+/k2t3C
ubNqs8p7EjKTjZrcv5xPXjhPboUQL57wfERl0+oE0CoV/4Qer4ieavb92Ip/lokUms8uIBwaoXBu
PzOIMJQe/iVTMEOWV8sEkffyIaj0ImeDvtd3mfte5BLktY3ZcpUsCXFwelIGL8foA4nNPg16aE6Y
jsQQMtF9hrXuXXvKxDxh5u55AjBjDU5ryBh21+Akaep+HieGjsDgUqTTRFHSSno2WU3rqjTAskQA
QbbDxFPv+q03PV4J9ZqorsxAqGA+nf3J7xQgK+byWTKXoDxWfb3/HdED+0/umtwgvIl4zT26tx4o
BnFlOLJ+7V4oepThf1Eeh5B4v5AtWFOTT7lc/bPSrW3Fc1QuXIdCHcAX3HXCMfxrjhQEQ/BTYCRn
9oV0qoKKvBDjYMpVbe6dtxYlUNwL89zwSizsL3IAES9OC+Uk2i6qEXqbA8IG9KAYhmywLa5hohT7
4ZAVNttTm/mUkYAPwSxkNIqqzrGQyyEUAqEcXbT79l85K6Eix3vje+joM7YF1uZeEEYuywakxWj/
GAu2ybrGwDKxHk3HCrdQq1t0nwZdXdAPz0eIx9uQ9vIOnf0wZI2OlFTFU4QcE+VATvZ8xTgOYu3J
Ny97qW71IXBvAFC+8wK+ALu5m67VfTPeGEMd/Rzfq0LDWqn2t7GRe1TzP1kVC30GKomKPpQPdqzn
anLcVXVWIFOhi7ashG/COEEyK94vfsp2UmnYoaE5sSR5yNQsPm3+bm7Ut/idkVy07U7tQeLnj4mv
CF47U7a8SMJgnSc4o+lypcXWiH7/CQRP0CVRMmnp0iNxWoy8nToiEolQXtUNoE3qf8bdczbme8LD
q9jYo1SFK4+SnfLVpKQIKmcY8iLPDzP1cg/7J2+vooOSOqYF06cTv8SoH6t14aaTi8yithO1rldG
HGE48Gf+mz0lEcNM/AmUAGjieilTD+Nag0wcN4cB+eh9FNw1SOkqsEIkUfI+WgvxPj8VL6qGzLLk
MoqQkguYLuEUpXWPNa5YiwH+nQw7+6C6tlaMod2bf3l7p4CeBbrSDhPvNiarjbHqQwjIWGH7zHqV
nLWqDiGES1hMsx3ZOWh5fJRKLc7fw8ImA8r6e+K8ADqmD7uLlNw65OSJK/ri/cjqUi9Zbk8gbCNe
dG/Lo9aOriDQPGHOVAhihAEfDXJ6cfLIr3AN8TezydFb+ogHwZOZKC8c6VR3DZghUXDUFzbZoJ/7
Jinw5xPIZWxBq8tXS2ijRD8jYPU17bCMXeD/452sQh5TbHXrH/2k5ddGIn1MUaAygMlKP77YjlIr
L/QQ6SSz1iZqFYwE3M4N5NzUjZyzcIJK2v5CBS+0JyI3l4P5NafGeVzUpj8DvujxrIzmccOB2muR
1FZhtWD1bVcMVveEqLx27nbQu4Y4E8rk2mDnVTXJIaKnbftN2fhXOKkhYLVcux3yWmmzjEez2kOF
bnzBM7ZfRZ7GCT0hWX1/KJNefvohkD6FEBlTbad+mQH8wWGsJjyn9qSnqN/HrLRDxX3G14j3TWKI
1HD3U4ZG6e48tokUK+1FpIhYXsRcPraU4FW9OKHs61VXFaUFapvimQTOeDKcmLzL5+2Kmt4zQb2Y
Q+rXZETQaFJZssdaCt22qfINrhdYp9pwbQGzSrC98m18beH5vw8j/4+4Sg8HnOwR26w6ovuJAIi+
pp5nPihxPy87WJypVXAEpTnK+wqHdO3YgmMp1hda+jhfulsvZZnrMud880Wun4JQdAspg8xw/Jxm
KaUiW3tj7ig4q/MXe0aRfAWDZgmgFrUsPiJnnKs0epa3fUl9glIQiXMkpL73ztT4MEjaRvCoPQyd
Gm2aCCnRQFm0heAVUKDZ3L4jHCTDQS0amZSNMEJOeqPocR679KRXNJatfYvHNg7SqLfH9VyH+9YX
t0f1nTGvctcPipLVsyP+OjxZBXCKKYawnS3lt2X7m+Er4TKpjYaxbBexVz6VyHvWeRF2COvJPHHY
J0kqU5G029PaphicuGtXiLe68Qirno0Up7Otl8GLXnPI70EB/knfRS7TG66iRvH5pXmMeuc6R7DR
IQzOrdwVArETYuUF4947lpa/sfaEjEJlUiw7mdvU1J/qPrqzKh/DeF/1mephmnHJ1vA/0aZD+G9Q
MhyeY4Eqqg2IAQN5fpDq9aYlJ+sFu9iMKRFX5qwvLo/oO5d3eyBEpQVeBtNL7txgoPg/K8qjJxPS
CRoFqemXaHxmHN+q8nly2B2ULiq+HZkwFcWrzxRgwZGIEPuKtTu4atp+0SJN3Mc9TSOPtTFCY6u8
j0dPmE9Ch98gyKGrFFXYSe616rxaaoKIz8yDOcAPfq+E3dMry6/9MuQOJmg4Xger5yR4wfSCzyRg
en5DFsT70kuyiAKq076Iy3N8o6EbJttrZxwGp8tnWdO70UZnKl1xev7+g5qRL1zlU1OPs/DLNEL4
lHOVUH7BYckSRRXfQvEA+CZdeOTItqSbdHnA1arxWkT7dnIeJFLVRJcR5E8xQlQHWLfIm5+IGLw8
AHRKPt8sqXc3Kq7WjKE0THd5jaitCdWy4lCCJ0Y2/yz5efhnpA/FRu+ICbNF3XGH6J5TZ51A8Ayr
HRGBV5+VxXw/0Qx3WeFccPElqZr4EXwpdqGfzyFu0e382RBYKl0GWikuHOyHnrwmXE64mGTHfdlX
8TdSs2JcIMPZXl0HWMzJEKbUGcS6D9r8jXZ5kNlEDDA6gsJBY1OhNcdja/ouiNDDp22/qsy7l0h2
wZLyzU3DWsLiXtuwoSMW3jhtERZtBpAL9zQEr6iQ4YMDsP9+DAsecJGSjtalO5pOh1okzAG7ICr1
gBpR4aHAEtd5C2Fcz7euKJpV1ta5Q+bvJ1tkXbE3UtFvx2iNagG/JeFY5xH4aq6Qm0Cdk1lH5JrL
h27/wWIefqCkAYTRA+vvW+OXOuLXJyy/MczRUEqaYFWz/XqqDQ/cfIdXNE3ACxYFR1nkrLt7Gmhf
VUHGwI5hCGXew6WXt5qz/MFhv7VJqk7TV0QRWe+7hmfz4nraKvgpVKRAhdUsqw8p7QbD7baEFEtc
/RE5kKR51xxHJ3xnDAMdmFaR9cndrC/cQCo/mbcH9tOO/y5odjYAewFNeSMowkUa4tnpjXHFWfyI
q4+JSazWa7n9vaYnrlHhG4hkcceYd7j53l4zkOTHiqIug3+j+dsB2ozEqGjH1LfBgKp7IsiMRvMV
yT6t8HKQj3OiB7z6fUDxgw2fY3bgJnqQyg0sVJaIyYvpXM8D4purcwKKn+YO1R1RAE8EVBjSw6Cv
+VjQLjKsxDzwt/Eg5pXD3j9zsxTqTxot+vxhwjaBnR9NZZhyQYQRtA7KXkw2dIu/DoY3c3AyWkWh
+rHS6IlJ5pbIxJ5nL0lelDsKZnkka3FSWSG1pcZNNjiUMT0jdKziMW6oWwB4uZo1O+SNyXcqU/1O
10nPfGLW9SWbX67DbixbyXgDR1/UJ7JEuajL/t28vadUo4hc6g1jyb5We1LgxtN/HHsT7/lkjiw9
6bLO2LKEQoWl3FlAa/c27zM3XSGD3XV7um7IxFdUxzd5oTUHDtDtnpkv2x6B4sJzA2EbHM0Dd4e3
uyuotJXJ+71TjhA/WZ1+LGcUbdiAbd+QHK3e4ENDDq6RpgTdOQqmUpV6JHkpxtG10yUm+zxOLF53
bu8Fp1jPJ1BGoDsVY7b9/OCggOdoicQzMPtK4GR8ltlwaliOiPev6Bo+Z76M1qdPKUfYyKBcOTZn
uPSejj97s6ishJzanyo+waM983gEuJK53hjN4QYs6cYZjIITNG074idPRu1MVSg1tnwN1ur58uBQ
L2nbIVNnVOEJUQyc41MAlCm3yDTQbBuSJpnM6D8+XqXHLGaUHsvhSzaHk3gzLITtBTApGbCxMDq4
ZYu3pKZsnbESBB9yb9gfsC/FV7PYQiL2Q/J517SoNcrSDcxceUXsV5UMajdHVUbK6/rcIlU5SVdj
ASRF0mfciJBYDy/Nba1p3bq6inDkj1yZymGM+Vo39JVukQLUTzz6CWqI2ozaGHkEv7PjdHGuv0OD
3zfQOETFpM3GjhnP3LGDFmH4msiAlgU3lcXlPsBRS5kEWhlWEBqNBIYiJaZ9iSmL1wD95zU7GM3P
5IyW2vR4J3TCqg15zirfoUFh/3GjmC93N7UtyT+Ac5xUk4C/k4bQMmoeTAThL56rrT2qGAfLI0bm
RWUR6iJiloN/1lrFORzC3xt+vqPMfB1Lsx6Cqc7eA7v5XBsPdVdiXcmcqyEV2MzE5H75zJpIN6ga
FrwevCxjI2KShxAwm+ymPNhSFzdfEt07K6PDS4/CuR3kB9FGlErrupxijPExQXGbCq3nVAHaFXn4
ZQsufdbyahdNcgUjzHzTDHq4VWXjg6m0OCfs0pzxAJMvxDt4ujn5MP4LVf86xrUH9i5rVuaDiZFj
30vcNHlGdtO5VizDdLwPhAVz0YIcXYU7KiEg4GE88eKPLJjkp3oheZFlJPFoYfDxR5AfjEXsLgOl
Y0eEnFQnN+cmjwHgNiHszds/JCvRD8/zd+3G/lgWFHgQ6w1iUAMtWyiWGna7UHGlRk82UAu3H3U/
28UporiIlk4WVBoWkewc2naXKZKJ6JS+tzkRXJdqnFIvW9ttXjjErBUFN1N53Vx+3hporhltTq35
LN6mUS5zIj8VcW3sXp7nY34o+/RKA9xWG+E5bQTZL4gl5udkdmwNln8j1T76skBGtZTxq07txmwQ
7jnI8Sbon3a5cvuA6e5ol6Ms7GKlqHae5WzSoDNn3XerAnPPjew63A2v+SaErtd/BW3vBn1L8d0P
m9jJrTeSSJuA0SIYNc9/BCJpob/edZEKMVefXc8Ui8JqVxF6KuqeuwQ7ZWrX7wfIPneXyDDjH3qt
Vp6ax2cvtv8g3tM2B/HdS0fTviJVVpQdmbe8iTn7hLY+iQHfbuDqbKjIjXpd1BfKTFcspTCI/aGW
vw68ZsDxQcRc2PePXXUshw5NcWz/5cIqY42aPmASVaU3Ck+h8dgQjY50CX0USMKe8hlDy4WZO5fl
oe7YY63ASGDpsqoC4mcJYaIp0T6zb8PLYNT1jNs03AXc0+qgbzcn9jQikwU862lhG6PiekIX2Eqz
0nN7chdZUxDm8leYumeh9GTGlv5BPjF89y/ZGnAJjab+7drucO6bEjfBW1JI4kFufsT+NNGGSdaP
dnOWVIPrJi98DQNWaXjJaOL1KII5PaOvcs/VHonHeE/fafxJxSLevlrarMhHlSwhr7yrPGZd5B0t
IrXR8ekFUy4FsXuBduPROgizLbAPf3Ci4Yw7oV6Lzm8DoPYRJbAbwf4woPrcP4C9C8ofIgKlZw+P
NBHmlciRmi9Ueme/F4kg1QnQThW8WgQxD5Q5MNuZIxNnFYc31/cZ4CWkLK7wte/YX15XzD7iUQw0
BHxGMkxFuF95xLXBHKJ+NaImjpQ2ptusAK8XEy5hdT0STdZ2wuYfVvOpzWnjOq9qhWB1LaGAEbnf
nVQwXxSlb9cvBucGDF0ufKcmQhYj7x8oGK8EucM+CZg0RqWnBLl2LFR758DOMGUy4yichawDvqEX
+nhQNTCjFUbmTtOJJVQy7y8Lh7qhXn9MDQY8sqOCYvGmqdZA/Ep0+D6dsfyP8TFQ8HK9nsIPUgDE
N7vsXHhPa3HbYzBScTDJSq1E5kuKWOuNF4nJUzGJyB+MYKJy0w/2K8AECo3g8U2BsKZo4Ar+Ngfj
2CNsNrY56wbgrx+tribPG97oteferr4kyRfiin8YMXSOQPAi7TsTMf4y3LLU7t1hYBSP+Tnm9XcG
QclP8POH/3rLsO3rfcCwozgraYM02zt4eTAgKoDd7ciFBEufL4GzutKdM2BmsczN1RR9yQ9jjeX5
EtfyCj91yMNqOCBLI8w6eit9RBcrtWpDTVh0nbclsOst7vnKiNSgWR9gTnx02zXg+B3YpLobGvMO
7dmJiE3JXiM2NZ1RiENLe6VGOQTbZDUTWoaknYKUgayW4Dc4S3pidGcDckRyzDTAucT0LPsTGoWG
nKVJADEpjkzgT4L7tIFSb1ERQ1i5Rtmb+Cp29dIDXCq8XfPQ3jFm3bQOlyVTdpnfRoPeUtKYc4pQ
jyO3mquHxTzV0TYAuwdvlE8wkLxavXuALiMiCdtVYbfOQDg9flsPSXLNR/LlFLQ3LSFkRIhmyYlV
lLFeZLsoYG2xxA2Ltos0K1CxHUt0cBEYu/R47onBNcKi/41kpayJKZ+wrLIc9msPj/AlevIr1Fm8
HeUf/e0E9cSMBlbSbdKtqlGfm4LBV/rnA6zDtgxBqtCcQGETvdLqf9rdaAtOE3XU9Jr4iD25M8NQ
9xuchRVtfipytu6JO+aW5Wxo2EeVHumWuNXeGWlIJsQ5zAK+S98gWYzRu+QIevD+qiSiR7Ihydpv
imev9aZBBdhJicEz9zMjGjs00BXs4CG3fynmX3iGo02j/SWLDPdWnx+N9h9UVMsBYEfXckC0zr5k
VGyjJsjK5I8WTQPAIIsvs73tQME59W/L0tVnI7KQ3yzLyaqYgKTvqezbW3z4Y4twRbDYqRXufia8
eRmvJeNdERwzPZV2x6RU/1ZCvbyCp4ZedRHJJ8VKGvsRoqLVkJLd1fY7dH+hYHtFQMBtaafa5Sxc
0zzFlqb6aNBJNVfIrzU2uwWVQP8VxXdkl2Gdlg+AX1LR9eC5zrt6eC2wbA3gODwfKnqanD7RJ6U2
dl3gX4+Ct1pyVfhfZYi0/FSTXZdvoifMYZs9FQgj4udk31BJ7bc1fK9a4SZttCY0O4zouWnhwC8w
JhXRY5ukJnV6vjzp2tQ02LsaClJc8KDLcGoTQMP92p68oYlk/KiIHKHplbpxYoAwvadZHGMHwzfD
n7WafdNeiMlEpXbvIAdWllHkQNLbDr5I22aeJ6ABUtghaY6p1U4qMZQNQYMLgjPaFG4fBuVbThTG
YP5MYEjYOj4sUVaO4Si7vOEdfgFZgArxDVEx76p6w290eCquKT2bZ8tzSUNe6zlsP+96LG2hkGwK
2Zmx8fX2yi2gGpoTo4sjdBVaswCiOjvUi/zh/RtTl2T3WAvypDasD4LovxIzbwN7Q9w59+teC1Xp
yDHB+cJME9cqUCeUDVBQ8TjU4FjZqe8dxgxg9JKJCSEt+ntUas5WsU1e8rppe0GtHwFotqWRfXoR
f0t38Zk/l4KCb5YG8Vx9E1PPQwTEI0RUir408sgAM/HSu52jWg/SF6Er7f67lDWVvkAEinuB8XRt
edWcyQi62fXJDcOGutyz5NSSQdKkanARJvLHz/EC3YwUuugMMOncMRjO6e134nR2900QJvWsRVU0
DX+P6dgqHXi5S/oshQZDEvZa+BhiplghokfKyNgsixzB7bMMolewEnHHvePmaEwfLwP69tQKYZgb
xC+zDt1Ytxu9py2TldX7XacyqGfrUSErX83w3uv+++6XHHV/zIQwxpO3cmgwEwtO/NMTsFSaMyKk
8G8MfAw7uE2vCktouSrkzeyKdrN5/he6qVncR3V0CsoLqTlJD3FxtXJLRLjpipH8i0rtJHmUONg+
y4MARiYkD6JxNuuS97Yb4lppqrJEk/nK8hAGACWet0ejSUhY+UMo9+JsVN9bICtsyO2YGM0CYsHH
ssKmy4BPJcT/bKLN1a8et9xN4hbS42Zij++ADvtvK1fBs3cmnnNDq1M9apfe9WmuJbkXZYcd25cl
nVpQYZoH1TGDyRiw54iEKySKibP8nI+Z1NygICiWN4EKQ03Oie6lhAFG2sW8vvNA//uxXTbDFE4W
0Ctz5toJJsbsXeU/KnqHM8InWe4AGdPbNx2hL5YAxucCbWbbEpWQnOjCti3XVVEoWc0ZOBNJaCRZ
XIOlUNRzplCxGfvS/PBd4RZa7QqrBhiAdmOpiGJmK/mVHsdQaiY77bdK0OOWz9yEqSt/Zy7cZL28
mqftfjVIHBWV4NENxC043/jUHG69NUSYe8oX/dCmp1/0G697JlWY9KxkulSKnNYeXa7XDSf4NfvN
y67fOaGIxsiijYB/KjzADOnhSsYLfORO7yh8hcBtpyBfuRfdAxqVjlXknAjuB3+ktFuCl5fDnoEr
6akjiKDRdjGPq+BryDQv7gVwdUYdkZmfAKbXM/OGIVz/218eiSzwPOfCY/guV2N0mYjrGsVd1CIn
lvh0/AL8KBlPnVyFALDPvWuj84NuTLWojnTTR/F2AczryHv+WepXP5/4un9NvQiYMaUFNGJxagZC
cmR/tkOSH0RoQ9OT2du3nvxyVrSBW3Kd9nBj+nvG/UWqzviH8r5fWxZ9AUA+Danhp0W6OiORdoRU
+7oUB2lPCfvWHPrk8TkXl9qNrnbkuPE+QDKMuzbCsPWBsXbWz/aGzAu5e1pG/ShFlUBzeg668Sg6
pwgeyxABLjm17BkIDcDhu0m/JYkE3ofFEh7te5mXtlrHOBZfnknxTn1JvpMcyLGdAtUIgAWB4doI
ttyyuUP0y1hm3pMdhqg1R7pcRV6A+cIj5+NVyHchszSyX8H43reFAovHuX9N61OcHp/3luQW+iN2
2ZOzJzKzwpGRYL4vbwBRR3GGFZtvabbJPjpjt0xjPTGz0K33DbUXIoWcJRmxf2wnA+4bGFbb3hyi
GAqYPZPZlbiRtN75yayi6PZ68eREIUfdVSeickgVTkAGDK+m1zd9RfjFRJTNVrX3Y0PcSs7p2gYv
dyfVk/+X9YLSPTfnxCQWeCKVXcUByBxLVrpPD7GKKSCXyE/hUE8iJR6XegX9ni+5hhqBiPIcw7TD
8NFdcdOVnk80uHrZLcvCjS6XiJZ/5/W237b+14y5wyb7MzGtSkUv6u8Ifj4CWBDgXU2tTZqUUCjb
e421PAcPApW3FhcWvTe1Aby/DCEygPgGChoQs/+DVzXYEQRWwdOV7l4dxw82mQ4nXqMz7P+g/0eS
U6fv9/h/hxw1z33VkSnyZt30HsVCxh3dMo5+0T39acHcuVk/DcOd43rXvuw31q38ybFWUOjxhKyW
I+2+0aUiX9Rn7vQiXiB8QslA8DH7fF4ayrxL2Sv9dEZnmrwwQdtd0r9oJDTfVlzPks+QN0tBxfUh
/NRe0tKaPwQIrEszcxo67+Z5ebN4HSITs5QQR6GJcrtT2dpxXAzIm0c+WGr3OVZQeY0XQhw+Aj/r
yusyEqBPn+oYME4u/7tjtNsAcVF8ZSdd7kWSrDfR2ud+Wv9ohX30MdcYWMvdJZ6BXADzl9EdCMmR
Mt7pfbTikASO/I19soCQIUNNetNkyKhwDz6/v4WIh2NzXhSGR5cILtDSHanUv8amFOU7s1ioZCTC
EjlL0xoD8pY6FL3QEG0KmJYhmjLUC7jjI3hi52NjNdOmQQJDFwZW9t83iEQYjP2AzM2eZQg/YXnb
t+qKF04dM8nPVdth9dUryj0rCBvF0KccRbUPiixmIM6AP7UVKGFxLBrQb87EntWfkNhLdFmP+sP5
3BUM8cGCZYNIOVRubVPsQXbVVvquiJX6dUwsH5BVXzWUs+UYazu6bWXeI8bYYDo5avILdQpDEemi
tYoN3NgYbPZ8UsyDlK+c+bC/yAKtiz5trJxjE/nIPQ90hz0QZXAZByElKxNmT3yeKqwsAnAGiSkI
EOMygjs1Ae349aANCMg0+R02OfGUJWS+LZeQtCHVyAwUr85AeSRbYMURQbDu/giKWLruVU/jO43u
zCTxMrdbibz9cgPhphfqit1UY+Hd2OIGtOaHx9TRbioBz3mFdBC6Ad4CCGkCHrp+WYCxeTasGTsj
kqs9lnSdccnWFC0XFknFw9j9eJLeWWuj/wGf0kvgTyC84C6yUfht4VAEAq0HWIzM5FQCafh0qBmV
WqnX8MaBIRFe+biKCY84FUgqXsvdb9czURJ/DfeQ7H6oJUt9XhmP8UHZfDnQofZrLptVw9y6LgLz
AIJomuXKQfalNhPjVW7RmjWXb5GlHKTq53160vEwcpvcKrb4hA63cqJRkR64uK4K5xC/N6zhp6yP
0yRTuj79lVoPnuQDCwmqICHhWhf6YQsrlHPJ3RC13eek/rNV9D4baJjpIk3X8kI9A6rJL+i34ftB
P7TJMegkaBbzbDDiRDLov+ZUSvCnhc0wA/VALcwo48RD0f7UVPmzx81VJbj1wcem4D93TXGV3t70
1ZWbtN511xW8Y9GsnBQpo+mMbn+HMkaQ8xPJ2JPWjmhRPOn/pszsB1ZQ24vJPPX98Z7h0xgQ1v71
rXE0bUX9qlbwnjhCRqkhkXTw9udz/Yihh+KNVDbyhmKCYFeJr0p14+jM7ayZcwNqKEDEulsKGUlt
X+K8lGb+r2uUiSRubrRSJX26iA3sWINEEhF8jda3/+V4U2HUhuVKJaWUM1cAPAdod2UgEtjqgOAD
qr/87CeqeN/63OC/JPslEcPSEJ0glKk/1CuO4NaP+REpix7oww97sp1bGIPCDtBWwxxuRZVJaP2Z
R8BJzWES8omVkDVw2AgDP2a0Ypn5e22HJoouXoHM8IF0D8ngsyjJDYJ5drrDO4SjU3AJ7EoRPVOw
BjC03vXK9bF9mxUhYEXWdg4wHm4SSonGfS8d/ywOKEC/NDxY5vcXHWmUaL9IiK05krjebzDit+ZL
nH28bwHfe3MU41yHcKyK2OAnefCP2HnyrACMKAK/Ai4D/z+2eud/uCrLLsTSqoHq8PFOwjb3b4i5
MYXu3BCuN8A6DNPgCpzsMOEUhAjrTTG+zJ3gb2vLa3FNH0ABRoYnrjcb9NLWic6wgDkf0odiiFwV
raf0HzyxaDYz1itQ3VJ85qAG/dhEhThy6aqfZod4y5RhryIdDz6fOOJgQDf/qL906LTfCJkgyBkx
o7vnGWiOScG2bjPrVZMQS6w01dFAJZxVpgdG8T/DIQTm+gkrkk3ydTasXs1NA7LOO1aNAzIQq0/Q
PMpkojm1o9eoZ2NBqhKjDdWA0NZzOgcwRc41AfZKQ6bm9rFPeGOXwYi06ugzEjHokBqfNSPzUKPm
mTRihoFCEg4BXOUd//DRWYtokGcX+MAV6dMfg2Y5zKkPdUBiHD8qBvGXudl5CGyr0vBDP0FjIPee
f/735hmtj+Iw6g5keQ0WLeCanih1UUDJkNS1RhDAqNZfcy/QyLTbKx1UxpRCkIZkMV+mYGoiCgKg
yXr3UrCxBnVP58Y8CNEr90G/2mSVVysWPBYRLIR/lDXoHGOtFsj7TbDnz5v9ZgWmspscVx0xiuwz
/LrmCaBHd9P1d2At1qi3ZiO+H8c2bet2HFDD/C8FnubT8rgC5+V0deVC6TcNTbEWJ0UOH3acZ2hB
mRhbs7r3Ayf/NKZaHcGgHjUtbPRWPvlQ/fVvkL5hh2oVei/BTQ8aqMuGKnf3aKPadBdFbfz6d8+Z
IAV0bqbjeflg/XAMtH4keFEHAUscaSUL0wpH+QYGBmaFsGG7OfPEwANjLxezDo9FSuk3sEpfjL0i
hn+YKgL1Fl9MVFswkVVlF+VEc5954WTzPoNzKqk8pSPZKLTT4mMoSEWamItByKFJC6YYrZAd/Yl9
Yzrl14iQ/RbjdwVl/NVm0IhPdZuxG9ZR7ON+NoyIhnbme9ss31uG7h9mX11x1V8NdXS0UB96z8GQ
KOfmU+89jGfNjpps0+hZ8uOwuM2fotz2ZbAu8XTif2Td+hwJAyEhDHAuB5mxE3XXzU8C+Zd1fZWm
U0BlKFyiyz6ngTVSIokWmzTrj+5xNpfNF4+eDlH0/4Nxh0jUfs7hnZrXldOaUiWeIJU4fiHv978n
y/VFU73QvumzN6GQS4RQzQfeVgHBtOJO48p9my7ZYiMj63IENSkVWqeBImonbRIgB/N7jq6CxBuK
LUOniYL50gFhHKY1JN1e047U/M0nH8fH7n3jBptdxUi7fx7pukdB9vSWlJ7Ur7UaHHKUVkyVhTuD
WzGLRMwkgAuqb0IF2xYK0xwhU+Y/KdPm6+eYLyyQ1iNaDAq3DRiHsqpUT1cAXVpaL1BoKLv9Hn4t
m1qJ6WnDBhVzblKT4IpaTZBkma5tNjByNiZXanAKjULs8qwzntfiyDmmQSZrf+N+81XggWfPnofU
IZwo+QfLwqUO8V6cwANZd83/jRtApAowz366E8VaUAPJ4mdFtm7Gx8PH7ghtp9Sn+D9XWmvj+ER4
OXMrzNz1fuzY3qYGSQuReaxn63smn2pVIcxTz4oivJMGs00xbrSxGEyzD7iXpwrEZnYaFQr41ITl
ll3GzT3yXJiKsmcb86922e8TtOlIi7RT7RtV+vsQ2bR4M95PQLSgnWIR7EpAowKlGDkl6jvZI5dl
yyIQmhXqnipV9VTbG1NcS35CXzEO87szKC8C2d8F/L9R17UdlEgC0niVAJfcX5SQFBC1PjkFGtod
4KJZxx3optqmskFdaK/44ltkYwhGLs2ssghwxtEOfBJFFuivQWToujD5J3dxkgsjKa/fQmy6PIeX
2+C1ytVJyTUdaIUy1UXeit22K7c1k+OAP2L0GFSA4ECvWFLLpBowmnEgugPVhAG9lxcswgKECq3u
AYPqsT6fksCWFqq6XKp/dqdub8mNVliRvKAz2GjuPoc6c8r1UOFX6JfgWecs0OQbt8Xqr3yDs2sp
pizsTHvYodzardHLJcRaWTEG3j2qozIY2kVEceegNxWPlPirtmxaPD+RpIE0I9gyqKWfsOH97MzD
orMlru8ktyE64gifaCLd/+wCSNeZJ4UJiP6NTxD2KqqsmdL/9E9cDnE1/vVogDCOlDgPMv2f2qdq
W+hHPXquPfRwqc/k/16v9lnkrtnlzi+0kk1JKsCJe+thkvvwyNEVCuJ++dw8c2uehcGHqa93l3G2
HihvyRdgBAQ4SFeZ7dOeyqIDhUQrdUhHBDyaOhZHjeQ6IKkg0Id8PVxw2VwiF0D67ZMuF8EZvuK5
h2izKMt/IAS0XwIDK/FObcifiKSgXzEuzgxafP4ERB9oTfHuV0uTwBlUcLsRv6OUZBREGCfluAUY
VVIWS6pEtxD95wFf6WXxKp0pyqrB3UA+T5u5RbDxOtuc3se8wF4Jxyrblr/DHt5vM/HTF40UgOpG
fiCpszrz56a5hLr340DsrhH8APpFtjIv1R5aEZPfk+hDfzoXwaNzmnYekwytknsykHnvtDDC4Ihf
Vf9ML2H1Mz/6I0pUewGkfG7h/5G+NCB7pciYjfRzGxVi4IzHWyOiJOPovV4/CgHENdZTOO/43S1e
GayH3yX7vs8LX45hZv5QQKpQEl9AkIcSx/1bXq/vw+NGZBY769jYgpr6QPvTMDJqgk9vp1ECdOES
ewqKPM3FMDjIJDMEGrNYMOKdwDcODYBk6dHVrAejzvEvsu4AdVcTtCDLJoDTsd8dQ1Z91WAhH4t4
Z0rGYkGRq3UmIKC1wQi3T+yRyHPwzKPjBBcT833Mib+0s3n4Ea+p26xXBbacUEpPMdAH4AdysKnL
Or0xvHUguNoG3hh/ucDyoonNLxvnvAm6oM6cCf0VdChdWfnbkAGGm25GLvBobeHtLZHjp5qMqFv4
xBh0XxsLzcMr1rAdACN0eEMKrkKPYXoe7lXBnwrmauAUXB7ZSS2OPK9l9TSZ8utc/vsF528BxZO8
yXx1rcdGTFMYR5zC2sTqz7Q0fMtiA9UmfpaS+pXEzmww9muZb9k/ym9pYzA+OCQy1MrbtgAYjcWb
RdaB1xPIRwKfnvTIigbso7m3+L/qGvMIMNIJNWYpjolhpzZDdIFavUI5WWHmZq7MNFU4P27vVJtd
PwZSClqhCfXqUkdMZxpHKJpFqTr55Bfduu1PJq96bb66K3eJ53rhfihcDIR59yoSxLfgC5+m74+k
XKT9c+q5zrAEO60qQjljrd8xrCsdbu1zNaYbWTOI/ewXkKVo0UMIhYvUUYvFPCu0Y0Fqbze6ahaO
ZPderfgSqORhNC32MBkeaBrFr2mr+SmUwLVCIPP0SXPqQWLqH8/Zl39b9BE3O1irKu2s+kAJKq+s
AT8ppcCrc8L5Nv2lqCYC1QgsJmlUoyGZ2EfmHCO1zWJg+hZd/rYyP0J4zlFMceuq8zMoA9dSsiK6
/27VJ3Aom/JZ3ma7tFt+OygbP5my+V1xCL3BvlWl2aGv1N15muyKXZvjGfIwThAIzXnLCjqMSebT
aIcu4T1GXAfWGRnrHcA4vbJ2/z3Inpd8EYEYuhre8tEKJIVfD1tUaw2BzKb5I/GoHbk0OLMIl/5R
Pt+yuPZ6iIruVA9JZF+B2uUiX9uN6pRsls3AUIS6fjjSzFC5YXMhRjWBA7d2O6nKHWPQS8cY4EC/
DJaEv5+jDd+kjY7VDca/WQXzqM0OtNH/rugp3dfmwZ7O7bj1CRyyySG9+Qdlc0v20087aM9QgXNA
HMDhdxcSm5jPhOs16SsNAOmLGi04Zr94TZ71XBTeFDc7n0PhRzduhRNuAlmtznOxh5eyUZ3mIyQt
QuHP9e8Hu1D8xT/2Se6zsGwKIN/szhg5OHKwQubus8+T0UpGGwWB4iyI8TAgi1m/K0hUWRN0bBWA
HL4XryVqDmnGfUINwD35DD4g8dNIz6OlFjZ7Wn45jftlRMxg7+l+AjEjoDVh/z0JxtVt8PjVUthz
X7K1OjZNOGAHL8pxYm87YVIFY8nGhunG/X4CXumWYBNGquXeb6rB2V8mXl+6+69MLCH/bURhEpoX
7bVSEupSFkRjHfnbV4NMakfBxreEacPcuc5i2sNOEd3lwIMwN7tz0pLXIYULvKTTisjY/2MXr8Sv
plcS0DRLzcS2VersTQ+6BcBehygY8PnC+o+puod9qiOS6yXzCY1Zyc6Yiw7pWnS3fSatymqL1cKO
X7uLeGBZQvwA622Zh4nhXas7IQtm8v1cxJ6ysq7lfTCNZntxTjlHmbNd9E3Pq6PPjgS8CSdzATSc
SuS5muKsHsdRmGCnmUp72tj0QgBJIg5U8uEqac4j7eFv2XZ4liCOMeKr4uZZBGwNLG8UalILI9x8
N1rpQiyIJ5CpEmP+y+Lp9f5npLPsopaSn5ESB8Z6+s6iRrMVb8X4gEpOurqRyZ9ENRcut5ZFRT/3
gj6ETgOKzTeWQswb/ANgkFc5R9WDnB7cV8Mb7B/tYl7faCAeStInrV9MCY0pznFeQovWtxe+iPuO
UvCzughdDf2/zKrtabruOiZ9pCr1v7gRz1XyApSDFlTJF66E1xLPOGdnfqd/WoEEUO+WnprOZrig
xl+ZA4LVmj/FRlUoquWiAxgk0qxQFMAm0coAd7y1SAxd9ZUMgQS9Wjte6CMezNUDBKYd9gMDzeIj
2xAh3cVRGO9MkKM9ciL+LnUq4W0y+joiBp0zJTga0KIRJKy/CW9GM32yveLQWjeiKjS6rUgUikgL
kQLHiWk0y9ifSA+UK+cMKeHVWMcPnH/Fj3PdUXK9gYjXmrfKITscnnFCbCoNdAnGeKeMMDon802l
dul0Zwl7gzeHOoQzFsyuq+9rI3+KPAkzJzeSaW4U7o23HEbfbszndTNr1Qe56UZ369ZHyPgJgR0y
EqV/Btkl5C4OE2Qw7nK1rPQcIMZ6GANph4IcbesTSpuMPpO45LqTaxSYvcHGlE5bEHDTi0Aufd9G
01M1rSsYqezMgQcxZ2+jA+AqsZ9vlr1IBNqpQ5qe0eZYcE2cWDKtgxgF4G67R/wTAcqolbc0Q+r1
5LOM778GiaTWjb6xZFXnEN0IojUVBcBuXnH2Fdoq9JnO6XEgQExnZUF/Scl5rC+nkX4WNBpszAkc
6nUpw5SJ6+0lQM/UY1/b07qyoz+BnJoM4xEQQUu69aesIzYl1nYpQFFQLh4PQV5+hTfZg5K2fWch
yvVdUYMP15zY+w9d/nhbOtyW+nC7Vj7VUXxft9Xcf4tqdNXveFhJMxjNgtXgBpSrWAXFFAuPPO5b
dU3wMPggNwmrQnhoLtJt7sBt1Wt2x03SeGLiwZbJDXMMk4lQlZpV/AunqxXkW6JHEET10xm/oF98
ownDc99KemHVktmVta9zfzEmnbLeS3oCsp/x2wyw2O2meXOEvNL9ee1mtilRASqbBTOHqA1DzCE8
uDV2jpgSOmzTjcQrULX3m3OME94BdSKVUiWHHZfaggnm69Y34u2pkmBaqYSVLVXsm29P4zGB0hmA
adLsbQDAb8V5VUSNQ+DeBqTf8BRFO/p+QHGjtL5J4Cm7qAJJxIB34hIqa3ADUquCMyC3CV1QEI7x
VNYIT0RxmVAQJ2SXfcYwr/xeLphNg+aaklaXQpgsf1hzGURjsBBYDa03hHb4ncRve61PFhaa5Z66
Mg01A2bW7ayfF5WFcyCEqUZD44NonNnFRFmroW8iktFiu2Em6gMJ4g9I+sASrOVqByGZoS6YW1kw
LOdc2IBiRhLnWh0WspOAut/w8pWizdTEh7wJa79asZtM2XAJKziLZ0fFgsPfn4snDuS1deotVwqh
Vzbmtc24QjhF6YsqiFqSJ0VF04LUbo+qeIj2IvKA2iJLzdjZ0hqEmkoR/Y5wCdtUpUiIi1rzEuR2
S24j8W8QB+1fO19zhvMF7T5Qd1Bzrdr+cxASKh8gr3WQTvstN99X55vfouJTNAkAXas4TdZehOxW
T3vErkuDSRf+3BtT3edDP6uzhlsjtc0htY5hnmbb0cQLGXrJoUe4QcXze9jtHAQFFME8NIBwnKlZ
vHqLQ7S3aUOncWSR9TowwdBJOqHFa1PyA7IhQWvysEFn2x+xQPPrLSUvHpYJmIpXJbGqcXvBhHwQ
5rtWxJieNS2QCd5tlcZ+LqdSzsXaOLumy1+iOmhqTIeodp+em1qBMNlVo2v+C/N7ZM1mfBtKsjES
o5AVLLKYmJWmV/gGXs+sKHx5PV3+0nzeFijPRgx5C1+++JTGU66Up6e6/oFbzq5X4N8shdTaa4b8
U8yeCPW/U4nBpsmdOcAer/7Rcf7rZxkGmVdrakmGDUr1oVQu0KKC+NY+oMvZcTNHpdoj1RE/Vc4u
9M1VwPqSZMPhpsjpFfXVbaCPE9kqo5xBiMFvUaUg+U+PR3AeGTeNYaPdjQWfW7nLfr8BoFr3PtCc
fw3hyoItgO/kAJZrrmnFww6niRg1pCPM0NTI7xbV3UdWLkj1Sx+meLQcOWp3jirN/gVZ9DXAXy5Y
CeeTzu9oiEKbG2ZPqoe5RJvaukd43i49jEZu/pQRy/U/nEHXfuxVT3Sa9rTp4B+LUgAlDHaShw+S
VbpChJ0HaWnRX33skiY0f0HizVxvIH1tHJccAJTUWPJuZqxvQQj62vSVqybwN+q4NqMVb73eQxAe
sxhLAoVQlQiFQ33hfA/6hW7Zk5OTw2fWvGxvj2Jiz/8GvdnO0sD3ZOQz/YE11Wb7Ew7kWW6GbWvv
3pAdDNfQYdNIWT8zzp4XVpaWKuWAa4So/vI8dbS/g8PbnIOa+7bGfhPe8akq5XYP1GL4xSitgUvF
8K1w2CtJYoZ6OvHUK5449fXoniPdvyMGbnb1bKZN7YbVkTtsxWyabG1LpIpZKJp0lu+Gr/TXnXgX
dbJs0si5poRa8Kaq2MBhsfhFo110Q29gYO69Ojnwf15KpEFrFIhL73x8Pv7Wr1V1zTwP1ijZW1YN
pm0Muyuk/oR5uTEPl04Xi5KmbeeXW49t7cJTDO3s5jklpWUPQWkMBloMbI9AqciibkEO5EszFtRV
6GrM3sZlC13NVtPTWNyDfmanyCwcmg8fPJozDy8TuK69tbeX4jX8Nq6l5yKbyElkxPyf4RTwudK6
2mi5YUs/0uQD+vd1nyiSw6b1iGHtuh43bDw9OGb0y7OMVM8l4jiFdA4UEe1l4Aq3jFZSdFiDltli
ibMAcEBxh89D54bBJzBhPfXCrgD/bO4v2M47xXLZNQ3doPkLOt6B7v7DstPRKk0+lIOFjixwFwMy
lmM8VenqlqV8Re+f8K/JI+YnqBU8EHOIhehRDOhVTUSq3Ql6PThSfCAoqg8mghI+iyIWa09RWD9f
X9JUB92gxVvTh+Z3XIUPyCvRqYOc2TwU9+RX1nSl6cQP6E1M9OlHRMUqhgPWmvhytJcItTRyGhyN
aYTa57UA6MTqO7Wykf9WUIjoNwl1vvuf76c83vtDjxHPeNyoNKKodVjkKKDJP/K8EhiYP15Drs+S
HRrcd5V9J1sb0jygWjt78ADg0JP5kF4a7pMhYJqiQcODWmpkRJGco1UIrHo1xNGzYzlvvpFPFYns
DRQPFkMwy6SwAu1QZQage5lkmja3eZr5g1zOVsmv8zHUXH1IdH+l6aUuFfxM1O+ehkGKKgivD3K6
bvPx3Nkb4FZatYUFF7E6rpM6hcBv1bg5Ps6sptV616rKOFjGEUvkKG0ZBd31xf/wpEVpImfp2hRP
ZAghCogrsPdDrXDYAOBlGzyWergymmldVhm8xQXsXAfRMFdBKP9GbVkLgdxFzLWTgLLHI2QTkqOF
Y/rkpHqS5PfKutC9c2DLAwyKbFv3ikmx9ST7JUzLuJvuxkYRW6UHfoOtfS9RBfT7aPwv8FDEl6lu
zaRi7NVq0NgBDeuH/f6tmd0o5kjsf7tbsq7aqm/tNl7ctCTwE1nGJV6SiR29FgqouyPwCYUc/TWb
8BEz9t4e1wxmFduDocbftJm5lB/53AhhNZU6nx8V2LmMOrqOwftzY5IcUwAeIkQM57e1AbnTtMWL
TB9PRqQAdMGFvHzGuBJq3OZSxex05rdnT9cCFYBGzoolVhgDYiHwca/GaiPtreSG263Wl+RS42Iz
ZNWYH70LtKvCW8eS5Vh3Kn3Z77Kw3g86iawJ26DOdEnOm0pDfTmLaTRvE9hAtdMoxjqFOBlK6QeB
zLjnoQI0RwusQZKdF3S6fFNTgmVDmYMFsXv0IKhnprHxOedd1CFW6JoBqSJTsQ8XaqJ9kQkGnT4T
sv+MTjfAB3k04uYokm7DySDF0CB8rMu1UxydWGEV0ePVy92JMWC/aZZkIQ6ECSlhICPhorF5MfED
1tSjtQrmXFzy54b6ri/Cz1v/omEl3Y3tfd83bUFeP2YFKDe2P6KjdZ9rBUkJuNxtjpFdR8fvvBYB
Eq/YY68kx8wiM4xV4FnaG9uJqDiTCVzD1O3Hw1xJtpRznAfUUmUbImP8j6ihpn6hTzXq6aoWclb1
AKCdT0y3i89Uq3mqhyRzWcGYmWYNaY1MypP/BdJzvlFCR8iE9VCtd9blX0tKhtNlwt8hgjZdqiEr
R6siGyP6amXKKbFLlXDd8LEei0y9JN9bTMM++zkQ56w+kaID5Q+wqK4MqYkD9BrhFl3uPh36GyLj
/fbsXb0nCtj6pyHEBQNdXJsNfJAiYv9UMNGF1MR9vBT3ol2Th6266pPRdwgHmGkVUPKsdOphumHf
VXkwG8LVSEX7lRbVCp/hFkL+vvP8Fs7sXB5o/5FWZUaOtEMPRd5ctotlK9aY57Aw3iTD4qamGZ5g
6jvykVKj3yuQxtSYVyXk+5gpOv2HCfJTWfJFbDIzV98ywjgAvraJY1BvicE9swEOdvQhIp326FtQ
GmgwTl0D+KS6tl3VktgY2HjIJdO5w51+GTGgPwg20CDquFPJIFvBmjd1zbmqXlECMWYKyn1OowL0
EOk0HJRVqT4Ub6xnwuZosExyUJFgelkfiqZOjqTHHBwhsSUYPz3zu33GDvO+M6z+oorqzg6m8Yqs
5+qOcCnmCu6gSZscrXzdVL01W+0uoHA0OYz6+Toq13m5sx7thqIxguxyCX2F/6MV9LjChQ8RAZ/Q
qZBNyIwr2z34WKWtDzde+IM62keGZEjoUzsFvacDacMJtTVcn9XgHQzJbQWS1dQs7y7N3eK2h9NY
XdMxLBOAGEVvv0QLT4l7yV7ZkYyqOuf9Lfx6akzKi6JtqyWYvxlW+iNxWhMnYYppf3wBpJC8ve4A
U7jWzr8fotJkiosZOojCC0LOlHupP5UmbDgJ7LwtvkPtmPjzZmNp7SKSWzklJL0Myd1I7VDnYkAg
6dUVIDFkKuQrYtazuQ9CT0J+EbyGB99Wfz9o3u5S1WrH0/Y1d67jfUhwdSNG+qdpwgUbExcMJ2KO
0m1Fw201XQ8aI6CcBRJCvEsryUX+uqfKja0xtLcmpLFeATEJY7KmrVCy0JyUvHE+Zk+DEGzgUfWn
dWDx72PJUm6I9jXL3NaaHeeXoaLRnrEdhcyGXvWaTVN4ofzMgOfAe4xRJC9TNSBzQDJE9copdMbo
UBg5IdgGPIoRaJvxiY7Hbs/6AN3dK3RevpFHuZYEoHPcjY4C+PoGU1amdcu3OtgNlEN/BK4PrK4H
8SpjEwm1k7cydET/eTKXLdQuIXQO+As5/OgnM1jlvGwm/O1aHtPyLjZfZCHawgRZbhHrdo61Lyx9
EEBLGVIezQLX4d+lLXKsIt63BjZ8jI1M+aA4PW+oRX51yytxY6P0roBtE+W5J6m+UZQMMLYn4KfJ
W9EEd+0UzsZArxHymGkmyU9jIg1bo2Mi6HBn8mQgkttWz51BirmciC6/dA37g+mlKl5m3XrYqqXD
y/DvCLHC9uO0EgshEFqnFEtyYJA7ulRscuPkqQSxHlJ1cndcVcLZbZvDx5aDkT/cZPqogf9zYkSz
Yi9IYUqB8xEoHVZcQJ3GBuQV3+SzhHxfYN/KRhVXby6VEuDXZYRIbIWk687laL4txL5PXmxJVEZV
WbyQIjsjqGP/qA2CFyOnEeGpRshVmbGNG6qw9aMiZfASFMb9sPIlyPbdQrl9R4qIAv1AqD/DB5fL
NaJOpfte7GMc9lk4jQYs2Rt1qHL8Q7tpzikUN5UEUeygIGeU0yqTPWNKA+rj3jHtIBGvAtQGe22O
YBhv+Z5HM3RR4tg5mrPv/99YC1a6R4+Ou/gxZ2tDvA8QTMwDpxft2Dlh1lbsc6VvNuqUA1Z32fs4
S6+kQR9jujllma72lqOZl6p1HMZMafeS8sO1ImaN0d9sWxOET2Fma3gdG8t/Zp4TKsLv7ZVM7F1D
rjJaJNE/SmegqIojd7mkePkiMvUPOn5DKj97T/Au3KIy75gO+vgBnh/xY60dRe/JJalG18XYS2hJ
z2JmzM7YVDj/OPXKAbS+aRbxTTbvQk4PVlWsXUiA5oS6f8fWvdqiEF0izGLilBaM0IV5XMhBxetZ
zww4R/V1Td4ydfKjV5djLc/RyxqGu7wya8xsmhPtVka8X+bSftWt9RouOzhi5dFwDdCDu7f2t/11
/Ir7152Z4pVL4Xr/ja+Gs7HO+Q0uAMpvHpoyqjf8hhlwRGvuan4Z3bDaNEW1PCTWdmHSsuKWtYHo
GKtJvThB8VziltcCKgMsUZRjlaK9yH7Arq6tcKuT0uucjv+UiK8jlPpObtgnlSQrCripzNy8QYw5
zFLeuRzxOXrepxgDsHkbvOW7uCBJ/En+W6IQoDTrnmANiGLvd4G+RvEL5WGC/ciyfsgxwLoW1gS0
ajbVqNJ2wC0brM2HweE4YNDosuhMMDKh77HjZGQ+IJnAjih2c40KGexZES9zjIDbxnAgW0MwF7Jk
v100i1JX5fK7t4NYthk7UdM37TpZ5jFuu8B4ZxnRJ5x/048iCiNRsZxh1jjzx9y7Q8DqXU9LCKne
MoOY+BhNvQF2CU+SvwzmUEkN6MBvUYOf4U6jOPEWmLm67pEECurkQRkq1LytFdNK/r+HcdCE8FlH
d++M2G53KLCkEvkDfl6jLwTogZtHWEW3T+B7UCHUuZD+NnU0BfCOMNanksf5gTKXgLhZtNk4VGTO
b/PRacaLoZv5y6zpWdG6qyUh4Rt+GWLysbq15hZjxqLDmuEGkZFPtBqpaKBH8OtJ6L69HSPcduq7
DSjNjisgrNJDSAdPi5tYDUY76p1Kg04i2ecE6eELlaEog0ZqLq6HX6m2bhMl5zlZI/k2hAOgnP0R
jFCzOkTziG9r3AKlNb5nB2otWZcAY7vyrQDmz5sfUviPzk9/nvPJYUHq3ffmuISSXrPZke5RINwV
rpC2llbvOEi1QX+XRrRqReF7893CX/LjWYTNfz8IZyZFlaC52YzucUvnchq0LvBwrJoejMhHDBeC
T6K8naQSHA488V1hCIvNuFaVEgr7TcX1fnkmNfW4yqR77FTpoQ9dPd9Hv/JBEWokmiqHnUSZeWbt
nmAQzkaDIAy9drn7/TEgkzP2ov8j0EOvL85nzl7+aD2zCIx0WRyidCwgsoFjRXpqH0XEQ1RoohgR
8NqI6f6f0JGjm1Z+BmMghoMhVmnNuTBn0kUoKJwqYRph752qsM5KfeXvn4WZdrO+PmeaA6+55Tg8
23nzGbn1sCROTF+RwIZ5BI/pR0XGO/dGPeKGiMQcm4vqXcnWWEUtLBWMZIIrzq6+w59CIB2lL1Iz
xbtyMdxb8H/VqCQTrxxPzyMxrc4VQ8yuL+Fakmyt35qnueoa4WzgSNEtYfQ4LRtIbjDdKXMneX8T
mZY8ylI7d2rAHhJg8Fy3EUVBPSnNkOU2BL5m34kFD45qyTMr1b2ng39lh4pSzYU42jRsrBnSlhet
n/vRhPLxFA/ndc19+ixcE3HCAvvjlOEetPhu3vHkFWZfJqOdrQV0aKwRi3Vr0HRqO6cipujeriP6
YnC9LMXJ3Fy02gni0EByHlKdT1W2wIWHrgujkl9M3uOYtp12u822frjcjT6Q5Yl4Z56twdVmFJHl
sSi7U3rQ+okrE6Q1Jpku8gpti2pf/r/+ryK6IcVtKvgao9vhKreqFmQMobp9Dpsap8dAJ9VdIZC8
oKA57AmR+vRo09g7NXj2VW0aFVR64wt2Nen5PnwPIoL+ZsJRSeJEgjgQ9Wn0zdkw8M/v5XqyBA1j
sOPUwnzRMp7esEUv+QV1FXRXcL0TrbhCh7Jz9bwVF5CHBMLgVmpJ0pCEnUB32GOy2Bmbe/vr2ivc
snmTtUnu6STX3b2l1mwYEZ8cRoONR1wq61aKULqWM0AHKVBymWNkwOIuGYPP5JlDxUXEtUgwV05o
J17WEKzamIjDFaA3JL31A+QDfNoUcRMXj4A0hoKokILfQm6B0BgWg/7+arvGJ++eKnwZBhLVu9Sr
jIYhlN0lUnEGoDgEx1EGPL+1td741ZncXfrrsHBvir0cbrg3E68fWCP/JgkOTXv+C7skCaykxFsd
c3lh+8RsDAhErcHx/r+KFZPYXVO+UzJjYn86ffbNt1Mr2sPDKT+qXicIKPLcL5F/V3aRLiPMqbj2
oKmPFcDL39Ei+PM2NY4GRziLYfQAxE2sNy3Qt0HfmSj/WkbIMqgVk0KKdqcRt2SWTeSRowHu5Hl8
sggUDVEBKH+BwUTTF8bMkFVdxnEDsvSQa2V0KccpSmXt933QkJUzeq6PRHEe90dRc13K5Dy3Z6sL
rCMI1RRv7ue5PAHhk3jbzsl8Z1Gf+e9TKxrkT00uguNKeGMOqSSRahE74yYmoNdwCgi/1txsggnY
YTHXXR8aWyO3c3X0pf1QsX2+DFKNjguM8YiH+znk+BhcGdOV5Rt1WdrgDLrK81t7lBBCl954Fgw7
UQUnozK7rDYYDTxkAUYzxy4AFnibnh2XExOos2kvSzMS3+43Qkf7Dp0hHDLyVpzzD+dx4kqHn0f3
gQRwuNdeNUoQ8GOT2HCX86xEookAMpQg8UKpg0c5sVGoH/IHcqZnVlzh9lyHM//bDngRzfWSraBJ
JOhJkl5Ka4dBuREEXzdh521xU25SYyb+3TKS1ywp7CwlgyGy+mJ+3qePTAuCb+i2qvy2JUeYTFpq
kpXD3Q8KGLXXuKF6av5Ba+3otPkS4XqRpH6Te/3BgnMXLmVryWxndoBgwCCeDqArltzyhwZVtspe
9wUGnGfCntlFkHrfDJqrFA4bhLdQiyST+9cMpEG6/dzloa1ugRcvhoxoe3lEgyyw3ylz7luHPZ33
p7l5XQJe/C0//y1wor+enprACyilIhgh92oCzWVB0Is9neLaJ9Y7VX6LRMzjlsRTxhMCCbcrjkSu
Q9o614YTWf8BHx0Y3IslsX3XbkoGoDSXlRc1FU6qiL3ctRyW84sr3Sib0/PJ7dCyIl+u/R/SyH1i
NXqegOJx+1Oo8vc4KG9aKspnz9reMrGGmcp5i0FAzG4c76NvKrtDjL77eyfskm1oC7lgFMQzwyRD
czzc0I9AF2alg7Kyug628ZTiHgaYuM86jVeNqgmUOqsRj0VtLoyHo15thDaGkfPuEDtJANh4utOo
C6heBWkfOPUARyGpOb1/jgGNGzJ39zH1XmMz3J7RNwzCOnrPKp17IaYhqXyut5DlhLTsezWpmeeV
oA9o4X2jNqxJnJnthoqARelTEtkpivGmPyDyIql+gjPvWjfFGfZzyq64Y+wDcie2bEMcV9u5PDXc
ELpyEUCGuQ2U6FGBEfSC1Z2ixYKxomAeedlRvXnjxSU+z/fStscr8XeVa6HinE9lNlyLHev6hWXm
aYTOq0/tThSAttaGj7SXLpns1+4pAA6jDt4oRoryydwj0ltpTXEpPXq3wFnbS87SrchX+73yYLL0
rLLMgZs9S1Vj18T2zZlpDDyWzjJbGAhk5JGz6gdVEuy9F3Yk+68wElXTnKxzv3S96dAV8PHXMOdS
UiBNZwwbjAiE4cQ5ws+PxCi8PrLNkNluGwQOjVT/l9H/8EQA+ysEcx6RAbjGsYHIXbMN9iSUpYtb
b2ihs+FAyB3QQKe5lPn6KZcdASzJejI/DVGgQgNspmLCvQThTu1wmQIAZk4315+lRaXub9DTG9Ru
DD8LHmRyEKk+gOEpF0NVMFpVH9Mcs27AP4IhbiFF96SC/qLSgmcYFPyVwdPFM2SvgZujQcrqzUDJ
kWkZwW08Ax6ZLrRECOEzJW8IyA6MhQo/9DhfLXJbnTfv/90zSa3M0ZFQ/iIUTehg1qEXVjn07hng
0EwXJI6j1JBDl91ykBKyXSdctGlKHQFHmYGIMtPOvJjymxvDOvak7h5mQPxmchNDhcZNL9ArIApd
2tulKTzNys0lX0tcWeO4QSHNuTLQ+ig1Lrr7TQzgKWKZ0IYsfjiRmtXaFc4Y91XhqgH8KnGRc6Ty
h6Ai8T+YXZSdFxGAW1xv10Xn8lyib/hMleoIuUxQQRXnJcCUcU9r8mEZtxbd1Ee+/th3g1hs4qzI
QUDiJgnLWig6mCofIyLd69HbWmNfwzPwbTMy8pl3sUKKDwVHJhYT9+56j1LbzRIXsSqqkz2laQqs
4fXr237r0qBj1EC3cJ0JgFiB0JAkrxF7A2o5CoUwXKM82xqEv3H4CHLQAfr0DkvX2zKBw0NTFHc8
Kce7JOD7QvHSydaH50dKZenV0aYm815aYRiCJ+9bXdNz/G0NKeNXQRKcLzrmb6CIqS2+RdCIBpFP
r9KLhJlpNtdXdYfP9Ovm11rCWC/cDgR8CjOu6UcMQKpM8PaoMRBwqtChBMvZVa7lKYI4x+h3iTQ3
5kSyTLjVfwkKnzHcXknm9FrYTva4AiaJrgeRCjZX3+jnyLGItXwm+KmMPMo4xl/k5difoOeZCgUQ
QS04xXgM0unFt6M89O4dkY3AwcCyc8ozRAu4MACnqfzwKaN7Tc8YW84+UyNqaGSORM9IF4f4Sp/E
STcBdqQegWtVGMJUER9cqCiZu/LBuGHBvtKG9EozMZbj6P6HHu9z5twXMhZv05grEacRDaM/eNv3
aWEOPao57WBH2m0kv7YfjJ5ZbiD6NEL1z12CD3zer+2j4eiq+QHwM1dAHBcTeKqHP47nNkt6PQi5
xEa2BCjNJ6/3tMRG4EMddWu5rRNQsLRse/rId70GO/KsHtUaBx9fz5Xx2AJX3TQrKyqHzb7WpjhH
WXAgo0B2MQeCVCDnx7s41Wal3TksL1bV016HkqrGPUI1im6SHH/6OmNxuBMss9W3aL3vSTPK9EL0
wnY/VfzEyxS2fke/zh2SOfn7qTqmvNAbm8MKCRUkkhN4B6yRPZNc5GHXm3cMQ3YRYJVwGzB7J9FP
jfyp1c2CWOmQEg0CbcjwfKdUzXEmRPhwaEOcRXDEnUbRMDvXoVBISe+CEXeZugZAcqwI6xtRkizg
bHisxLB5ZvasgFOT+BeLMsQiuvhDb7Eiw1pOkUjkMpazawspbiT1iu7TyoN0hJ4ITIBQawtluZxY
I7W90FGWFpxs4Y1IT34ybdJfNN1tUL5Un2rjMOl9cqdAILUwjGv4gJRs347YsU83SymnU/AGwi8Y
a8uYssQOaa+WPGGM510ZB4NWCOkR2hUpT/Zl0elSrKb3DYIXzgYYK5CwJ5kg+cPnlalgjl6aYRQc
mS/vaehc9P6JF8uVxj+GrQQv6j4EpfgPDvcgPMUMmDMZ9SpVAqedEtYTWExYdz1zQGeMqjgsfGJn
DzAwzh1uRKG/P1k9recaT31v8bpswZiu1Abbk6LGDMHjW/6A8b8lnF71HLFz8dWOqFFtxgHO4G40
lO71S0DaiJDD/RwYDpX09knZONSJD+51MsWAhIAnjUEE2/i1z25xSXn19OtQijI3MWbmExUcoOU9
PwxHo3eA/Tck1Wmvi/6QXMP1ynT2c//v6VH9bG/gvAE4/cPMLl5RXZ1Uhh8M7f4WD432NizK8aHX
z9zwr389fr6xSolX4nYSSitVJ79MmGQARPIQyfOli+PQUklClQOlq0Ccn1rG1nk1lQWTGojwddpH
pUg1OMLOe+ACTerVbGL4I46Zr2gdJsmPo3r3flhId9MHRuE+I8+/2ZblaBUdPNIxzXnl+7zJa3fU
Ii31m0kicGC08wHxRBVtxyDS5g+4EaggeZwnWKd7JeFEzdFZBXqFv86Gq4CHAhJdKbTMblez8M8p
DLtJ3iSoDURRJkJR44R6VG9loG87sTHTpXEESSPwz0InoCWy1Prx0eT79IDqXFCxOlRD3Ii8VI48
r8Bdi7nW0TEnOn43uPcuWRMsNFIWwUUfIZSERcEQqFyEvwqF7GOjSbLJILnb4X7QIXYFEUiiytrS
3deYHcH8ER9QT8jKdoOIvPgyf83tGFknh4GrQNY+ylZ2BP3b+aV3oqdc+A7C3NCuF5OtMGbS14qS
uhIvHuqG+/gSpZCoQSQHPuhrkApiczfVv9oNkL8zNEXNeC2CUHJw+qA0kg1x4sa4Ri7ozoUtzPyU
XLGgGEE5WvPBssLqVazF9CG+ZU2bspHQ7Iz/UVtUVt0Q1/iyqb28U5nGNmNqUadoKwasNRhyu8mg
vakCWa7D9QhXNDhK0V9VPF+1LrYSExu8gzirDwxkRbMIgnartBhRh+UTePBo5yJjEK2XotFQR9g2
0k98PQEQ5qL5I12UUPzzYSTBGQsXY+uVJMWQRNkBSdrI8ZwflQKEUC9oJE9AY9++lNlWKX+Ma3AF
8bxyVZ7ek2v/6Q8N5jXCpHYbdVIVpgHAkGzayYymSGrvJgroEZP/hSSzILCqx33HCxp69qQYDW0b
b291oHgSukXZJWYFXXNiXVCT+YMg9TG3KhchPSrVRL+c4KPETTazoTnRaphCOWrW7W5IhDMH87gB
eSapTKmTAmUdi7dAqcyjWL31wighx/kpQSGvWEbPHZsze247y1WB+UPZYlsxYv+yslHg4AeBDleF
JjubReBuDpb2vUpv2feFzZszGTI5Wkt/pN9w2kATYncQmEqKFPUsZeKqB6vWQJrktl/qbYBitTgm
FYzjWO2U+ArnsaeCo8mPbckYpl5tXfKgq0/T1xaenrftpgyvNiHPxxv1XyHT+ashcrmVT1G0i7w2
NvAcQoXHUSMZyTZdRE92s1XqPKyMSogyFPkaXtpssOszOSweeepsPd5NhL8udv7D+89PW2/WMID4
d+oxJpAlsDUVrE/NT5w0k7MgzZAyw/xBrtmXwyfJyqtJJOQDGvyz9J+/kghuJqPmXEXucKCe+AO0
V2I73neV8s2u5R6g5YuzxTj5Zbp3Bp4zUZK5Jj/KyUKrUS0LfhrqSAu+6yBWc2kf976xqk3tTpV6
uixjaFG7/1DGy9Dxw2L4rc9qCl+FN/tg0zvViNptxP2qbe59s2pH3FuFy6s7Yg6pXXvzaznGyICM
SvA8Akm4kGPnCMMORbMZ+PAXJjGkm0klanYzVd+XlOSLHHj4fJierkaNIah6KJTfTRBlXrFeGsAe
ktB+pd3KPHdpFoYcJHQen0xG/SQqpMnFHAWZkIvvNmuwzQmjbyi+DSwjfFzQrQCZxQv5qThklKgg
VPYpc17xY6xdrzt4HziSU/+/3GR48sfY2F8TAOjmYURxjLmh485Fm+aLO/WeCfimuf5rRJaNweML
N6V9aHWQ6/qsFHZguXOfX8lWqor0dZn0mEYL/oC3iVdGN2omVRlux4RRTYxdhEX63x7SYeIOpXCo
aJOA+uDH+/CHD1pOc4wsC554Euey81iSMdS5jqX9gqDYNULBdVRHcFI8uy4/PT5qcDx84pI4Qmat
JBlU4o+n/pPiHVGwNbXbnX1XVETd5cMN9z+02N6RtfDwG6F8Zn0ZgNRapArRjeqG1Yf93A10sR/z
PpEgwFY+66VgBwrv4CXwzq2QYrnAwHk8pD2xdHXVpi6x8kjVb8eyYnCe+6AB/V0Yon66JM6Abn5x
eKWJB3ihTgWyj9Pqz9oNql42JtO/Ygtutp2F4MrpVpLoIwiiMiDNSX+XeRMcq7GZ7/32F4zfl5cq
OjUXRcVHZQI8uwlTSI3vFHaizxUg2ou2grioy/nU0udjxN8E7qhmpOBtoI2QYHFpIGzPLULJU+Qy
1Zxmv5EQC1vdFvgrHtLwA8N1mWZV0K06hRwueAkpjXFxJu3aCarZSqlN5dZl7pWRqBCi/UfuEjvX
haE5sw5uTWqFIMfJMUNoFhUo46OzLelogjTAafMuupvZLdrd4J8u/aSKbo/fKOjMYyOwII7H2nwN
aiHBWfcLqvH84REPk93HhD/wYd5HznOYRZMQy2O/r3bLyn5UFa5EfN6/Tnx3ZQ/9sep/lxPCmfuY
C9H7WfdQAC1mg9BE4NegN+TMdd2+e8fzE8P4+dMPoNuVJPHXdURbkHq3IzYNlRtRZM0zAznB069Z
rChEa2UwFX3SLewF00uJbJAX7Eqo0EwLdlkuCdeIOAb27HX4yrrx0RQkDKrs+xiHy1d2OdePBfIw
9jyO4oOt2SMfw2QQt0tSfuT/5HTsNdXhGEWzpBvuvE1ylaG9Fu6hyPL9iO2YcJlsa+5qe8FA5P1o
cdXcKBkJYIJTjH0/I/Avlhfemw5LA4y5kd2HKOoFZp7ng8Qf/NoDL9xEVpNOnWjJL6qH+y2RFa+m
j+Z/+ZOguP+xuvjq5jAPAgGe3QlJCaOQX/SpYL90MA32dI+qAXVV/QjSUNpLuyiO82sJO11m5Gmn
J70YUkB8DD16x9SPjLuA7kkz4pqLR7w8n9QR8q59rNyliHfUavmCACiDgeKaWXKAM6ICqcNcpJOQ
DEfu0idDctfUpHZNb9Apu5uHaNDxaV0Pelc2mlOYbgQC/RhUuSIR9oUE0FopTs3LUzs7Axug7xEH
equ3H/m8Q3vaLFmp9i2rdTmRlpiDpbpnE4I0RFvK+NRiDhW70AKaCeBVXIwllxJXSlFsFzj0N09E
cedimU7zOdLy0E7e6BHbTt9un2rQZRkkvBH7ZHM0bxI8S+7KAWVo6wtY1tp2beG7QDPAWb+KaQ7y
+ULmIOJhP7029hdIwMJqXh9t1f+JptAPvIn3mZCFVlHMOGtw9tcIvK++cog+6JpatHaK1uJvNe62
Ji4FjNpSLUrO8kMAua4bbTgzNMtMB5V5fEWdFvbj1hRK4Cr3b+3UfdHn801N6PlbL8i+hDl52jMC
GGuojhHeLrNpU/AEWs8PqWVsNSn38j9PxjI7LYnpMEPTMI2vdWUwQqqF16JT6lAza4c/5OYxX22E
aJiMwWcg1783pvD6qF+fvYb+fmDcionpIq4E8X84733CFVbnAgp07H37abIViX6onKjV/4gmTDEG
eCvxWBdAaFpuRibgUJkQ/7dfID+wYEbb0tDev14q2SfT/0opFI96uShKzfFOTxYkLjp/ULEH+3Cr
oZTjWt2IuYQKEv9vuRbQ09joHhBLjaG6yXKs3B4gxnnVRkckQ5dDwwdDEqE2oUhEL8a8tgl4go35
RVAh8Tf+nAhJoCVGeIi0NO4RC9lfZLaKYhGxB+nUK9bLRylV8VBNGC/DV2qW73Q8WKDEuIpa3Q5G
uimVe6Rbioe5/W87ejYi5cPCsOyW+FhOyUstPeBfWMlg5K+S4URgDuslTe1U4c/1FT0dv2oNu05Q
tgNGDqqI567XktROEHS0xfqUx8tJPGaUQHd6HuC4/8AaySSxi0R8nwd3OBObIP4YwLbeOkKqgI8Y
T56fSzeUW1SSMTHPsQmFo7RbJO/cRghRLHxMDXSm+Se7At0+j0VKv5kQCKfEwCmZLyAK0g/galw7
pv66JEmhrwP9NiFXgvSd20Ytkvu/WlFV/H5S38+s15vd5WaJiZ7nP5kHvj6blIzUqFr4K7JmAhPq
jNJK4q9/kPe7r7AU7oUxsqfs4QXROxygNT8C+yWtx3iHKdelZ2d7gb9/KnTE2WhniDHOPQ995J7w
s/S5+ZSBqajbFz5DMHnNoyvKbwgSd8BZG1QvKeYupQViXqK8R5i91ZNndNPoqSFNa9ghqC/LXdV/
czfk6CcZ/SGVAlLdi58lh+1RZgL4cKcnl1XCIs6G/PDcugapbLU69GILhkOgohZKv3ygB1a9osQ7
0g45IHpJzupLZ4CLNs4heQgnSfSu6+PVSuzQx9UXyMHRjcQ0NiIJRu0L1Z78wMrK5anjfKy+YTRT
rQ3SDuTYm6u+J7fmpxxfbOopZNCTcyaAE1Jf5q+6dkojQCHppkImfu2FncVCsl9Hu/Mt3f7qWRVh
kpeaWncgwvfy9z+pn04VRTSchJyFQrCrmjVCuLf5IWd93ova4D/TKRTVjQYHUA4PtUSwDxyZwHkL
Fszzz5zQZ1EX7FDow3t/hj074PYDsZhV6NiFfWlZEqtf9xhRa79NIa//qv7eIZx56yklfVEzf58a
ax4dyRjGqfZxZxXLZWJYtBIEtG9bNSjyIf9/884L7jm7lJ/XPWanjMjRN3uk3DpMwx69zShODnv4
ysQV1h7Aaaa1QVh+u6BLX/WOVzpQE5W9ihbE/pjjTl2Xjly3NbIOFzkZ0qVZWBXdwqPDf8+THMes
P/SNe9vzLJKlV664vwWup1L4VEyWzL74iFjOPVSWBf/4hMml9zk/hmrmJTYvvVrnrMOWSn9C1eKf
Be/fkr9ZJkHmH3DS1eWomrOzpQ64gWeqMIadt/ZU+BQLCbEjF+pZ14M6BVEamyOrMeOZeYT7Rfkv
Ig76ke26doI7NWx9BDjsDvPOblpS2vCrEyUnjeka2jRWeR038X3Y23aKdgPdjjVnkfARAYr9YHpE
n0s8mFZiAjNydTdLwdfy7IlixwhbBM/hfCSTKoTHmHHtnyBoaEcq14VFDOWRleQzFuB+lJW0q5Nd
Ez5HKfKt951AdB3Cgc3lVwo4QgutwSYj9/o0ZM+07I8u+khgHMK9Reqr5HdHtEphTBEKBQUiEn27
fqTcTCpRfeHUeB0tWq4yUbqSHZFJ0nb/+nDAspG7FVxEnMs61eBa1eF3ycO2WIzu9lc8iVjpsMPi
Rl7AN+fM5+SkNccK/lkiuP44L0WEbADXNSl2gMJdPmWi1du7Tn0Ko46K8eVvYIhQ4JqWfhhzW9Yf
X43sPHICvtSffbzWgOXyz5Re4HCG3YunCh9oSkiJw7rkM8PJe75I4/cinw6Bkio7B5KsyaLo6Tjq
Awt5hJ9FWrPAVDEaY+6pU2nI8L7xbgMXViTGBiGUiDlHrzOa+P11ZE0HzxvMC/SAkgTMXAxgv/4D
fdtE8jX6eGXFKYAeIhaWA04hA4BWIY+jiFJQMWjBlf7o0UUFHvcudTcSs1Zk2Reh76nRlqT0u8Tj
eTsTuJegG/D6xpsen81d08ugZY97hDgZeBs+e9P8JPU37DLpaFEmdXsLub9oYljCYHObZrgtFHsd
WCAtTqNrcR7cd+FMEgC7GMtC89fRiO9KdTeRTXknSuuqlugbZ/elGiQMG3PauQshZ3+OLxrgLshM
adV/uKki23AGGt83KrSZScZZEOyLhG7fNXsWeU/CN/edsCusYcm0LUZx4pJvg3B5vIXw7jBMYDkA
gaREXiBgIAeIW9ZgKpIMsojjlhy2WBaX+yeayqDx1Olsd+cv6vfdARaWFU9gefvN2FzI3y64R0Br
1oujA+fyWG5STDtnuLobMIE0O1zzznsQszB7mlnknhyk/2UWsksiB+rJjOOIVMC/4Vo+yUIw6BKi
/gNZxA92Xvso9pHHUjTyMLRhVP0RHJMTi7HI4+NLBYceRnJqmarpJGMt/5jFR+EKHBjmYSbS8mvn
tHHXSvkPDFQsicx82gVsWutovq48061WONhY+HmyeW0WGoJ64o34K6zRrkzzVYYVmg9k+jHtkrzO
VMpepfeE/fSKxV9zhXGl8xy/OAjSCJ2zRQt4dWyy0OALreUb/xehg0f+6FxEpe5awp3mvM3nmctc
fDqhDKlhMGfzD7/YTde681kIrJ2w0cEtfhuKREqG133JgDUYquxXnWt3Sl7OAWpxpSznD5az++sY
neC3vXiGJ5C/wOoHvUkC30kpX7naC7Dsfnn58ta/xchht0kFVqpvKS5FP8LDgu/+okTtf8XSkieq
Q73Yt8M3YTj2lhQ60l5BQSK9KWE/8l0jAdCIn0TiqH2qsub7/I6Q+HzHwTz5o/p2WixoBEMNCG5W
0D+OkAUNsS8eiipd3YiK0+arP3ouzgjvBnadk3F+Vh3T7cYA/soYlO0ij20rGZIt/EQ/v4R8GshE
mfK0iwYJ9sG0XoXz4BMbjwW+KdO7V7amffAS9TX5Kyw6TEsyOoYUorbJ5kr92KNDOcAjIa5pUNq4
nvRkLstOEFpmFBowZYpfpzs/mpQjMuW/Z9+5hSgGOdXBHsEbXDAUq+sZg5KiAqpSp+43k1DcJMRC
w7yxtAog9rAH8xRhfLO2iS/cQOReiFO9YRBOT+zYXML51Vz9buGOUG7AYXi2HBg+yEycr0QaKYIc
9FfdmqUe3YQSQCDWSbCwFRA0gMH4XwfHxTjoEdQK1yHkIY8eD9J3oMFg6cS/T+Mw7ez1soeKSDMX
Ke6Eq6ow1Z7MCy/uIAZ1fOGs8yvcnF8b8ityx5wKyHsg7m4We3QpLbT405Km5YJJwiyQbnjRstFM
xNZNpE1SKhRf7Qdo75+5QtckRN/dhQQjEaSQ/G/TRLjeH65ZtYwxOBOXzRGzhN4PpCOj8GCt44Xg
Xq2nCBmVU7eCLQm7RFhpgqyZ1ILBVKHLRu1B+ZDam7I5QAK/915CTjHe5wQEokhmkvGTKh6LcGWy
lvt7fgc0HkJPELu4gi39D09/iqqLxoHdnd6qHxo2U+zMrTOAGS+WpPvoObFcfDG5nktLnLk03d3H
amJHzpWwZG9jvM2857qaJWvoODl7MxRE7phGgbYpmiw+EgueYsUC4Q9cVQ0OF84tRLkqkQ5+f5AK
7ITL4VeWKbsSdieYZ4ucqELovcnAe00CFuGdAtvOXEROhZrNMxBfzVyspFnFMBJqCsHEcnq8hk9x
fE+qRFRrtirIGr9Ld1GnhhfPifUso3+q3ug+zExO3pqCjXt21Pm7b5syzSST9GGx6IWSc4PFcx1b
hAxcvNhcEf8d+fT7P8FJn3j4ygBlvlXemNctPDFIYTY5tkswK4Impr1Ita1F+GtZ73akK1WxJkQT
ed7p6fjJsHqqorPCmynCk+ifg2dhsuJ6YBJmAD57XHv3/IYAgiOkr7zqHnwkWopzDtCd0auR8V+c
SCtx2xW22HZNl3q7jiBJRJLKUWn+kF+4s6QJYrnwyHOQuhpNNm7dL+e4tkKIXy1/NfkGRhDp9wjk
N+6O08TM32i4XcUi0c+BCojsmr77yqwFjkpbYqhd13kVc7MliTC4whqvB+ns7+bNexeQ02Ku/8Op
Jf0VPZ9jkLPFaQiHrycKj+3b7GhwP+wbdGOoM/UeslmCYYwmRRA+sSIPntdjJJu6SHLjbGwFAzqj
IPFngmFgzsWIUg4EonqZSAcRb5+ivrI8hllhtgEAHuwEV8QK6IOdoasdLylb+1io/rz2B3HsIiFh
n3zU6IpFC7BQeDM0goXndNQKWS78Ojv7G/tVupOU12g2wnmLdbc0LMYp4iVSxJGwVdEcXSdPVsAA
tV/8aO+WYdOkVCZac5JkBWpwTKDmQmXhEspJ/6kFiJ1CQwNVg7hBGzZIRLXX1p5IzJogEMnXan1s
l9bk1zNPFCSlx2nBo7uJHNO5fY9M2rGW2G+4G8LxDHfRPExIiJ41Xib87hK2+TOZH979ARa3b9p7
sRkuH7xe9gKfqsYi+UStxcv1NGk1l+dSysUroPmCGAAgGfLV22EtMC+fQCoi5cvKWzWNymtps8l9
w6gbpy0pzm/NiCnWNugv1flDIhfWFuyImZaWAqwMr8D940FE5CGfS++Jx4/VJVnnjkW+7a687v8X
XucSPvWp8TpJPQiAm/Jk4q7vtwOVZd5tjMlcQccpGUaBsNu0HNi426tk411ASWOrxUTNOTaqYu3P
w6YYULaSlhatxCUVCPlut4ZHsDzekslDPLSo8ke3r34Aq68rjRPOGj94upFt/qCYIZ8KVeLz+Gil
8WQj7HFBeFoWnJ/CYJIy0mgFgk9KrCN/S1F+jbJP+Um3sJndJlt1S/d/ebUILhViNUeYz/cWHh+G
oQD4Xy09i+hBjtTYCFr3JLBpbX6+yaAfU8AWHbVSeT/xr61ATk+f72xUAvSYqmo8LUCkeLzOjuzP
3jmfORbf6Gx0/MQOI+9F/xDiii2A1aEoeRPK20DNzqnZ6qbVQKUPpiRvIgf2buYenuXSJYbGpKH4
+cKWl2T4jrhr4BTDNoe2dKxtfWgi/dzmmMoE0Z3CualMQzVAd/HjRSDuIB0PUhaXxjaRGW+c2pDQ
TGgydhE3/lATGZaw6kd+zr1JaGduldgdhmCo82dht5CbXmAfiuBsScOdWgHwVeTtUa0UveBl3egC
d0M26g6BU033+2qdaSEQ2aFgCJIyoIn2YeTuB2KctT42xI8EPyIqS2lo009l2kyhx9T1WyMPc+4P
In52CSbck0Hdbb5/i04USUMfc+/m7bjpvzDLKelTEFwNUzXVcgyFO41tfgVShAIlPR7S/Vkzr3FY
4T640vw/gEZa+ijyfVt93epDdmanA5NtJVb8TYmwXwFAoKBZNvGH1grnljDQHcYS16P2XxW6PKkz
gJV6keD8R4aQAgnVN8P+8szCNbzv22hr9sWBqZbSkL9zQcxXkBYmn6jtj6lCKg3AvnS9jfy5CZDV
l99AzFs+Bv+Cx5wuJ57ioshOZc9eqZ9N13mjA9A7FAtxhwEklHGQi7ZA0Pc4X1+B+SKnPDqOIXtc
o7vraReunqUn6It/7LHQ9YSKLdflFvmZo4ykhlkuxTLXpZH9Fu1eEwvgm0o+FapClW8TxvhY1yZ7
3o0unbzs91OWE3pIATKGQtDMAHMY16aWTrEWtIoi8IHwc7QKS9mprQ98nblyeSaakZ4mI3YVVrqh
vmo1PYApTy2H0chN4rEAqAw4K+qUNrpIG8eTcgoTpg58VHaM92oe+HVvgdO550gWX55yTix24Pfr
hO2ADCWwzAi9OR3WiBP+qVcdQzCJB58mp4/bMgK2xRgrg3aO4K2nETFN7uu0NRhgO0mju1O09cq/
AOj0a7kJFQPZ5rvPVY9WdMMT7GY68mCE2+m8kJTMtfk2YPxXV+WdCIDvTyZTcecfG5bnEcjwJDa6
V0cJSIREDfrB//G7kpIe3uuJFm2YcZl8DR9wlXzT1ypgUbVz+JDVWZun7ARmN2pIbZiviQViNdPr
JVkpJhJqM4KkPw+wy1tR6DvwUfSqayiPtZ8Z7feOwlQ2lOCk4ofzbz4qKygp7h2HDNquPkMarDqu
hQ0GAuOd2kOt4Im2aPmKOph01auJ15Ln6I4xff4g5rZ4c1k9yc3bd4YlSqt2Svwx2bRY6yoRTC6j
vfoMWOo5kHML7o4BcrhSsAd/pl5Q2FA1ZLEzn0RFaPNPnLh+mEqKtCF6u8SFy99VP8yVF2SVIsKP
SGNvCQPeTUVP7kdVq91gorIGbsxacFTNKE+7VvFSzK8Lm1qBDScbnP3IrC7pr1rtAbD339D+14Ts
dTPd/vpmKeG8S21N+rEQ9Fe1v8a3DYqeo3eHzuBsslMogPIcn3w1BRljON1g8WFLdsL1lyCX+99Z
yEhWzYDkjUYcrCX0ZKFxWSm5O4JxNDEYGLPLltqwCvqiIznP5K3ZPpshbfVy9cGWI88exiflu3Ot
BdUEuxOz+9JyuQk4RofUVo+HnhwDXUNN7nUd/jwS9e+vIN3GLfXWyZYa81g2lFvYn7ybqUwMqvUJ
WsO1gDdbrAFMBFw3M45fULTmkxIt6RKs3yJ9yEvoxSLWmH7gbX4FY3V9vhbueNLs+wUt7N/u6Eal
zadeaqiSrs4CliIoL0sOpJIq4TDHIitifc53NlgqM/GbnO/wuVdYbmCu29tkWw/7pRpg08Rhjcji
6H3KhmjkwLc7a1/Qr6sADW2rSpD5J43JcfePCXB3Sl130+RNL5ZwbKV+Vf968WX7B5MdEdRE6fzW
Fhf8EtkPKhYRrfjGXBpy07PeWtup50FZ4aV2poIRQEYgQwnHeGdfPYZXzYgpcwy1oH6ZWQgXgE09
MGhpjaezqvPNKNhuHgeOLq8vDup4x+C/HxeXtAiwbNjjcqr/F4g43XI2IknfTJqiOccxxk5z61FI
suQTQ6Lgip1PJ5uZT67vVqIBBn6auYy3F9q/LEtKQYDqg1lFgKVrpDw/Xkql81MvIOCQGBydVm6C
u7D27/jpZXgzvlv+ftqSGCgsoJMPbXgvGGz0Ge8J13xNHxF3Ue+zY7srqtw856wJZ6jl5Xq3y2t4
vnhIRfrkdUdD1rIWHeSbNeYUMOm6ZUGH/qCCMgrJ3Tzz5zAvZHBISvgEgq+OQlv25RmbaPlRs81E
zpQNls3s37kzfvasoGWFwCvXPgF/HPzE/wpci0ZSP4HK+gL7uAnwIUAHNYp6sZXkt6MTosjpXzjo
ALQWJ6WgAbZQ+YAK4u14XzFkKxbjRf24j7sFlrxxe+c8xbttIWxRfwGoS4oP4TfWdegSmOdcHvyY
rNYVAYOJkbDMrZjGeDn3Vm1WW1ksbz1u5pu8rmmL9Q3XLX4LNBO/PU+txLhB+WL1SfPyqXQjDisj
Sh8jKAUgGUDA+5cDAtIetHybyzHHseBRiGpaUYh3Xi4DQ8xmYmlDCIZiliN95bWiinuAHRlaeZen
7VQxY6aWXFe5NCw5I+f+NtHT43K1pZgcVXSolm7n04bjvVTWpJfhbigMhr1AydMN0aXfaArVzJ5a
yIit2AydkPgwn0OpbNHhBD8Z6aI//5uxjh2lM+zgArqgh7XcPbzikZOa2Wr35xCQgA0VDU8U4tze
XlzAFmmM0yS3j+L/+XJErcdAoXqmIkP/VOLc31bDTL5fBqA6V5U31QpG8CP42beYjaJX6ZT31C6L
slZP2vt7b5MTQApTuiwLjOr+ALSPTvfa5b1hHV1YRE8imBwbaR0jWxeBZ6DdDj91FuOV0OdjpejS
yWB/WV7IT0l6pRy9IdZT6TX0Az4XJ8Xmj4HiNX1Lguv1MGI+z+itoTWcMNnxA41XyxCXgwSiQ9Cf
DgsMEr6HTomvKQy4j/02xY8/IXAwX0v+TLwQxCVKvTuuoiJiX3QrOq2qDNrgmwela6V23Cidc4LN
V90eM9J+HzUcLs9M416DLMBZdXfYpkD8SK5tt/tteZrSo9Q64C34nWDqn1IV4I7WzusLRn+SfmPR
MB8pHngGzBDS7zC2A5b0UvcP8qQjCIQweR2O6XYQ8BKJ51WHXwCt7Sjw7uLUgKYLqnBVusR4IzdM
QRIBhpc0vNfNI3xH41MqQnYuzOxgoYkBcQdcmTIQ+v2ERYp4molOYGZQf7aiBXKSoTp/J4HPN9ky
QA0pwxbaoJ/TtEXw2cvv+3mr6XriY/Uk392tup/5iIcG0fLgGD6n1VZNCc/SbIn3lfOHLaWwOWSy
o6LQYgMTA8LKgP4wzejIpL/+ltkHb/ec5ioa3oK8aj8rs38Eos1CP05b6j4GhTKYMFVvKNEgt4cb
JrMZOO29NeoQJsqTQsMxuxWFZ81rmoqXQ9UEPrQPJdi5/qAMm07Z/WSqWywicgNxxjDefe+jPjeD
i08542aLrs2ALf3Z7yVBn+RE66/aAE+xu7GYU17JwhGGyJDDmL7T1TVidr9RNgaDGjO0G94D0una
l9JpOhIFYYtPgPcUiBBkqRy4py52hbntulmTH9l3TEoMtOM3nt2nGp3wJIT6Zk0wxI33xl+/WooT
WS0bniCkbm5FD4UTOXSb3KxtV112tk0e62TFqb0MS3MUp8XbjoaGsJokRYb/4mTdDT2w/zOIymnH
jBZh0A8/DW6X8sDchmRGGUJVInE2ZDoOT+Kc8TYLnWn3Qz3UKE28xWvajSMDb4qFwrZa2Q0M+B0Z
HBupHJ/+apP/IcJMd0SZNhl4rgq79dEIROcbnSGGX5v4mq/6beRA6848YbaSu6BMhhC65Mkvr65m
anLsDJea0ZEi2drbBCxS+TohH2JjcwnGWmiCt5t2i1G5ms7UEZNompY4qC2DNIIv/1+aqPd0DOrp
ZDCZnFSHAsE4Z3UtqaJkWvLCFr3NpZHIL9TxlzEOdYRicLWunaMJaDM0C/BO6pJbeYSr1yYZjtKK
ALr+eGlPl0U8LXzMuvLrIgOBRh9ozZaZmi7VcoZvo7LrhI1qdbGdzEUbnA3IDJB81hdYal4pRZtl
7Xva9tHqixsrqWqISGJcXjouBVZ888BDlaO8N4isanOi1nfMggKp34NvLvEZpLbodiw8Q/G+W67B
Pq6zDAVMRpJQekQekcNeI77OghdPkEX1/Qb7BSoYQqcsiq+Nabv4C1Krr7GunalJr0bVLEWg/+gZ
1bqLQtCcb3Q3lWzgJuAdn/ChEbgzmdK8zC3VnbMOymkek2ZCiYfh9fJmEtFYQpKMrJ4hXDxGBvQL
LsnZqPAg0YFdH92V+fO7aMDJBErJlDb/xf+j6RugYUm8Lh1zSUf3NIRPxd9uZQsP+ZsFH46Zgp0m
nldK5AXqk9DdNXU5IAUp+O+qZDNXy/af34pzIh7D+vcP+nnrnrOI50OzxYkQ6SGEzrGo53CbB4nq
28I40pYO1eu6sSwD0VOuGx94feVZDijEiBAOYf3DoTEOxyzouzCFezIc6GHRB7c6jQoE5j+zpl2W
7z62QkOTcroZ715Ht/+aK4dp4RTMQ2+vEvL/SPqEUPJXqKG4Kw/XsvUrhOKsh4JJU2980+zVgL2t
5XjXNdEYEnc6bJMD9H3Rd+uMflInKbiFYHHhrzCsZH8NxRnwcH0XXcrVRWVDmui0QU+dfgMffZ/G
n897oYoLaIc4Srq0r3OWlh7oo+CtcN2nTgPLyKxmoD1lJuPZ1Hk6gT4sa0jd7pBzbx9MmJ2zP4Et
avEhYNrW/zAfid6UAADFQUWH8mPJRYtaYbLNk0pt+LxI9YUUSWANGxb2NCS6TmWu588yfM6x5LNf
j77liJ7KFfur0t1Vu88BTTEv2JHb1knrWY5p1bpQe9zdjLPC11fjRhgsvNVtHEu1Y4GobOK9L2/I
1KrGMqX+5RYSNyiMCoQS3xdEOazEk1rhZV4PBVWFIFNipGBTiO/pA1gvz3KN8SeoLhZ2V4Ebvdiz
SvXT/h/grDxs2/thRipSB9IJErYnPQV1rBIatCQ9Z61Pkaw7Tdb0p2J34NEoI6yE5DtgIzxL1ggp
EWCR7bs/wgmMJfHkR4DeW7wB4V63nGsPubPmvw+yOt/jL/SJDYrPczslD3PpsQxPq2T/upWVjGLc
9mYqihKxx4sm4IQJkwtUivyd9ZdRuK0HlaZygtM+A+d8BaqxPXCA4jvSuwJnk5/J7eskGPW7VAQi
bzntDgvluL3ZZkW83/uU0Pfc7nHvw57gHBV8Xsep3+zTxBdGB2a+YD8+OfE4KWiQvb3YIPHePKpX
y5ohDzrNNpGFSEHe8NPLIuWZi+Ah3Gbn9Fpcf1a49L+vrmWn/2rnGrkGh88jt+B776Fi9CxB8Snc
LKM26DL+aJUhQSM2/yaTOpLG2JaEluawxvf+Fsl4k3DdTXIR6esV4pDrl+nE1NiZ6Vd41Qwhx31X
Jvhw4+hp8sso7arP9+175tY5xwBR4OCZt/KATOgSXRdWihPxN0ywtJiVWSbhcZHycrSZlhP3PHPZ
N0T04OEuATZ59ZpeIXMDqtgwyAAyujwk4kFqi9ivbzXRoCyoegt1M8hIrZbjYXc7rtHbovREeRZY
+t8XBr3ZVEKM1UxHXz4AE/t+PbRrR+BwwMhu67NbmXAzrkKTD+2qcg/2tO7WJIuifRPlhRasaCNt
lEmy3mwQemXMtOmheaNMXmzJMY3ZiOzMIGdXZ9AmXvEtb5nqsV0Y5L2NdIDEMouc0R9FP8tqH2M4
HLK+5LbHL4FLb+ynXIOp+upWQtcYo6wCjc8BNO/pfhrLT1ZHNNwIAtY8AUBb0xrvmzzgIjYkybCP
MFgQsvQT5HdiM0AeEKmpHo6M9DCnWKVx2OSgDHYUqwI2GN1Io2T5Xh8FcgB/o6dj2/1cAZH3+VQQ
8kObGot83mSZ/2UylwkRPSNAAfKrVXM0U35FIm7jzXRewpon3JZ2Vyu5kX9xHmNtCfW3c2JxhMfl
0Vo3vrAF576lRNJtWmn6j8OdRYNBd/FUG69UJIXfT4Pi45K27UpYm0GfyUV5iJ/ologEK42cn8xl
sm+HlWp3lDY7Z0pQ6/26n1+H3R1vFSciozx2JHgD1ZQhCkeBL+8PKnDC7WT6NJm8uHu6IOmsODL/
JFAw9TbyUSJVTX4+Ng3I+sIA25052KgLNAQTUs9HTda35AUnbHPWVoGHxRcG8t2u3hIgM7J1uZQ+
EviamzX/P5lWhF2QYqEhQKbfVQMTmtt6aOMNFYpAB/Ukc2n+FehePmVeOU1l8vGh64dUo5MZf3It
7XzVb4WnkOxfnOkGKgivclqt8J5dCUGIlBUvKoQNVtlFFbQ8qCmgBvDuFcIi2uZCckZ2Ays8gFJ1
RUfPecPUtA4aaVUpDAHdkkd6SVJjQwjCxrpvyVHWMbJoxFMy/Jx0zcEX81tdFj5XmhiqsXpnjri6
BvNHH9ZsQD42J6zbRRPG+aWKOz9dyOBtWbEPWDr4K800AXyGz7pcq+spFjWv5JSA6HL8ajzEsLMr
Gln5PAVlskW9l/fZQrnl5I9tj6vp9410QzL3+u2Hr1RjT4SwyBPGPKOheL8jIyfZ3/jKABpuD8YI
YRq5qRy4Gk3Q21fM0viHXSXPlDdPDCkXzIOW75ETOyy1gl4DhTFJk8C+5amonaW064Lf9znPec0M
0iAQaoHqLMB9Fnws1tktyjRNaCn58u8lv8Fe6bq5HnzCEwPRGfjNkprBqLD4KzBdRlAisCviwmxQ
l8w2AQJ+TBM7UjWdThMojFU6qC7gDhVuc7eOa1BTJ5HM8Nfj7BVFz/PlnLRciy+uY/G2U5frfS1Q
g9HZGVyXolYS8Zsr+l48yua5/msDMKA+P4Geg7dzp7Pn5Y7Bmi8kSceQ5n3SOqiFRAggKWem+kKM
eiD0VKRO8bbMl6Bwcolf7pOu8TBLenDr5EYUL3JrTb3EKd66SR1SAl11F2zttNl1XRWOs64qtPMJ
6H2fUCDDTILAsmXeEZTpUpPYJebSScTx2ax4AQIddKgABS7YGXqmPXU5jzDSKbtDN1aO0+NuOwpk
TW2ZVibxA8V+fqcge4Rr2WOzaWXXOuv8EGp80YYrTr8/X9B1aAltjutGZ9MnlLh6UAPqQVBWTv0i
tvwKqYExkZulggfrVA79FuvMD7oz7OHOmC3KIq80OCvF9OP/sXU3ce3BFzW5uYWURvlf4x3D9Ock
U0e16ZYOCT6Fhv9rSNsyX/LnA4Tj2/rw+WreMTljKw7+TZjfeVPdiyJkVIQQyztKBSrofEO/O56K
mGqCWTV5zT17FR+D/9CiQTPIuZ/UaDltIkVKgfMTGi599GgUw+919wTsD1F8sdBaIzcDlT8HxBjf
x1P1WCn20kKJEHROiUd3M2gUZfEWPPDGDqF9ThJpYC8S2cnA53U44lNb8Iz9OzCt17klY1QxzEt2
flfiNkn+AfO0dtEqpluver25BX7kfUWy39RyHAlv35ESe/qmHwH/EApVAkKhPrwmVBlykEcjMelu
fLCFEK7RaV/FPeUhwiMb1E66Sy87gV2HKEzr+XgUWZ+M/P0RYs47YCemV+KLlduSaeKzzKNm3sXw
yxbSf0P3kJsBcx5MXFwxzagqcSUxlyW9yLDy1Eix+U3rwZCt03IdgYSqsEMdI5PQBo+vtWKyGqzK
vnT2+WmbFPPd0hdwS4L65ofKxB8PnLSdvDsrYMCn+v1NKs0vKtZ6RPvugUIdhoPVL/UYDwBTMW4m
K/bgtd72ob1Jmvf3dHGMrbdUy4h/ebgnfZQXTzcxtvuKqvOvW7Z37mebBYzjVuS9z3X2Htc54xQ/
fnHRFKxOy0gcJ65TvAc/U/WMv24+/ZZtS3y+3N8rSDAQd0DKFJWnn9sVH2O5+NFn6TZdNytt4k8B
qZxLZ8Lote3L75KZUf8gvZfKt4Jv/XaF+82VNJgEs8/FI/CK25Mq82Ab2+FEoZfs/K6GJVr3OAZZ
Z1c9rToBFG52oM2H36H1Nn6d9saLs8kDAuoZplzUhz+ZqIx6Zx2Dr+sXu9Cs0AHgpI7fRqwTIEyA
vHtjPaihLMvCl/WxV4qzdBJ+SQCkx8Rtg5g/2pLLV1SDaV+kbgVMW+jBw+03AL9M8zgjiw+f1wUT
dJwJxWth9PCK3GS+prxVbr44QuJupCnNa/fHsc6N2wImp58pl39gOsLoilZScO261ohIIRd2ikIU
j4YdFLqzb2UQHq93LK4vVcZxcsDIvLq5HU3YUO0BTjwYB5YMNUUe4dopPF5cogOzcAr/U/qJ2o3x
r58De+1bwzl25tfAnT1LUcSFxq0lj9kwWSaWLIy0AH6gw0LE5+6HcksdAdFFTedq6ut2d4dIOgSQ
yO4+fqRFIZEmVNyPeSEWgJQYYM8UNJYoySxG4OcF7tTt3v5TlEA6bloifZZE3DR50MEqe6F3NAIx
fS+HcuR803BqrUdBxY+6UV0t37CiRFoHT/ZzVki35sKIqTZQOeMJRSNy2ivYUQQp1A1F75HMPsiU
WzOyNyss4+9ok5aFkWSw+WZoHGBYZBvV5JUtNNgK9xt8uCOcVzms2SVSCry9PNIXE4YvKiTwkEmF
08GaSRENH8DDiJElZozoCOJ4kL84lPDphVQ+MOEwrkI83Uyk06kjcp9roMFeANIPD3cSjE29aQ6S
PE+uyFmqKLnDLtfgUmaKKqEV7MFgSDAzBmNCBfya+frZtt0n7j2PTD5yHveldvaYNQfyN6BE5Ec+
xPsr2DJJp9XfHzV/c5V3Q/spXEmSnCAz975KbJofPcUBB2BG0TpSImF8lp6FrT4s2oR+GH5905UR
n55pSIXmjZeSyL7SeTqMqi5ikEQfNFlBKUwCqKn3j6WPJDvhc+FqyqxmrfTAwcpwZGSsrquS3GW6
fYOEr7O8mpkvuQZ5orXOYlGYBi+0yQqhw81udVjhoxvutk8NIdiGQr+Ks5Mu3qDZWabwm0BeCoUg
VpsCQSqhV8ob1MnNhb7tUUATtXpB9y3MSEB/aoNZqDS3kaaDZRk3J9RSZTHX8ven+9xXvC+31rQ/
Qjtan3cjqWqVqjVO/x+wY2NBB4XmYKiO2BZ9h/N7V+E6qRlj3jnDWN+mZfH3Kvd4+mvpKcCfFe7l
oM/Gs64W9AxXbXeSMzLrT96gitM0uztdItW0NGHoH/J1LyfI4GXM2y6965lyNSwkeetaWGCF+0Xa
BZWv70Zy10sdjTguYFGIDgT0DRDuIB8FnaxihiwNGq7vL0rmbFFWto5S+YYuIBBQYRvOZgsrqtNA
nF9HBiIamXOgKx6HAEGz4TJS7r83G29Zjqv7dlIY3shT71jOSNRe5d5gejFh3E/G72AMLLQjFiF+
i1JqNyJ1+8BVKKKygGCUXAsXL1Y1qcO/opi3+eAW11/8KCrrV00CFy9HMu5GEdQ1nGVwIBbutgcD
YFgc11KuH+2UXKjLkNR43jAhlL4O7K+q3yUk38gLghdA7fC3VeE7SN3k1+P91jQ1CDsSmcCJCpiN
1mXCFeQZx1+6pyvE55E5ytiVefpxXwDZdpmw9Mg7lGe7ti8Zl2o6rJ8Uuz8VfVW7MSPcjCR4UaDT
rdDaLfAskLIoQiHTwozWrL53M6V3fBgdISDuq7MU/Kgj3WDfEq2rSojQmpUMfs6qKEe8idCKI5JP
CTtM1VtLsVUCjOf5mRSyttE7hEl1hYbJd3jM1H+QH5WpfxygTRW/N1KuUTooFLXOgxzlsxqCr53u
eeRgROceVCkDmNSgqsefATUOqiF0B46RGbJgOCoaxVGNlw9DR/so6RNuhr0jpT70M//AuF8IEguR
yqZpFKGICSU/p2nr+2jH1YBq4wLJxj6HH/jQ+RTdao2E/gmC97wY3NsEkltpJUYqYzbVrbplLsB1
5axMMmzc9UMOPa45M+N0CKAdQsPRgGxBcdnmW02YWebRSC64I7aDg11J4fNvRWDEitY42CJasgcU
FblsPUSj0QfD4GQCGbgvI+/EIhzxQN/PUcZAlHpXhUjWmXNRjIBHpit5YKFbTzHR5lKc9VnTdR5S
4yUx3JH76z3Y81Y53GusI+xv5kCHoAIZr6FL0Av4YyA2NhQLeuAhnkRmVJAwLWcBnxj6ByHWX/AH
Jovbe3KPKvzQ7YkV1TS+/+zToUftC6rx4LoPaouW8uMNnvvDWF0aUopyQebvp5vufvSXwn3/yuOO
PAnYFxp+puF2QENTUguEJqTQHsUmTvElyLCimnl4naMJRFHP6vzbsBCOWUz3wqjqB6IWeY63mds0
jXvPo29CLhpxCvdoTfpcqRpmDqUqVi05j+eLk2EOKq68s2MMz9gbrpw2cYFuM2Yz3HRhvty6wLiw
T4WAXYD6Vs4byW+2Ir6axdMs0BUchgy0rgZf4M+qREecqQIAsXCy+82960JW5iNQeY/FxWPQGlHV
Z+Qp5nsTJFHH4B+oRP/56KgNtdk/x3Icp+bv7cyeQWDaM7Zvzn2Ri3Lx2fWFzTvF3jsl/B67j9mi
xVTXy5ccNVaLFRGCDGeKFKDI2udmE9Tuq+itwZX9tBHu2f1/7TeMo6fJnB0OJCsTYo9oA31BLqqL
vuZmXKNd2uK3SsBSLGdQx7UI5kqGxXzKADQUik+VkIceSY3yQBDpnUhF79jp6fuXca6Nv6Io3oZj
7edYCeygFzTMrbc2cCLr5hyBtQEpGqQG7rCGifCIPgMRi3Ebik+f+7DU0sBfqcWx+fujdZM5w64U
n37csb+DDmYxqRh9g9HHnlPFWBBj78pgvuSeoDsD2gsTUSeyQABj2kzP19wFK8fivsIXhVOBo8E4
5v+5RfPAapNosUYmISnH04pB+ZO3VwKcR3VHnY5HA1Dtez9hdtN5mG4unmMazieX42z/YjFuwDLt
MDyRf5Xp0Zmm8ybQpx8XDsKjCwlml91zy3JRnwzTZOCzy9CxQeNWap7SJLKaczwRuexcw1vZ3il5
hJGkDyGrLxCxhORWasGF02egxuBpBM/jgwrtIg5YpHDUF/wQTHkF+0TouE/LdGYkqjdDPyfVH8k8
p3S00gXUxbl8NIJX6OhcW4qj0mnrguw9iUys1YIHlKwOR+f/+4F3BIoWfUsd47eFwCYypdkLDHfO
kSioIkCCkKlXVTQsLM9fNlXk4brPZyRLi1dSn1z7Al+EvAc6oKoDUiUTfAkRBGW3V3rruSGr53Zc
6DLa4DYmvWc4vSw+VirJDvBVW0taaEaoMdGirIgcW3NZFEzX9cg7eSOUpXx2NCeaMh+ggpa1K92h
9QsD5MJLI/z1X6pMTuWasHkd3LHNXB22QhP5PAzyJaRmBvq6DEIbHxDC5xApw2XdduRBbppf6gih
8WOepsIfrGewfrvtikDPM0RBd9aR3vdB3K0CcjVf7FsMbJBUJB/krmm1aobLnmoiyPf1f8QX1R34
clnSVuhmQec39CP/ulKHz201jfT9bpi3vCX5+EZYk/mdzI7JZzvUXnd+SEupQ3Ye9LbTabuft0lH
QLqpfZP4Y4TyUlpOxt10n3qDSIW2h+X1iJb34sJFZGrXF7KD2dYQFfMHi1u4nqKnjY0EXY+pPepe
ydx2GV5upxJIqOh9IndMYyS3gXNn3TowO6hhDUIZkOg9BiOICxDXS3zcQtRxpHugNx67ezSbpsFH
DClVqESubXvwU9vIX0wfmeeH3DQ42Lu/yNwrBj210ihiya/7VmOxsZgNuTGFpRWex0FVF1RAMH2a
QPf2dhpkRGGW10gRHqoOpZNivdIK9chcpvh6uFIzFoShlGIM0ZeGhuXw142XFCMdLAVUOtuiVguy
gC07lFq3N0fWqx2x2VMvKhrCYtBrgKA3bMwK1BD8qdv2bjCXXN6LWa6mWA9wtNjdmZNhobKhhHQn
5nbNEg5EcB88gAF1ERa17/EERQjc9uZJAJ+6TQK0m3UaxplhRaCi4qzra8KRWKKur0HyHIzlYIgU
glVtkqTS0j/NaZDb9PktNsEGOt+omh/SkS7NLMZa6ax2TWkhGatiTamvuP9BLE2Imamcf+iT5QS+
Nf95yaiU7zRgjcZHLHy28oO2of2VJm+2d7SguUwowL0rcV+VevFIw32aGE9vRtosDdq2POzD8RZe
bR4sO6I5qpt8fT/ODKWJrlxtJpJbf4yn2XbcwB4n04sQKYjqC3yTLv1bPG/y8C9s3dHZOOBXTFLN
SzgYz1FyIFBnDc8iprucl7pyaT7tGnNopQPK/2jMmfvqSdhTUrY7py6fDWaBX2T/by0la5wKKjwF
oK8WacbuVFvk7g9ccQ/58UsJK1RI404/2DmnNmHxs46c6nDh+1o3ezo8guqiH/FLmzYDKHwqKp5m
5VtwjsTx2zwuh75E+RiuNXJm+wQX+EGT7uiPsku7aeF3JqxD6luj0H88viQXXwxBmBCRtfzwOO0S
hVvuTY03xc7gfLAHMq0Ut/pg5Jc/Ubw9NT903NdjWL5LOwAsqVoClkDxGKm5L31dFcySa/jDRb7H
8vVXahq1hbAdCJFcOPLKJVnt+6oPOEQfOtx1r8C+oDwV9rXR3fwMMwaGwA5jdL6/x9RPwmGoOul5
qGyzmRSbUdMlCun+uMKEOwpP2yMgMSL/vJfiXNo5WdB36QL4ME4ZVyAtA7T3ine4fHBJMub9/7yt
z8M/hPbwPqZ+Jeiu12CGs0R3nPs6OlhmIpRaELNtMQXJ9ho0INEu31+WrJUKrx+sGI0HwQ+mHfhZ
roDExepsQeiIXOwoAU8oStU3KJv5QfsOcFtfoyffA2btbO9r8c2n46QgceQ2Zu7yWH1ZtHOth+zt
59PS3OIeZXmMTUOst84bYfE3ZIMFklOzdyjZwzkOoUqQl/IpkAIVVkeRbLPdtx08pVE0J9/OSkdq
hj42ux1WGSO0rV1ycHZ9806lmPZ211N2eV6yBOydCpI9+qbZSttrXXXT3B4z/CGYL3U6eLyR68oQ
QKUX0moKGUHnT6YMTCnir2pxWarPAKSEAlLsHobT6sJIgUw20hdAUDEl7obbH5uzol4MFvb3f4m1
mrFe+ESe8pQQXHqeYl1VkV+3vcLETAA4CbxPX/oLdcFsEvKolx773mXDwhbIFlrm+B+THPRVeU8j
aEWsid0H/AfYNF4yGT0/eRUjMPU1t8hTZzS/O0MnJ8p5rBNOx0kBWod9rhYWnW04lEoR7A0scZNi
sFyD5UkFMAGlLYtX3hOgNIXPiBtuXoFpqnFMeMFlBS0ASUeIjX3M3nyF+mbMjzqeQfCrbPi6CisV
ybjJD2kb8fcQC8LeWxKO3d371YEueGFTS6XFC141mw+6OamGteaBLa6BbjCIaHOWtqHaCPCobDba
y0xOx8I7gFQIewAYLrvVtwc+rA3AjR8gMURAqL+oBDLuV7R0equBb2JuepxbEhDIYasz5q0nPy5r
egxYLc/aMsWxDcBv2kzwerP1fy4UEp4oS62L9LTcDIYuZWJxHvvauVvv8+H4lek7vweuce18PAbU
NN93opoWzLD5ezsmddyooWq+JDdpX9cz3fexRRJX+4GX9qQDAwRVy0HIcSzH1wSjgiZW/Mz7oFKL
0kCfkME9LuFsmde/arTtaydAaw8YF6WdwG6+7wT+EyZCy5v/N/rNQk1/IOnZo7gZOeeHjghCnZUe
7uMsOiduCrk/WoWkMnN8yOQTgqzgwRendUv/Y6tPiwDQONFzkeSISFCx5NGV0fErWwVVBey/wUQ5
c/Ww9bZoxSBchR99c5OmOdyfjHNsZcep/dFIJe6zX8G8rlh9LwYsLJS6jTtjO4GYe4HFg37uNP3x
BAiDVmh1tuzRM3P22Yyv0PZetDi5JcYDm6rr0sSya9AOX1Q/7T8ZAUegd1j9Q9jjVTMWi9EFC2LR
/8RS8vwFpT2tunOeCwih2gtLmSqVxwkY0LXVW68oYPD4TA+7maJejxs1t6l33LrKyNFGwWfpqpR4
4aEfBIVf85M1iwSfMI+rPQp4zhZ/AjsPdoLwxH6/TNuZeVLgbWB+Dw5IkMRphX1UHOQbQwUALXyI
RF8BS3/PvfnFNoqVR1Zi27f7sMNc5QX65omlYiwAcEz/KYMoqgYjav9+TUmshH/QCtigjV8XWOW+
1FrUnQa2/VccwQnJ0YaDUQz9bB4fiT4YG8aVif9olVVyEHPloA87iiuGxtIk0p/hasXSy3BkCF2W
SfucP/hSIz3NhCjWKcskoTf0J6T3bSvrGLl7onpBrqVyFK4QZ+I8pZlKkICqbNNxO353kdWIVUpn
SILtcMHtvCIEvPCxiHSAyovlIbJR7cNfmyZ1kQebgK9lYHZf/ldnIABv1Mym8GpCouo3HguPbCRG
3R8FAdEnPm36lWNRdDrjALzpr+Vo9/RSTGXtYTTXd3MTIVX7qDZQngJYH0syx/G2NcqfSDYeX/9F
/xVb/W/+TCcCNzzV3gsp9c1Q6Yzw9iHCHgxybHPKXlTQgcZB4mDk+0f0UkDAf9RFWQtQLDKxuJoJ
9oA0BaIZvXSgq60DcmDusBS6u7JDvq6nKEwQDZoLDvd+Zf+91f2kOOWwb1mCAh4EA9fkyW2RABcd
uKWBJOKc3TgD5XP1a+zjeVGhSHEJIOQ7h5YjO/OCXXd9jz/qzT2PwGtslc7/vB/szMI/2x7BLkur
SH46KbuCueKQcCy4aU/Fpm+3OB3dJsLBwNZEjOd9FthyJAc+joC9P+3+AuD/hj1oliSNIj04W3wa
8jXI+C8xcubUzU35G/XWJEX8dnEtUxn6MZeCr6QKixze4T+CbYEaEhsNPEpIQLyKRxAfFE1MqQQh
o9TGhCFVAvMWPDLUY94wFx1kKFt9Egtu3rXzezF1iYoJA0leDo+dKt7IG4bvdNsGns9FN1Gc447v
mWEzyYyXYdCB6muFBCVB0juEzbRlH0xSToYeGHLH6WuH5VM6bziZOvK3EOZButXEQT6wvFbTy3/g
8THEP6Mqx6VTxnV46Nfr0ZN37f/0ucG+4+rOEIGRgXaGce0QpatWeMJVT9iQofE2fZbxIsI8WS26
or4NfMPQdmwLX/o+xOrnJ/YkAfhI6StlD5YRt9a1KyjznII2ofcgWT9nDQZIyqBoyWPnjEu8aNAa
8jrm+SIorKTMaNgWTR0qb6bPi1NBP+HGEHqefUJEDPBS1VKfLuLdqV/oyWrZEYM2075CNkAluboi
KI1ADkgL5s+BQ/LVgNS8S6JzRlOr8y2VEf1ixrf51Bs7RXb+m0Yqkn9pqWzHa7BgqR3pMmJue2Wv
l7ppE8i+bWhCkPz7zqgYLBBsotzonpODJBwrZpBqPDc2vLpSGmLaPMWBfHnxEOdssmvn8n+SmE9F
KLR6OGED6NAjUbaX3hm89+c+CvbV8B0iYM4p9wX2UOH0FvMZzptqGjbpjXeSbXA6v9DbN8z/ZYrN
fma+bWOudHMwj2grLc6SMwTpn4oTKsyo96bzpHMi6K92eayP6w2OrTgmdJ/eUr/uVVnpf3pQzDG4
WR7Gq/42FhfM4biuzQOMPPj9ez4b1pbExF4M0vbswu8FRFhpqOF4VssSvekkVYS/FhgPC4XPDpcO
m7e6XVFkpmA7kDj37MvuxtM6Ng/ECyTBK0/AFdrt1uMj4uWzXTqmDT2XI1/q60tn3cXC8J74hBC9
88cDnvbDU8hLESRW0HP2q24E5eNjRNGS5sQ6fLa/EZM+js8jdi5rNde+FBGlzf7ATPTFp7RDJ+U0
/I6eNX4l835AGgRfz6rX/J5ihNsQWVC+0FATs+6evsPVFY9Swo1QMYyiKDRhhhFw0X5qhEPfEL1x
GJLDq/iRs2N8+Z8014Gf5Ou5RnmY7X9JtR4xv0PsYUN7Px7g3D2X5uLr5rQC/RZILRUnr8xRqKWA
vrbZRyPcFN/LSkeWmr6GiGVy1Ar5Rc/8r2EIFI7tMc65rpDKt4jN3u1oIBMK9uUJ8jaL+lNFxOpj
KpPiuoQIb7C0LbOMSDfvmxDQ0KO5c/1LBewd0K8axR6IcWLqNzmFlEXqjMLqSIN8Sp5cYreeLE9J
HxdvgD592yLzn9iaoP/9BA6x323xDyOjczTqWcwz1QqQGoJVDDPWfP58GuwiUjIFZ4jaPdyfpIQJ
/Jn/LlZNoeLiMVvfkfdMFFcGSMu5AfiBTDS0uzOnlAwlx2E5qguxWWF0V+FwN27PRkBFioxUVm8j
qa1pXnyb1Udv6cDoLlhc9G4dnSW2CJJTgedbPJCzygAKOEPU6ksTcUgKqAzr+n32NKwKMnOI6iL1
CyG8pQenPb0UVEwRldpOjWxUxVsQu3Q5GIu3JBl35RuJ+xayvJtykoRDM7hoIyZXDcPQdlhx/4nt
rCrATfNwZ2/H37iT1wCyQQjy/bK1yHA10u+vEmnMzxeSXXn64fWMBoAnH8fDF6MqeM3aEv1YKz6k
V9GVej7CvK+735qRLzPiDQ63ygkwmYZJ09B0KbMa6qmGhRrnviDFp/VdkWtoIVLyOyL520N4yb4Q
mmxZnR4xCJMtKn805Y0Kc3OnLSQhPT4U5o/UFxk4x344kFMmTA2s6VHuJdqvwqESLvvUWjHeCF6H
BqEE3jdK6cJsEJm2ctm6k3RDt+DaoWTCSjaOYRA1+zyY+PBC8gidvPIDeWXO0uYRe21fGXszI+xc
iP09YUtHQmOuXXBjVtwF8O1AvV3e1QQRAqtngPRbbr97Kcydb9h/toqDlgDOm14CqNB2iwj7ZuI9
qxfdjfuLD9t8/d1UyvWSzs4HNK2Pl1xl0wmMYFyXHlkVFw3Dbfefw0Pvr7CkFnEhnG9VQTP66tbY
yWcO8OMCyjfAQvePish6VuDKszJX6EuwYSpTgjXalPokmkkSE+cH68jyaZQFQ3hWOcTmObtusSc1
f1LcYlCptN2g+VHizEIbRRdwZuegCKGcgnKDfA83ImNkMHB6DpUyDoq6qvjxee5ErGsItkEiyT/A
YH8Rdicm0nOSozae2Fb58CX3PfXY3W2xty6hhNbCVD0/v6Jp6Q/cli/ZYUp81PY0PoChCypspiMj
taG38CybKdPTcQu7jrjhe82N/FAS7FumwdOvB2+CctoG6DSOvH0ddcAICC4S9/4g12wXhbVuG/NI
l7y9dVQoUE1O4Of+9ghAC8EZOMZScYi3abxYUwVCwC966/6mEaw7KlnH8HNzPzoC4KR2WB53NG8D
/8T1ZQMfwiycDO9bxjE8MuAy1mexO1st/uOvqQng6NJ7WwVmcA25QoLYJ2l8xnRsNh1VSXScRad1
X91ciiIyVsOryilm6t+LNqWhkRvjusq2wfF7RJ0XUEnkrlSmk7G4SqiiwujBbtENR8KbZS+oks9P
MzNF3h+sUEEe7f+jFQzSM8DSrwmaYL+rYEWDK1tYAhBk0fcv1lDWCWWv5z3rpTcYYbhRnXKAh8Ez
Sk2QtdI8+XvY23dAqHCaqj2s6GOQJ+mygwtY/TE3lQbobiIO19xsViLRzdvc9TR8oud2jvqaJwxW
/mkYYGakbnJbm7JOVGQ9fFvVidwK1ikMwLgvC1qES5hbQYBtrj2jfrGvq8FdnXpDcrwc5QNaE60z
yl2kq5Hy2mhcbhBcqAzJ7kbdmfpU2epylYMFRtSDMMF9NynBskVAuFPcprvftOHU1Q7ndTg47mWt
VzyeSV8aWSmgQqNGg89JWpH5wbl2t0f2Oy3eYFz2vlEAVqKmRHCyXR6oNTGqVErsRBPGOUopbYPD
Oh+BikLhYJsMd+BHHOqIFL79UsapuDMwWDcFYtNmYAxACpA1wPSJZlIYezsL6W9N53PNv1BCkMxd
ChmvOpfhMKO4z92gjfhsHauKcjHyV5IbmDEHvj2DMV0aLFkZPGdIZf5q4G2AG29w1pcyz8/UPIUK
3UG1mCOe8oY0x2uba427lpMgpjiJ29FAtaSS0yUP+IhmvXgVU6eu+1TyF+nlzHyR7l55bszck2iX
a076C8eeycEwPDXGRrAbkj4C/7+n6sdKP95wBdB5HpyYYbEhRgilGm+qUL5qepZdrAiiP3dEiVI/
O7PTLOW7/kcgAYy6egNfsHqf02D6CtUHmqBy0a+k9RMLNr6r9tZjeCMO0HGm3A3jhNyNp3kfstJi
f/Yg0Q4OpuGMlCdHvUSvz7mD0z71UOUKVIFVEQ2Xeb15+H14/RYtjVbFgfqnFJVdC+E5phYzIYxO
D+GSGResYklLqWkM2KeMdCjujtYIN4ToVufwvwaffGuMN3eh2ChKD4wQfh5hWWJcxruwKrJJaQhj
+gtx+2qgVCPasvoPZoJjJJSPlSylHJGYZ2emcKg/nFqWrsgLQcG2aWFoLbaq5z7QfiIm2KJmqCYD
iZvMitxVuYYLlPRIX1wqD6dmLZAkT4QcCdW2eaZ7y16HCqMugfVMXMxKivMkNnbOYehsNgNI6l0f
BKVk83STFiY96ZdkkWpCT6iANKRnjxs9eeZp77KXNGsnMF/TW/KRQIGQML2YsMYI+es9OxC66dgg
JWebNJSr05yiQGcYEB2DgaUbjgS9oy8oeFLud8/ui4qoqEKYGI87249v6wPl0Q3BjfjldmSX02AS
piUIqV3diMrWevXDQK/gs5/caExMt0lD99+vLfJQt4cKiZv75ucJrR699UIIEcHn0hfXID4/f8V4
B1zrdBAJi717OXe56Y352vUxXimLbsbAsZu8Why/HLGANxVjkFOjEvUyw5gJMc+YkzXt/3hesd27
66JiH6mhPs1wXxZ5v0nswQMR+t46JGfA4dxbKvZJMebk/60ezr6a1Oc5a1KTOvhijIBh+QLJTJ2a
ErT7fsqXKv1J8mfe3u0UQw8GalA8fAlt5EZuRtmWNKfENJJLcZjv2cFv15yhtTsVuZIGTtq/SY5F
Hr7RzZP0UPk6XI5eBKukAuKj6zw5YEcGBzrRry3CzPfB+BZficvVbvK52hIAtOWD3DSJIDff3O7R
/iOZHZXmDFoo8c6uqk7iqeUKzCKecdKWtZDOpSqphpjPi8VrUIU1SphwPlfZnyiU3Kv0vxCVW+EY
mJGz5XxwIamVVPzhxuyhgxUxacP9YegqO1/OMorDKSapFX2J0r12ipaT2eDbfgQM37vZ3548aCzl
b3hbxFbqwmhAQoxXFcVA3STXiTR3RuZRIsBKBnMusGptta5BLD5iOx+IvizoDGioJFAK02h6fe+w
wyk73fXcMHTvuPZsseTO52OVCSc7EDNbXThB4Wm5FmjDazHILOJY/7Yrr+83j5fJTRtLLNL3vM/Q
PLRMz+okBjiHuFOvCac9T6FMNStwQqTxfb365kF8wA6r33TQvlHCbaQGN4n76+jqoOprnGDynsDX
UNlBPsGyLIoUeRNEYQVRNkDJ27KYQMLUkmQOL+7bSDhzYGameonLNWEJLsw9ThdYNRgiIsbvxZea
Att2jz8bsrLnABuePVOA9HG0Ta/+6uI4QkTZZLNL+dMDS6yZULQk1kql+P4eyQrYruajjmWwIibc
007Y+SKAwDSe7gJ/5sxEIXuOxvyWWMssFxBP/305R6/h0fDxmOVXYznDi+L/IYU/XdLUpJqyxBdq
szNo9QPQdmM5ckN+hrII76NuT4/ZjbPSye4BIywAbxAJoG5QE145MqTukxK45Tf16GC/+6AsJY1D
HUYre3YZWdt2ga2vtqwyqEfVU6qP2kE3KFmAgtf0ovS3cvL6Zj+QSpg3BFuM17cm9DQTYL/mrMys
8xkpoSOghHa8ZGJ9aW/5cNIkSR1iw+H1pCpDmWiaLWMKqSaWW4MQ7V/WYJXADz9fVI9/LbxXCE7R
6ZuMaY7DRNNEVKhRpaals+JagBkdqgDYNUrNTd4kS5SitrjwnRSHSoakC/6eTV11HC+4eO+tcyxC
yLFNuD8txkYc9xA0d9KrkQGB6mm3YG+9qpBllEJRkXeIpOCdtH7wTIHHLDI5RO552yAw9vNpHOjX
oZ3fK79W0kaAnEPWM5fKYzBBZx0NwELuasvSko9ruuZ37zsQGqkhMOUhdGRbSZMgRc5s6Mm5L4Va
icwr5R6xyqjVJp/eZLcR1pOLJSABnCMOzE9QEx60S+qF5Yh4M1MQelKknWwGY8KwpGmyxkyzmHdo
GZBUwDvYradp3nkhjTjc0M8AWs2FsWfn8iqNNXg332O6H3ZG7rNoSYYnbE5FzqhElSJaILV3f/nX
eKgGZLS6etIiqnEGrsTGpKbCxajTqu3QVdyt4zp9k0JdLzzjezzvpfwQoWBi0fAIoXwev/3Qu6U/
GQENyOY0rspceYM6d2KgFtGmKzpRVHTBCt4KF6oMf/7rQbbv4DB8xKnlFNEIigF598IBIaLkkjO9
xDzGYtea1E5JDyi/ISJwOYjYWOReV9E/okbPoeSsa8T1wW79eROp8rPOuP9FC/gQ8L+cmfJXLmwt
pE5aUeGbt/+zdas12LfXp/4KNGOKLavGkon+QmlvIu9KLR1C55dXi09/BN/1ckWVJe120FG1R0bO
YUXuTvDkpM8DNm6vrEUSqDzFMPyhy9Sz0ALW2dpGnKTGUfaZOvsU5Mo5ai6QOxBz/zWR2CfMq5JR
04wZw1knj3txuUXeh3Ep7nu8KcVAQQxQUASPV/f6g0kveKBncZtUf2mkQOYPsW8kJG9PotrDJ1Yk
Iy+/tPxmjNnd44LtgMOK3m9vH0h+bBnt7IYoV+etwNMOI3jbtWjv1EM9G/RXleKejgblsfb+cRgR
MM5639JxmGZyfd5QQGm3U/cufdTJn8qeFr72Ij2tYT2ARUiArwYDhUiVjiaEb7NsN0JKJD5HnA3S
XMDa5QcbjnEt0FBxLgROoxmrv975q/9ItJYhvuuPXSWIkE1vCPI9mIw5XUy55/ofQSY3xuL0UubG
joFvaTpMPy9S01IBXSDyfXeiyV0soqpOACrDJXn8/PMfsuxrvz9GXtuc6xl0tSacUWi73DNo7Nsl
8ePv9Bj0BcZ5mSm1DOuwlfRX6KMNB9plJdgLgOW3EqPAlg31K8R7YcZhkuitiNUgPGAOl9x4vIxh
3/uu6NpoZfVFdpJ7taSXYhby8eXNOs9xKgQItWZaXTNj1HT939yUv4wxtgm56xwPT33hACQcdwvo
FPSkbjNFIhC9JroHs0lOj2/6dKiq4/YSvwyFXXuJ1z8+a6rxfpY18IFBzW8Q4nrL6cP2lP41yaxl
QexCeX/NxJlsS/rtWU/PTuZDUPjaaxU+Qn9/L1xAKB2wIP289xdtLJIQKvEzCLU0P+QdFefJ0e8S
e2idwpxCs4sZW/D+FAv6B+wXDeSVZsf1dhYieCTsfYI0rusFG8OwONJ+pVF5HT6NG8G2j2V5+s8r
Ng0Uq5k4kU6n8w/aVv/USPKF+XEiaWZ+3Nw/Acj1gENavD0IJSBPD8J4pLWZ8LmBYcwIQXjinYfp
SnNHjyPEf0BysBrjwK/egwmHR86mbKzrA1XZJPjBUSf/4XocZ9oGYbY7zJ3gC2aF8MdOu/AFHYU1
/RIwXz9gS04eEwif1FF4AJkB2O8fxA6wpjk72z3N8ftRBG8GUgv+9lAUcbJeebl5qXYpR0em10Fm
aigEM5TpdLi/AE/OTG/q6UW+xIjCVea3mCAvCoIkClKEMvAJWHIW4K3tzlrs9Jm/u3KxK2Tqwp1R
Ox1xHCniK/Kv8czng7/csQC9HnRbcBswZCNj1+MPkeYKQ5y2LD29/2ToBd9wXkDqpK4JVja8Wgck
oaKMk68xATIipGG1Px4Iy5/q5JnEKLJYM3VYEKJRPJSj4hEYGvpUZU3rpFSyXVgR59SUzUeNDFIT
5eb0MR8k+74tEkPHW8hXeei4a0ltmsZp6xAgrY/zCsOYYPqXwSuF94BS4Q6EkyLCtslIvRhH9Ijq
8CzvfjByYTlRJgFKgfL6JBjXLWLBPZX+rOx6uvDthOwa8kjYuDI75p15xP/mlMKHP4inNEVT1CD4
N5uDVbgrHOdcyFuC71pDIlQ3keJFLv4M8FTJNKBbAPQ/uo3fBp5QrP4WAthJoFHrbHQgd2NV76nB
d8ZeFdezrEgYOBHy36ea+Tchq9hK05r4y443sgQ757pesdKrZTG/3PLm+iN7ChcByJd7B4ALWLKf
mhZX+gw7h2wpQNrdlf62CsRauzpNzCWtc5DSOJ8BpHz0mguO+NBkFf/NsADtYuegZIDwzSp6yt5K
oUDaGW0KwhhUmxdQZZ596jlj2YgDRtL5PgFHplk71tDw47KTWG9j7AkZOBrN493DSVvWfL/LlMGe
UF9xa16AfPnJtXYl+r3pOG4E6YQ6BiQMXKVzWNrZCeDdNto1EjjPAFXkdecvNWMcuykPhJYMjtH5
Od7khG5lcJyja1yH/dP1XhSi7K3fnULD9Jas20NcQx8KcpfE2LPoH08ZuJXMKtjZ6jKB8s+VjA6A
6WHej7fAZGMNkogclh9wGKlIO5i2eW4lBefY5orNM9CYGt2T1BTc5xy9JyM+mW9SKaVfNhpcP4ke
sEdyT55TjXJA11lHOt18UwkU1m5SG6TX5SN/SYh+epHl+Z+gn0NjUrhK4rOVWPAI6tC2qzplXA68
i1dvsr7+Xjrp4fOqg+kc4uffqYGwqt8yEC44uL2hq3r5yxy2bAYUGRVA7Uv0xK4B4tVc2xNfcnQv
xJGBcQOssrnN7XbNbzadvAn1KfYsL0KlRWsedt7VTkmekT2yqnJKsmdMoRhQkRXu+KCV7xIGqHN8
7n4Dr8EMRYCeqoudIQBdl5+ap3FMYiqaCuvI0k5Wvz6CjEye5IfbpA3qJLgCANN5BXJ/rog9F35H
ZKm+fSLYpDfDSvbcMpGadwigeaciHT4AeXQyzOlhjl9Nm715nMfiw9+dQm/pFtCpKcgz4ejvutmy
4Q3yLh8MkA5OvoNJsfL4FLWuqH4AT3amKfecoJF95YkhXxBjJQrD4iWHOU+s9r4iV/Qc/3wdfbaH
bpPNMofOsSGUCOrZjxVHlxuoGcvnLZtb14yPM9nF7jKOhnfy30Cdq0m4oY8X6LAVVEGdrpo1h6M0
LqgiYAX+Y7vDk4LJrjQfQssnMW65aqQHIqeMrDdQ2viQDTnarWGb92w2tHsrEA2bsxRm8zASEsEO
HR2T/RL2r/Zg7TnC7wkTvdzehgYzkzXfIxQcynROmJnU9e6NHRIzScb0gc8tmcLvIK9kDQkpFnYI
gIYmZUtY6R3WzvDA87NWGZaHMRFjE5TTsZb2PWbKOCaBzdKJCYtu9QBnyUNQz9s/DQroPbDaDf+/
BixQ3eL/yNJhLQQTlJQ1jE3PezOZ8eQVKUfsmiTNlDn06KxOBXZRlwVu0nBLJwGbdn4oQUsaxR68
kO/36g+muloPRo5c8Y04cndqiMGW4iIeMHT6AB4goJw6o9EywTJ640pzulF4Jd/gLcohjW0r7FCS
l+yUKHSWyDJ3p3nw5ig4qLtVEpbRXXOcliVBZO4SZECTOHIcgTQkkeF6lzFAJxM/DLZs0y1XqQ2j
LRmTNRLAgMMI8Wle4tNQM7eIsJH8hyitO/FvQO5601uh9EhreFqrE69r3M0W9K/iysxl91lYp29c
3jVuCWxWaL14MvWSGqNL5sd/71bMZwEfJfCOEGLyenTm3lbcKctN+zA431Ng6OTHPR2cnKHBVMj2
jzvLzeqPREDzfSU5Zd8wYNDloHQPgSRM8k4VbvOzfH7cKx2jyngzND0nn0cMgtI0HGVbeB3syrCm
zXTdPssQzr2rnfrtTpo8YN5xvL3Lv+GatOV8A98aVT2a/nLzy+H3C3bbnAMmUARHeepQP8bMNgjE
w0+W3Vz7Ej1SlfZrZJArpWL8kYnOisJtbU+F5+TuLEUwMEJFqpepsWrGAgF3uANRBKww7rGNd9Zv
TkUOIuDdrybqq4Orx3+EGL8nr045Ev+UowESMn6l/4aLrfPo7Ie1PyPYy43kCaEv0U1I/b3u8lVj
KvS+aiAI7hrrdUjh45ASIGp4L4JaIChaDalcQ5NZrSpz3NR7BSBIC+l1vO2EaqC/AjtaaVswejqU
VKRSUs4Megwp0FlV27RykmVCDPa9LsGefonR0TRJGoPN2nm/W1Y4XPXWC0cd21QVB0a2tWCIk3n2
AWvtRX91lQJP22KsoaNZwGmc9Rv4Wam4VvgsiC6ZJri1xGDXjSVzpDow/idhyzymxMrBVxQ38Tu4
U+ocCsN+HImJodlHB0NqEiUm7vNi7DCmq/57suHhDQvpnZUTiKLCcO4Vgp413lJI1HBCnAfeITl4
oknw4iOjQs5ICe9qpNzDKfWe6yF4nMM347Uuv4IqchZn7JD0leMpsScdQutzqjjJrzRWpyl0+FjA
qfF0AC9jTbaOs5gux1I/l90Mx1ObkTL288CuBXZldcCLvnP5AGpGUNOCcV4JHCYV4e/NDox7gV7g
LI5SWqSDPtALPPLFN5I948L7Kj5i3xZMVEg08Yh1UPpNG1xWN+rOOJMrSv0WYHfWFljls4BduH9F
kvw09J8MAj2gUZTECNuqcDJc/OpVLVGDkSg/VYq+TOkb92MZE4jEop8+HEr65Z/Ee7lPdwMxD+9N
hodAGQVnPq3U5w8HG18Bvp8G8QAE9abxUNATsLi0LBeW5enisqgXK+yzEc7for2VheRCpASctcZL
fnwLQW7ahS8oLy6SueCZJma/veNPcN4/+cUaKKacsbcjepboNy06TPgXfHH6H+AhkaNgllh32RTe
NT8P0coOCq/2KxD0SbtWv+4xNnsRzYBOn080wOt4tXiFeeRkZzw7wAz8mDgWpWoOranhrhLlz5VG
NUrYMghOg797wJ8jmv+KZ39t3k/Ri/DtTfjjdqqoe4cid/yj01gawgpASXbzbgPe/klIcm/c+kVV
gVYzyslURjy6Dwm/I4vTMKcuW9KNjiDEMr1ese6pI7g3pUcSvNAjhx0+lexHbGogCkvfYk3RIOaU
MOeivX7MS6TGIFl6kQ0NJnTEVY0B4lEjiZ+1HNdMIG9as2JmN7F/aGA5gFZ6zyVlWE+9sjWiKW1n
pbVvwLDPW/YQFxJ6C04l3ctFEG8uD67kt7KVVIur1rMRI8WXCrYpUYirFYk/RUVSSz00XeTbXaFV
Ny4r0quAXVI/CR49p/Wk69SlqdxphmYRLukENy3T6ZNjP2H1B6chkVMRB5GAevuc2S8SpysyvARy
U0eBE4ibyeTsGGfPC3VQFi5JJrAPdIIYlgkLUeeBVdYQXSJ/bNcubR6rSrbUOEE7kMXySMlpu6e5
Px9SxtBBaXLJKouiiSCGrYkJ8tQljyLVPqyTMUzBidoSVsW3AebIRIEtg92m6WZ2fJXk8k4XIMIT
HEnYbxI2BZGI9njNbP3qUxWjPQABhpNcNw4oLgVSz88f2qR52ZEVRj0RPWICjfXs9JVOYx8lmrUC
ic/DddN5y6jmW9B1C3Kn83xHxqDqz1vkGVjUKU2blzVOtJodkTHIL+t5/dfKmnYRZsivTyuWGtTs
fxS2/kf59qkcGXAZn3kwjITcvp4mNSgnEoCiQGl9pNGq1OikU8BwoF65EZ1WEE3yJ5KzBi28Mc7i
IRK1vE/rA/iiwOy276saqkS6gZcH6tZWFHW3JZSP9YGA9ANXLHy5muQ9OKYeEUJMGvlku/y3/NiV
hjT2T9iirRN6ZN88t6xJSXkQO55dy0FYqrvzFC5xNHeFGVICf3SsYaCYGUWpciCiYUuTV0uMlsNV
cxh68FLbGFT5w9ExSn1cGZDVh4dtz/rYMiAlZtsDF49QUO4ey5RTK1Vx/oHvwCdqg3GuLQCOAh2P
Mp1WZNE1MGIKTVwBFwi+hYjGAPgyosezx1ST7mbugaQhYJbqQxRNLhBT5pGoEYoka6qHairrxb60
8uxtnmZ82U6Ux4nrCrzXwqk/wgwHaZu2V6iIhE3NGhY+bZPX/1RPXnFlDRfVIGCW/4KVbLcsG4+l
KPOwnQpj5l9RCMCzYeU4jLbwivbYxdZFKN5vA/CsMq5rWc5H9tdRn7jh00l0acFA4vF+2NiOlksJ
pI6oqCKh42unEGPlxQHWiLNnzZdPnxjgPWK2nGU7HimbM0Voscn3JSStBz/P3ZwJc+Pcc2lv7Xbu
Z4SDYnT7BmFEx7uA5CtOQAOg3TaoaEhEbKjK9QaY9KaRUJM+hKrAC9VfLXsbc1+XBV7cg5dCWV6O
acJePNpl+DwHoXlhz8bi1lR/P7GENE8T1oYFRnITbASSLBO1BJ4a9PAPe4/uWeYLKK9sZ4zPxauI
PsLBOE9h3uYPYoikFhozUgIMx3br+yF3yOUfldHsyZ3hLx4TtHtRxGJLb7iyK+rCjrHnW38ovGHj
/M5vaOc7X3GaLJfxcIwwt0nwUKawKQAIWN0e+5SX7Kv/Ik+F7brewjo98V3xDBwm7GffMlKsFe0d
TorK6AGBctD2izfvTYhagjmVWkcT8anjpYt2VV0X5GtKGdOWTktgma0UxsYddVn4YNWpQNNcHMwy
Qtd3GH7WK0OyIr9z/5G9l2XROfG5p0Cdg8BXLAQthg80/DkXrRjiRJi5zR40BBEJNc0Lehz1IYvm
d95l4wKLCSCFRbn8XacFKbPrJhDV+BvrbU0u1pnWBNjPvPMMkfb3HaysODMKYDDK/qq1TXXgiUi6
93c8eD/vrERXbfMHD99bTzcRXgZIof9t8N1kXp8aZdIjDpjddB9Ziqd2Zw/A8IiRV7aWdLol+vif
LOVkaot5UaFNbX6Oau4VLoJGVe10D0N9mG1uYqYAdTHq2pKNC+2q0lL96z1SPnJBmNkO92bzbh81
u9BfTy7W631iDEgKbQZ16oJd5YM+mNr1mf9hq4/l0bJcgHDLldlfhAa0E+VgfjzB8L90OdXodVYW
rqXVj/F3a5JT9q+oyuUB0NbFCBS7BG3wfYdj6T/MIC1gU1AdPQYY6tS2tDyu5gLGtbf8O1W0uI86
Y5Ott/s5FU5sdSn5xvN6lGovXuOrxqBrz4e1YMucwx78uOUDGDvpBSsS7/fcfLgEMsIK7LbHhg4L
CmWHaAVZnNSOJgEXCKRQxhtnFJ+dikzt0k82pKs4x6YgfAMC+wF3KAhR+LyXJqI5vZ2X2iv5hlez
IQ6AhEDsOjOREQ2ggYdSApISZ+ujmqq82tTwJUkCGJ+b+4RwoKUni0oje/pXisv7Sz5WqlLXF2To
Sa+fUixrn0BNgP4AEqMGY3UnomOE9ayQOaClIfrv9T8SUrNMbVFjhSAReJYNXp/7Q88WhHXpC5uU
3iapReBhpSh4Dpo3kKUtlQdeePzAhCEZW9mMdNdsfA1VieIR09zSYjUP5P5Q7+vk9lmxzFbyBHbZ
UO6PVeB1MvyZprivNJ7rhEhS97+nvNsiTwpuqlM4RzqF1esrhcryItxYPf+AQZOaN7JwIDofhj4f
gg3rB0rWQ9CGfm7RQ40P9V8yzviSRjk5nKvcdhO9DhTCj4qh0WJe/hBwLqH21+Qff/vAVDbWzMdk
gkYQJ7oLKgcT0NBS9OgJPVN/m61AyD8mwnHXgCk9PJQCxvJFKjAAcilWer7vrE1Fuol+0++HDH4D
McAIcNRcAfNFqCPPrRlDc0FhucXxdbXFQZ0jJuFhEZPBdlLjN8kei6qLuyU4qviYKBEPUmtCbhoK
RgAjGp5eFpNPLOedRtW6HXO73nE/kQ3S7fBVfDejVb5kg7OHtMpjg4g08avLIzV83Xb/8O80nE2Q
GDp1ovVvilBt4MXYz/0FV8qrhtktgIqd/OKtigjl1Z+sAzyb88sOnVUuW7wIr5f1pZWETreZZqrn
g/kJLFAJFl67K8rIRoMY7LUdW4DYSv8pEgP22i8M13dG40CYuZcw4z6JaHRbFUGIOmJjpSj+rund
B4XZQomlRULtuQ1gUN6tWIbflBZX9KVvCujN42CPROB2Q9wZP9XtG0msJxzMCIuhzQp+0GliSjdQ
0nvQODf0/3VXA3q2SiyaEws9XaNwTrMuQOAowiKAISjY+o6hgwlXJU9OkD9rb0IVi0+8yc1eekx5
yGroBpYQkpiCBB2rtv62Rik3eowKwAl33nBhpoCttuChRSunVnFIiop+ZAduqsGyZ7V/UYTWyn7Y
zO7e0NYIMlO9DBRhiKb/sEu/DxP7PH6U+cOtIcxofZ/5twQwvbsmYnktUjBdnWoF7Ocu3D+m00Nz
S7wuQt8POXZblA1sQ+XrmgHOXL7CDdt/f/kUnqvVHENCJDEC6cekhOY+/S4keHvV2TkJrK5iJLeQ
ULVsRHyPDGcIxRX/XgF7sPYPtzw7SZRSKaNf99tIAFcLg9H84YWwcUmb40+Xq8I1dpEuS2E/yrge
vqF9K8KXQsyhpl9v1DD+mjIzba1rPzh8g1SdqHWZaZLPfgv+iNAM1PKJKv7vCqPmvhG/cHKfnZXb
bcU8cfGk8paO+FoEU1i0rRG/ODYdIM7al2xF+J0l9dA7/hhykIIBxu8ohmcNFgKbT5d69AIh9XY7
cRHxo6zw9E6dl4bd+URLSy7UkyqHv3XsNUdk5CKHHYjfpkMaDFDPZoSSpPhPWXRRPHkzT+cqSILh
pHKsO9ncEDXl6lcdfMyiYhMbQ24mpdU7w7/dv6EmVwz5KruRyF28hAwLhia7SgSd60ZNlq1kUNRF
ctWYpEit2l4/iTO3gZXkaNWNJ8gsQMr1Llu40ZMKakPylZGYA5/tHwSnlCAeHvg89j0OfPjP6EXo
YmGwvAmdj5dtbYgZtliiCqgiPiKNCs9dSzZjBX/cZySx1Fgztd2nH9Yvj8ZN+18swZhQEA2bILnr
1ZpEOBhNRDOH+HXZ5q0wJ1SK/4Guj1xiAiS8K1p+KXU+7dEdrXekQFx1sITdfVMKqBsZSdxXfWGK
/igcw+7Xg9OlmwUp20X/BOadYXX2frHE7HXTQ2/Y4+aBI14sogc10Y0B3y0/5AQLPn3fR2Z4EQZc
QFBq61Inr93DAjHBXQ2KL3CoxwEqcT4m6F0UNe9SXMzbpmJtkoMvsxP8b4Y/8R3u0OMkfTA+x13W
3n02+lM0IXMxzariTBf4Hiiup4Uh4kYQ5HMS4hUQLRTjHu1pWEbQQHZOvVa/a/PKK3uMdrZ0O5Tz
ZQrjZC7mfe+621EWz1gZa1uBThqQqSZ/v3cTYpnxmiWYqAlzwvkMjhSlrK6U39A1Xxjyr2jyX71W
xaLSU5YqlIC9Qn1AdMO+OGOciTaTm9uB4lNEhhMyn81Uq0Ie568cm914l0+wgRF6f9dSx9UZ78V6
5XXeXenrt3qDxeQN/cnPO7XtlNN1gnTfzO96hgcLXIk44cC43WVqTSVajJBv/312Ik0pb5vXXC9e
1dJ8HwLlLBEYhFr41+m6amb+Zkqnv6r3MAn8oyv4wAOla5asWAk/fWHG95RNBGRkVwmZloiRV5lz
OnB7mlshAk652xyM4gGsDFA6Ib6q0RDoXja1dKqaDiirK/z7SvJpI6VCHMeNU79j1KJUBoA8BP9J
j5yAIekT9UmOF3DwSJEAp6zJF+AlLm4DpEhRzOO2yC07xWbD5vcx37YUUA8xUj0OYeg0fGksv710
NX/7hC7mz7B2GXVWHqI9YvUNNI7TMpbsVVURS2uX+Nb4ogKRkliCToyQyrxxdYxYwrPSxj/t6P5k
VS43p8FCR3us18YyhXQVIWcmZU8M3aJDteYOorkIU+2bCsjPYnfrrrFuzqJZaMRhazEbdMaHKZeV
Si6y52V8/CG5XXAAbfg8/fIM3dimpgfeIoT0uPomGrlMt+enpuIXJ99YtkqxM0l6ZSBKhlQ89PlI
T2hMTJF7ETQiBJNg32RTOFc1bzOO+gysN+Xpvem3rZKAOWQRWIcF4KAUyX+ugbF8b7HBEHLeZ4oD
+b8s6l6yYwFxD8bFUY8kd24OIUH9ezHqoaY3Isz+e0j65r9qiELM0pAXCaBvBkrEiHsZdG3ZQIdK
Aayk5+TiRU00PkKDCnWN9KU4CKOghmZ2ZOuIWAWGxe/tPHT3wnTlI1RfHjRupeefQ17IFvYXA2M5
Xq+ENh64US/ORn4BipSjroSb/pGnQsQ4ZZMW7JEjb9B3vjIvVL9WOZ6DmQDE/1emDh7B6V4ocwW6
SShGnPif4zFMYS7NmK7VImcwhqgcrxyreDj5mhvyKZcZkLOI7MaXe2oNVpML4aobveClIu2C8n3g
BAx3Jh+LkLajRGDdocQBQxbxIAxPEnBjgm2lFHkXisgyfB3oJf0NJEXtCeZh0F/Umhfo+VWEkjLb
+3c6+6pgU1TiegmJpt3J4upww3I/XgV5lrobzrGUsrY/jChWVWeWvXQrZ71FyrhYSUQRlpAHcwzu
F0mhNY6d5XWQxMwnyI2H7TjiosRmJmaqxE5pp/HnU6j9Umk0SJi0fJdKBi7HMexMb6wjxqkIi0ft
ZiHJ4t7dbJeo9meM0IIN7zanj94o1324FQIzdjiqFE6i0x4aGFkyk+SdbQGVjeAGTnDb2TeBeo6+
oMJQACo0BTECCDILfRPRv9P/s/7TdFOPrSUjiGTh8FHc0qlbaFvyYp/t/E9T9K1eE5Dki7V9gTZh
ei3JIEHpAKuv323BXGJjRLi21wvcrFHF+UeG7fCmMc8RFeMn0C86PQ7QAEEMurd4OVKzJp2D/ALm
9tf8RtPSEhmMHe0jpOWTq9vRtmFOixkT+vePYpBnoh55uqh7agdTnKKyQrzrrwk5w5IISIZbjepw
PPawLkWVe1JbjvIV7YjaXbYoxS1wL+9cIwMK79t/AgVDAnJtkhk8pHLS7xcmFJ7sv9474WIAdjNf
wq0IuyfmhJMpJTiBgNJKaGbQcHP6Far52R9b+e9g21sE3sswjqHihccz5UMF/9AIjMGoFPgS/LbN
qz1IREdLfgQHaOa0DAjVkOcN9f9StQBEce9uL8IQofxdPAL7PrAPZX9RpLqrb5URkjXDb177PsK8
rQ5GF6mWUk+vrs7zzWyx0FBj/3NhvXqqimRo/TNPfoYnTrwmCU5W+NWGJz2iCrUgf708dSHcxIm+
+zN4UpfbgnXOxxby0FKjT7UnPVuz6l0Zc8OsOE9XHd4lU9X26vRQzGDAh+FJULNoUuGYKnriigB0
kA9o2rZROpUoDGJn+1CSSETTPq/3rphaqixd/0Fv5tEGPItWhzwpvX3JvTRQ1Grk+jQnpvsbRR0B
uDliN63b4EDMMlz2daJrNwf7T45epvJ2LZEAZRzGIhRvGg192nNaazq40HoBLEFY1e4Z4NotWFTL
JnrjvWIoFryhqeLzrXYaOjrJrHlaRRfEDvPU+0WgCYUQ8Xo1kV62V4j0D15m7c+rKmKzUMC64r+g
SRUKmWRaDmJpErUfpGPQhlxMoax2AL5ubrOphr3lwFH87tR+mZ8XExdMQDm6OMAzyPPqlu9xH+NX
7LjoF5WRaV5arVYLML+jCNAU+zVqbcO8rec6Ne4rXMsCd1+wQ7arhw4S4Zku+PFT4NfhcH3MqwWE
B32sJyzf+n1ygtRVHSz/zNv+H/RrwdHQrM681efeNgE2VavS13PW29cRx+wkrRwTlxMOihMw0GV9
lQ1XUZ853z9Au8QgR3++umcxydNpKgq5tZY6YR8zFHKEIk8/KPjwC8SZyy/Y1kyM87AxtOQzzE0B
SrNibm0KebbdYX79iBjETF58Rg5EPXGUlt/r+lEjvqHhMjEuQ41c2gBbuFhrJgoIdzKgDjpcltDz
4vpuvmHjPM8pdoyOexscBDYiyybqBcuI1CXkEbCZjjdtq0OLhFct2ikjpilsnXLdScQOUeBqQpg3
HH20bdSVMYJtl5qaAsUQ9R5bm/mNU9Ppx8f9ukQn+tGIVdem6VMMvLSyCAyOFin1P1b0GQFYdLTO
+EonOMYMSGRREFa+oHhHBbKvp7BmTFJ1Y8iFuRETy7uUAwvtRP/GBXa7glyHT46ZniJ6aUYoh9Hs
K+ud6m5v98L/UrN10+piGkbn2/PU5NamgkYfPeWLU9eaI5LQ1pmolg9dtN3eB85eL3e8fH1RdOsp
fMyLkD6RhpvqxyjCEe+R6VmW/osSN/aNw75OgssxXoshACuuSHtNgA/hTcndvJnY2cDfLDcwKfPO
My7lyvNWvNNKVDj4JX27lDUNf52Vqn2furLm/CZcUcPKfODr4FYYaObAWkWrTkcAzVdI8MzW0/1l
37dkT5ys1eNGhk/dHI2YdHClnrtKC82VOjRzRVPsq6PinsX9pUpUADlhfP220HlBih0kflFPY6uu
N4lveJvKG0TvzrsgAonZe6zmUY/yMc3opUajkazuYBRlnneahR3zz7HYHbewhyEemqlKLIU4gcLf
yKIo5F3szWqdLCbZ/AHz7f/K/+8gDI9262O/1vtE0bZcJKKSx2V64JnP0B+Y7u9kzlc+e8KFb2a0
dLHXmnd98ShTN6hEmQrEpA+j5oqI5Y07po9crYoGfY8HZKUjn7rnuUyefrYUaI0cOuNFjyj8o5Yi
eV3PUm/Yn8/SM6z+mvEbhwEv8M0DDHByf207b9UiUdx7/keuou80jatP+B2tTedImJWp9aYcMMOJ
auWdOAO/k/a5ZFwasOTfuSHPJNy/b0ocXql+dY9faLPx0wEY/ZbKYh6F54g2EhAP8Nd5gsyFc4jM
4BZIAFXXvTF9gpBBMMq+o4cuPb/dg6dfYkh5KBEOFxetJGgFjm/rG3ftvuN88HdsvRhk3hUiJ9zZ
SRZGVvSix3zVzKNqdzmY8p4nwlDjPqoj6FFFJ522v5bsOrDkvGfC2x8ijDks0SIqdikoEWp1RFme
PwI3zrvNLDHz7L1BpoGuQ5voauNTL7rvCyC0Bainvf3NHeoAofAym15eNfW6vnf3WURqiC2SJr6+
ESdvSXx6eOhLCrxUzZ5uMUpnI7KhroZ7XqqsbOZCqZO0He2YMT+ea5CCYhPgL3K8yx2VXEvNMT4S
hzflOgXgl9Vw3AqnxmtFoJWDyognRIf+7843gQocIYL0WRaW6vB0Epxhf/drSLbxZqhAobbwbBWG
hFAy8Os1r5NsbjMbRZXpM6BFo+yaSUXPoZnkuGKUL9uZJ2A6sHcM+RNAOFG0QRmdeZV7x9011GzR
W2D46GbwDUftsJuUzWmGOWD1Zsz/4d+LO5MemIWv18BiZoMboKv/8W+Pa3puuFehogHPIxoE8L5T
drVE0uAlU2cVdbSrgHJU4n2adCc4dwUplckEcmtkG9YU26h5c0fg/1D2EiX3pD3wWK59uYkJrFW7
k4Q5IKLeX9btZy7C3Wb4Qte9GImMqXseDPg9RWff2N0F5QLBTwRkQIGQ+on8+NG1TtP5/urA0NCL
JBIfVJUTjIMXqmvLy6aSCpz518L9Uif1+EEMTPV77Jvi0L+FhCLF5r0c13u7AQYz+ef7Wdme9Nse
FSZXM073K9Mz7i90dvq4Y6PsglFGU8dMuJkTd9CE3w8uxsX7z9q40v0qYAhEx8J65iAaonLxwbPU
cEbHzAWdKtmomMPZMA9B7f5FGnRUizDU6X6rNCjTGQcLP5nrrhLs8dw3bYDRwrvLigv4p8qmqmVl
cuUz553wm2+5HZHY8sa1by3H0L8Eu1vgjXPrmQXcNSTtCSAFfsmhXuAQiRE71kLEBWjqubp0xVVF
Fx7hJkoAY7dXdOtrUk+Zi0NU4VvV6nNobXeQggOvvcE/Mmyhu1z0sIJPsV5vNtseotu9RcpRHvjc
6Mw1xxgOctzqlnHcNufjBHCzlcXfjWCn8xqqfZOcPpVlT/n7XevcSHW4izUvY85SY9qvA/2Lh0en
9BSc+crMn+EAhraQ5FOoNOHIM0GCgIE8OfXmgR4P6bWrKC3HKlGpH4B2LJ/98ovGV9bTuWSkfCMX
Y7K3qqFSbjsPKvO4Ypvzrq8tEc5/Ai1qoJeQZIxSgGVY0ucylziLRGzJRuGmEtQAEMwbYoB8vsst
W9nqpDUffYUrDJmaTdkVkz0/xSYeZXP6kkTNuGYnQJMkerDeRbdnjMCqkfl9Ki+1+02hV//dEipw
95jFAxcSc2OcA+ZoBDCUcJvvLuB/o9zTca2lr6iBbfICKCKnQ32sm9ugf1RlmaoVAb8cCuW6msKR
oBRTywHDAnrHYHyoYeVDgBKOvGroqys/EvR+aP3cTMV/YSI2OTrzYL6CIdyqA9/3QBZWQHctOLRt
cxnxR52R5/cFqhogKmmWCnm1EMIsD48qyfx4yotaSsrgkup33yGL5k0irM34012MSZ0LZ9IcEXTs
IDnMTj8qLKJbfu+6/QcdZ6PywhnR0vv1kNj40HWhXK3/RA8nxCat5bFDcvNBUCIVnpBfvYJ3PYKo
OwNbUMU+3YaEXGQfm+FRUaKaeAElBhZEDOuFGlkCMRyv4s1jeZ3M7IikVB8Hxy1UgGQK5FQ2gyrH
i3uaBuSWov+BlGXcLSapyd0cvkCDZGKVSICp6aFbg766xHwysH1fEx8urgi3dyI1plBmE+NWZZA3
rU1Sa9VfZOts0wiCkmxZTuGP7M4JOpCq0O5kL6Hy5E81tJ7v+QfPOaM317KlEllZLMCrVZW02z0e
QXPoxf9XwyOIRi3RiypkkWD7qcPLW3Uilp/4yiNNVZUsMbFTvE4WxyVM90wrIOVjSuTT31GaX+J/
FfVspkyBg3rbGK5mKWT7wn31aGJ7y3b6fnDf6vRkFrXrZz1VBHWkKbKDPf4GwSxvUywYXN0jho38
K84dcvtaVTFcF9wjQcguIfyQCR1bHg3Sh7jlx6ZWY2OT9dkNZKjt/2URS/8RPtz57QKVKRBHL+Ff
ZJoT0bPVnLrqPN0sctwkoRQHcnWMuDeY82LwT2VBkcuT+XjiqtXiqytraOCi9wzypG4M/NWiyRc1
IdM8rID98q2+K5dtjNfMZEXWXloWOzBZm3La0Nqoh8kQhU3lcoeRbj2Pf/BCXAhJt8BzjVBTDQ2M
YpJAOyBn8m8ux3cUV72tL9u7rfHxSPzcxFSecu0lNNP0yv91wCy/kqmFbs2PCcqc2onxshS1MFWQ
QiSiGoDVc5tbhnkf88D2A+SjaWKzMuZw6tHVIrHwQe0NmWwhESXQer1PKfmI4vwTp9r4V41mufPq
G4/UNncXb8IFPGfnRwnLvbeYGiuYkZ5nwCSytnZpFFgBcfo0SY5Khqr9V38U20EqAKAjkVJSZONI
TnwxwWlG27MoN5YtuBSDVXzTOycw3oJAljzBA7fStJkt+1eGbfiKm8Tibcm2jJKiblHZy6cGd+gI
X+NadhX1gq4jrXDY5r5aDy0oHWIYyKVT+QK8zIUp4mMuU1LWdczjv2r6CoFI7f4CX+/0HRZI+dph
wmntBpgerPseNB5UZD1xE2NSqTY+ZLrghnWPpmLjDDZriMBPv9C3iaoHYdzDQ8lvnszqUvxw9HuL
yfUOQKCHZ/JEAqIAIIGepTpejRWpq/5XJotaEcTWfBnPDeKilPdbqcgzNKjle8jKBA0l0NW5FgEz
V9AT7SZLXIFWheUhDFfs6Q81FoklG8YYvlwCrguYH4EGqP0sAz/pjvIHL8PYFiQg2ZDCozYk5zjU
LugPmH+6BlLOU0xOczOyxFrqCWrK87xupxlAoee+yn2IFiavSISi7erVIk2AeBcAa7qOz23PQ5NK
5HIWteB3lYhH5XSUNEn77ZqJNjvQ+5eSxGqUu8O1Mz1dUXWhpLBEcDywWsHCOltd9slU9t5KVfbF
8RNWsIkAc9qA5AxLW94ECOcIp/fcduSRFbG0rQ0rqm1qA9V3Xj5hMDKv41EufVFB0YwMyHakV6T9
ZwwEm3dfQCci5926vCxFdDFFt3k6fpzKembj0b4XWOY8gyXzLBphTNE83pGQzKEuZe985P62R/gM
FFIdS2n9UY323lwUkXYhEcR6Hfocl7mEtFc0WbrtkKVLPH7PyIUywzmwQamuWxwaLqryhLe9cfCD
j/LFpr4LIswUmNoawncyI+wnJWmJauosyhe1AnXQa4bWe9oiAHzC5yC3XnGPQmhgKKJhxdjbAI4b
+ZZVmFHu4rdgQ9RqYF8BnQjbZiOpo4QqHFfwgWp1uKJIXW5GVbnVEFZ+sg26gx7Ig/2WdTb07FJO
c4ckaSplu1rTvJkbnWlHt8bQ05XjPBLqPlAjax6dtTSGwauznwD89f3rA9LNTGy4cuUfZ6B6JmJ4
GZu7B84+H6tl9jHF7GJ+wfQMIoMD8QK+VNRTfis495bBetvG41qwW8HmpONRicAdgtBqm3EMxSrI
9vN/Zlazqm9EfajHMYsZKPCkAzHEQDF/A68LPU1gQkosDOkaaR9mPXBtFzC5GkXA9ULXrfdvzA2J
R2KuduQ8L/0153Fs+a4qF+xlzPL+hh+4jaDu/71TAsbZxsSzpOZx3W81yeKFt3pXsxPXFydGj9CV
lIf8B2Pw2G1IqEoyXYqUTUpBT+VzzkvxZTWuphRnYM/ZAp/JpPHqfHSkmsk55SKzBaDPJ3GyvxhW
QPveqmahOMioS5K/qmBwU15fD/h+oSgR6/1jcz8+I7g8SdLfju7JNShtAL/mhXiz43MOYIph5Fi+
wGg79jZo6X+ot/dj/ArQq9ioJm4mr+phXDwT1HQfxZ0KT8bt3OiO9cEnvUd35zEuwbOWQQORBQPu
8JTDDaFwCRvVyvXkf0JkSKziFjjYU6SDmHvUWmtDavIU2MbW+WShvmpATmQPorssUvBK3ND4MdZK
d0MuccTh2KdkkfephVl9/qSj95GA1SibudkBIQOpAIpXfBuZmsqCzqZbgJaj3yUxbiW1HYtFSfwB
laJ6hxUJz4gQgAEnnUUTzynYtGMjRhoxHIqBV9vgyqtapL23wPFVmecSVKJeZubFi6janl+6u+lU
jFn2nTBylXqcjbcckyw4NYK21D2ek4MmSviXLgLmA/AR4w/XgCxQK1uhRyz4YQlTVxkGzD6pyoQT
61ZauH341MsEGxSels7v3f+9rq9gqjCZpuaLag+Z62WFagcrQqXp8274qr0kornsd5UB0fDT7Pl7
ldYZXU00bncVMgpxz4ADIrGE8WrbYtfEH76wkLyL3HRqlPnJTDAlNT7uC3J+eQ11uujatgrsylww
YSs9H//QaFABDtnmLNz4JDPq22IP/dZizM6CWEWotVBMkCyxJvWhUr1udu1WEgANn8B867Urr4CY
OB9qwJ2CTlg5tYzYPEXn/Ddth90ug9rAdh+LHlXy+nUbLNcRA6igvbzwKqr7N3C/gh4kJDUSW2hV
aFEXkMVl4z2bZFWdDpmbsJVgMasEv897Oc9+j0lhjFD5he1+XtJOpCdRM2qM4XWWhYXlO6lQYEp9
jnvGAwV/0E77KEQ0OHzj8lWoewY4LrS2EWihGWq/U7NLKaWsSBSYgvq/X9QyM6yhftjnUSwHj7bw
U1xrwVj6xWQ1u2i+1ETIv40TtplwvtO+sckVOL7DDhYWYK0YBz1g/UYpA+tGFZ93r15tVIjxJagq
Dn01RtELwL2ozSJY4lH5F8WAxVi+ooUDNEhQObZJU/RPPU/UiQNmmyIRn+6qYHy32c9Vxuv57+Og
dg2B6qr2N6PvRj5RrlMfb+ZLm7KC+m9Pg+6SfJGGZgnzqTYevM97MRb6yBNXbiYkzUgq3eshQJ59
S3jNClGORsEWZSKJM6IY/VYK8pTBGq60ER/X4lmhtXua940QSYPGPEsXEW0jJM/pYQbfphK5W8uz
ddBvb1/urCJwS3hwCq2GYQJQ44cfEKwVjKBcxiAmkKUFkwyAE3Goi1P3wxIDb9EVx9CbE4OyVjvW
3I3N3sCVywOOAokPhKVOQ1kOMayyYfnJE0mTEQF3Fu+ohRHo3G/XFhT8hozf4kInbWKASXDx4tWM
zJ9bw93A4/HcgrBfCf1YBmFaikEUGWb0XQ0gpRUIQkXGwreOksehDxHj14QlBXRchxWY7GjQb4Jl
aLTslufIHvawtq966/J7IgFd7znYfT5ON6glpw4jt+nsuWYghm2Jwk64jAWvGYkG/rto7Mx+th/w
0ZyvwXJOrHq9Wbj1V00Ro3ujjPx2vtqOg74Q+8O5cb/J/LXuY3VpGNa6FwG4NTDRzpmOZPM5CTBE
c1yONQUBjVSG6eGocUnFre2BYqV7QuoUYxtpHVHl8WEumWgmzCPjl3R2Q6udOfeFsYq8j76cFfU1
sLoR01+A/+iFJonDHZa9YJbvxHgjtaEdKo27u/U75kIGEEJVq7NKJWrLW8hl8Bt5xRw/WkTCE0tb
V16/dlz3uwLFHvy/b3BWuLzh3bLVfaUAfXecXJtZorIRmrsMQfqaO2xsGH2I99X/Myvioo7/jp5G
Y9mPejxBQywGdZVpHw0bDW6zX+XbPLbEhGAX10z+D8x/eIdf2Q4grWpUxDz2sgvejqG+n7nNxjN6
+apbgz/B8iUAluXQCCS8M33+mixbnRV8bQ7UzZSmebs90Oth+ygraErwy/Ls9Rc5unwQM6gYcoVr
aaDF6QTO7HN4B/kMYOV6AhLKEiteVj6dAy58luYImNT0dsRLw5SS2+1VkI2/r5ADqqLg+PLVN7rG
VsQQmRbc3h21upFQtSsvI8QJ2uWRyy3412h2REy4ONXk9KQAMxzpl7AyYXiPRqnc3YPbOLI5/uvI
oGlPE7YRPItcSh2zbbfAAE+ocL8EJ9LZRtWWwAUOSHRTi9R2tytgcICgv8EIbv85W0hoFKXEFUvp
jSzh/tADNNvL79g/9hHILAAb+zhQAn45l1pvomVO5AE+RAWZ77Ql4JHFRto+bE9vIT7slDomMUFM
BupzlJDQ9G5McKKB+bOi1C+08cHyijgStwxDkuBxzBNPweeZi5E4fyMi8l+YCHR8aVwdIrpGgpNu
czx2fZ9hiKtQEJCQlEG4lW/KO3FL66Yoz4oHEFbuxho2REmbtjN7QEV8SJ90/4jbQEORtTVFX937
OQ2feQ/USOJXHrmuKJNaJY2yu9Rh6AWZnRSamOmkxNshrCRbeTdSEG4k1EQGDBvmVFyjg+Bp37TJ
mAzBAp+6RdXnLQOyHLg5V6iQcxKdHzJ4H/2Fj7qK9CMrWypqYhnu6m2ZRNOv2/I2vLBV4S7CcSzf
mqLX/j72GIM5p84J1jMXfR1wJTLTChX8sU1scezpHlkUVS4H8PENAP4r0ZKxLe6HbgSSf/weeAQu
+KseICnadMk8gQ68yRfWyFz0mqGO835vWKzT4chalv5Yw26d73YPjDECanR0L5qJVIHhuLvwxMRv
Oyq9s/W7e6f9kF1FBtGY4A93tGf4uNQORG9uRO2FinUysJNklby8NzfaXyVTQhaynum+sUOEaDw9
QIQbvuEUzvN94hL44ToIiNv33vQqtZcnQ9YVzp/z41xX0ftiPVBfH7XUaOp5L2Bon0zWVXo17sxN
RbGjIF6UO812WmHesSzlbvWUOfg5VMWYAM0I8XYNuO974XTBqkqsbhC81J4PE9iUvNZxm/TnjczJ
uxiQZRsYdL5n+aKk7LMgMAPZjtTlZoI9jnD//YfiOSK1t/1LqMRkWH6sRHqk1L4HYlpGMXkZz1+t
Y10DqMDXRacYzRrhcUOSCDlf0XmScyunDJwa7yJO6smZt8Nhb+Ia0vV8G3UbWNHiQDGZNPPLTdoy
V6RVjodbXmifK/ibuR2PBUpNG/jd9IJv/KuentS85l0+5K/QfgBfUIDJFdzPW3sN/u4Zuj4Mtx+m
op1BWOE6LO6wiVQHnQN+QOJtFNx1VXXXFi2PVAdIIswrhXTdxACS8j9nARhyRg9LmGZmDM4/znw3
1Gj6sC1f/RJ+x0YPuV5MpUDDN2sVNrYablquV2XL0LMgqc7QSnsNg3vM1l3Nm3SLpKN95X00wvvK
UmAHWGy+AedFygZiaHnJSRYbTVjxsiTGny3h2a+qijxrse02xlcG+qOvhOt5lH5AQ4+XpHYdl16N
YS5jRcO4z1S9ZKLHcNhdh05Zz41Ssi3MATvbzwlYoxV6fZjAs2zd5lXWtoNLweci6NSJfI9DkkmQ
CCLKT8btjOF67n0H84A6z73G275xewx+k+S7mOcR0Gorp9dsqTnQpKP/K6fgC0cLtd16IB21RrOg
9howlHlrye7O4yH8n2gJrAjOshzSVOd/R+g8Y5vYDS3KL0ohgNK5npwsRAkZaUtbKvBRoCxtwXDK
SmMNq8tObF9RiSgpWPhXU48QgKFKFZB+/JsNVdTPlejNak/OPqy54Vs2gdZDEPsHFDKb3ILQkRmL
RtsCmVVfnEDmCPl4Vu38UZH9oyoy6KSZ+msZvAmyfUDtYDEGm8ftFnSXznXq5Yk99GuA45rQcrW+
Eipi4LsuLV6Y/ewEbWNa2s0PqsWin7QWOydy7TM/sl1gS6y92wb+aDwOg3q5ptwncZiFQF2IyJi5
3osvMtvvN3M1Hcu8vwNjflcLA4GK1tkRz9CEAm0btZfFIG1ifnSPs7fWlMjgTD4QwjklfxTcXBuP
/3Q6dMSxWqxMBmH6HoSCYTzyUu49qSOHZCp1IHlE5279YdwwOFQYJww8n6BHdhyOirOyxvs9CUbR
f+e0QDJ3CXrmHLqsR+/cx748UEeTb34dOAxnu96iHjl2X1bodKQh6zaOW8OQR0R1kh/uEKGyEdx1
x/w6AKDZUPnzeh/oo84qjUsFZeA4u3XwbRkgThpEAkFLUE/nOO6jRwj80VPFh/t4IRE1i8k0zOgE
tBG+wp2GHJvSJCWxbxSHIIreuWoZosKaHWrS9aLybHNrAs/0gJbYLmjnwosPO23S7AHdylQSJlsN
XxmgF/Wl0lhKkkVw6Fyom4oHQPv7mmRGmk8I/jv8NUjUgdW3lgwHUapCrQp04H6TWfDHjfJIpBi1
IchFe7DaIJexeeOzKsVVACISPCYL8wvjc9XyhsEW8jpWiHn197NOHD2fTDV9MLiT06dPhOgpgC+c
jrxzBHM7qGX+D9SQIC+SRHR9OvJfLupdADdymhqbZ09Dmn7zSdvGKHKIYFogvdG2H8ouViqemXci
ycYmKbmpxl3dM0ednA5eWJXveRSC/Jrt0wUrpV+cLSR8g/kRH/AJh8gh17z/98vWl1rXV7NmzpKr
HqlM04i+tcm47+vRgEyE6DyQQ1Ro7OB2C3fsfyWcuammCg9p74glgbBroxYNdMCLaeG+IAPv4SET
DiTz+4gZGDw44+8Oyo8LjS+Z0QGY1bX0WBc0ss6Ps5VCPXtrbuXAta21x1S1YmqBXKkc6zgf7y/U
X9ihv1sjxMnbcKEz1KfKQgbZB0UUXnCILJb7BtUk9hflXC1XRl5U2NvqXZr0Z6bwCUr/7LbIixaW
iHC3UGx44HhifbWMioXeSSJOuAlHw8xK0dpcrzestpfdByTgMRbVPCUQP3M8A0aTS8uLATPrb6Xr
RhFlC3IhnPXzz29400yLIpCM5Ic8bNLA4Gq10dQhgFGX+ID75uYtMqiIywh9z+oiZgdpQ9TDy2zY
/HXBCcG0LFlQVcmWHODUY+H8IgX5N9BYmo1TrGOzMrPd/z5lUOobjabJWi6Mf7l7K2GzMbR9XZOq
jjI7EPkIHOdtifwJKZcyzSRCUsS2mBa/dhP0/CI1XwlFFfoSj5jY0b1OTy4f/2RVnOv+d8JcPu6f
xI5dujgOycWFnHqtyMZimeS/EX5dDBL40jutsmpk2B6KwB+Zl4+gm4Xsim7A7LTkGYOef7ipknkD
AbdRctFnnA9vDiE+yo18yjXGHcdDusoKyzHdwrnp8H/s9QlIy6tYR2qsnnaCHc+Q6bNefAdTKZlt
5QconhyNZArQNiGRELKGsnkV1sgtBVZA0B0rIRbwT0CK74LAuB+5Q1k+je+PSOjFpgmI+FxSHwfz
3kxjM8C6yaMie9X5dziZ0ugvIFAYlr4WjJfBcbY2mTu5erHtWQmwyuyS1aN4ANI1Jy+Nn9xPVyC2
eCqx/bzonhNG68dU4uOwPPTduLPmuf71NmgUB4ObGT0w751dacfieYPJxz++Xuo6bFTZ1YZkI0N/
Vs+h7PkOpAk/yBHKf9y5FADhIjEZn6WQc0LAq6CntyDo4SamPToOlkURm1R01NzXG32y7M+PlqTD
2xS0752ackCpIJ0CR8Fuihk+hjIx2ggZsd2pHeeTg5LVXSjjcoNr6HYJIRP+SRQt11GCddAcMNH6
Vni2+QOKpW09r83GyMP5wmq2rVTqiRJmAijuWd7/KU6N2VYT9/4TTotHPwnzHk3kkB1Xl40VW07i
+cCk7oypUn2t9YuBdUoGvwCl2qu8pH9itiqJ2TMT9x/fQXUG9F7mkODStI8afOuHp6bZhekExb36
jHuWgcMjzjZmkYHW3YwsP88PyD2xmeekCthMKOio0lvN9Y4yzz0+sM79cnUXf8f08znlW6kIOdZR
EJTPePba+FKEalMdmuQae/Gt/ZaeGtHhZkxpRfBYBGDL5mMSjH4Rvd5PI9xzDChv95ULqbBd+baW
Blm4F+bF+aiYOcAKslJeaVlw3KYPAkM50sSTqCCcxl+5LzhYQdUkD4/lzpmPvIEhJy1iD66yJldU
sbnyaZLSR0L477kFXO+OP1xdXyKb4y2Chiyd4aF0LPIPzGJTLbCu2lFWZcjEEPr/b4nau4KJjKcA
LV4mefvKe6pkMEjNJyKlyHrTauKbf7T+enbYPnam0fdKAdfV32lJREloMDONnIw3rW8rxCenlHD4
7a/uxgs+5kMgK2bwMmlE/Lz4ZpVfrXi2FevBzGOA4W3mWdYwnTqJCuo8Psb53usxC23UIWdGoBnq
wRtq12xGU5peI43kPF6LfweLG1MJLDXu2UW6vrItpwHUB5DMmDSOgFw1fz9/5FO6jO7LIYiBbHTB
mWehRx6QTpQDHNCV7Njqw1bwpeyHftPxPRWuCRS7YpH04KS4MIAfs4biRDzIZtxYj+ttSABNALA2
xS245GgxjxMZnfePQR+lEUkOCmExexMBUJa5O4+/0c5TetECST22cbUdNm1G9q6A+csJKcfvTZO8
HraqPfHdn6mcr36SVG9JThVfnQ/f2QZxo6FfTzX3tijZLTV5p67JSztq0LuFaiRL87ni1oVKTKzO
Flix4PKkicjorDGGK4y/quhHkvbmQ3twDLqdClBFPCqfNCQtQnLAXX5AJsUqbGY5I4a4DzxfzjzM
5pu6Db1B+BiMcYkCsRiDTJfz1DglaMQBaRG74wqyTowAai+FgQlJ/gcXR/+ERDWh4ldqVWQbM+/y
7/sJIi7b0jDCyU5U2ZYVlAu/DD6hz3F3sR74VLjRWoKQNKIIQx6klHMuXnYWuJHF/XgKaHJp0tlt
EI8UInOTQT2VJYQlvLHJX0UAMcOzvKneQBtw/sZErlHViexyGUic1XTs8lksYekSFVG9phRdS/Ll
uSkG90eSZFuAvQml+UWF16xpUwIfMn6dRcW2T/beZMzj0NVeP6LIq63OUqhzc37Z9ZO/yS2GFwI5
D6k8KO14Pk5QiJ0IwTbcifJ8r4UdHoCl5f8bOQNjrT1mqDUn7Z9syMacgAJFPSKU5e5qM37u1XBT
byLw8klEkpPDguTiZVRRO7QpkcrYBu+yWFmP3bDsKdzJ9eCXdozApcGDGMcfBfkmxUexouXBh7SJ
gxBsbgTF6wLHDaptpfA1JfJlDmrcvS025CQ5ovKCbbC4AnlBUjQlQ6xUzwfWyFgSN78u/PQFieje
j5hRZVSwKKRpokXiPxdUmfX3EiLIJMlzFd/U3txn9ygoSFKDOlIMG9o2CT6aKDwNsCYI3z/rRx4V
RPkLN2a3v+1l98r1Uf9XQowVfdMp8FNwAuYAr75uJ3am8a9lCPOmi+F/IOTb/gYoZSylQqoywAR+
obApm0O+KvVCbhyJtPRg+N7gqUa7Bydhog+vsR0COXSmqr3n36jQ3oThKMTAfFHtrloVtPmidVZL
vmDu6jzFBW0ZzdeAk7ZrIMv4CHlFoEFIhtlqR0rlv2h5Hhzk/QIAYIUnqHrfvhBNYqMF8JSJ33Vd
a+ZPzhg6SGlmkfRYv8fWqCq/1TrwbrQLQTeC3xgB7ni7FSfosrJNFi9XGbojeMHsohF8mvyEzRt2
h74tAGUjjMRVDIfgSugqDuf29OZ1zP4mCytRv/kNGb+EsgJst3aF3aNQHi0eFhj+JAWpGHteHGp+
KlHPmLquiHyj+ARTlbSXXlw4E+f5ZmTQ5si2MQYTZ5hgGBEGJeT64m4m/Pxb7BMPa5IAX77v4XM6
Q1aG9w5NpqgeRrj0bRXc0Si6sXFIzAyMTolFd27nfYm7rp1xMtN8SwHkqlHZELvNsrtkAtq6N5ua
/fH3R/DIoY/D35WXJVApUEdperAlaHUSVxw5laLSsX8soqh6M7qee/sZjcrS8IWAXScsszDG7aS3
P11QjmNRnrjwccvLGBbWERoBmdGu5cq3HfxAoAfjve+G8Cl0nfIAX17d9/e0bM/a92l1NkvpseOO
2PbtlXEEWkuZAuIeHsJMy/ZdaZCJkGIp2wDwifiUNiCijAIaCklVRBdpWy0iKwmB+gVYTWiYTooo
/ggORrE14XHTix2h3CzCpjBk5eZsqkaI5eBfSj59KSU3FvN556dx5PFtOK9sMczRHSsVHI2M4vyy
uayfK/AWTBNDLVl8Hr3wLrsF5whm6lk+VSLpK8IaUGkA7rD/8ns/yNb1pF4XYtjVwAqLRi0qdgb/
Y/qsj7Tj+qoOob24WvbVHWW+ojHQkrC6e0ky+L1exTp08WhgtLV/VZfKjIlLAwLZWJC81Soy75ZP
NkkkUV0uJ8oxYKuHwg4dSJhvEG4SioMyNCGU0TgiTXSMDgRaE5xI8x+eYmQpdOu8eL9Kb1KsiA/T
BJ3CfnBcLQhUcoT8O8nKbuGo4jn70Z0a/G6H8PWc1m2dTfFkk5foqlkZfKdm+SfcGMkz8zXQeYMs
UayoBidnzxnkvb2N8eE2791jUYqMWvCo1+tg64zKxzcXYHrF+fX3tkFW8gbvoXQkeevfo7G383ZX
M0hYOH2Dycwt+B6O51cWbVY6BlNqnfoDD51BXspCvmUi5KixffKngaX0+RcpWfqd1zQpU5vQtPun
LtCEjs9drr+NIeYLH2QNbQUcw6WZ/mkrnzopj/JouEgaMW04IhAqfMJqg7JCpoLXvKREA4+D+4D2
IqSCf8TzX8yRAKqGyQxIn2uTxFiF+X1PMsV84neZspt0/ARiiQC0LSB/CjZJVTg2OEeDvkmlsZka
EMPzBGsTo5JwfruylWiklxMz5pzg7dS4CuXkd1TxUiODsAXlRtEh3YNiMg4H6r5DSIxg/VOZYkby
tddBilUBzOh6eCV4BvT4o9B/bO8836BIcSOPbwXC/7NDAb7JgmQ8AikrTnO3ZsTwHjvB2ShEOUgN
vB03RenmZAS7KyLXLfBcySX2wg71yGOG7IW25pHPXa828DN0WviNMpdO1Y6EitlHZrKQ6KFPzd/F
MNr8ihDeYo6jMKeJ6Xd5UHlO2KleZ5CR9G0AyM4cduNKktVdepwUJw26iNqfKEjtolhJh5s7oXxi
Qf5mevcug82nJsXgyuWWUruYa4ZJtBBgbqQVt97CIu88XfVS57SJ7dT2otkE1cT4lJrUEtRVhHsZ
FDXEVD3js3LpHqWXbbdJBwxKfsnzNDwezyBxhf98BwjlJd9bMQRZDNYo5MVJN/THeayGNqp4vvWX
7cbxeRk69I3nZDGV45a5BZVQheZV5ONUaIPoqtCE3LiGV6uj47XVqB/okbkLSC4//82QYaDnvGHZ
TmVHgn5W03GbB5y81cVxXXCcMLf1Qd6eMxThgI97jh9aP08GLk9x+QVRnh7DdxxA4JyggA/qPyOy
+FxBpMfBME3F1CxDJxRqm/KRYn/n9zttVksj9GkBkqZOMDNK4JKqKRXAMmVwcpHvBezOONnhQdSp
9nBDXNHrT7zsF1+v3Ym2FugohwQ6bE97mJ/BDd5nBdRqSnS2Eskk3yHsZJvfV+0Un7fUJDXJko7f
8PQ1LxeueycjVRv2+5JNi7VVRIU6YhbhGNlA+pFAZFSEG8RcZ9KvwueKLQjiowB+ACzztBM5YrSo
1Y59gVUG+p5FgZUbjgtUI2DxwE+o8zkdbBjG5k71XVKKZaEcL+RW11eOYFHfKPOrv0wlBEF+pDh9
oCyEcGejK+Y+JHvJ1oKq8VnTmYkc57BcvdLRF7VrVFeNCNLNQ7G5/qQBC36ZK3coe7V8EEu8tPTT
ZKueQYAfNCMbUcsp+xmNj6y8GuhSwPdrrPP9nxnDw+D3ni00aWexzT+UzljH3w9x1Z9ucYRyDnTu
VTztWndfPgkY9dG12O/foOHth4fWC6L+VWHCbUh/7GF25ZCJB/F44gcmBexXODE0SFV4fIJN1faB
BfGgXYgL0ifYdQZ52ZmRxJd5A3u97r3VT4lCGH9drpte+tso3uaSMPGhUYoRv+Cbn0KAXIMgsnLN
q8mFJtXE8T/ZX8IqE89a0B5AvcTi1w9+rRw3PDktBY+FiQcg6HJhygGFR36R1b1pOrTziqQjA7Iw
Pcyu5Vy6CQar+I5OhXwipoJ6aI9nzTljmVXhbmWDopCh8ZepXa/URMNVJgvYpPqC1PUB65Y84Q3H
sPWdSCvwM0bFP118ZopZQITmNI1MLhR998SXdxuQ6LtiHeujPXVfMVVxwiG5wzyf7TnzJj4bOeBs
nubin+wNrN6wUopGMLn9G1xgf+lXivXYkqLOmXrdGEoyJaW9VWXZQYNjy5N0u+svyMd9nhktkSrr
RfvqflBbZZePm+1fmcUzgBRFmLV4H3RLgkAnpNia5gZSM6yYaOzRSuHoQTdA+mDKRAIYLfs2Pmho
vbPgfE4kij3vqAtcLEHn6QL6IL/bqJSXtMX5W/aoyGVxe7G3R6YS2pTybJpVFICv848O0oTaHht3
LdBW84PkVSeaRo39nf0dIV5XjdB4vZOzmcr+FW1U3R0AgSQLBHsLSbHHCOtkuHKgu0Ui+/LyNErG
ezgQGNak1Sl/n6TFnXD4ip2OzrX6oqVqUzwO5Y8LIZsKIXAfAbGmWbvzSMXHKUM0nzjrAGP4aFRS
Y4qqbgIG+rKbR443BVshr5O98cpq7mtJLAOg829wHTsvrwd5Qd4JntuJqZZ7lpzxkom352SG9zsG
MOeKQv4uEg7AuRWdFOJNxPPsxnCnxsglVgktM4eBMw0QSVE+MNiZ5zgPGqxzBSXdTYtLJ5qewGKP
twFjx+8ySbdB79S+ZYndxIqhqyaPY37/SZZEWylSLgfj5sTZsQb2fShXPToi5UzFAow5sJETvK8D
VgtTj7wyRDAlsgIwl4LGfZBkO5adKGtdCzqA0nbItcfzTqob08tziLQuWTZKcTF0m8lO/vGBW9bs
i6PdrJyAtDC4BCQM/DG5a4LZPQdwymE5Fh1RFP37+uQAChD4OudX4DHD2DqLXTrYPPwx0Q6TNYcZ
1G8LYS5T5OhShFLiE21P1kI7sP4+KkIOoFJLTW8rdafif1jIC9YJdjHUFvKz1KUPcorn7t7ZwdYL
CTWdA9ig/1f6D7oR2UXq5GYQ2JILuGw22VWj/UqCDJnGoEimOY7u/bWtUbvhVwj/41e9oBQk3L/+
W9tDxlGBUAu1xJr8cD4hwYqO4EI9LcLsIes35Lzb+MmIfKgvhpkqNbssYVPSxuzTrwye0c1+icZ+
BDVFW9KdaJOMzMflmcrOYyrhOvMrmmuKReJyI46lkMSeiIptPUKFhFhofBY8pUNk9wg9OR52ZrMx
zh57t+QtUNfNMlxB8IEPZ0ok89IGFlmc6C6NHekfQ6TeJeyLvubuAY+gj9S1AUfsGikdSXqnn8G6
M4uLvEjk7QxH62JgTJDyzcujOgQKNapga2nLg9wWSdol49+2FSmmgDAm5oHe0ia2UJoeQEHtfaVF
IORvJGvI7mjSqEEhvkk13N35UkAK0Wgf5Ef2QAvDP60KjIWfcTJD/KOsqda3ZKGROEUIdsvmUpSL
iJYte15SfnU+BMOwzAYLAaiN+cnQRb12BfkIjmJg5eNNe059HRBU1WqprnnExLwbsQ3ghmLJsPd2
W4h++gtqxijxnA97tnhK0XdbaNBySzNFOjOMzUlVpYL7ZyXs7937dVqcl3XIYI/ByL69yAHeObDd
3hmVrrU7XhO0C0N1kH4EoX9zwvyEEUWSEwAEQOdmUCDtZOO0G769XqVpr8EwYESlH07olWCbnWy4
vaM2+giOR+5nLT2Oh/42n0J9JKlaGCf8ZSR9w7+R7U3h67yvYoqtCIxeEq0np4sovuFexw8Eozj8
uU9zZHFqikUr4kuHVhzyMg4JoKYZXzxWLjOr9Rys0rhCSpp5xpE7jEpuWB0cX4TM8dW2bhnVsA8p
4amGbYNmF5BbkFWCMrwnSGe4BotxyYO07BuVhf82p3DikxeoSWOMpCcBEbB2m/diSIQYiSopexQN
uC2roKShSxGUNgM7dlNCwGSyD7uzKHAVZfRcWNkDQREmbsSmiS9ZEBO3E4STjoywJjisyoHkAKMP
RQv3p/4vgI5MRLNCvd+IHWHeBGDbZPgq+UbhXH4gLTr5OTqh0a+8rtJ9vIG6QlzvIMwgvdS1MXM2
KaaIHGKEsOsk81xGobKf2kVTqQe45bEW+o08Ml5MF82CAMfPqoawi/W8ooolOcBeAkGo/DqhTBFz
L3DtEAeVljtaeI93hTudbEAUVG/qvPSNctmsjmD9y21XU5dIdbUTzxYprO6pTgSaKQbNglOi6oBl
0ZWhJj2P7CrrS/ZcrBaFZPCOmSOmZ+qaxF0EfbE5oNmk6SeyfW37jchefbKB+3L4J8koeeTHzoYO
PKNzRonIAbxrDLXYdkGc+0CVjowEC81pRamZ3PXYOxplrPW9bIQFNdONbh5bO+zIjv4+QVnqri7K
Vpmm8DDSkd1jD4SSEjJDe8olWhOFIS6NcHTfb7hvIZYt+NTK7V6IlHbydzKpYFBVuEBHZtQwWzXs
+AhPj3RnW7Ou7OGlEdlG6ZrgJ4PFBst6ohxmJ/wGg6iLWLsXutBWVvfU0MjfPzvFj3VwUfw82jp5
89RNoc0TSstP+zxa65MOx01IN+mUVZ0gTfM6QRAOhkg4+qWh5k/pfy+IWaYLbfFiVa/H1JQ3ap7V
vIaVodg/0BGGox8Oz0bmO/pEeNG/zXItZRbIszzDzJ/c0QG2q6LTdbrwopX010gIZ0MuLFgbmsRa
MND9lBgc8F7EhyOXGaWfGjsUO8iyaZ/NaY9kHk9RcyTd39p9uf42PJlKm89ja3DTeOF/9ZHAZxtb
s6QGTdcokBAyFHeb2v2uZyImgAXSMlcLYEGkMnFM0aUh+cX2Y28VIJJB9eAsvnH0i8WYZFsg9jcb
tfbAb8RZ4AQTQzZby1XMB6yFRZofN4RSE4Oa6XCh0s8s1HZZaCQsR5z1onewePPnp+JwTpw8U99w
WS6lpbvuFRqAWSWglAIM3SpelQKpiZoM6zjJYiD4igzxP8ygWtYcqkolwc/1qWflD+jvx+Jy8bpE
Swz/WLqYJ67qPbuW+j/mRPzo3Mb7rKHAZCBw0p6VkpllZMnWwTabXmw6ZuS9YViM4Ob15wzONj1N
d+PZSOI7/MjmLP7ysuyZ4oRcqDjvswQJdaoGdWXXVqTVXw3QqpFPQ4hy+gr+xgs4Bm7m/ggoItZD
37k/riKvNia0WT4Vkws1rKWJZkhLzh7ALoHY8htxnFeAdReQUswuJWqVZiQZG/tW1neudDLYE9HO
H0dQIiYK3HybuiDfD26as5cxMMSSIVu4Ga68orVvtyVpAMoqI5Xf9f/QrJ8KI5+GJMYxUusqSVuo
+Q4BoPCdjPJMqBiM4LmpQ/T3ShmKXUnJRTGqfrmx4LrQm8uO1TQ9ybntJII3DyKx6OozaTft8jZ1
2hdyvFV/zQhrpttwcl8CdTtWFWE2Ubp/0Z9UGyUCYbW5a0R7EkgDeU9bsNPA79cSo1HmB7bjYP29
oSy2TKIuwP/Emm10F7aO0qQ4pR/SzPP7j/dWYwfhkutIP6UVzvDhOIch9pkRlNQdwNpECTipz1Q3
7pHajehEnTsAtkOBng1yExlRiOxcgufq5sgnRsSJHnD3iAp/6PUqU0Ne/p/rRSVzUeXev9PliG06
wlLauQ0fydZdkpFElh/R7nE5lPDZDHbjVoSj440cGtmAHCTb9EoUoS4wl/moQI9FJhnj95xEKW/K
PqAlSUKUDqrnOxeKkFqhrlnSAkejQGkdzkSDkBAN/SpeCu+fMpmb8gPCW/HIKWyesQ2fI1DHN7z8
GSXblZaixtbsUSl0Lqz4fE01/eogL1m4FYIaEndl287P+zoCiHFjaU4RDORQo7UyCcGWAh9kql7E
+iKPOKoRRSA86gUoAfUrp3UDZcSLuFtje7gyIITFgUxWbj0mVBb+9RyaanBO1HF5enyOb57uC/mK
5XuXcSjcR7eMqEa5gkD9sCgIP4zWPnQgYC5AmYz5yV4bvkJuieegyWzYXpROFZYa6NV7tME+8mcb
17fy8sLhLZSY6cl+9l38SEKbu6F6Qa3ipWiCcnTPJVIwL+H+U+S7yZnD8Qzpph68fVsedYfxskkO
pl9w4cAoJWl5xlY6Z6zpX02Ys0QouFnwdC6oh90EmpVxdwnCUaznRbaYDpr+68m7xV/+BUIcs6Y1
heD92WSWGoAQvRh581pE6AohvW1oxvo9CRd2ipQW2Vstk4K6A2R2wPaYM+p3dDgJaVV0CCC7/P7q
Cs7HBfnWxxuNtOYUaF6u74hJTnFgjjk7XTef+uN0AG4nOq2b0Lfmq3dzOhEHy0imOWw0lsAwtXTO
4gXSfsDTmGale7s43bx00oZN5FxDhXW9EkMAGL0Ep2HGOCMU6qhwinpCVHwAby6UVsiGcLQjVjd9
Q4wY5vELJ8ycbhUzfLHu9bzWPJEflVl5KNx6Ffjt2xfyPfhhGl0ZuWOn5zLo82YYeWXl8a+r2TU0
R0dba/o42mGf2ieZ/CM6Oq6EirbvmZOhHI+rG7kDw0rHKzR/RzUe+vAZ5DMt2TBuKhH3AO1w28Hf
m+6KzTB3jbpoRhs83R7k2WtJsotP1qhLf1k18W/vnkgImvuhmAH7cDTvxYjeOF84miQOhuBtWwlg
df2wQ4P53D565v1l1q3zSY9qi4SjGgUtU6t91vlHcAlACDOmaaJ3mx+V7oXHygAXeXV4e+DTEl4N
paoTUZNSvI1sbwrzXs1/k3HH46wZ2BEO3JlwXrUs527rZzDXrQHl361z5Kccs/5A9LG7uL/RX/tx
h4RafSD2DNYqFl69r6+u9eHCOYvv3Sd1gToL1Uk2KDZd6X/gKo75gV9/Svkk7A7KFV/lPa62gFye
qRMhxeyy+PH/OuW2O7ZqSrh/RqGyrUmsV/s6bVIcZ5Vej115kUq6/GX7M/haeep3evwWzT1tJ92s
OpWL8UyX3W2f/IqQhXNFmmR87mvZ4Ca5uZjqeIfTNvuEl6oyXJbLLRFWZZWPGaNGwOBxCInFC+tL
sz+BR2/Z1AvCFghImmlaVE/1wL6kxMuu/GddtVv2RPkcJXTyBhWgdgsp/fMr1lAUZQNHNdqOXV5K
0LnSb/3NWnV4aD/JV58s/IB6yjge5LDfjwwzV4PDOVbyt+OrllniIKwXMERquOd71jMBKL4LJdw/
9jllfIpgWZRVv1FSLUdsR7EWy2/zdzADUhxHGfFTjoJfu/yr4NFBVkLILoN8qXh54bqweInBoJFA
BGZvCjC04cD4NSP5IBrjOLNlSzHvBoNydSZypbUYWuEr3KpXpfN6cJfDZoty2ZMSDRt6Lfu+Lewg
mQoXgVaFNYkgrwDwGTTsvGw6ztaxd/EJpgbAFakSxpIyRdh/das/ToISFFHKHo5p/YBO+rk0cXTt
bUnoHiSEon6V7IpKj9HSF/9F7/2T6THLh0mMjfOaizUbEc56WvGHzBnnaWWwOSMIGVJbUBv3kp8y
NabvVnjtwoq1MkW2mbvslvkPx0N8FtsjxFoX7blmHJC0CWtf6/KG4GCTpul1r/ZQPn3jAqAfUVO1
njIPLOAEch8zTTyureEfjiWlhIcgiP97pAlfxYYxk3mZfLuKGYgUFTjZZAy4Z8f5xMg/XKkkkU0w
jIA4MAiLAKqrSSHoFbk+4rO+IIp4z3AHQaAt+2EBgHWOGhtRLzpdMfNgnUz1F684TOi2Hunf7A51
e34UUrjVVWADNO6M8paY0QXjTqK9VZNTkwHpeYzmhn9SOFkv70KWPkv/zlyS7FjIc4+4FXqGP+Oq
1LHfcCIgoMMCJwz/9JcBcUwjnnpYWOSROoP2H13WanP32pNzdo0PdU9qOtmYjw7UqFA4LhhQ94cZ
eOHfpTz+YAGntLETRaQHxL3h9gjRjv3VMTdA3WbFGlGqakQZJRzGp+8vVgp/ahPVupKNXsm5LXAM
qmX4Ue2A1f8BFbnSQxgEMnv7z/XVgNHGvwvD/bOHYyNcEZJMUBoL4LSsm7IWhPVGJ/nvU4XMwu24
v1UahPO7tbSZ6HEL7+D/y/1NOWA4A1dmWIU7JJY8ohFIZ4zXCWRPs/jnG2wAEz4VRlz2c8+6aLtQ
XswLScZHFs2UrjgLTCDUhT9AFWdEXuyb4lPJR2jEWFd3yFbkgtnBT0Acfw46qsyR3kzPchHHk0/7
BrAVobQh2GlgMntVHahWT7TBgC3pdlvIYikYf1Y5QMlv6R2cB0wj90JhPguLGeegdOGOHaEeGW8a
LFAXkLCjAgzEonC5QrjnR1bl7ouEI8EXeISwGrULa47zoXH7ihkJKA0BH8Bsx8gX4NW/IkLp7kUr
WKfXUdDGw9ROoFle87OfxAxTGW6ULV7eQlDH8jqM2RhMVbRiFn/+Ct6oU6I2cV+/DObsqkh0g5bM
2YXVPiba/jH1kRWdiON83JUX6H+vOBzzVWe0jDHDv3Af1SqQPMTz+US7bHbUXQncyONY9dTc311Q
NzAkqi9ABweslsSJEPwI9EWZDe0/YAIiQIa/AjAwu+cEL/B8Vi9/CLrG8c/nKqnTmwosrZbYJuG0
EUQYdspvfXqc5AGhVbl3lf+WySeJGu+LyPMLnapi1PUC7Mzt6uDGFEdnMg8/WdqUOc8glL1Az3Uj
lABR1StLT7zsdyIueloXdw07jZRpO2glGqz/mpSpKfW3zMLnJoUKonN7rS6+Z9Ianr35PR4wIytZ
LQ8JW1DJlsa11Iike21gKJOPFqO1aIwPITaxrJnlYAFD8aA3Xe0whDt2NCCgyDEyMkd9pRbjUKJa
cHU8RgHiohkavMVS6YKvFGBgudGOJhQMaMimZaAS76Nwwhb0MQ4fyzJyV9NG/bOerourgyJtjETG
kQmk6N+c8MjMAT67bVtIiw2mQtaU7CtOVRPqyJ+PBZyfXpmifRryTcshd4b1lN1tXAeL81AHp9q8
iyHnYAecmybzFB/vFTgADLaOMv3/Fp5nFtAiBSVYTzQdBuqHS5jnzhNeDbOekbXQe2Dv23jvc+B6
Y5M7s+zA5etcv4vgxS8OfDL7Ghlqd4Bu4y5OX6xCrxbJEZrik9wD3kfId3fedv/mGCYRP/vlIUXS
rH5pnA3Ou71IbxA3AaPVrMcXQui2tPUvQwMXCQkvDr1grPV+AXIrRayKJsP8INqgFF28RarYKbiI
FHoEL5aUPv6dyfGovKnY3XveNydY3rwVrG7ujUGUAHix6uZ4OOf1xZTUUVSIXfVJmxHVtr8BA2WB
PiOnesQ08j8xcWqGkxWndZuaGq5p27XOYRU/H3lixW7Z013uHp3UKOq05D35CdxVCYFVdXRz4FHu
Tv888O/RDbSOI+IezGa8JD6nuc5wwz3uVrCGnNobXrREUlJ8gCPgJeYAnQats/yKuvMQ1JTTOeE+
hXLtfKrhVGHDQSEVK4K6hDOLflnJrbmRzYnUcITcAe2cZDKXxjat/znqV1DN2zlVEcQv47eKPo9y
xol7aojeIJMogZFXkLuYjjHaGA8K0Bl/Vcl0VW3WStV1+c02sHxsORS8rXZUH9TdISYvbRcyqsJU
xEWo8GmBTUaagcMQCO093XGWl7EfIpSw6bZnMmaJ6n3ifxYx8lv0QS6EXj0GvgJGU3oDdehcmKQr
YQrKO4lWAqgCQ334ZGaA3YJehq3E5697i7Qurdp+CvCvCMEUe84igjhAJA+rvuOszW0OPSvcmMSa
BewPzWhfu5Z3ZMOMo36weTdDMgRjIpKx7kPt5rb/aopacUWSKtaAoP46ZpIHImUSQM62tl/pQw1l
YVb7XjJbUJu+IvagwgMyj+dFTWPqqvRp1UsFlH9yk/7BhZP/7LAbGQwxehThq2RRe110vQ9vIiUu
eQHCPKlSrp0MH8iLsWKHUPpirG64A2IuvTQx8k4GbtMBpptK1SoMh5M0wWQbVWXrJSs7QptrPvij
PMuoRh60xIjG/+ADKJhIHCHDAPqQn02eqPwCmtjZw9/liyX2JUxNIPHpQAGao7ujwzEsd2VtwcZU
to7Pqe78pVIijE+QVAIW4vsdVpDnACG8t6po8a9WnOUAD/JbSOyHZCoVJzabfi50otbmQXe8N7dJ
hA4PTzg/m/l4RUOAl2u2nha7iwdID7Z1yth912yarOLq7cp8g7LFxfL6n7fCLpV3kbiH8VY2r/nC
sj1bMkDtwG3bIdBivC4l90Q6wpNwjiJLJ7zYT+8u3AzopMfr3AA/661AU8YRgQHV14ceFGRMrE3P
dX7qMfdWn/QvTKBiN2jYCtAPPQzoYSx197NEcOdTc7AyTjmfsTJZzVQt6hUoImWd93UKxN90tY1g
ttQ9+mzdvEX0ztLUxzqPoTG/4V/8IGb70/IasZXpB9hIuYpBomXqBYpdmGFpudUtb3KWXeBhAFD4
CBMf5Wgj8UMlCIGJuaroL6yQlKIYUvLhvkRDjuaC3jp6Gx14eUZ59X+CSmZaor9am1ITteyYQv7C
N9fYrgXR4o/tdGfABuXQIMuWzwGSkJz4LHiMKHCEedgDuGbTK3xz5hOIqAECk7srEU7Jb4QZ4TMq
8aVZL7aNsllD55g6hyqkajzaakd7AQvGPl5hNo9VZecSa5NgYGUJdazB08c5L7prlmjphWXoieIr
AOBw5RqqzBrNgE5iABYAohOCLxIZUCpui+s8M5Km4oJeg280Mkl0nwdK2KS23B1M1azVSS0BbFb3
ipoN51KiePVktNdAGoWNrfGU1UiP4ZnEDd/XK/hNm9gL71QYPmoqWmcKEUJA2ETKnK7CreU+8Qcu
0wAS5KbzIJ3Wjrp0x1ezdbQ3LpG3OMLGyLmvCvcR17g0+JIj4U4ZnVocEZLeJozCTIZgOtN/Zdrn
U/8jMatkrcoZyRcDTT244KBGaoOTIV0GtPQ4UgXuU+U44SOGq6Pk1SaCsDOkPIB9XF/2ILhVEfVR
4dK+Jeu1fUH6IHWbjanAkonelPZJ6BdVhV0nJm7x/ISsooFsPn6QNfamY6gRR2IHb2datmtJgJ7P
NyKaNWczf8qLMpoieQVG+YomWChhr2J5z7OoMADuEJrI6etv1cEPahu2hm9Vf6b2UO/eRCpgl6Rc
/SGVH0nrFdn/HmM7ZDyPvcznokNhi2J3cq+iycYiQHcEvvVvibkkK147qW196/fXDzEAjwzEjjeW
aVYj4qEp+kQHYj1TnLACQZt7d7A12M016lA2sxIR7/kQmqesNQn6wE8TuguJ2wspCQSWFv1jHb/w
tzjCRjhIIQ1kaQgkpZtP7MkMhEMQfjcbp4RD4sQtWCy9noDPK1izvJFhQBnoHbiIUInFOss2MRlU
6toQ2pl//HBlU/4XDSJ2qUXqWPb+/RSGys3IpSGbJBuKISEfIbn99930hvk98i49eZMIxOtutlFN
BLsuMGS5rWpUwPQGEOGPsUqDmlWu+PB1dNzntCv27WOG0myfA8n0hkNPDZRVuL51Vw/7A4ilB70s
Bre4O7rVB2HFV/nkzxJZUbihHm4Vdg5RQcQp9MgT6YNPlMQs+9KcjwupIeI6HC09D/PPClES5RKK
Y5EI0DHSktkaKVQbSclx+/Y3IpyFMz4r3tALpX5P75UaLaCVm6UI3DLbL8Rdxb2np1lUmKSoyiny
DLySlS1UKjwtNol1QY2ndSr7kCBg9DKqEe1oDqYP+hR+x5pVkYdBWfToNdi4n+1BTDMl2EzxupE8
hwkYBA+VaU53TYhgd1ePZxfvr6kZ/Q3NhEhg8tS9AD2Y9S9pXYDpFobYx5ztbKLGJ5lcRY2vV/b2
IweAxHdPrHnE+glq3Ig+qa22Cq+EKG+J609qdEaM+TAcMXJCIB7FGACnwonSGO1+/iUCnoXOUR5/
b2MBoa2YJww+51z5XGnfMq+c0OXJgjY2u2M9vFZUZprAJzF81NV7fAo2d6BKXrZLppkf7eEBK30w
IAW5xa3kzLoCn8Bu69v///4boD8JdEK0IJVgG2I6geDi97gUh+LxgEoZ5V5nKJ3wdBnZwnpuN/LJ
7TtmahkTPxa5y8npyWflwk61lg7ZDV6rboZ1MxOS9nMMuIvIgZKx18/dDZ5UGV3rnlbU36qZNogY
wtwOIoTmtrcjWm4Cc9xboiyIrsO90B4Koy2VKX446FmmGb3Bu9Pih0rIsRWJP0d7trpsz2LcWXx5
a7bj4WSWOZcHB7yLgjQXSCI6dZHTLxoFNiVAe6NrV0QifiD6fR/7PjjBRKL3l4J1GSxQPY50YnKQ
hc6K9f+YONTv8o/lykB57RVzDMwWI+UB+90P1st3GDKCo7bledO2u9LVI/oOVVktfSu2Mub41BQz
w/zidPe2UtgilurYx5RdUxKdp1zmPd4uds46fPvwQnT2OHBHU1lPydHpswmUiTDjWsQu1GbyZWdt
sBfXWGhcjXWsPutIYnkgYyiYxP2EcRyDRRHqLvOhWvFhv3RJgqNjvzs4HokI0wirZfKOpKrtCJ+y
/VaHprDIWMClZyux8+T4xKmpFQcVFNeb7cR0yyx2QSxbi0y7nuFbrqAfnANjBu3gzONRwgRKQzXr
gN2trW7ryydKINJrtAoY27PjfXoggm5ufhaIAn0znoMYDhm6AsSNxM7MsASHPow8mHxDs7Ob6mu/
xGHK0sHCq7K0CdXqdWd7K6g2TMOp+5iJCc9ZcV5332oAkTYfh9febM8ZfSkqSc+ZZVHgQMYlOxBt
b0N6O1SU8P/lThQ/xcPMUledbdQeSjfFzFhQ43++R2bFEpMSYvw7lVzSmyR92Ic2IX8zxPCwJ91d
pIInSY+bwwlpUu113lbujhz/zBNhFRyk1uN2eEVeZr21///khFOZUTmjH8aWA+B5Sml8ph9/5/lS
P8Dv6SESj+iKGeFekj4x7YCSGcLF0ZlBgJG37/bS62Q14xWh7CaZdtzu39ituKrNRirjUmIyGlgj
w9lu/B0Zv9rOfiuvMWi1bxNneuva13UYjcHlIf2BOM04fGe5qMzypBR1Uk2cPJQrMF3SYE0suUTn
0fy0WeNw8x7qZ4OU1So5L/n3nnvB35EUboDcIUArs74JoBFon5VfexKx/Qi0xblxJA7NLNLujz7U
pm4Y4aqxL21FehK92mZhrcBmkg9ucH3/yxgYig/KPvYdGTbXKOHfC4sRQoI1t4oqzJFU+Svx8FHg
UmJCz/3fYA1vta3cV1P7EovG7POLcmnX9oUBnarN4kEiRGTUTLzxCHSCQirMRY7PCkmNyjlUODRM
nfMaRnVcrBDIB/wOZqCQ1zVErCQqc4Zus0ZR9rRFTHdlCoqcmVU0Er2GF7vfXC1ejkoDz85iXnD1
6rrhwrIQiU8BPFAQj41QPrUJrg/Vdh8uTE6uzHPJEGZuoYJh9x3Bad3uaH2E0LuhL7wFj4YHoebX
L5it5kHSW2EBPt7DykQLNqscqUuDNsOAF/U9tCVXOfyry+ZbiBiH/CQETrmKT2VmXTM6ilJ7/TTM
Aoy3Hshr/7YI8AMTSGqD4hCeRUT2wZp6U+RAprzh7CcFy5Ct6AoLEhdxgO/5oSGqgvOQelsVzh6F
3EQm3NJrUJN0dLlPm6YRLma7zWOVwXvT2fU5zE5mRElCIFoL//0jXB2vNsAQGbHRfQVNOgqYABjF
Jnw0HqMUjUtFGo9Ir4JN2n4uFD4yVa6Vl9p0gWTx3rjQnqLOrpLRchdf/xBBcuo78hF4L4/MWAho
uvcBIYOOqWVaNW6Qak65oPxj4WaVDmkaSstG6/MRJbjRsX/L0H/B9EpOhfnY0Vsolbn4cGc4KvUW
oCLEUzd/SCo0ZARQQ+4VSFyq+GJrs3ZqKOTsD7Iva80cOEYX5+IhUPcL3GXMgznaxzO8MHyv7gv/
8637eIBEUSx18RN8iKamemiMSPaOuRlNe1J8H7yRqaI0Hk+/ufj8XaZnIql89UoDU3mvXDv/8Moi
z2iCbB8mRg26A082Mab+XZsItxK4fKegcuOtbawYphPiL9+BEQB0faubK9rglRJbxMQYgYNFKb5U
D0nbENRZxv+VC1xtNV84iqUe6C2EzaJ/cz4Aff8/MsU4763oVPqjTrywbvh1o4etgdaxbcHEysA7
3SDrM1dk0nj2g3Zux0aIv8UjJ3cmq/80zrEbUEWK1vIwYjb0x39P76yX0dN9NrG92tv9DYWdeD4A
DNPqHeMuQN7pyAVb34CRMR07onP/XwhKbDjOFWvdFSe5L0nMFJoaJZABY3dkw/t8iBhgBwMfxuKJ
4pPlg37DTXc0SX77+coN1SjfQ1mMZRRrymxnLqneMglZ4Pg4aLJqYoYT4hamcZSE4v777h4KPv+S
rlPWNOYaj5Gmy0ERwkKwYAqfJHJL/+C0ajaoVE9bBF1HyASInJ5D95itQ2sp+3NnPnje60f9Q4Xk
+WTzwrzjSw1iWSoICvN+dywvY0a/q3FtsFUO+HHJLPiOXRw0CxUA09KHI4PS2NcefYpExAKB/90z
yUguALDBYy/sziRwuo1JaYW2Sphie7zo6qJjUvPiw8pt8m0npulugxg5r+24l9asRgEwNX8OQP/D
0QetT1wfrzSNh/u3q3gZCnpZ8tpOtO77vzShh7/5Ttn8vc2N/+WjVqAxnDkOEu4umJrjGLFLaOqJ
IuYEVSlFjw4sWeI1wSFnGHWl3LmDufckFPW6tbTeCAd7AN3CoDXmsCVGLECVP0OlDd0tpzBvVTIp
QgBCb6PLOQxOwmNeNbgY+530a3n/JGTGT7R+yhNnwiiyXCaq2Y29+EmK/CU5CQULJ2Mmw1qdAzJV
Dirwvhq8DuI3Q5YW/4sHSxVZdeQtpluflbOiZ0KDSNUwqH3k2Htjxa7lG5EdFvUzN63klQy4FTO7
F+taWNj9ppeLobB9KPNULqUIFKsdQd4ObccEnIk1BCbYb6s+IzJBb5XI5Be2D2huD2VoxR+UmOIj
KVa7AFSFGklG/DSHZHQ9v6piEkNYBf+K37nenhUnGUJvtGKj0+nHKZWv9jIiW2sUsHFfG4Q8ooJC
yoZq0YfRmwEyTNXcONtrDaJn44d3uBzAG16Dw/CbQNiWXxsKUlWrNcI95xDW62uw/FSWf3l9vu6y
Fm/0f8BlfWV+9kKaHqkKcYOsaxXfHwSKH/y8N6qk5y5QYg+AZ8BHK0criKnHqZf9i9ZOF0I140vo
oWKamCw+//jDsNkVYZjh7CNIgBDEoV6c18UzwX9cZHIUEqqp7kvpX+WyWoRQ0/Y32t29hjXQ76TD
Tv4RCeTUcm7wvYswQCSLUtsHIL9RHiej6hQF1EMzEbJQQTHLYOZ1Whag3jbnTkn75PHqXVGrRNwc
h/ncfyhFihvrReYE4WXIYkM+jnYl3h5XN94FNUE97D3mr8AFAa4uuhvghaEpw1JxvU57MtCLw3z9
sfKPdZkvcq8SKxjxWxVen8okOCjkrXnWvOqwx8g3gLb2BTOaQNWPCloDnDKoFz5urII9svZ0+Yfn
byj63l6wbTPLf8R3AQzFgt9wCtyjyP6x3y2JvgLRDohEkWRvHxtrrSVTn31oGCTwCDWEqLN5qOp/
J0sJoQcrRDpWoC072VBfKlojYEywqJDPQNyvjRR6vHXbN5+ddRqEvpqv2DspZyiRuWs+gwKFQ6Do
FE0GVWEObB5KrFwMGjRVgaE8GvO53RBV4ThCxGcoPG1zNLQW8iSgeA7mRbDn5Q6VmwkiN7zKH3d7
SGo5Bd0z+YHli3XSaEOe6IcH/XRhheQUqlbywiCuoHpfEhYnJ6AqkV7ex7CXdXafTMWZgT6xP56V
hZWZAqcH2e3CWyHrjCBbKyd60suDrzQXXIwKqWpzA7C+5coU1lE7zoe7R2ezdqDip4EzevOeBf6H
uPAkgZLhJUhUl5szl4NhQe1X8eF3/K0mrF0Q7uGB5G3aZiWZgswOg9ekL6zFHtRZ9ydAZN4YzJhy
dxOSDkJdVfpFyQjZ20978//f+L6Xf13WuS1RSW6I6+hGM/1VXaUdkmkFT5j/fKDo9om+qUuGZcp7
6K+Ox2fBW/iB7awLUqvZSh5qjYqBIRwC/dVOTPX8QBeufUuQGO50aGyiBCXz8IYqHq23c/V9R2TW
iAIndfYMHl1abinHyocbUmA9oPP74J2DB8DxDKodOUToW00vguy+hOWPUmqLfjSeYh6fOX4nUJlI
Heo/6xA+xeOjjH5UmQSuZR4H0kRxyRsopYm78uXxIrRds2IK5YM3ZkAb5/PxwsMaLccVW5Nx1tAs
1a7KQjH56UD4sRgJsPmeTEZnqJcEJ2eVmieUm1VnCaJlzVNTKFzaLfe8Z9B9vblkmr8HnOBBB2k5
xctpfhRd4Fkn5D+Sv9QYpWIIK45aYBfNw34bcV0RWkEUhhGkaMrFX1EVqNWkGBHSiPXIpu7OJ0G0
wtk3UORB2Fl6G2tBkXqZwVLEWMXUeo0fKTzUJ44+f+G68HI7Wg2OMZshJQdnMBIa1h/8ha9tNjrg
H/I4U33FFxB3F4N2Drmmt/VlQ4viXWosyA5vs8rian//NMV0VlQ33ui0htUYFtvm3KgbRo2Ii4fx
9pjOle7wSNOQlkqS82x8ZY+EliGZ6bvpqCgHeIEuNIAUwSusw9+BEknW0f1LmrOgWZRLwDowEca/
wC1N8IPlKieYZEvOm0E8zEazJZ8dIlbjfTPwvzpIc7HaviExmwgJkhb8L7QeUSC6UUXUXi9TMjWZ
1iwgaCe78kKT7RkEqLtYY43klVIlm1fJug79nnOSgwHNCJNlZZoM4pnDpOUhSvtds9b3QXkV5V9i
qSKGHmuwOSCZUIoGKhcrIHnPxx+Hh3ngcleKJIMjgAdtdvAMXqco10RB4dcDhtIJMzYX6s4YSP4/
0/WNzyntGeG0h7wRGRZuK6gK3zy6PeUJR7vBnfU6NImvwOqcjur8kZYNiF09XTpEw7jYImGSVVOt
qUG0sv8mYc6cooXEapIYMwZhXHJNyL2j3XYMld9ZZPoOmCFaNTSppF/9s+imY0pHi8stm11u935X
cOZfmr3z/JxL7m5ZVsBH4Eq41tHG9haC4J8UH9Zq6fExhENhIy4TPIRrKUMy1UrcKJubon6PD7Gv
nHf3Jx19+2ecv5zNC2bKcQS6qbS0IMatd8VrTfxEtoDdu3Wc+sIcN/TjkvSwh06QNl9FhCIcnvkd
gphiIoTEVM8vvDMHWRItwyXa4708yGPiZRrCbuytBfSXRmIiftT4iKw7JO6vffi0GGA1/fNBKkdh
rr4jB+ZEdxiFAeD67xIYsdFGwN6vNdbOuypt9Irft1y+XirDzw1w8IIhXJHgRgdLSLuYi7IZg0eP
cynh1mTaf7CQ72PuVAmH3OLdCq98nWJkdClRckhnZKw3dKV/YnACuR2RcFcIkHJSPZBUO1TJjLO2
6VCZudU7MvRGmvoNOgwbPN4J/h4cOJ8HoUeGKNxL02WsYdoxM2pImts6EqzN3aYIfgb0cwE/aHG7
W+RbyBL/cjYhB5GR3bLuf20Vb38q0ZRXPhrR/n/mwZmsCwiWJOXHJCIr6DZIyDnE1E9AI5EQQb/R
+wIctSYZGgnH9m8xHNMuxbfI52+rh1xWK9yoFpbWxxCuPvlP/y1gxY7srpFqUVckcJcDPwtweaye
fC/w4sIpLlApgOzJuz/gtDhwLLU/trp731i1r1ctqvIYR+qPgQT2owOo6ksShHrfGHJVlo7y6bpC
MTrzC4sWdnVI9Gew8cXDHUj0n0suq6PEP/K1XIhw4pi+8bnahl1yaXv8NfxsGd6UYPQN9t2zXKGr
rECjd1h3rsOeNgCbCVBBvLhYvotOd/UE70h8KhUABOlFaH4i/7V3OigGg3fUtgg6EcGIu4rRX3HD
fGTPOIaJHWsRHT3JAJpJ/uxfqO79RxRrxh/u0S5lTXLsfnKIa9N8M1y0qjYzxIBt12pXL5XdI0jz
xSq5FAKkMNEHjr0KGjefiGRSy1n6JkA7PFVW0Tmzy+5Ag/BOToeysdHJ624YGbWL/PDXUVe7RIHN
DP1p10bKg+S2xg5YSg5EKumK9k58dRv2VlzdaVkoq0cfny857/OIbdAjUxDg6XQpZ4xTBE8yRYwd
YhMgXP7M7wTlZ9/FitiLDB2CFvKBxQ+YZJkAuyZA+n1U//17BaOJxR5y3BjxWJ0tCCThnzH8YfH8
3ShwJK1AmwbIafpYK2q7c22M3j1j/cCS+6bkNO69H0xeosCPViJMVIhXqXu4pexlP/7AyJCorS9U
rLvWRP7KLUIlQXlkE8oV2MbOekZ9j+NOazlEwxY8KjDCPj1Qyk3OSAznrUTNtiY3xM9nyTbV3QZD
kgqHmjt3m9Kt1C9AvGhJ+5BKTBWzFAY676vBAH8lT3t3fmeB0J8pMYaCMB+JNf6oAQWoUFGhnFVf
nclkV7ffdREnJDc9cR2iL9EBLrblssrspd9CSbGvyPvpxkwheNXAce49/QUharS72EIx+s1HD4b3
8F1vp6+zy9/BjI9jyCCLPMSxGPSAUsxUJohYPMwc+NxKCj0xhwzV0arG23tG267orwfehs5Su9jb
n81euVOC08bnm5+CFEGohwkIUQx4xWzATem91AajiIFilrhLnYjkj06m9QxSiC3C4ixW0YFqi6Xr
F8rjYEmdAxMROQ47ONcGNUCFhKFFSAYjKT+FcfeUZpJCfHaDikCf/9Fi0cn7+7n7LSatQKWbbNmK
wAGJJ9jJxat/hqydUAdvVKSjJVHnMsy0tMtwGH2ogo+AeVwogAo+VrgPc6aoMXY2kPSl5MRhqDc4
qoeycasguwXTD0tq3ot/J1gWrkk9Ym6I8IwYlXLpkR3Dr7KIROv2JKG3jAkhnbB+8Wmx/cFiyWkM
Yz1ZrNMtNgDIHvDAEPzfwEoIgrrFo6qWeQTKzprec4LgaEQ0MN2PkpcLMZw5JAKxrqclgaVreWCl
QPT5Pv8NEdoUCkAEjyrGq+b0d6OFdJHv8sOXFe2eqAbCzxB5vcfBxmUwB71cj4s0stPVb0x0niWr
d89aT3QcHIrCZYGDkwubH/dyIIVLQjV7ffRBrb9mWIyGHDnspnP5N+y3vK+R9PB/KBDaYkw87smV
YF1s+whqGfuQlNNgO946q+Uia/LdSn/xl0P69CjE03HfwmLoMiYEeU82Pe+636Qbce5jbg69e6Js
1MdmTnU38b2nn0hIxdE1KYj256tV1Xzf24yJaHXt33jqvTADkik0KAO/4VnrqdHCS2TWT2HVRCuI
nCh9930l+04BJylMU7g48jgL6OU+epQ/0BO2njgpp9px+uHExMR4DC3NAuT+V26ZCZgkOkCoQb9n
nVxyzYhWUjwjcdtTRDVGHZ3zgmOdChmtQUdESptuURloaxKlZ99Kx+Xc+gAW9xHb7T/UiUHc8tfI
dkbxb7R2NhWEN5zEbb+h4ggsUYGzAT1zcbQmu2sIZEM+G2p9//5/X7RYAMFSHXesO7c7VJ00rDlN
ftRNz1hNbI7p4qkY6DkY92aQqTPB2M9uTrUXu8ynWGbcAw+RG+T4SmY/9+paRvhCZA06t+CEU6WU
NsT1bDJJ9IYe59KKVQB/cDnWjn0dOTWkIuNAzLY+BVfaJb/dJG0O+TtxWFAg5ukqrQ/8ePt8OE/A
dcoRYCVmZfHQNx8hpVUsnqrQTEgfBEiItIg+qpU9SZrOuDxAgPM9Havkwr4or09Os4csoO10PHb1
DnpTGz9RXr6xNZhBm0snL/3yfBKKL9ICAoy3Czlb5AOiBJ2/no0M78xIclGoK5mOried7i8GtdFl
w/dgILJ8roNj8R3Oxczlzq2UxTRQeh0x5MKQMWDCIgvMqUzngW9qG5e4H0ThcwS0kTp122ZPflop
NNy1VdV0bLwz8C/f32N6KJOlU9D0BBkD2Y5DMoFWwf5Vn9NweECWmBPEaKgMp7KZku/yn2/EfPVk
LrG20vPfFuTRn0x4HGbg08iGILe66gmvE4/JU5rD0/0G6asa1aYZZWc/aHWYB0RIDj3sKmP+t5yP
ymccmtbtp5Ipc+2vCDHQDt2o2MONhqtmyc/mo4+ueRZlxWy3yuWEN+huQqTWtiYaViVsm+HfpooH
wYoEQY9dhhKYep11f26qzgBBQPlvWm/Vm4EdZxEh9a4bjA63dUR8e5rPRmhGsScTLTVgX7maS88o
aFOBTbkLQSgxRlUCaqZLGOo+ovxnmms/y2cKFXLhrfNL+k3KAH/3OzWYi2xRrET+HO3gJmFy7FCj
kerNM4rJMPvePLy0UiCqI0xj1hSvoPDRAtZMn1uNZ58CBF98yrHSkmgP8p3oHVWZrvGc7LfWkFEz
CpGdR0EzGVvFXf4llBQeVelH4hueDqhF5SQDaNMBJmTA7Mc1ng53CTATpsl5EnYCJFylLbV1VkmN
DMtHVKeY2x21BD39vO6JfL0rg6dO9fPIfOT/ZHKAh0j+XFXTWb6szxkCmHNv3x6jIsRL7k9srr0l
vjo/J1Xw9/5MoLn4D+VvC89v6nwUEZri3Bz0r53WWwIfwpVvRzW87kA1/nQWOW1UlssXthatx4JQ
IhfYRH4t/PnmXl8XeNfa2sr9zRpL+nBmMLVjdDjnQ+ORJ/CjxJ8+ZHOdJ6yr2N6z/lWNiB0Xe+1X
7RD0x8d9a0kPlRw1N31vcHcUGulu6HuodPd/xnGSccgc8R/8SS2qfHJEXQmAnknVV6nVvpgGj+rx
R8VaRtXOU5EPpR278YIDx6/urq09HnvxQI+8PrRhZo8w7GGSnGiSAYlXlWzcwg81RFTKtxAnxIYo
0OTC6TzDjf4XwzWnxMHOjBbuk5LT2+E2tS3jaAw3ac8qL8fRYiWxB7y4trP2bzDSF2CpjjB//xmd
gDfXKIa+XsD+fOugfOrWqhHokVf9IAqJ2q5Fow6l7ciirrf7MiJqDWyWywBr45/jDYO9xpJUp16s
XY3O94GOD/XHZ2/ZjlNLvbPVbpCAAFiaghPDdvZ8DS3PFYWamwFI/cgXsoVRvi30ooow3MqyLguv
26YCteoY6OT1JnurTfbUbGym/T/6Ut41/96yPY0AZTXk5PdvvR5X/Hamliu4UhUWHx0JibiH7dcH
BmsJk9TF54JEiOWI+M9kUx3a7D/JEP26CTRh0A5JcEIDUNUiFurZukKAuH1jvCdlDVL8qH9NcGDo
M+cjngQUjdfHs20Q4Z2jlkKnarrSdRRB4jZ9lQo/qow7/drhLYq7b7RxO5ieE5Qz87zQux/F9isU
kb5xs2lFwMApNtGFu/oHg6QGWgDK2Q6bcY96L9IU4om6yUntXSRrC3M5WdkEhO4BMtSGPjn58Pxj
HQ1bXS70IR2Pi/dD4DTxjYGWFEQUDYL37pZa2S5cOvxMLYKDjvoHI8GyUZ98DojN/ixBRBqKFIyW
W8ogdRa5tAfcwlIp7uUqoDJMHtbRn/1Edd0STuR/f8ITRI8UJLJkOcidc3OoDatjuEK3H0+13NB6
nX7InMyV1f4bvXP59dttF35bMmzYVV4TQ+3GgNfqIVrXIB7fkAhfFtlncJz9CWo22ssHuSHlorIB
a1G6YXWQe4E2suAHWi6ADma3I6OB2k0CkksRL5fyvlzxSg4fLRN6/78+tfmqWY0DgUPSNsVpLCj1
dYIJC6k+uGDrReGwoXE++N06eMIdxaxkfa6RgYAiz80LYPe3nGqxAjjMohJY1DmY2eGwWsXuu9vE
F2jW9pyfz2MvhX3ZH2HcBbLbcRbI5ITNLrZoNbx4f/bfLh7ySbMpG5pOLZwjTUBmI2ePl9km3t1M
W/nWXMCT6en+TrImKg6/3zmqmnSAu2Xv/Gryc/nNYt02ErVBAyICPjcKkcslaSxTw449wN6ZzLs4
/uIB+9PkxYdI7oNr3g+4lHqqrYcHiHq6jvjgzWOzMypQkqP6qrYQpgLCeJT7WO0kbbLpQED28yxj
Pd5W+ILy79aKBUPDtv01r8gaPGsWLgJVvMNPxhExyjzYWyTM/79k0/skOz8Gop8gkWeCj5NfltPT
IXlAcypL9xHlgA32M3c1g5wJqPPgfg14rYxQM5vLjrAI5daQWSvBE/aNHOo+TXg1Lm9cuxug6dKZ
saDKIWwMBJWzODRSOyzX5RhjiH8J7jGfMnAyIcPeS4qGufgNLY5Kfv1/NiK4FAJKN2UEMSBPLliu
s/iDk9sR2UrZBW1jq/jw/sNbQPw7Ex38kZNOd2JwR/1103B7fxtG3XaQ8wgI3MW8q8ID8mo05Xdq
xp01v4QiMQo2pTYNaDFD5mmZ5Y68603YeTOlLp4Ja3/zxVyFRSO2FErc0e4gOVYRxcV8maNxOV3F
/JxyNM+jldOwmrTpYgbvxdB44YvHSXnbC4PrvPcrvwKTIDUJWkoaBKBNyBzEVWQ4nDKpqwczC8Mo
YQaxWbOld8loHXmxN40BBP0Ekk+mA1krFFzVpJ1u54I+ixOcFlPBe1ka2/q6Qs1+5MMwLAQRAOc6
gW80oCbTe5sZG6P+GT5brb3ZdDolbrVZPJ+ykeaO+62uNrN5uLQtHQhAmCfn7gqeyDg8Du6BbPJB
ihd977+cKPe9QTTxMEcakYAmWzyHA9QojmtDx/S2RftFUOaoBRKBOHTV1Nrw1YyX5FQof4qBMHs7
4P/aD/6O6CIduP2e3Crgd6GwYOhLmtI6ULd3PiCGaqamFTBf3vhGIasq+XV4wOvxkS0abZqL3llu
KUQm+aNjQAlq5PaSyo2hkpq008YSQxa1tvlFvm9UZ4XRu8xUjo0MOeU+AQS5E3KWCpvq6SrajUhY
DVaH3mkuOiR8HvvIClqFaxQt5s5WLLVk5phFe1uttVzqduD4QHAzRFup79Uo8BMUZnmj4SjWkCgj
GT/0iFBpbm3TDAdpbCYXX3nsDY6Ef/mNrNS3eJa9XIXChwIyfVedX9puG5BvAANwOHIWq+e7nTAE
OQsQWOwdC/uymov3+m4FYovRxnnTqQQzRa5HJuIKAaOo/LM4Zdvu2tMgIBRSYmw82zd/gchUocQs
hbYMS++I95ajoBMAlsS2Xaxvk2ZjQSW3H6NGmoMmYgevOA07wDdOtzb1feszPR+fnqRMf/oatMnq
O5nWI/4wQFe+c7XofhnbsaVIarqSWly64euKhDr5mDBiae8upOlpsm6V/DS9Txgj5QyiZ/chpl1o
v9/RnURvQMroHqVmC+xkAIaf5bUJAnExqe9pjFs6j6ejft0y0rEjJaYWKPOW6lSDxCNaovv5Lnd7
SIB7PHjKazde+dN4eDMLVSeYjpBAEEvtxejRbw0wIgMhhD6rsnZBFVGoFuHqpcdCYCQhZPG87jBs
0nSvoj2YCyzys/OyGNxiEWv8IeICdCEvUEmQQ+QYbjIfdZ0ganqNccXtLE1mf5BNik/KJ/GE2l6L
qDhA82CMJfGvy830kPmk27W/X/diONIUGWw1HX0mxe+m1gDxdFpfXLJCEWsrQn2bXoZgWnp1JXhx
INDw5vCdh+F3OGVysVsIYZU3ng8HVUq5e4bjSwYz7KT8OiUyO+h3iLDRYxYm9/snF0NIONh39FvK
+QNHrNmK+PucRdIXgi8oTNNqoqPrKpecBgG8fpF3yI2A0dwUCOV+OQhuwvr8yURpGZTehbfZI6e9
JfSsw4ipULLyYwsCn5eARKhmoD6AOtZz5CEqP8mIxS8du0k9OZlyDbheosUtnGRCo1SfxZxpUh6B
CmZmw8XsJNYgBSmWzopiwGmiefM+zdERmrXkJ+eZdeOEovsF+otGOP7kQ6dDb+g5mdZujrc5ycmo
5/IjAS18eWIRGia13q+eBSx1YT35btXKTLnQbMHcsGiU6FcVswWm+UKBv/Nz5j2kd+aM9TS1J1QK
R/ZsfG77T7EuSjXPoUfUZtgAj2vCaSi0FpsGaBteyWM4bbwUYLAPrb12SkWGiWhXHjxnop7oitae
X7YwrjddDthfG/xXx/8JVYzT7Y7OzylLCyHuVpVNzJIwDcLJipL9J4oQynbfx39sxlrOavP5Mhsb
Te8+lBHOHx7Cw8KbZJUHlFA38d78/t1VMomBtWnDVADj4WJCFo76XEGDVfPYIKZzGeEPpMAUarLg
xXKvOa8vY656MydqW3H2293mVvUTd25EOl0aVFOGzwJIuaexKSRxTyhfpNpPh8tIsr2DG08WsKvc
ehmsD1GxXBRD+xF1X5ImSLjR+Z+PLfpVNv/EeqOEGTcXsSOS2IPv/zLYBJFKk48CtD89JFS0mJBA
inA2K4tvFOglJt95gAKHxQO/TNBw9oH5RiiaAqRGMdOFC2TnaM1Aci42uOdzR2FTaVJ3BZAjb0B6
xub7DD7GTPAZ1Jr2XX67+wLIFPc+9RbqVTP+tMohaAK/0YJiEcrL3p1BWNdy9XlE1tKXtOZVk3QM
HF36UqvoHWbf9x7o0XYUzfCK9sVbYC6PYYCgJqdH2ZGwGd7dvmvmC8j/ohj+952Bz9gx8eNdENKk
WPPRkXjLyeawuMc0xMYh+6eYVHPtkyntbO9UFxxwDdVren/y9lgEx/vtL7HwhHH2eoGr11P5D7B0
TmTvHnwR9i0A0Vc8Ooiow0e4piQkoOQpIjZZdRXM6wB6yDFcKEEjnTlX5yLHpwmDRf3EoqdRUiJ2
o0CvZpFXNA3PepBCU0cupfH5eqpOz5v081u6JLHCIHwiuA9y+v1iMzxjxseQ6ztHCFyCjlxdt5pj
7x4g+htClrRM4mqOWVysXGawCPVCMKIiEXMQBoHYVYfYB+kSEO5m7jiUlqsdF2stgNUjoEO3V8n2
pphbbO4y1+wUjJzCdpieO0hRl31AcCHbVX+G3N+sFTzEC/vI+fH9kRTRi010X+bNFstpq+mwjHcs
Law3JNgVjoxxSA5Q8wld2bZmJHgMAJDkH8BuDqoQV4kTnacdqa+whV/c8PhkeBzFciZQz33BA8LY
QZM3ZNx3JMddYpRYSBLKv1ozETmTF58/zkvdmj3BGMnI6ZVBxj6MU1gef5YZa8K7eZySU2qBqZ82
j2uZd5/Mr+IXVqS3U0mA24lBirhq2gWg1jBZUiAM2ZP+yptFYFHkQXUB96puJTAeldOdf3LCJ6da
akPQyI4p+R9DSAfm8MyK3Weqfg8p9eg4ud18/d1byxrOQ5bES6nAVzDgroL5fWzDlM1oXrWhDxLr
fIBdgjKQKIo2tsMkWj7JNRmYAruqbcf+wiz7wN1CV5flGezC6jMOVYewNGk5i1w1vEVJouJRBUCd
CJRDUAy0huMX9erD5lwDIHMhAjkNZwcNbugWn4XhS+HrJIAtVuS9qvAIFU9LKQA5GJewNpnrUA1U
2d2ND8+WdS5D/D4Db41IvfbQSyzKSGIAYCYjPUdvqwMJkKhwt9raqogqG93jxnwX/QFwONYDYznt
bDtVN4yoolnp/OdC1CIGx0DrVb+5LhSCYG1/pAH0C22/tFR3rmhDyMdQqFh+LQXJRGXomqMPYnfj
fsesDK/lygVaukN83zyhLKH30B/pco4nLR5GTCzCZA916NvcGn19xcWK1RJsmuTu0flnj+mdKsJ7
B0VC53uL5QTKw9opHIkqbi+ChnLY8MFuQn1ITO8ox7HfI/X/MqI5nZk4l0TWXdBJUl1EsP7MFhGl
gg2PRW+hXP7Olnba37W133A5Tvm/Z8St9A70Wp9HM3ZYM4mvelwY7swgQKIUml6jmCuVhQhbOVDs
1g2z5HrbQZE93rZHtuZUT4HEZks0yvKM2aV+oqJt256EM1PuD/EJ4kt00Kl579200qyylurMJsVJ
JsiCyDCeodf6JN8HrACZOSc9M2xogBrO7GfjHRcZvt74eVTv43v+Unqop2iKi7OwD9HLH5dNndsO
kLkpVEbxNFmFvT2cMRZ1TzcbST9gg+O9DTW274Btbjl6tFqaoZo3gvzmwbln1smaHZm2SG3o8/aL
jb16Mb0zZ75bgDkYi7FQO5H1xyCfQyyDqMz2L5DaiMLPNESwi/6h50VXaYy/uaguUZOKHLPNhczs
8l7UJ2SUFy6EkCqYtCFB7N3j+9JjMJTMwmL/qM4Cd/Q6VxocN9vDhduaPmFfyWZUfg8AfzeIpeS6
hf0txWmOBHbwm8FEZYXJZpSKcBtRpzWH5ec6cQhW3Qln8pdq0QWCS+2v13BrORQzKNNtk6SL9wDs
W1nIOIAmZ81rMyuuaNpPMuJkYEbDdIylBFmTzZpVqv3gXR50ONwUc+1r77tze9J9kmFRzH3OVZ9M
Ir6AtJdcrnrN7hPqvNONlGdaEcS00q/wQOUJBOPs9on2qBdCs7QNBq8pxjdck+7nqXt4Tf4BAoyT
JRdZnluKJhNQfOLqXG5kOx9m2gsxxDc16AjTfWS71cmNcpOATd4a/OIkBFFUYEHCxRpGiQqzmdQx
6E/qGsPLDE9Wf32Bl5VXPe4smwEiQrqrQwakRVZlwLbIFkLRpRr8eVp41H5Io7r2N7Z8+F0ApP4G
Uyia3i7JLbIefXUhrtfor64Hd5YVikfI7uIpHB5VXYPlNJI+CTh2XDy6YbZdVsvcppLcmiPRabQj
oDCH9huJjmBdXzDPQkD44d3OYAIz03UmcyKbQeDSilUFA86c8DEfjNsEl1QfemZCDamYPD6AxNbm
e8tdVOcn4tTtEy+BnOOchrFWeNItv8asX9Gq92rJW3WeHNWXJK7HuO4G4J071snZBa0z+dKlE4PO
i4JAkMsu5AIFkKgridARBGfoGyWPfeFiP3UQd61wyHixhUIC3DUINNau46Appvoe5JAYWlg9eDEm
XYVcoNjF2Z6MJXJY77lirar9jLxdQpD564MuKoRyX2nn1G4bj+zSqwHOOadsqKs223vCkJP7a2Fa
M3nclsSQmHq7Onpx3onvhBpRYDmHT8yBwH5kUXWUmJqf88HG0+sptbmaY+QOYNMnaxvk6kdnLM4s
ODe5vyRbt8VRpGYXDZtm2khoAeKnM0wv8mYFUObZTpj8UnlARvOBaIQ2QjQ73hwjO1I/admzIXoY
xz7C5ePJJnBqaQNmP8JQUO0r1haIyOYVeXXFdZGKlFsH/7NMTaKhj6ckyNjmLkPCEBGTDBOmRhYn
9ty47JzsPZJ4+5E9RkIefOewxaWzRsX8JccewSGw/WAvKXc9wACJz9Qn70MW4+xsgYbqUvUKGGem
f4v2c8hfL2bwM+p0YRGRSaRGjf+po1MScTzE1CvGErgw/SzFe7ntG5jIsvLkqOJGtmmV245/0CGg
Fa9+Z9CFoA6faXTxN1owR1MqMLfVE2vovCdcPY5m+UHzrQgwQLTaiyjNF6x7Pav059dQKbze3Jit
DZNYZAR9fHXalI+izy4Op0WdplXVwdqhEwdyd9yzBl58v/a/TIVYGzmHTwnBOiBJp89RjY9ppwgN
Dn6n80sG8zEoLKt0mF4Nr1UvN0OHAhKhzUwuA1cpd371NUbFoImke+st9CDydqpFvT2X+zyIxxl1
K3Cts6Og4JSFwRLIOegXvDITT3gTQPMrdRf4MigfxfT+qzpv41yGab0GHY04lPG4p8HSHfJitLDW
m9BtsmYHn30IsJHWko3BoTPk4pSc1cpv3wlkQN7m3RbbCyqgW4A9m4b7NJhvUJ7beO/wuFQx7Laq
jt0N/EeUYzqTJSUGz9Ppf0R80OiiDRp3fNd3UhHEjdATb62ZQseNTJc6P7FYU2HIO7ieq6hPXXGB
pNcKhx2UwEchKugsMyq8ftcD8WZpGajSO5tpqi8MRLdxTNMDoCArRBiZUVch4u5KNlztNJZJv/zW
ngjQTqb5NGQS4JmPl3GszRNAMTMgohfz9rO0rDXmRXPrYMYJ4XNMCQ0foOJ6oplE3aGak9o/3m2Y
6/V8bDy/K3kikBMv1jmPQq5ZKl3VZ0+y05dF0gxOvW/Fm/7Z5Ap0wP29RXhA77zFvPV8jyQnuBm1
YzWjsJkFI+NvgSZbcz049AOhlhdD/AbyEMVicinDwUgR69faUv/8s4FPHPm5pnDcut1BR8JI4SiG
BAaaGGbm6uIjMcvlQWbp8QcW+WLoUyihy4AafuE/7tA7+8cvN2ZujMAH5vlWaeqoxL1VCgUajObg
6vJBDI0pCu5+aPzO1Y/h7KwddXDJj9e40KPkN80o2ViZVDUR7lBieBZR0gxdxxa5RKCpUF6Hta9Z
SbX2BWkTSR3lXGsTTX7VZAoB1Uxj7RmefltIA1wqgKCRDLDdxOS70nYpnq9KeyBrCty7YRwcGEPT
4/C4ONZudOXdHjTVr7WQy1oSsJWFJucp7KO1DjY4EiQ90i6QL/YNzfNgtSjoM5TehbTqj6Ovokeh
wWdqvoCQjFuUZ+nyVy9Byxsx7nP8BusL3Z39sdD9Yg8Xx5hIlb+I2Hf2VPpoVni2Hwt3i6lfqd1y
bL0vbTa8J2zcYO2ZW6lpOKGroPv/VmGMdK0WTjbmUavlf26oHHKyBRjEeu9VUDBdyeK5S6oumNSY
ELPVngy4lZQWgWiNjzPnBtFfpYce+Qu8EiI/ur+aKYk/6agLI5G/ghNd1j50q5jNZcS2ZwZhEUqd
NEkjo3joRKcKCspTHdouqyr8OcltlDDjNP7CYIpz3tQW+T2fSdv2VYdgEDufmJu3i5fmgAMxWew4
dX2X6fdVujzhIyXKzQSQS4mW8EZQZEZuxwQooCBM9uLADVeSbde8cSz5qW+MKOgSZi8V4sxhra/T
SylWCHBrIT+ZcAOQe9661AsSK3qDLDR5Dmf32wQUIcB3EKN3USUTqpnl4XzLQ36frt1bwx1Ig7ys
Y3ngiS+4NsXOaMST26fV7MFc6I5OKkEqbfNiODT4rI2FNAuSjIac3+He00Kxi0BZOR9CdPPenAhi
L4Z8IzHI2wYVuf/w+oLQ2Dgwe4klv8/2F1YJOgEeKo/x9+I9p3MafGoAbLqufh0NRoGwy2Hu/8LT
12J58ouCZ5CuLRrhWNxTz8zBQnFiHST3EsrR/DB15JRFDJRF5qnYoo2It/dupkeZGDKSt9EGzL/o
QsnRgl1RDhFBSWWnpFe9YphygYSYeeBYo2zu68twh6C4wIVjDRlQYzOQVAe3Sdx6Evr+SjgwaNzZ
zDyrJ2aTWhFHyn7gVlSJGOEXDQubYz+q1Ln1OKIsEcmaewtHMi9v/opa/n9WByc8f9fSfiM7Hm/O
Ao8UUl3PDtw53SVNaK+XpLxEuQ7qQhxr8hZDgri7a/O96XPzHNENAk0dt11CqznhYpsDyzTZVSHJ
XkQpD8PjZZwl6vBxzB00kork/5+pW1cosX5f/IAA3j4ptLnfrO8Vm08vxEADXMDNbnj61gE+hzIw
suPmJY1OSI/PD2CCSAwxyDY6zB+hhc62zK/R5bluHlj4k+7MZ9tLS9USdvNT9GrHwc4qqmoVsf7f
FtEP/tzy9NQTCMnIhpT4fjYyCVqjmkvNJ8I6LIqo/qVGZV0P/pyTZs94WGasS2hhWaB6dB8CgGhT
IVWbD0PNT8wiNMvXgmiWWwQaJtM1G2r9TQebx/cedzAHT6N2lnhwKRjPq2FGDJhvM0dpaxpnPXPf
6FQkOPPrUrWoHxXRLK5RdixlJGlHbPDOZ44ny4+cfFFtvz5cMVJ+Azu/6jHd+vuXb/xjfswo8Tqo
EX41yI/KZpiEQtClwrOZ5nKNXoQt2yvDbyWV4DjZZ5nRK1JjcaP4sqfyJWJRwTcjrYDgLP8jZrax
z9nCvrd/q4JNd0b6Qyi8anK8K+cyKJ1Uhsks22G22SG0LtWycbdrmuaFjk5piur/85JKLbiZ0LJw
x+ONeX2atfpAnGB6R4JNFgD2dwAGtOmKrVg1sgsh8ZkLViK65ljERsv157EBkcPtZGNXNMKoOL6G
AUbs49NDqnSTEJ7KF9D32EDzDNi4zSy4LAjqFbhFZnjllC2hCGX/7PmS4hBG29ds2emRsxSW2wob
oK+mkIJ3gDY/ieoDwglp0o1ioE47x7kKtWGNh0YT1a7TMbDHu8Z7gjWAxuQReYXJ937XUegJsE1V
hnzQyGiefex4ODkdHfrCZ6hRChOFiqmkrnjasVjg4mg+/isPN6DDWcGsGGBTmyddtEHFNlcDJRi3
7CSGnt3gpBaxvsQCzxu9AZzOBGdWn43P+IdHZ+aJym7ApSIP2NNTWNoh43VSseIrupxb9bGVBlMD
Iv9leEz5e2/mlIsaxNuzncwPNUBQciOTuInHVTkc5OhX/ou3esEnIMAy/CiKmLbKBPOG/zQtGY7c
ny3LOsJfAzPBt20dPOYtaevMvwt7DeerOwUO1rhRrj38hWvCZFV8i66snk+6xuGLR+rTMfVxCQsA
cxVAXQXhHgDcmUZeQAKpIEWtTr8T367cWr6GvyD7rNLzHZpyY7K9eQ+F1YKh3fSWdIbusgqON4U7
o0Tth7M5tDmB4K6sPFyygO+VnwU/gtPJ1zPrxcKILvfT0ZtK2F7jpMJMjEDzdy6ojewYJkFnMjMJ
0GXQ2V82p85YVaTrzMbtBdfcW2DTiBMAot3H7oOsziVIUdcY9jVMXO5wxU7fFOa3SbZo2qXU1e8o
9PaYFwCWl9L3F1spC+/dxXbc7BonMg/dGX68XfTXpupztxg3Qn9Ml7pW+zN2l2zVR4O4S8dEtd+q
1v2bLFVUlBwdKy8NAlgN5T/Im3rALLEa0dDGc2b+LlICE1BaMXMRci3wc2MxuKSsiqYLfZ/6vPUI
jMqMCqmB5XsX+k2ZuJmDa704LMCn/n2rK3tu909in9eb2C2LYX22Szkq8bm11bLOU5o8cpJUewEm
jvkoAYD8Xi5+2bhy/uFkB2h3j+ltO7eajJlihfxwYyGYBgN9eyc64XZaanoXGgXWdPMKCPaoQBuY
p9D5FTeN9xZ2/UnXnSJWleEpxJAtARMFuSwMgS8LtHR9YTQIyk6O4pxa37WLNVJSwCiBNVQiDQoH
eZDZtNmvSXKg9kGhrNdjQK6TPDjZZeyCzLAEVvkYFKptwRgL+ucNmOxIPKEzuMjb8VcJntdC13/W
Z6ERGR3q6JC6+SvsxMmEYp8cgvNPp0NPW/z1xDMgksP2MbF3jA+ELJyaAWnlfDQfT9YVtGjmf0gM
VyBJfoAOZ+65u9Msi6ewpvdXEMFPlHv/83Nd1sty5M2aNpeRXrMiD5wrMV5t/svvQ0VMnbYg29Vz
zIrUI0SBzPTOlkXRebgotKjh3OPu7KbQPkqOZSdGk8m0bS6yLWB6oqmdACFRzHRttb74P0V/DTG4
gParhsihnh6wFzNHs9Z3jAbdxIjwVdR99R3p6IVtDEg9IgbA6nQbiWBCWVdbcHTsmwH2v7tuOae7
DvtEauDfm5E33sEYGOFFaAcYz9INZprwUo+2NYKtYEq5k4x+P9LGe+QL91A+9c/AnEXY2BHhpRcQ
gJvVfmFZfKK4mmjfpJf7jhh9uMMifPX+7/aPy5M3YtgDAsloMdJ5uqWbbJ7VqwJ4tVWpWosZ0tna
he7MXbW/KEnrdFCnpWRQbLIU1DrxIp1psu4t/4sWlIlolANgqy4RiLryVCRUlOXGMM8KLu3Xu4gM
PGqhIWZkyDox35WC/btGDyI/wSb1od7mcjWWGxV7lvjqiLDTRkdzytLoFOy+MmH0e17TC2J0VCis
im2CXlG3jTvygCGFdzqEtRu/zY4XsoPWLNWzwI+v4dLDk2dQQe9SLVrzWr3QlxpKHO0Dbu1AnOg+
lL9t5Yoa38oKFKfkA/+lF1kqbN82i2zxr1Xt9NHwhqnl8m9VDlPQpMY5FC+0bsPOj8grjVQXx8xc
TBKRqIe0w/j3V0QgWtq4uhXKq1QX3xNxPYRR8VjXo9ideOU/L3s3oqeWjnDH5NEj8YSS2v3MJXkA
1Zl9YkVcTj5QWboNq6TX09cJu4JxQZjL9N7ZL5PINYPTJrYKMhNgen6F7YFFcx1oSDGdFhmNd627
aWCBYTSWG+zq2ozy0973H8Ge/0psHUOt8Z9H2mvc9w/RTpyHss3JLbN1mxfaxPoKgWCIxNhtKm4L
6EMQxrgsONciCrllzYQi1k8mPJFcrIIkoK/fao97y/iRRpvJIXp8rinE8jG4eMsz/fofPiF4xwaz
D50sJHvHj83EiDGeNZe1U/H/D4hwrgin8w3FGK9xswU9GGXbLc7P+r85Lq59Ro+q5fEsvqEWOtuK
A0Pb9KqdC4iXhAJkuVqWQySuLeBK4jtUXnHnf3hGs0FVAFSoxtAfA3BN6kPO4nVZSkp9jk7gDdSM
ESyZQCiMOSP414I23ViA/Q2JkooI1yys5M9iB8AI2KFHLqF8JcC44jYqYZ1bA0dpQkRrfPT+O62q
l1tGkmckXNHVqc2Yo49PVqr3039DsFpFi4II6tq9jZW3N4gKlFV/0aOTkDfCL7d0ZKJLOsPV1bYl
JcmwL8g6MLAFWOriYnkhXdx4GepYS/7vh4I0QQk0FiCBteJfhR6Hdkux6D4czgQ2DNxCoHd7aXzb
H/oDXltrm8zx0quY5lZBntPH0u1kKAmFIak723plgO+ba4+4ttvcpDLwRyPsX1f2j7E+irlXGvPE
NzHzZdYUf3WMb0N6RWKLIhOYOk8bP4RWcPOM+MrXYyVweoP8/syl9nZXpOfJzLRprcKAM2FaGxxZ
H8NgzXXfhUkIr8EDU7EVd4i4v9QFmMRMG9PmN1H6ZtU7chFvrHVA0ttTpFbc+zksLt+K28cOViOc
QAiV9tiM+EpFrO1/UYZT+fgqiU7u7N6ej3FW99/PpwBgWIYLelSvIzW1dxtpESkoo5yEfJNRjV0v
vEQ6czwZe8rDpXWqLqa0IN5Oywwv8tgtLDcGzYvqVcYDUqWc71XmkYuGCHFw9aGpUCOxbOobR4Jm
JuIjBjzAz/2uhBrM4sci1OuWDQjommRu/M468QLPLSHcMQ1tcbqeXASwZwdTtCQGqjfj8UI7EpjW
TV+EqVk0gDj/0gZ/sCqotVOw/A+wog57i3ELLJO47e9x6cwvoazDZYr6AUCaGIIoPfAW6RiwnLrC
nE6CuvRU1KUAEm5IApnwFOkhckDcKNWWlWEJJdXrzGc0LaJhugaCxw3ww+cSMFpng4Tfs/kG3QRp
8t74vgZjLvPJtaRreRu597n6Bz1jIggwOcfNM/oob47A9ddoPN2LMvBdLeveydDC1IdZ/oAsJn3m
3Jq1+PNaUULiwPgMIHb/avDtnqXCIcM6IAbbNUZjdJA5FhFLSLpNMSYe/p3cEnzqJu/ccQLFlHYu
TkLm7E5NbrgaHjfBZ6bVuselpPpkdk/keIBfV3YC2TzN5BAL2vpxC3cWhpeO6A3rPnNycovIxr6z
ox4GzXGB8O7Ua5JCzLLaY9ihzXGyc8QdJgPzOk6ZclDhdEXkTSvYwbg1prmoM1Oi54fjVJ12yFIb
1F1tgtq34+c13RR0FB0nMReU1IGdEAiCTEYqfJjxYAm4p/bJJBeJZ78vmjeXSakd2Xj+S9990wKU
szribaawV9InsoI8OclpZHXuza7Ff0+x/0W0iAEjPMpF6gKLkzAJ3e/hBDcr5Z2Hvg+Ts86S76lW
08XW8XVz1bXJm7kzfg0N/kRjfAQ2eHRCPFLCnAFhDtusVYEsb8vEr6f3SlRnb5RZXRv/MVqWgCoP
558iGuw55z3ZDEAEhGZMwkUfUblSwR236cm79ZtzBJARq9cgUI+eqXXQRLMUUb8FiKTl259Wgt+x
Kx/Gzty17k6Toegw6OvBEJehdhgjhrtpMRzIsrvKxYjJ07UjeljFD439V/d2iLLAA22BaIa/9Acx
gv0S/72eJxTwrVtbLAw7bLs5mLS2+78zHRDTsM0qHvoFApu9yacjaJXRcF03WOzu5a2EuqaA6MjC
lHdNuqiRw4ZZMrPLLZmnf/c7SpTg44vG61xli0t8ADwro4aRB1G8L3zXhSJCMgJGJJY3Y0nYH2JQ
oj3jYpkhtGm6x3GAcPBTU+VDJQOiWcpUFsYoXVxRUrAQ5MAmy/hZtBw0jkWqWGU5zaAJSUapFtr/
t4uZJW/rkJ7TtCs/XKIQwyla+GVNknEannSC2x1k6b/TKGXPRnNkVx8D2IRYR1VxYJajOoi4rj2U
mWmNnKR/RtHqr54QVCLinIZkg/LK4P4u7MxHy4JAUMkK28W7JMkTVxJ56Z2Q/rxZpeHAry9CPF8Q
UzUw5dO14t5WY6SPuTJ0tRMgR4gsNefT6UxKKY5pKXa/aDfHoOm5zUPPSkGKdiIc5YX+Cz68mU02
CDVDNZRHjSfLzucKlcCRlXT+tnKAxx44e4dXWq2np5KiGwb21dF4vUtphqwdycBX5H0nEx0Klf/4
grHdzz5eHwNLAnI2Umw/9XvOYEV4Mj9d92Dza2od3mYxpTBfWNRqKd1K0xL7V1rGppnkVjXIHRGx
CFh+htAO3dq6cME5lzgLoacLTeen8pB8Wgz4YIxVSLrfLFlXXlCTGLiffGhYzdikuKTAM8x/1hyZ
JhCbQVpeGRsNWHnSMud7gehJQNVXP+4o0rUH60xbNMVPiHtlWgubm7mh1kCnsGM2ZuK9QocC1yyz
vx1apBHj+UHV58IWfbkd34Fu49WcYp1oTySOZcUQwbCh4Jk9JNFYl7aGOOOUPXrleXpG6TKu3pTY
DfrQyXmV7KxdSIQbA5uqADU0zK3JTiN7b3mykh3J9oUicwp35wWxlYyiDujZsI5ZTLfpK1Tsqs+k
4yBMBV/XdxRm9Tvu2DgjAxmHR8922YDK3jIz/YCzgfLdnUrNlPy+MProa30tj29Tf6SSSgTugpoU
FeOrFFXK33UATPF9+KmdHlI1AqY7AJZiiRyAY5k1NPa4wF6NCKuOAWXk6P1bStbdt9SzcdCxVjLi
ba7nJIQ8CEUYaD+W6Tqx9NKXUW0Z/YYrbRZVedunoiBsyMxvBS6rypdiaFK2WJ9jL1uWQgAVxVba
77OwnRXmSzB1r3or7NnU7UytSu1xxoF/BfSg4cCnXkru0Mx86Hwo6qi96pqlrlDBg6z8gjkQ7W79
2hsY1oPeu4g0scA4sxs282iL6vpIqL/tgMWhk3WsnrsjZuj0wAJdBUP3p6Q2wI9My2zbKPSvZm+i
/pjI5xyz7cNU62hSLBI7/YS0dFsBwaRqDd69QrbI/VT0IkMkHyLEanQwTNWMMvdZW6yuYAH8QwAZ
sorRzFIhkKqFFGzJYyyTcyumUmsF7wVk0x4Phg9AvqY0deJ4Y6bB/FhA/YbYpRCsdWvGlRpOOvXV
DpYHIPQPjwZhtKDn699aKNKS/pbfYiulb9zLFK+47ouWrZ6UqWhiHO4sLjE9HeP9e5xoAEsEFAPX
yEGzIW5GPEVFsSk9syKYGFoQnIo//EXbn3X4nV6tPN6MNRV90KfY4gXJu0Ybh+bnQfZ8JY7f65Qf
0g7yHTKKmD7ZQp4ovc4U8CiBIjf/auronFIbHle0SZ/rAPjYnhK1QEotd3J9xZ7gyJ5G0R820JKm
O67tzbZnEFzQY8825ktImK1MyI74cX3UcigWLOO37WizSJajyL8LKxg13atNCldsnSYPbZLYPPhu
qPGlz1PeF9iI0ycOWaVcHEkMlVQyUY9hH2H7bQnonMnOLohX+l/hULW//A3sJUrPE/UUbZvNLj2T
5kJAL2Ffo1h2tAAnMb1pxuSa2snlvRYYhACzX2x7J5KZtZIrlC3rveuuIXCl8bKwvdDVneJ6q0UF
ohP6XwRWinBYb2mzShKPm+fPo+HTf59TH4uF/zPuYHebMIcqBVLDVx3JXGo9eHs5neP3QiHfWteZ
0xxJZudiU37M6+dK9ZbB4yMc4vMUba0uFRZvrPHHEmLLG0sANEn+BhsCk/17htljhfLejDwfhC1G
o0Hgxb4vQujIXUdsQ9RVS+BrWm6Ssy3nb+EORu9/YZh0XDeOykyeD3uPBayE5XZbpIWQahi2yUE3
RIIS3gQqCiYYJBm54LpMZ2m6bTVvEOGRaBZXrjlMpSEpOwt7ZkSqBCquQEA8m09mHt5la4TOSwVC
/wbipDBKN9CC55fBFJewwl9Y5Jad0yfvOM9wjpy06f5y8riSwBnx2SA5YI3lUwD7izCZ7G4sIIqG
jqkp0EsfUj3UOgqoNmCWxl5+6VNMDIzpuiH2wmbmtnBzMT3iqMTd1GbuFORA6xzKzmzUoSAlKJ8l
/ZAm68p2fo//U0KoSQA2+P897BcY7YNBgPjpZ3ea2Zh6IAcOx/OCkmxlzBk7/pIF1bDO7JyVephh
Oc4rEegh7VN+rhaXftm5gtywB58TaRLtaRc8sZqoNxGf0Waf3vwEb7BL21Zw6LHGWHNos+kPPSAK
aPtsRySNTyjr+HGJCAkG70phIYyQtYlfLbVsu++4utbcMTsB9TKOOktICldLD0kQEzHAECB+Grr4
Ge2WPd3imcUR5fSeCMooUp96RW0ep/UEUgE2OmY053irdQcwidYLHhQP1ZhjIBIIJMENYO/3UxRP
FwcWLx1mgVS5CBQrjWrhivUZFutl5ubkP455UyQSZAIvdwbD/TuE2zQo8LD+hC4pTv0tpPfRce5b
6Dz32rqpsH2UByy1UIfcv0ULBJ41L5eC9pPHzyKqqlrHh41aa1iT3p6ZjWPzbiKOEmpZrt9+pJTi
MLYTrv/c1ZG5aPbtLPswi2CraaaAXWXvk4xXaHe4bvCIOynO0gt5tEa3Alm6NDIUd7ua6yFFuima
ondkQkSIGUvKPiCp3Y25EACVv2j9UaL2mG+aaIr7OwEQf2qAyGBWBS5zEUxVZxzZL4/hcL4I5JO7
b8k3TM0ZKv4iTU5xYXdioUHbgsqvRk9vBe3DJE/VTQcvQQDT7SIMGtI4w+GEnOcqX7GJDPltoaCC
y2otIO/l3KyM9m8aPus4rZ5pXC3EP9LhkUNGt21eSIpB+WnyFYAwjBQBqEo9pq5wReCVC9rtc+9B
T8cj8lIFQ7r547VTw0z/xL4oB1kuS42tv1UP8HxElNVQAWdEPS0+ro3HB1P+3Awf2bur/o71/Qwd
tYJaavW/gAEMopio/3cCfZblIcTmkcTSl9oWMM1GslxpxvBg3KewXYF1nLB9OgcQvb1zfj8NlF1o
cGFDHyIlkx7B91feGoH2bE+o3IH6dcZEY4XfTr82yhs+zWXJA0i5dlvxOKgUe/FvHw+jATET+YIA
fDPJ2gCkIk9/f8SUiIp3FnV3CJ3Qdnq8hEpY7xLzfyrXM3jDRBz4x9BjCu0JsRS+wbK8rOn7R6t0
AzTH23Hw8dlrhvUQaBxwNsTYAfAXL/TAbQH0geaHnEPQoPlRpqRqgCWuA9zELTEDR4vJg1y70WNE
f2l5/ngTkPiAFb9h3BnTBmKkmv0kAtgI4pun35Wdj7jxbtrOsvHnS6bBcKGhsSvlOJMBaUaQ9mV2
h3a2CyEqwrwv4l864+O3wRKMtfWtH95Tsi7ENArmnnSeIPdfIsVpVsykdQOmIB3BON+7ugh2NTm9
bc8z+l3AiBPeVrvFCwewyczdhE43yGzBNe/w6PTKu+Cb7CFuJ11CyBePv/R+0Votj8zcvJBNANLe
VXnkWHaj5bfVzYFhZqHelvk08d36k6tscKHpC992ebK8v5y4gcJ7Cy5dE/uXEtd+90x9q11jLD0S
tWQowza1QwwQgJp6WlptFWdyCxFsHVUdWLnbGbn7+06Fie6GCcvmtUN1aoDtvwbH61XT8Vs5Ue75
gbvCrn5KnfDHS0EnWcpotYS1Sgv5W8V5YqF45NWguZpw/ngIeCa1IfGa+5mAEhxEADGiLV8082MI
8jI6oWE9aErRkHuwOwnVJkIltDYTF479NjHv88MNcG5WyTiHMwR072ynM/+Z5HXfPx1dIxsd7J5x
cGlEpdgLtfZhrcgreS6HqZxb4GVuI7maVJrg1NgE7uBtlKmaFr0RQsGXRzh3yXAYwF/Ok1RyJc3A
OyPLFMNvpcsMTJhCu8cPTQAZHaJ0xMOrXroG2auF62RvTafvRh/0Q4sdY2k3LtsJlNieFQTEfvi6
TPSaoIVwlDrJwnos2eDAwJJM2O6BfmYKTXviGOkIY5yUO8xPRz82s8ASkZsUSMtveLRlVSOtk+qP
gB7TctsrNfFREXRKiG8EUiX8Mhzi9SCZvKBZbnCHumn2z4jS2c4J+yADrb2QDphcuUnRYFr0FiL7
EQM9jz7DclMX/wQ2Lq6HPfCqwmaTFg3vPAAdMFrECNoWpOEZ/BB4NC3yogWDJH4O7DQVhlCHweBK
dptJ4InS+GmcxFZjffoUk1xAQvG2WI2jryunWAlM72XIHucq/Ico/YNWod7YlsqoD7dsvzb8ZH34
KGRsuJ+B/nZfCZ/A5ZZ9FOcKTyTkJ/VauIIy8keQtGuIL7gguUN7wCuMG2kJSeMZWRujYLyRu2xp
WHbgarvJ1YZ2rcveKa1UZ85w+Ff+E6PTrU8+irxRgtUpra95JFO6kB8jQdUVDNTQ6A77s4kcT0Sv
4K/7NLj9FLHzdNJOTLwVPhW0GrkGxX4Nr0921wi6BbSvLT7OpHzyxqQbLRH20oc0J7TkojbXKrGd
2T2GvH3kai94UmCiEBDuNP+uQxLfW7oC7GAdBC64gzGh29rSecvEtBul0az1S87jPd/OeUWacG0k
40CobV8V20wFdrqSWt//+eLGjf293tqxz/3g2wFJHjW/+AI6ebwINfuXJC4jnzqXsCaY3jkFtsYn
P6LuXMlodHC2cyPlL89RcXevNo1UMIAPG7wApF4X9v1oa4fj3HJpoeSty7yBTLvmBQujF8I63g/m
5cUpFCxfOs6TvQdXrkNeyxcrwR9hoovcN6rmfNAoUKLjalL2OPEQVyaLygf8DupJ2nbaoHfNJzMt
SVvT+FJTgAEPtzri+k65K7YVL2R9EYRjSqlltKdc5zi00rrjOs0iq1QDw77IruPI9DMPaYzwGLsb
wVDXE+c81bZEOgn8siT0RPZz4lsDcOSAzNFGgkPLriB/V4yhmMJhemWK1ciGeScxdYRTnVfWQeRn
puEmditxSuqhnLw8Lf45RndgFuir6DBirJDBXOlu7cmPXU38XQGiHVvKG/xvycFw261eZgl4aY92
QkwTkGpMdZPjdclEcuXTA63EHDrMl9JlCqmrUhpY02BlqKg/TH/UuR64QAeGU1/sQNIYHz+/XuNA
5oMgpYpjnINM83CEB7yiB4ltzfnb0YBVG/Xl5adsMwbgN03UwEb6JhN0n/ev8bzsk6qMwNfi4BIy
ISYHkHeYRrAhKR0y7QvXai4i7CfNIEIMBE1jKUHuDpqILCbX05g9r4O+KWu/0DvHnnxMyqNGxfRt
3IzKEfckjgzkQbtXnDVANOztZCMHJCvixBLpPoIDQPqZlFsA8Ueqg6kM4JYcg14+mcnc4ibUPr8p
4l6DpwEJmgiwj7w9tM6gv+SeL3ORjTNYtCymrPzlvx5tlYhMNLy4R3N4CSQ2nLWYvxrUc448HOw4
l0jB1aoFAROz2HkJoAnyUPolX2br65QNNqQyP973K10WgH5kdP9M4ax6LWLHRb85H0ZmH469hazg
ef5QKmSv49HLpu7DBf8kO915aFdf6JPLiZUU9Q5fXXc2R6Ab2O5i8XEyUVKZIOm5b5QiOzLEQ4/W
bJMAQjuXKRzs6tVYrWM/7c7sZdzHfQwVKBZfZbqnLxHbY/XZKwzZtIRU5gA4IoqgiNNEN8iY0F9M
twr62batsyxKzleC6GoW+0fxc/nCeYNAQiAR8yS/bc0AWRBGIiCk8ngdWwdIZ5ceRDZzIQyM0BlE
M3y2NayVYpjtrLqdt05EiZaLB06K5/2PhPkMjwAn0cPj550k13uNDFoEGPbtxRUuzUnpQU9qWHSO
w5ScqWuqZ3KqS4REC7Zbxe9XGJNs69St88S4upAQ7aVlotXF5KgOZ+B7/jmq2bbJ72LWZHEEuO8m
2JH0OJ1m0ebYnKKJ9cts4lMt3KTYLJ9mMbhDpfCNLjONUTjYfs4H24noXASMVpIbQCtTNNWt+5jG
pGFRJ4li+lLyT/uEOclOlF4xj86TbanpMK2MnRKpVe8TXZfJfmf0WaLbEe2cyflWa6rybhGOWy8s
K1dQNb3A28BYEdKsVZ2VHl7a4dxcScpQmsZ1Tx6yIv4VSjdMNMgdD+b50oyA5Ryq1/q+L2v815x2
JdfMoKyUpFEvY1OQ7XrOqqhApAp+95S6aYBFu0eeiOP1PVFNvJN8XZEuElnQx+zvIpcjdnDy+dKg
svyRR7q2agcexNMN1gKrsHfEC6/J4Eyxo+3cRQoaon4MSTYScHfD3yCg/2BhaCxGjbUR0Ffymp1+
vHIltTS29S89miGubTDWogc26WXnPSTN74i3Q77SboIrn3BYoOYEME65mRpHOyBf79ZLIzzLoN8a
j0yYADtUVfe09ijKD1N+eFI++L8rJIKub4Mp+gRJVAl7t0GvFOcxOPqGyBZKzzohwo96eEgLDrRC
aC40a2JykURZRbIJqLQ80I7+Q/Cq3NEsg421ODtAmN/LP/HsFUy++B5F7zfFQiIiHf/yH86dg04l
ZXvzJxWwpvvoWfGLWvYh5FALvgC10eC/RdM7HE5tjHjbMUVzXMIAclEzGv2zFF0MmqFfgTbYAd4x
5xtsXt0Rt8tDjJbu3E7mfxDTTaamEOhqe9pTBnIyf+lp9ORAo7C4o/EGJn+Tbm6ZDqSjrNXI41AX
OUyNgeq0ZRkwGfbxfFUGIbPUND2FgQdR9JCuOe6kI5N7LSayIIdYvbzdC9TTZs0G73NT62Rud0E6
4DTBMw8lZLHN+glso8QkPIE50Jb4E6BsRhsUBVqAAZym9Ojwq3qe24lrYNQ/kQaw8yBeCFqZ/d6L
LTQALfvWCqmaDjt6v2ovLwr3RtNPhT+CQCN9ZlVu+mciTEgaCI/PhdYOCq8EukUEACOhZcKsaQiv
MeoujYLx1+9do3h4cRWre5fCMtQ3kFO4aDHvppGaIbbg8Ka1KWXsGomYxm28NAsZR+Y6xR/PGQDM
53I85MsOVuVm+Zzz9xPICib/vNF3YuAOD4KGf1tUEoPEd2Iw09YG6s4brGmACzB33a4CAivjjzYo
LWpPrNhuV68gIX2UfRww8krfDFR7HaNP7GKlIIdQ25Y2wT1GcIc9UgZdVnvjHD1Ze1FBhQaBmZmV
/Lfh5j5+3NtO7L6nXKCTbocXe+a22RenFIUJ6ZWMCDaI+6/txlXy6J1P0w2U4wsCZSpOyIMKjO1z
+0/hF/Q0p68XGN2iBhNIuP8UG0zwkg+pUyQD5xjyhZwLD/O/mB9+tp2g5VuWNm76tg2m7h9hKYUP
kvkJDxx3XMzv/Qkurz6dfD1MwC769Gc4BEsiDx5Fwegmz8s3Ui5zci4phE5jVhK+mjGGVu5UDUm8
YTkc/q7ahEGwSjkchTKdO7GGg5eac1H6csCAzlIHUicOY0oqi0LRLEkGKqFOLMWZ0pOmxm0jncVv
t2b66S8y7rDNsPcsTVAaslkRyJrs83oJq2ywDBH4JkRG7iCwlsduR927ud1qSwWqO6QjBZHb4btD
IKiH6CxBeFIFe/nws3L/5JW7M1StfhdRcTWpSx50LcFHv/0t2ZOKxNsCiJp78A5RcwYrdE3lJ/aE
toEooVo1xOERyuvYyhGEzqFXtd3g+johMjLWna33utxfdLkxfZkG5XvJNIa6YXAJjweuMcsZdLw/
YNW2E4UYgQ9DwUQ5HrQWCvmf9vLp2KjZkAXgh0GBsn4R5z8/QQ6tl7939ZuMhNyByrrFyMAQGrni
PLsCprubd0xv4hTzYYxZKqE+gDVvTBcQnaHVzky2gMaRrb52FqS4TlJhg2m9Pah/nfSukx1tBq15
tHDHQTEq4Nq+v39rHMe8CJvhBNi+KffV7vXecT54SWKDwBJ3Kn4iNi1tPgQDEmxzoEO9maatKSMw
SuiNk9lzhosoM1FR3V601CrX3vN6vo7AiWq9BWIBaSnboV0ojzn9zh0kAcWhQYHRYqQUK4rkK1wD
yB22PjbwhrTAcqDUCjVTKFxL1K/u/2YzluA6JcAQA4PI1ZyABVUoT8uf7KCTdr5zwdBoHEpu17hK
DLsTPahdviErHP9PCz+h6EeHvrt9mdjWkEcgJqdzEuj8zys5S3/waBMjazg9gKHQZxyszzdLEmJB
K9vzuGs1k5yYRtxT7bgC8HXMVAsr3Nplp6oiA/jsWuXLNlbN3Izk/iu3fwYNGGTRlvv0aL0BugEv
gSWHp0IcBe3d4NmF5nZkzzdnwcieIp7l9Z0goIdSSjE/QwNIwXn79rxBG6wZE/bxjKf3n0BQcOHm
8+awOpPL7MYa3XCSfaRLR+g/r2WeWtB8nRVKw7EpNnIHeDRKQ/sfV/LOxvC2R4hTm9uAxhyPpqrS
m9EjDwDeeDAaUGcidetHwMiprJluzZVud+vgQ5RepuTZr48EvyBi29dK7YTouo94bfUbCnwIwvXf
vQoftri3CYhNhbTxVjU0Sn8h6VJNpiH/9bUAJCThTuwTnA7Jg8c7X9Mj4W7TClRQkvT1oVQMcLRx
06iPuayQQ048d0GGdrr1TX7B/FpQs9aHesh+nG4Z/hW5oMdLTdv/wV2ZuVdzO2su16BZPlFnDqqQ
6CFrPzIGHMfQf/fkEM9rIrUT3X57f8xZEC84mbAKuyZQRUTHkuQIERMthJxhVsPXHbB3b60/SAxd
B1J7RAXNxrx5XzmyNWvDXOdVnH3aB+QRkrbtmiou9J/hGz4JXSqBTpVvgxcTArQop14y56oQGuWR
w5gYS4SFe9bQdzDWHDKFieQTw1Ldgs/hheMZ1FqOJSqa/N0ZOADgAiNzozUseegeFcDqQ/OikwL8
Ali7+nGRJMMAZRfQSHIJPb88xX+P8R/QTCkrcFf48LxTSqC/jcFDPPfY3tm+vTTtkPk969RNmA7V
1wcoBm6NvKAabHBQcxs/jocS0ScCRGMarU8GAdtC75OrupquYX+VKyZYRbyfFq0lMxWbRabSSwLe
b1gzhKz5XhJO0jJJX2OVwq/86jkVzrcpDGn0aiKxhloqXmPFJF2FjyMUk4L5gTY1VV/31nQ6Qw4c
uSo41Z67mJwocyll1HTPatvqAKwJXrX7OO4vOyetF1QbAhJFXsNadKL3+0LU/stuIhvfcRgEwtNw
/bt8X0tTOKrcFueMMh7J35AFnG/T2MHzsBgvKkX05S5JV9WSjtgWGhbDCbqUIHggVbt6sbJaM9MO
aqCFtjsyYhHR4pWW+kK49X271XdM/6WAkLI5QDGeY+MsFwCpWKyElj/2l7CBnqfFSU71mkVI6bvA
ku+vaZaZPklWLyiGwcLD7iYEjucw+Jo8gQGJJagV7FfWONF1/FBRwYnYe1AmAlhh8266fFXzHsMT
kbQ9oK71GEqo7jBA4YpVWQLUeCfVhcnBMFwlhzbQ/+Xp6I3XYa0FhKhYOGzisFcip+vhA49OKZIH
ExhAYDu0mSmV/BhoSTQernlZ/koq+tf7GU8kXARcp+p+ycPwymu+VFJnR/F77UIxnPuTKjHHWHWx
7F6AGQm15+hcRrXpilPywVSoTmdR9tIeInm57B/luAw1w1GrmO1QpPz24Gvo+iGkW36RYyknkYng
jxFY8bBS1nBsKy983XE7VhVcN6BYktYr3+ofPkaOZg3l81xagn0QdXRf6gCJrtjGPvQDpRJu9QZ5
SS3GOfP+uPkPYZn0hUqdtrRMUg2suK2yOLzjKmzuKbdPqngvyW6Nw9gQ5QdDTQTHQx9hg6WSX28e
jWQwPIPVGUXcRZwUI8GCj4KcGeV711SUXcrSOMxhhot8P34LtrYKr1vLH2MDPUV0ChWsYp/RqH8T
EvtouJP6bIfvr87a7WKG0HgvFMPBru5U2lba8WR6xVmq/l7REgXyxWN9tHy5aZUdPe/YwdildsUz
0VHIKaOpa2IQALDpvJbNTXIIeX3Hldefx4av5QPJwJceAC+JBJKV7CUlp7huK/hcwnKbNVy5e9Zj
yqLeYD4vZ5mGMk8QG++Dz2UG8nzSUHVhxtgxT184Tst5eNTLFa/fAAjKdHN21Txcu9I8AEZfj+Vg
1/s4eD71/NWtE/88hGpqGMcvK9ShaN8StkHTOXjwli/VLBBAkFouO8puz25RnPEurPOtZYo9ChGc
T9Hk8i8fsiUMu2+XSPur+QTeLqdip75EiWO4qntJRSBAARDkbCOffLOvfZjEboQp29kk1/9Ny9OW
rd/D6boX26ZS1XiuyBPtebLmfWYasTgMQ8xb8PHTlrBccv2myUGp8+PjlaQfyor9w8wjtYQv45tk
IoaNXHb5/hQ0v/XaSI+qksZpw/OFv9ewDcnqKmrTsIUryS66kjEGYZIxqmFfNOArakbBlfRvVq8c
F+sW44pyehTrkgMA41f7+FjJ4eASRe7X0nyFN5CcxdoJkVf5TmvZbTeQ2f/rB3aQ95zl4/+jJ6u1
b/WHRkDudHvWXPKrKunZQVHDOLETRzqvItJ05EMAXqe7fBLo5+RhoDgy2dth/f9QLBSnd8G/OuhW
aY+YLr/46bzfeQ8mvgdoEF4IW00d2eCsEnj3PDSrzjvCnZY/MSbRS0wJLm5NPnVunqt5g9k80D9S
GvIHDyE/vVXX4/OEPyUOgaYgIFSvIaRUY4XHojMjgrW9mgG61JKBK61altdCgnWJVD0kGTRNqi6N
7cGSwhKq/ssiPRutp64SX/I0gI6TVSFIn0MFmECInNXhDJBDxHMUe00PAlE5XrWQhsUv2OIEHvIS
te9+s9Gtbc7dJjVSUwvaOLvhl7v/UKoRbzfzgDtLdwnBW+qS/mfEDKMrEh+lKCcmeuTmwuy8bqR7
tw6xy9xoXSfZB1Z8XO4OwVJa0tA3FJx9oKk9zH4/ofbHtnTLWRrA8lj6ynWKmIEvcTikiiz5ugZm
ojUtWNFUA/t4TRsfQtQA9XeIbi9spZgJ3UZwmHWz8MxES4eKtcLWzBB2YEdpws+nn7aUUunbq4jc
S/4n4vgikZgOYMH4GGqUkrfzFAvfXP7WJ/JCLnlxXj2EFJLcyqArgm6217d/DKt4TNxQJW+pz8RF
0jqNa5Wwhb9DWLrPdENQ1e7HVIodMSaz+/GsmqOfiI616B/JEwhxpq8WDklr7kT1CKM7clfgl7tI
2zfoGy7d590ZaqterJOvJvIqw0E2rObQxAuoFbGcEn5RdfmVpKeRUWgSJxz5FpiDcMYQpjgDKiB+
y7aO5YFUiKpn64ZrQlMx4RfwLEoPwWWTGMVnBl2qaPH+NbWgGdHlE0HNSSnKWii33QzwKYlMErhM
17SZYWV7bqUpdOFpTdohEIi5lg7dqOmVdnaku45ybtcK0J0QqkEvdZSRCPFTZQ9tvqUE74aBwiDI
kN/k4E5/B9FUNIPlw+D4BhCUDuCFBj0NaaVPs3SaGI/XeS7wtB+vjyT9ytHkI+Dse+zPUhFwQsMk
P8LBu5PGyiSo0DMA+FjBIo4GcWbTs9w9gVAwuoAEdw/ahdZAbldSlfb4lRDU/BfaxnjNwcgreJ3h
o06dnao9NbUnfL9Fc0vfnigJPF5WT9dXQyj60Y5kkh+edxTYj3uU+G9qiH4sNVm0WhEGUC25zZqO
qRnVybcMVAeRb+4pXwAMscQaB+27+ma44Z4SIEnt1sXmnLBHA+voU0wfiEQQvn9X+nB9BrpmhVFb
UumrK3x6PBfg+2U+6jb+MSFpmzlY1ln4nvbgI51bYpH2WkBkc/gj0hyY3K70M6avTZg7tnli2xvt
c4p2umOazjXkScfCanFZ6B8rHeUy8l0K7bohpunRW0AGWGtDGRMFxNEmBMbgdsZ5kKXhtmwPjUm9
nQ77azOdMmVUiAG4X196odhBGs02li1EeJuQ/gn7yhPufY3wOknCHwjOuR9IMY/S3edmeStJ+fuM
Q3OG5h1+WfnnFPpxxFa4+ErAU7jy+Eyo6Ht44tqSdfQ3iaNzHvsoyP3Yl4yOPy6TX2+IRB2b8BmU
+liXXtG533oSKbYdyTEVGuKiCWNXftLMiTbG4nW2lnKv9j/dVaScAURLZkJW7AAE2oLJqPmjaM9e
mjRtco3jtkfTNHsmQiZuezogB5FbjZOHgHVK0j9dJfowF2vmumu68hR7l81jMVvkACFvVV9EUruw
qQ8miLuR0tZe7sUTe67hlkFBIsMU0hN/NeA49fLMGWiiyShkCmEi6q2UXRaCKOgHRUBxxa6DlQ5i
8JwOlIMwh4G3uJsqb1Z18EqZeHept2tD6H+yhGqNL0StHhwkKbSAy8Joon96PUzYVyZlNWjiW1pz
02pqvdUrZjx/ATd5N3yfMJn7P+DoMsRDv1nJfYj2cDC2FSsKYlAxvREuqQZNEe5WtEgZq6jC0m+N
BhLLzIT3VOKfjbr9E78oB51uTBHuR+h85vRtJqKrinpaWQ0jogjfekqG4IJd1fa9WUCuaMrRjl8t
Suh35YKCWQ1lFiNtEuZ+w3zs/M0Qh4V3Qbq/BKgZO27Zsz2cuFZ+Gf1gR1bBeyXE8InECpCR4plN
DYTVvSMtT0besfHLZgzaQPOb4h1QhJsZfqCtndtb+r05zQWc8kvQAmGSpAeP3zhk5vp03cqiUZ7Q
N7kiKj90j78g9oJPVVayPuDRBTH2qSXETA4HVMKCg2+iMY4JuVg1VvfdAUn+4HEW9562xE1HKyaW
nQdK6rTI5xmJe2tTN7pza7tujdM8jiyjaGRcPzBCpxh9BgJCYJM4VYy4Ft+Tn1b0jMvsDg3SDVb7
Xny5yyJrHAXszWxOSskux0BFLp5BRp0PHc86tLjuJ/pISPbh/fe/pRkLxkKwD7g2ddjL+uouYjPi
4cEXXgC1qVhDrEU3wwqS6zCJG7gYndxNG2Re42Cj5q+mqpwGUi/rlOlmQCDih73TK9S46J9656Rz
hhcrEnjLolaJTSsX/NDrSnAevDuVNZsBp1Nc0Ifv7LfPqLaD6k6IsQpLuVkV0v9BP2np5xvNK80t
I9Pq0lEW45u8OHwlaK74mbMu3bUZs0KV63wCDDodgCxcs2UAQQbBYbb3cy1IymLyRjDHfYQ8+fpP
F+jjaepVrEYjI8vLcZA0etNe6g7jAF47uUvT3lPZuJC2ejEAoOCn1v+PZoFUjnDE7lG7ht0kBKNO
QtF4qWCr0bWYzDAtb+4QjS+wibJiBQcjGXqznwQynvfdYXnfEUMbOXz9z4GYOck2W3IOz4tgY/Yp
bIHMtRk5GSD099DF1Zfy4nx4QIgGR9TlMvJZLRIn0xjzmkDk++XC1xuzCzEYi5W2vD8RehB7tFWE
KIiy4JEu+aADVT3uwJnE2qg1qHgfDdAk63qLLtAIgmWV2uSB6tSVdUjoR8xvzOK7VGHI/UcArKaF
E7zxH/O70ffgXIZz9AzSR9aiM5oWRBi9Dtau6Oed/LBN4jMhz6rSgRMcw93n9x4HW7ZD/WfyEQII
b0I8PQuILtxS5+gLtlxv6dGo125jdbn/9LHYQGKk+RNUS/Y56aqp1Ys3Xg0t+YkXBJXWnl0jD58/
IRCgn21bNeE9JzWM5Jym9KTeiQ5FBCK2CTSSn89tpdTRuIwcH3mFjBEb9ETIWybNO3WYQv79GpcA
DPUtf9zAoe1XWal9CQkZKVm97yjYm1nJ7hAmrtkMN1cPt7VVtVu130NzFksWfT/sgAnqFS29kX2y
AIp2miSlJxSNM8aMzLw+/h4T+paLewofq7KtBv82bA3342r2SIHVuTqXwf3WJvFk5ovMc4I0zwWc
Qbl+CYKrEw2AgGY2uVfHTuNdHnnehQCRUCwi0owMNhWnUW3rNbgu/ccZycwN305GK02V5WFX9on4
oYYRgsFXgHyVpoAbsdG3eQAbvfoJJBtgPeSe4WUZOaGErdOWtiW+VzyJwl+aSX9+S0RNiSGjBUQw
C6if5WdnIhsGGqpRV5CEcX0PFFj+o4owVZG6QqhJM3+8nw4OpTdlePsTAU/Z25bi16WsQJ/niFnZ
GSLAG0JGMXQGwv4fuyz2+9MwZCXu0IU2UiZ164Zbdv2jceOfOz+8c6v5+FHUeovGFpPoeI+EB5Jt
AKvS03dtmZe9gGTFfEpY2D6A8gMabTvPmdc4D40XyPgrrAmDn308L8RZTAk2ODEV/Pl/TU+1hu1X
ZEoXbgL6Dmbu+eoYH35EHtnTnOc9O2GMwnvgU/mt8pMndn9FixmM9LlJR4ewwlUfgHpfwwYPudYi
jJGlTKXYKSbUspwBoeBNw+nQ7rZwSgvA7kNsrFlPW0GWpSBr2McazVsvr0I77/G09Na3Es2KM7kZ
/jR78a7bvLKQQADdz5mrs4PHMrhPWeVx1bOcp8h6Mga3PTd14cM9swHubCwqvjGdiDrKaQR7HGqH
A8bhMggCCbppVgygl7/7Vv0bGdzrl9a8qeSAlLZoq0oeYPMD0nmgzQbNjQ+657fntDzRqak5mV0i
Zab7n0587ZV2w4UtX3ks/VF1qlSwrhG3sXCWqDrTyhFdfU/w8BpmiWuW0UIJPCny+6rEjScDp8UE
yBGXjZ71vu9bKedkN0ys469jTtCQrYLEK/O0yLelO2hEUQPu4jwWhD3BPipwUTyxhk5qL769k4Vm
AXLWqskNFQNUZ2ZKZLzWhRJxeYK4QqJfh+/sRP1gczsIIg8gx5zshe9Nbwx2mV8cKb5qkTeE+Aix
hU4nviifxwChyIGetCl2g9DPpv2JqkjJNM/nef8qn+8qFKZfa88KbJz3bvq2akIfxNYKcGtUIZYm
cSJJE+q+KJnIKx/lZaAwIjrtdEA3encCp7hNkmWltWFKb8CphnarnfOCc2JdYPPETK9EfBG5KzhI
Rh2rTcsI37pNv/yJPU1AbmDrB1ijgbyHXEEx70P5owHuWrJOSOpqRS6oPearKbtZ/DWNMMClB/yz
MAR2qR0Xgmul/Tbk3TwcR2mJNPhYyN4R1VXK9V1ezo5pL7+a2FuQ/ymg45b/HiquxkiAumzK8x+/
I4RDj6wjB6jyrOgCrKKR25gRH50/mhCUmj1DBi3k/tmyHIqO2mVnXpabeihmEm7M7OL1c3oZptKD
BOaDMtm57oY5i7f+BZwLqUP5jBtJU2pH/o00Q5/WfRC1xo08CnTfaaci94/h0ojfyAQCmAxxnBj5
//bnBjbgmcvFMr8dCfNW53/gpYFKYsFKw9xO6mtzauFIPlfe12JCuHRlcw8C9wnWOWEIq4Dahisu
k8IGU9Nk3KXBIO1lxGyZaq9E2yWSzAjcGoQvUq3PqIf4vQDv1cCwmzBEy5h8+5ESL9HyLOvZzoVi
CmkiXkv3mdOseFFnTMm/Qn8tXrtLyq0M0va6nycBOSQQEDcX6PjDRzFQOP6Sl38qNvQ4FuO3DOyK
ieiCdJ1a8ErBoE8O3xE5LG7pBt57F+j99UCCT63Ex3Q6brbFVqj52xOeetpDgqVjYFojDR2uQBEW
OkSEaWbrb0WuqtKZJL5dnCkJephtiaZUV7es+LSURBSjcIM0TkOeaRPF8jgJvBsvXc7ZA5hJPDH4
clgK4PimsfG8h80SNK6pBJ8Nd12qhjJOIhzTAE2cCdFG5X7UaGrjx/88+8fK8W51r/0wbEGRy067
yg9sj7qk4AYXljH83MtTRO/uUVret/Nc+NScDXeiudeKCuq5l0ngE5KOP1Ge0dv6Kdv1pyuOW0Ne
2XVyguOSKc+miSuN7qJuMAoNoUqI13948yeNVSw6Q2CAm6dJLLcyOEIws7VkELGVhAcZtQi2P7+P
NHrWSzqyBkfIh79h4iyX8Ba2a80otSd7415rjB3pu4QKn//nZSLAodv8G6YH7RY9VKkpD9IGMmbn
QvuPtyfq7lIerPGOQC6UKR1jvVhv8RGwkcxdhIz2vXdexjo2UpzvmPGZQjVZq9f2MbLRh5780AoB
cW+fDaD2c64H12dG6d6WOgQUGJJHCRDbqKRzE+IL48W1UmvIPnosKNSuDv/xbIv9LTjQXhmNcJAc
C/3w8D2IGzPBGQtzFCC+R70JuVr+HfL4O+PrNv9g6u4068e1HgBoaVBr2CoIsDY7U9/5IquLP+7E
nAp1YhXmHM9FWCNJHfdnDWGe3hQps5nP6bHxmCuSa9g8APX9SyipI+giDstQIyAcH58F+zfFgDbd
R1IrH0DVLj9YkuNMbJpVtT8SaPvh0nxrnJBvZG6Ut3cb/+jVWnlEx0l5j/ohEp2VqKoDraXWngkF
sGvqWM/VX7NiP/K78rdakakAgyd5ssFDaUWnPNUUsL7QGEuKOJpJa3rQ3Zm7p4SARyOOyRAps4CQ
+YdTb9aL/uoAGiCrbVesL33eMbt7Emgx1Agbs2Z7TLJ+zmj2sjcWOBHW5gv0HjypCzznJ3CrK40w
yxDrOPR9Dvj+KQw2rIxmJP5fkGypL7BhnKauL53igm1N5RZA6ax44CiF53taV5JAmgivIqhLuOcP
ccmt/3t8Xd+dfxI9c6omlQaL7CrtQ2wL7DI7W0SOY3mV1nng2eKjGp5OlqmF84eegQrlhq9jEpU3
O+UxAGVuDqsC/B2v/A7MOCCrHPvRKRjjPIgEYi9tZZRs0h+ChR85TgwfLsGx7ckFG7PsOlVcHGsv
NU31ZSZWj83No3wMrnR1UNaIFKtcrwhf4FO4PsH67IMJT1H8XgEQAFBR8NiiO4yaDDuffpP4pT17
kegT5N6jV9brkG12ZNk2HD1RZNboBFLed0jLludUR0k9/50+9spkcuSajglQpQcRdAfCJVTK0alh
griEyWsE3S2b3oPfSXUnUSjgdfs/vtIX0klbB6Ugbt1QpaOEstu6LvrhHF0WXWGXS7qJ0ZcKW7Dr
ZqJANcV96iqaLwNz6lNBKjMoTl2CNfuVD8/SdKLQ0PIkHawahBs4oC10KPMLowuuWYg4nu9Z1SUg
Mw8pxUN77bgOOKT/aiQ2K4mhcm2NFuwLr+NYrL2fCgR1/Ckpot2A+0rmBDXUMfhartadolFwgRAI
OW8A/G0ieRKbfKfnmrCgVSrxTZoLC+fwWYmyh6kvLv0XDmVcZOvEsK764K+wNZNvqtN6bVrBZgji
2d/xyGe5HVb8uH7Q7jFPxa2Y/k2LkBhy/bodGOIRe9Ek4vtyF655KrmeqdHK0YtGfFtIrd1Xbnga
8SgXvobDjcWoquEnx922Dq+rqBu0Ay90Wc8jT4+xQDgWgKtYm/Nckz4yyH3R5nOkQuzzCTkZEWen
oAZfqfxC3c5irKeXxfhGI5KB0szdqLpixwX1Lgt+2io1hzupzZrFUbQw3/X6QCxflkO2xowuVbVA
pS8StuIAh8ZHqBosKGC9otg6ZZvEgPt17hz7SOMb5eAaBHXTjS4mfMxlKDwKylUR+V+q54JMhbTK
/FY4XAMuHGpYVFvziaiCYFuRaIwerWzKtGwrJcpsTvE9xGLaOE5DNYCxlimlza/RsX+5x979yMPi
ODH+bWVaBG2qh+p/qmoDQlC+KMSsrKwhf8HSgTCeUK4jbOVRebIpbk28G81VQ/BDmLN3FZMTLCAW
ZAfDUto4sv0yzu2XxaAJTUbdI1+O1jXWxau5B0F5Y7+FHFWF+VH/1t9ZPb8+w3sUni6xPZggdkru
UEchjFBjj+m7qW/NP2mOiPMZ8d4oOpsydBFPR313uNdvZMld9iJegHU74YbOFxaVr611jybFz/j2
P3qpd7dS2eTald2DFWRuqRRw5ZufmN00Uqtg2p3Wt/TTYdgSAPwoHKEloYyt6nKaXXF/aefFGzO2
Kv5LLjJf474TqiouMj8UMap4nzRYsEFJ03Qpd147NuprEdf1W4RgDCqRYQcZ4Ss0JlXuoiph5ef1
JluDcLhg3cTm52ZlsGlGOXycvMYT4WTJ5XJYAYRocZhD5gtl+o4Y5xdRlcvP9c9AvPuhaKcKvOaK
nXxAW17sFAJztQbM7pljnoBtR6X6vEdo1qe9cirs7A0Eit+hvSJk0vmzuuR/9NmtzWX5xp7OWpj1
vzy1bCa/OPaKtuvBMMxrEoYnS1/wgc3KnXIJsAsY6SnRKOtme1zwcttpCmW4uYw9pBorMlqxTbJM
mrYMVF/prUuPzLz1npF0Lurie1vtgWn6WeLmb+SpdA9GVDTx083tkE9lk7jtopsV9ydzg7JQ+87q
k4dYZKmIENo1IZr7N1deDfpQmBY99jCBiF1YVl+zuwu0HdXFAoB4HsFyRG0+z3Vt3lrwDAyUcrit
R2ZDSLxooWaEr5lYE1MZyraq1KWUtJ3Ekx9D393kWZNnhjwkmuydjKJqFF6dqe3T0VqMs94bFacU
CJdJIiNaf5ZPBY89p2gZ/DeS7MZ2WHBRLsabZWEBvcflhUMNTj/8XeCHg05ttaS3LQLmhqAAUDym
W55lBUAR+KfP/cgvRaD2hFgATZgntu95bQBESpS+WR/xcaa1pXYc5tTMFa8ZUrh/68cDHKodEVzA
xbyBSbmEt/gMnmioIqqPn3ccZvfhEItaeMPB3v5mjD6mL3JlZMcU88RnX6hB3BO6c5+ib1jacLbH
A+abHh0z6ejtRXaXeZoX8qsynJT+GOp3YewKM89G6ZlRZzXDlgfpiKVIpxV5pugZob1JChV05tQi
hMR93mMLM6ZQc8uorrouK9/HIdidxbgp8dfqhyTUJRpt0VFwacIwzTkgkg6GFdTwqgaAp+W3J9zG
7SeQWA9g9EhNdo2gh/Hb0+IW88JNzh1ba0t09BAFKiXxFAqYRybN13YJKoZatvZ4nNSVAhd6Xi9e
q7WnTinpCVAcIQstLj7q5R3TzXNDJuRPuQ4qhZMpYbUGTu3ysyjM4s13ReYrO7lmJScmstjEL3l2
LhbKd9lPIpoHiSQXRIUaSa2drOzT5Z2PdsXxwp85SHarMV48FI3Sfhe24GU8llnQUK+evbtrsk2f
J1OHxVj5Qt2PORGaoYPvz99EEdPhQgaagXEP/OtiaTaCgSW+isK3UFrjJBawnDhGy929Bh9Wonld
kYkfumiF+kn5ynWXtNPB+bLLGl5QHoMyEMUWblGDWGX+bvLtwjX455t3XyiX4UNCpWxNmEeGhqXL
Q/pD/Txi39DflfNYv7cF7Nd3GK7lPKeBU+elGpuxEP43ce2R40RIGZartHxin/gXa3v7j6xA1lrF
JpBgBKup5N/3MfoPCCLOOTPAQIk6XNw7MkIo6HjVi0XSMv5U7fvVeor+wI4qZMXFq29NwsloXgTI
dUb6mjvzUelG8hf8MbCtXxRVHvZrQx8G9VpeQ6cADwGDq18SOaI/5ogX76VemTbzgF1akl8dCgaM
+hjqAHm9XHMYY68aNGBLUS3DWboQDhqFRjkS8Mj2mcjaAmpkmXtw7wdCUzzhtN+lIm61RV4H9vvg
SaAza3ygQufZpnKjxNbg7eE/lAGvzGsCE9XQz7kuczvtuTcddb3cO1femq2Wy/mtp2eZVzVyuNsZ
7P+JD0VUanSCawUF5g1XA0lR/AcXOKDJESHH3+THaK5eYFhxMwHuDh6DjKMIarhpRkCr0CufXz8b
Kg7JeQ/XxZCdJVVyd4yvcRSmDskzPWpfZYDji4SA6WaDHSza0OCksMTfco7ZCa3SulqkCrJ5yQcW
XNeM6MMvwrhK7xcFpPbX2MwaNNuoCcJ289Kpo6Zv8TIiygEBhnXRNNawn/gTMTGqjyu1qi7dggjc
z6lTLp//Z4+PMPrJQmeDHzLQIFkJqxWyWQf6/AqRiAOG+nuBx+n424L4WwWRny5nQekR9GNym541
K3UCi8B1pryBrLTLTn0DxsgyeRqfpk+sfMfS1VhWd62epfw4/tVUT6V9rY3KldKda/hJPFD9Asve
uVGVPkduPNwFOOZd3mABHbNVWYzPP8K80ewGJ8rqV+E3iR0kaQXlx/XZItyDX5XHZf2Hdpin4Eaf
Sb4p0yOXruQjXNDAHQ0uQoyOHW1Y983kI2aNuOioAY1PnGTYsm5UX/gg0pv7LdfARhXOZPNGPHF8
XZ5k8V1SbQeD1MOpkeuti9XSZZanRMeRULHpvpaUdBLpJTGmSR7SD2Iozv5lQ5JerRw2hz4F++xk
WpvdayXCjYFwfEuAZot4OroPV2FUxsV4mjTfYcdYOigp74Zv8PgcxDUI3FirOZ4WWBbhDhalwHwG
hi+5mLoz8GokILFfZ04zFMfiOlZtjHgW34cMyTSE0/pknxlPWobtBh67bIWKebJ9sfzx0ctAcOfE
1B9lKYkkZ0GWf7HsTvCSLfxYo/EDS/OmV93K9e4CFjs+lgEGOEnh49RU4w2xzKb+KKB2KBzyBca2
i8GaLNxGVphTDsVhBNGUPEQAQq+EgZ+s5FManer9kDuC814jl34VscueLSD6YCH6emXiVqAktnbA
RjgwNafWzfAHap1GjYedag4xS+S5P/rhbbdsNXGV5sC3Lx3OiPN6NaTbjfuZVXu43nqDkYPpN8Cu
Je2VO0FRUbTrUwbhmwGK//bGJTB8lEYV70zhKnFJ8HwLXKQFuWa5EesXK24huN80lYNejgadW0Nd
VBjZK/1udnCrRrrnrRZblXBYffZINWKkar211gVKzg5LRwpBD83RaPgNo6DPUdzRXMChxxlC4tfB
fq2shpPfxQyLRcAGPcukuCqeghqP+sxD6qTCGJEwcPxHR2d1CWMB4V/bWR6UNjBdd6z7NSlCsLg6
EoQ44bglvRMahepqe/5SKFbeu4BtD1V7r6EwfTd03b5HPBs65CiQticQXgXwmBrxMfVZ5oWqQZF4
PUjAaMPA+OUw6dW2TQgfUM0cyXZ2XW4jOvWJ6c/VDM0aio1fXGkeuIN4c35s6flgXsyGDqf2/bMo
exzecWeAx21a8eHUCef2I8IElUXe6kPLvX/k56PuD4QGn1Mg6rLWv0rx0KZlJDCi3IMNqqFwILgv
lzztd/k4S24WCcq/O+MlRlx7uYnMxGLjKTcCQyWEKNQleUI6Z8stFL5yyughQfjSLVFv0IBOzGXn
XxWClLCFxXKBdPNcn+XTgNe/WltkD4zZ3jFAccg4Szy+yf8P912C9+zfitNpJi5+Yt3o2C0r7zWV
aaAogRAQONzRjeLxfIdIR6+mqkLkPegRe75VHzPmUFSZ1k0jmHNOnYhIYmYN43wqmiArB1Wp6E4Q
PaqvfcnTDgp9+v2K4DTzhM/WLi6tlC60WYSfQQkMVOVzJJeN7U7au93PEH9zN9Zkrst6qyqQJk5c
6gQbbL10vVTxB73rybeCSJZQZWAIfuzfA4e9bHiBhDoYZmZ0axiG5MvXhV9/CBiaPb2c8SaYMPAH
PhU8EZlSa57LWbinwYOX23U7bPseivQwNYmTP3dDLr3katnomVIqr0UCtKTmltD0S34SoTu58TUF
ZpDBddZ4NVCaevsth91p8F1HL+f2hKQui/pG8jxXM6/GS8AqzZqnJBLYQGHTJK+KQfpNyr7+zlA1
9smovgf6GCVhVxd5NxCw+xJeePZ11r4JnsrXIwHDvk6O1mi8kAGFJnnysX1HIgjNGRejPJM+Pq8R
nH6SjRqfwgO9n7EeFjakC3MzInVT5Khcb6fugx9jEjIdEhi1SdpXPlV7olPT48j2/KYR2Cv2LyrS
PB/4Aq/YF3OOdWdJ0gCgXEx9OtTgxAdK7uX93Y7xbwh87h5fQDMduUl+3e44vj+qOZpjGyP8USIc
gMLZ43iLChPlpLPFGvoHUTN0zrrKfi+Cnhn/qvaTtcJrdHLSy69giRZPIITSQ0g0pD8zYmrnfD0K
wJ3uHVGeANOHeJ75F1Yyb02SigsiftJLpw2aF0Rbm6qYkHMvzO/C9heqVdmL0lKqf2NO8Ri5eGiu
mlKnpCVzZgQsazoCJORYebTNqWCfjyxfFk2ta/II25FVj8dwr7FEW5fkOJdt2fxJ3UdQeC0HJlrY
wlT9ln1lHMmS2dtkOTfCnPb+RhvRN3G5RN1oOH8znMOHnkLUDRmCfxCGsT36oJwqvCoidfkA0hM8
lgl5fNKjsAcsXKcv2HVu58rLl54yS8QBslKsCFrV/dD0KX1UCOkCTEOCzy/1628+AcHBXTbF+59d
S2qv02N2cZGpk6B5PuKu0rJQZ3iq2PrJZmtxeEWAym1oa911JuZRHWkzHe+XjHAWPos5EJJjskBM
1i2pGYrC0Va5q4HhKuCrPPxVwsNlc0UOtHupsdKSx7qeBQtAP4udQkAnv+XSr50fh6ohHYVKhTn9
E2iR2pFEt9Gbn9/DTSzVWPBnxOtWBEwDzKb+CeQm5TZCPOpokBYSanr/qIq9kCKoqO1LFWGDifTI
7V4eWuPNh4hO7D1tqe88qQWkZ+AtU/R+Y3wmA6IDrtK9UA2ku2jrl2NKEyexuBLKBOopXgXT3zIo
Chcp7j/6v9mSCyGfXZK5hS69+1B/+QtFodGEMlAU/snBw8azCnvWPurweooAyP5ne9jd8IREB5SZ
slZ14zRRBwIUs5h+UjbOUNiPop97nsVahtPMgMdWo07ieTXxhSlzJkqiF9ngfgfPcqaUr1knUlZw
uFk1c/CX4R8gLNlhB2q6+YVsDWHn5qNH1WwUsHDxd+AiDUoOcaELeOmWgH2J8SWqyMtiR41fsI3b
zuRNAbDcezb5k2nLcnBcSeY+9s2mWRqNTo7RnU9rEaZxHyEr4+G4YCMH0TIFd6DqRjqtN5DuAfq1
LpOOmk5CvEGzpCPpbvK32cVW6SID/FJ6ti35BkM3s4FBk/uv6NW4YOWw5YmAvjsb/AambSp1jU0I
Y16JsVVJyP0fZ3hLzKYCNMUOqlHaSLWlZzW91RLtLyODSGAkH2ZgorjPwisjjNNkmLPFEdibmUh+
L8egqqJtXPHLORBvW5BlH/h3K+gpiczGVWA0rwSLitDrnT2vKo0EPW2pYCrK2bvYiPpfYpky8XS6
cqfl/gKh5tThMCpdcPYCPhNZFpsQ3PS6dy/3hi7qJ2q1x/zZooU+cns3KAlyQm8PcFYlKT/hfM/h
Hec/gMxsu6N5nP9WNksdKqO2PYfoACXiSrvfo+Xl/lPiXZGl0Jl0pFbQW7zSZ2Gz8WTVTTJzqxod
n5QvGrqJS0nX31H23/ryemPhg0l2/ImIDe07grzlztx+hfoIp8zNIsXt/yoBgnin8P8a/Lc93eks
qaFOoqxE4hdjyYQ02B+RqRj+Axw0EXuL4D2Cs3jsqEJn0e8LmmVORLXzPVGd65rUhX7qK/T/u3dw
rfc18kK9zyTsPvPMT10jTB7fkZXyxfcGFLvYDUTgsf90+UkSuKOGoYqcoYSj1RXxmObEXhoBvxgc
jTGlSii9A9nP4JTqLd5xp3C/SQYAEes8mUDijmPTug1MehQam8R/RnDGfFY0hoEckDP1gImgXEfR
RJF9287sufsLSMU8C0TlmqFa+jZLGXpgBLixR7uvWjnjSgI0chmAYtMFiC8txVl+VZmXkk/wngto
l4QgzEGorRBGqBNrM6QYz8YkGT8OfV/sR9I/DV4FPr6VrISu+M0N3PTlTmde9KRSo7UW0I50cl3J
oxRhGXc42rIeG9nazXnwHt0nZmLSaiayCWgnsPncayTWGb9hdWyZRB83e/QGmeFxoEtrTzytFvEK
x9iAHzoW/BoNU1DCbopFrhLtiqIz9XHE2xtmjKWgZ5v3EpL+Zurjn2LRP3Ak7Vcw7ncIU6SL2/aQ
/hAubULy/WGf9wabeJ/aEX/GkM51G+TK8qBDqHu74z18wGU1jYcaiziwarDl967a7yl+ItruQvC7
0Wi2l29nuY0DAb9AFEwA+V3tTwApP5t27Wj5Ru14ZbUuLppOOrRZXh8RZMGBXS6tV1X48mQymJkc
ZovihCi2/5Hwc5fwy+uvU97MC/sd3pMl7mMMTZ1V3D+TUlCeN7U6916o5J+3/HTn/OXCO/cJS77e
mvU+9jE8nP1rwK6ZRh0ibiGBLSFMbdQ3bOEAxYYyTuDa2wq9cDUXFQnIt3qK6PF/Dsf8cNGIzE1c
YjJSEutfgwMngHUtMf7BtMnawzzwDIhDT9siSSQ2XpIOFXbZBx4sMHzoL6T4lSDhtAw+Qp5WOa0r
vJzfen/QdMh/ja/m4WR2K3KN3oBUwq9fRpE9Hq+9hrxl4+zWysYIMJSfXq1wxsbkEDtTI6QS4Dyl
w4p3debEir4PRkymsNeCxIH71eztMw5v4zmwmpRJE2f92laOQk6VVV0VrrlwQ0Ktfmm2P0Ym80CD
wo3jQV4tF2m9ftVgveLdA941zgrgp4RQqK24BjFeX2yfaPqvL4mMyT7VJFeNAm00RHL07MynxeRH
e1oziQyhHQPw/FXLcfuQZyI/Hb5VvgPJDMHYuqf6toG14/wcAOkJpWlJM95xFHdJBU3UrVBkiJKN
j5O4+gVkoTwsWFm0Z72ycG1jCqkzvqtirFBOffuyu/MZPzwzfkOpehYvgunB1aLluQDW5nzKVMRU
H+ej0OvnLd5KXxQTBLopP7Q3sXaHLGS3m3HFNla5lx+JygLXGSXVIwQNZBxi+ip4nHGL4dYRd5SU
g45caWt3HjyJ8dHP5SF8rvQYrNXf94UVLzgK+eP5lZ2nYHS3krj9hGW5Q6pwL7tNPuGyLvT7BMi7
leNbX09SArCBXtbhx4UXlB7dEiIOyVtUkKPnyv44Cnf3SPlmrE0IoY3dxpUrw3Cj+evjDClWXeaQ
JSicwf3EpYjtC/OrMvfxnij9ogd/eYNXiXFu1iWhEux04KSpOyNMHwquu5DnxXQ1EDCjIdLsN40J
kL+/8VMPQnnNqwOLnKbtB5BuRjRp8LSyyefXWTBGqbKyuLY6sz0rg5hgNtiRgZ3M7sPE/IULxUf8
PdhBBJNNVrCpXMXAdYEeiTUK34ns0xCOZyW5QkdpKawxLuOwQOsiGXP+YZvEt35FxpaZ3c7mYvOr
1Ty8urqxc8ASHeROJmLdgncbDkGvnjYytHkTq1GreawT9lgjSTHA0npdtlGp8pyG2MZF5rxXfFK3
/cJwzC8PXX++oWTnePNLq8TKPh9UDzyJLDIPCnDL6fspGyekojg59kXWNp/dYC0c+q1AvrgrP2G7
k0VLJKjZXjkWdOvkT6lTjhwR0d082McTUbxjNWSDBgeKV5HfvamiyjecFvLU3azDjsMajg/GT632
/04BLyZoywEun2u1xfn6AstMlf6e2CNCmJmBmrtf2v4qz0PLqJZ/X4BLprbfeKuziW9cItlaLFaQ
MFSNaVVxJvb2ij+hIYD9tyRjNXkLsl73KpUoJ36MrHdWp9T54DJRLQUrqLqBLfdQGMWrnzm4i/Rl
2bCqZn+jRL6mXJC+WZ91oY9KBxw5evn8fXGCOOMTGxzbnx996bsXMfEd8ahWDyqBhU8i7v/Jg7pD
8Mnq55+ZpQSrlOQ0PuDIQitPJ5Oc/9WOQ0dObRGiu9LSqefh5/gXXFmIP/wUVv1NXpAz1XOP9jX7
XB4chSLPVtgVMYodR+XbsX6slPOyMpFdOo990sJrtMp7D74u8Z8osAso4pQGKezumpLf7VyHPc5T
3Wm9ycE0ceV68zDGdjygIoG+NP8Cc1CEnREp+qqlz2BnkzsHMcnIOKJjlY0bAcieputoxVmTImw+
lU5r0B5C0hEApiNCClKxon1cTPwMquu55/o7DcHnLQwfsdN91XuuGzv/S5PbXqLu7QziOxETDTaO
DokXkOF4pYZvhUSrtWYLFu3g6bWvp3t6CNjAigiUzoSk5NX9QzlAbSSMazXLKk/phGl7qJ454ZFx
5bxlJtFeUrBrzytf0prlJC+LK6JtILXcGJGMillh/8ew9HIz/XTQQvVjs8FGn6JVYlE36x6dGJfR
0rcuACltJLvn+LOmZ18ZKlFwUwirv5NBDO4AgJYA9MH6vFBl6Jv56uN9TmrROsiay2PHoYoDrwff
IEeC035Xnu5iDQpsyHLA3kATFQk979/jeF8oEWb9pW1YbGmKFhvH04gp23E4xrueDrRhzaxmdTyM
TxDNxHpLlQvYmNDSbxgw+CVMoM6SaSVJ/s/K3tGde7OWdivdf8W/hni2Q+bVijTG/p3srGtBbE4c
5VT5X28ni5liySXRAcEvfTwQyzZP4RsMZDpIijoPm0DhoZYnkwVKmqo3reYSZvsHzGM3I6yxOvqy
gbrFJirJRDqB0r68MF099+ATM+72JTOYuk69zkn06RjzmwnfSTZ/vXpJt/w0PikfObxbEZAy8Ens
ZegZofLe5bDbUfRgO93cBD4uQAh/4Naz3asm4EL8lDWnPT13TemVIcbuOMBoMYfd3FrtBiN9SAge
WcBLATSheoXmStbt+gKoNZrqtRQZ7x5YsbQvjUHAw3xScT95OYj8jkrHd77WKsCAm1KAfi7TzFES
mniY9SXCj5QGximPDqwUXOHAU/79Wws+XsHSJPpFwYMkDiP31sWyVvO/wwiBVtOV0h4hY6IvhW6y
6S5Ny5ZBjfMx5dwA3TV8DiWp6MRl/ZgfiYrhmFUiOvqcB8/ISYSrIjiIzabB0Y4xwebNePZhHJie
dp1j1VOPqQ0M/OntoFdGEBL2vQX1ZPZVGsSCKQu8brZIw0OD4RMZ6e0CTy5h22T4cW6nKPxi76Cl
jRfuqcdWnMjuugdl6iFWs3fznjO4Ww9jkPALSe+NVYwjyv8ahgFIB4xVH6h6ygaa+nXYyHX63WFO
LNJwZZ6eIDMIWlO6XuTQQr7gp3c2Sbp4z4CHOTORlTq17uhtjXZIQ356hEalbzHk0yog3hd1f0ic
LUpcM6UdtBb250O0fR1Of7bpZk9ne+O+Nu/LXRToXgowYaIQfPUQoZ1mnHusbA1Vd2ZqUOYrdE5z
CQU2wu58fUDdob7eb3wXT04+BdhOWHAvnKiiYuDlFf5clHlIb/0LqJlfUpGLCaU7SGCENngoe59T
kfS6a32udnC6OOrfRfvhe17Hmw1uw08DHM8tcD0p7efyMq3L+6RUBVDqxVGq2Tmm2eEcUHReb7Nz
Xf4BXEJ6i3Vu6L51Ldsu/WKzKjIfYIMhob/5NvewT6nr9u9fxj/DpQ1pTItgHB1sc/FYz88XRA6t
xnLDxn8xgfoXlrlKUPxBD99VjDT4qpgMTLVIhrxdPj1NbWuuID9g8C1rRU8sFcQWn1/818d6x1G4
wvNh9gymphyKN2fxoUBnjkMbcG3zb/MFK++S+CoaW5SEDUQFeQTWUdqLlEOxksHR5LD5Uxjqymze
voFQOjvwsMTk8ynz7nJgBFwavano6xPzSQzzKmwkGHnsrpYXHQfhMTyoImXgd+BHJleTll8+QYdF
sTi1grqvpc8yVHXmIMa4T4+qr4MzkF9h/RWpMgFkTOpxQmGQtJZ4aXhZToVfL0w4I7Mvat9Zjin4
0CgF1JkctFOwBAm5S+4yrxG1OpIRcJTpR7YZWW/5IdNEOaeHv+hpPwb/kCoZDGdhSaoixm1Vzeml
2FgluuIsBGfvaQWpANYcqP1mQG+TKTynza10CYABLlUFiVvXmSBCyjCOrzAeYOojyi9COi4hE0Hg
rLFkqFG7zETgbkBMYubelUWi40/iF7wtpZDGVO5HJe4lZWc4sZquqBRQC7zDOFe5ZF7QuRQhCy28
5jPZf/d7E1g8KGOf349rSNcALhnmjKuMQ0RInySwyTL3ab58Hbauuo3gVCCAUVCEAHVK+IR8muHc
aK62G1WYlXlXWMf1HWOG1aVbdBvK2ecYQAfXdqAhfvjZRD57JmfYVA1C/PxDN/FF/KzU5qJQqYZu
TF0TLRQRnZ3gQzsLSa6bRuZLEYO+2bs4NM2XAf+H/MxYBjIZDqZhECoPslR7N+iTKxR21G7SVfrL
8GQrloegcwWtDnqt39fsXzLU8sen41jnRMiUT8xgUgdQy3GaDLoGWdX2OqGQgEy/ak0GmMmxdOB4
IeXQa2gek3p5wZM/IuY52eCMxeU5KYdMI4B4WkoLxWA5yuWtjen3//1shRMm8RQ29HZhz7wwOFtj
dKPxYmEV1n8MUV3E5fgYBbJ/hCTvpXW95LtTCPCCqCoaBoVWbrwOVdnjJVfyfqDLzHopNcvSpptm
bl4p8IWg53ZuVMuR69f637UPLO5cJm7wAEjIoT7FiV6wcjj9gZ0B01z122Vy4vSYTYPbG9qpEw0p
2guNfFWVBlf2SxjybzEwFfleuZtILyhT92LT9FSgrY4ofEpJhgfabT+fUaMlJbCHuwwReaZwLVLH
DzW+uZWTqTHdYMfmXgCcxJwxNxyroZACreKl1uYGGuX3rP9vk3mdAMrUhgWPWEH/R97C4p+dCu+2
EJtSCrZlvSIjB3x3ZPHWhD4U00O7VzZYoWf/P0aJDXyaeSD+Oww3yJanwFzvyxyetwd3fRHucbRF
sPXpzQOS7WACXrhv86b8QNreHg2jePk2uXYkoBLiAx+K/+c1l+Soxr6pcuQ54E6hIIwxo5Z/6ksn
RYU45YyW9Q5NirPhyJFKZ97AbSjCDPD8x5nx3FL+XaTpw3p3Oui8bt/IFlLPcS9equkqGBsPOnqe
VUtuZDOUl37CRzAcwpiPCQ/b9wMAeCXUKDJiQlCRMZu7BitPI78idQ+D8dIRrB0hUYTjDSpxfMJV
o3dT0bZ5b4UQ7zF2nDCgmtmyilD0zRSnTZFwt2g/LlbvHtJ8WY2hpst0g8/ahVejwtbuhMUSxCVK
J8IO2+C4oyyA3RKNpXH4wfADpZfgTvNicHnnPB+QUNbASZnv5xAQ7KBjXG3pyY9qE/Dx3aIbvSNO
nDqATCIf8Ab2P8baT5Hlv/39muPNouKud4ZqUh3mTV05DZGCVHmefZZDpZ4wVV6hZL0XrT1UUknY
LJAJN7JLHlEIDJL7+ToR49pVyxkWX25ghl5Ffb3SUwy8GGHdn7VfzqaKsWDcpw0Nb5Nm+9f2+VjU
I8t7wi/HEZJmU6tw70TZdGKeBeyQydHhdlNJh+KOteNr1OlFOlXqhFPW5Tjz6klejmN6aTize15e
5KI3KGzIBpgEs/Vz7ctR9U8a1QL68RvGR/mbykrgbdUlWKW+V8qvCyl7B2ScJGQ+tBi0ZulGTzAj
1siJvYekgey2JpsX4Mecw23WhfOX4n+R/CQpC83q9RKJCURfhUMtGhDoti7T8zlewv59XQWT2q15
vkaMSb8dV4gWNl90nR0ay9wlfWMEnEq42uU7iFNMU5pU0wpkl1vi5PVQMy0X6a1CLyPs9M8zo6AY
baW5fNf4NG9zbuTD2h0IegYddkgf6iVSh6JK4++F/uL+boXVTWG49jCYFMsIJS5dFTv2yJzLXO5D
uQxLRyt437AXq+lasTZaOt5UqRf2FvGB/YnmdZqsahP01uIwyapwyZT+kVUXAWrYUXuo4xIWxk6v
ECaolxG6UUy0JjbukJK+iXabD8UMIfTtb4KKlkGHj1D6ftsbgLBNer5UsatcolHb5NI4hnl5eQCN
kpYjLarNMSgBOfK5bTcRyXfz86Mi6h1vfbIMYrmLRPuFluzyxkeA3pyEkPmDqZsLKXN3qcfZuu7X
AP3cCir5Oy0Pf2pGgNx0temeTl46rf2S7taYhMAR+UetDgiSNgPVnnlJXfvNKDR4qmJhAwCW+Prx
g5KQMunkhDtniLJFDWor5VZP9dQjulJpDKR/AmR5w2CyqQUDAHXocRDiIusoTcB2Qmyxik7jiyD4
OF6OUOiwPzxBykpSXaS9B2Qj18ZjOY+Fvgi02cLdGr8ekDepu/a87DElAQWODeW/baotSi9e7nOn
KMNHa1foNEfIvqWkK8DNoLbgqYrSNGF64QXF68al4/wMZf95bFP4Z2gK43zrHTKstWmFJVjkzO9H
le6ZYS/D/4LDrNvQZ98mZ/lRteXr9PdcwxozlxM2uJTZkAgYDyqXMp/JFn/hW+EHpDLyuu7OVbho
1vZooAIDy3l3EMdv9m9pRq8vS+4vFKVgtEa6oPMwN9GGYWvkUihKzmbygMD1Rzrdk5cSivAMu0O6
lZFKjs/WeHvfbk9p6aCxjtC1etHyAMtlR0u2q5MJCn116L35h//W9d4a55xb7vYkQb+zKjUWPoXO
n/zgjcl9MOSWDXly7JSrzrlP0Mdw1fAwOLgxk41guWrXAqwLW/fA52HzjSSEZbXTCAIEsI0b/z8o
NV5SNJzYzJtFFdJLESHmnzV8ynCQdDQm0WH50RxPj7IJ2+aJPfO5xOfPE8skBkQb3RbFebLS3vuB
8zVDPPu2X6zC6r4j9E1U8KSlM3iwbO8/IC3Mu8x5h/y9iUfywc11TmXCPamO8KF8rUCM9LDo7oxS
XQOvqBpMU9iyNAjvs2J45fMgzE30wLL5BvjP3X2/qxB9pyUzfAUd4V8y84VVa8xAnTqQtHAcHUxc
b5JMgUAJPAiNVmo2dgW1MULdVzQz5EOmtHuM8NWOaXo34GuWwg9PKTGrMzMCG43MO1rUTGA1LslC
lSZaJB7tSziAGVU053D3/Y4EJf/9ztTX/iKWOADjh3B8kalhfNV2alxvuyybZ5kmjkRY+NHknbAH
RpkjfTNp5JFTXNoOhEqJLK37bTJAQmgKqJpK57VHIp3HBv76QLnrqcUUnhUtMEsZxJ+1C9Bdv8gL
KksyxyT5MCyjtHmQJDgE3Wo1dzb+tvv7W0ALyj9ObcwyM8nNSiFVl07Dr2A0eUoCR+42tI+CPbtJ
LDQDAiwSJivdSXhj51KeB2yqRtss3/7L91SczsZa4MNxHsDP8u7pV6MwbtB4ABP5HV2li57C182D
tuIUlcZlN2+yduHuyHd/VaH3G35ay5Tkk2oUnjIIePydtolWQ+ERM95ru5I/1jd1+b0Hu3cyYaol
hQkrTX1uwy+VWgyZxn7iqqpLaaXLruPXHXhZ9f0x1uOM7JLqmiHj0aeRCPOH2rrFWsMbWMKlMXzh
QEOlYAjfmqHFyPNiaea6MDN3NNvJMz37yYjnTF6dLjgMSqKy9kn5TJgYMdJakSbA+NPVoaUMKP60
TxPWc6H6YA0AjmUbBqOxiFzJkd4ULuNXZcPqrV4HHqJUJaGIEjCZyyxctDWwrpOb6fYuzklNNf0u
VSNPuHmOWv8RbqrOjsGrSZU0Q5R8mPcbcsgX38qE3QMR9pUbUXm2FxN7HtsGoslmkjzXqmHJS+Iw
9YUsOjfPddwryY+Bo2prHEHwkgiy66iFdY1hApcvR6M0Cepw2VfxQVSJEOJwV0gR00zjiPh/GSZy
+FkgzJQ9vx0gLJ9qW81L2FN8mYbL1xD2OK3P6KCHEVHksFSMJqtRQ6b9vR/f0OoamxcHo+OAxHNB
z7oyjDg1JQQ2lM0zxF4mfX/kgPpBGFx0EL3NPFDqAsTenNk5YswxYq7pkLzkvH8QlFan1pQbFDNQ
u/u5dSOnYIb4GRsJa0gDl1iskX1OTCToYQcmwPUPhPs+fABSE2bv5AL90FlA06faZG6HrezaIXeP
75DdBdSooD8gmDjtbyiDs53ddXbdrElaqBnsbiOeH8xrfJHxtYfDK3YzYFl9EjOMoVoi7LrnBRBD
NrRh6a2D9TBUZhnNovHiAxMCN7c7ajzWg1T4uDU+Jmd3p6XyVU1U2z67KgOZwTuMltz53Umz9Geo
hdCAzjJHYh/v/Zc9B7NDVYf0lU6vYsp3C1YQMOzUgWWHawGKr2BApKE0zSkBqtQiJExvjiZVZJsu
2R+ptf/2tA91hspCe6OtrKsc/+CwGuPYdxrnAiQsIUfLoQC+25PeasXkBVgOC4K6kPOzwJR6IUzy
TvkhUkw9p38EpGWOPPcjLSNYG0PbCraxIbtx0hspSCeNuLfQs2cOTwUGSpGFC+ixntnJB9nCoIyV
hS/rYx0rID9Co/NPNRPz8brZ8/Ulyu5f4rqMgce+QXY9jlhym4NLZ0P3U48jYKHEMLleSAsE4uDD
0WgusDitiYh5zaP9Xo61N0nJxjZAZDL6ZYTAcW2tV0P7UC46WJ1JksaiiXNKpPPUp7ata1NVJz7e
L+w+uERhKZqpdeMotiVkNHOhAUF7fYJ+Cr48HF3g0g9eHZ4XzyvU34MjACr0gpAW1TgWtwJ1/R60
aBxWj/IK3Es0KGCg5vW9dtzIZZM4LfTnFbT6FwAfCJJlJkdAsRfWMV6fULc9Nmkl/pUrrQ1xjEfy
UOP7CD0gguUkD2GdoLRaNxL8eSxRv8A2f+WHc6XNU3molPPmR3x2YE+wOY9YXX38DMjap5BBxDYq
uBDRAv4TpachxryTq5QIcFdj+WBx4HAy3/qGARVYvMrz7xKmeloXCdlJemT3fS11ZfJjK9f2MawH
34QOMHKr/JtvIrIc8m5FQpnIs1Eo4ouKOvZhFzJpfVLU3ZYLrJsx/Gp6KZES7S6uNezsgz/Xj8JH
5P0sCcFTNzuCkpmB+vfOYD3MKal0SCjUHTPAER2XAdrZKCx8hlluOyIwgCD7SBYYdDNo/ZkUrue9
y9vx4SuOE07eb/CWNUmhRg3wqNfpaoi0eIWeWH+QWi4SLOYl7DpF4GGowHjP7LtDVPJ1WZ1NbY+4
v+eV8/ufcQKZgC5CKNll6Z2L81jtqHJ3IsN0304rylkUIOOvX2lGD5OMJ6CUYDMLHPlR/ZS0TGnG
4kRqbLaKVQpYAUMRwusUE+PZp87W6jGnH6mOWIYRau8Og98oOeFs5DtI7AqITkILJI+93LQJroxS
R37wSMIZHPst1k8lRVQYgJsvPGuPqGEGqNJSFP/B4hZPt0p26af0rFygbyyfV/Q8LAaxhzyyWQJ0
disTkSMdJvvV5RPf58Aj/dcKVW1YksuUlpd3heIPY9QERw3Lbkwyr9sYRMf04uke8dWAS1WsgkP1
ZupUxAzGDHJgQ2DK+EUSOdp7QCRP5W+s8dvzPDvVtT9QpcxeKUpZf1fBb5Zo3MF5SW5TxPdJMS0I
m3uA1vHMd5lDFpxjbasjorHmcPyNDXIfrqWWzrRVi4nXQR3i5UBAW/XK9KZdarnOz1MKRmcVH7Vr
dDwhdSB5OIbx1CbRbLNP8SeTLlR9zZVfTWvILLalhJatuJDC5K7ClxESS/fUIaup0Iq1m+fq6jiE
DdHnwlu+Tz7GBoy3Q4cBiJGe5M7YrTi275YtX8u0ZAZZOOtcljRi7HPec3dKYyK39h57bZwdrc4R
TFxo9GqQJMxBDSI+90ppfJHXNi8iQN1KT9ohKY/E0EyOcCFWO8jLw6iHQkF1SaeAeimde+ZYyXYw
E9gs79kF1XhEBW50rIZKJqT9gEZcDen7jK6G+WAoWlrbTo0BbFzfwMhDBcA+ZXuLPaAWsL0TlB4o
OkxJiWkTS/NhIa6sHdN67gIg1LRskLJvdsGiQGs3sUl/gAgO/UJdDlQws95qAUqJeR1fsZhb7SU6
8VNYJjfiL4ShJXMnOBLCyYeTM6jIdXvp/RU/zdml1mv2SyfjpGAytWpbbDGjP1KBlTGnr+wSShDK
zRhgyWWoKJ0pR5CTKKRA9BnObtkZHHR3DJOFcP+xWKdx6MLfKyeMv5ps26luwS42LZogNgKEFKME
cuW/jJjRsGk8ERLZXw/W1waBXgvXA/KxKoqhh2efB9k0xHVpzqqWOIHXlG0xMyqt5cGFQ1Gc6Oze
AlBpiOZRIUzAX2wCWchrIkrTWga0Nftmk1tm4CTAbJhIs/zluWcrCZVvqF1wPKg4Dm/iX4pyCh5H
uLoTCvuA5gFNXc1mrLucBDB/7+mxf+IZIlIti/nkFfjwSJf8FyBHZMge0OUcitWbVetqMRDzuoo8
UiJyhCTulndFmH/9ct8qi8zXM5ECTUtz2l9VT6fsYFHpQUQRY2SjLWy4gKgq01eScA2mEzk1j39d
7sY7spvTxKtXLeBehzgXncj8B8V7G9Sb4tPlJ4c5nA1MMMxeD5xYEDgslQR0z/EaIvQz/1u5MH9b
YfJtLIuT2Vk//MWlHg2ZpTHmttm/NcV8jwzwPnRBafCSV4PMWLCNlc/zcjmHaGkFg/GG1vIugf5H
+o9iJ1h2Eufd75WwfCMCx4h8xMrqjCp8nfUB4cTsPxkYasutBosYf+Yb15KbdZjA0cpF+w9DSPx3
/a+bW4XAxRT70TnNUlKEwhhwuuH7XUiMUkL2MPC948Wgbtae/ylvcz28sgDlfW35R4cNjfSl+j3x
OlRlAiMwXivZLejNGlcP0HQlF4kNheNWI9W3GK67W0xKqm9FWf4LKLu5Ew2OTKFU87A1Ca1QAsxj
QR0HABNgrhldpDXPbf5B55hqh4hR90sFEcPXFTgmgirDnibGI+grrPmswFiQaxjwRATKskNqFRI3
cOEYNHWCjxaCmxT6G2w41W0mq5q78kJcGcuJajiuvJtqJU5YyJPz53OQcU7VR24Em5SPesKzcGKe
Kuo5oKLmH1BU8krIj4Xw3xexTqqAk6TuzcEKmGeFrtRi+F+9MXLf3DJp9M01Y4xsdF3Bi3qombHe
udvfm5LMMDn/Mvjdvz6hTobvJcckLA2GnVtT+1gHDn/SnE0+7IFIEtvPBam+jx5dNsuHhorRWyKB
kkdNeP6BU8d01MksLRwRvAJx/GiUhc2aEBZ/vbynA+rOoEgseuHA98zHRuc7jQU9gT83KoyIVBCG
87QD5mjjtS9IH7WB0DwbX+O9jTICAQO8lo0jM7h/xi4WZ2aVqKyKUiBUB6BfTvJ1mgUnzx06UZ6d
JfzW9e0gaTACia6wc54A2Ohgz3GxZwsD2zcm6sbqgxQrTyqpo2WT1YeZmkU02FoBgl3mSItt6AoA
S+cQKu9/pFphGQSxyQ0w2zzVdl6Ntt/lQt/YxXYujdOh/rB2nHm9klH6xNQSDsGFLvjSLBs7RNZd
qK+bCp5Xww+uTRuBCrLPS+HNO7n9mLBKmche1zwsPWiFOJeQ9DWfhFAsZBJdQHh9DK3Uygp9Hc5U
JrPaltictZRMT+Q+rwdxdg8sCuEvoj2NdiwMoJpeKwT9UsgwrUU2smsZMb2cM1jP6z6pSBz/4mOQ
reOtWTudm0zXR0L+tiO+2EQm4RsazZ14bF1wl5MDqB2jXsnycrsNGUxMJoz+f90ITIL1qfV2YKVd
J/+FTxEVRKHtdQYFD5AeW03eSqvBzzEz0fCGbaZZTNFS6vKOUYTpPJZ5UlAafSwH2B61Nn3G0Q3j
6qM9eW8+7d+P4tKJs1aLd4Nf7Igu/V8RxahttUulzaOvbvsk69a/Y58JU99B9rvM3SrIpUW1TznW
zXJS1iVQcYs+KvMwhlga/4RRyvavRAfzsz+NNO5SRHrkGNzBHOzEciCT24BRWB/3OWF0yv0nExik
Vh2SIOznUDV+/HxVHN+M3wHWAqmy1DQdkAX2uoawV9F2EYUd5pggyaljOz+nKy2+MRP+0PwiqF+0
oyGvkJ5OD+FWjvUqqXv4l90hYUYlQcTuywUdqPcFnMXMCTrKCEPY7eH41gpCZYwjRhPFDg6Y8a3H
mwNilt5ltGttrGskqLGVckiWkhW00JokJSzumhocVP2bpUzVD/RbPt3I90I+lh33HOrfJ651bpnI
d33aCo3RMkNotQImUBK1dQ52fIDyRTNucntF+xHMbhQHM2V2k3OXLlyGDDwldULhs5lyq0sdx6Lt
tzOURXPNjO0r79P6NEZxBN9TkQUukINhzDYnaHflfl8kH3/V8X/d+HldHF662PAXIf8gGocpqCSZ
PNE4VQN3VZfxBA62DYcJgBHMGKlDz+yrxZkPzcA1c6hYR61RfCeROXmcO4IIsNk1xVXocfPGI5xf
bSDNFObyFn4eiVpqMeMHLJuVtmvfnb4LAaORqBbL96DLCNksoukDLUropnptjMX29/bH3BrVkNyE
NdUAmcbmO5SS8FVygJXL5NbB0Ka0G6e4ADWHQcpGPrkIePn/Ecn3tqoMB2uPfTfOva4WaEqvdbC/
ZMKbnoAhKYGLaUMk/CzgfedEpiq0oSjGx+RCkDZL73tzP69IBFV2SVktWW7il0JxylajgAhT+kBw
SNt2h7UFnQRsn483UwinKGJdbBAUf4OruS1Nljn4CzRdvTWHhIzvekmHS6qcdsr5GFtAg0KnpUa+
d7S8thGD0f1fAhHa0vKKztyz8jVC3p8j6FsPHM0ZG/2myLttHwofh/yNzdPOAPfQdLC1euHY0J5d
UkmRd7Df1t9RFCopyBMeIxPF+TNFvmI5rHYgvEcSo/4HiUV5N+i93V+0aiJ4yvQgKw2BtI8DzfYo
+Xa+JbvoJdl0rMyZex+hek2Kkkr29+wIZHQla+XiFti7y6RPWyzMoNYb/76U8ko1n3lmmTmYqbYx
r+NiZClw9wK5trz1rzMuxh+91+BJc0ROZQNYkKDqAxSgO/COlap5PBoqJ7M6Uzfwtal7turtiEEl
65t/9RJLPwvw/HGRxlrqVTzEgskcd3gQ+ZiW6SXBI/O2btDfNpjzJEwOFg6CMP36eDCiQL4ZHFfg
Mv509vKnrJVcvVgeQrNi1FGMv2CgtKdZZ599bAE6zuPY8QYkJbJJaT9kILKO1EM0HD95aAVB+WT9
JthVbAQta5FGj9V82aIp8dLeX2+E3C+hQ0SsVrYzGD9f2mPbggbC0DIIu660OOEPo20JDR+VUdHs
BeShlqguTzlOQIe0D7dNYTmrUbNY8xjZToezRWq0KhOS2foGv442byslAccT6FnG1T9r14txPocZ
AB9l7ZGlLuXjNr9sd0YralMkYFCBA/TQIrt8vmgMvV/ne0RGW1lVbfJAe0rtQeTYwQ1fwaluK6/b
UDP4j/wH0hDk3p4u2TC9LLSZ1iAGFO/M5cJc1djEzPZLs+0YYDAYh4TiBcYh9aF71s5bHg/cdJe2
UYYQO6d4msfA71+HkOq/oZXqK5kO7dr6Sq2QSXlGNp8UyzVQFJui0ADQlSTYH8vUQAoc0Wb2m+fz
zKBU0SRCPWF8s6WOCIE2yF/d6o3tBHoH8j5xKkjqbrfirQsvHuf9gD0AVWrCGkHXfTxJLo5RUr4K
rfVRjmMd7Isl+MSD5ImaOu9SDuud3a3x3KymQYzXj248SCbhZUU26IpfedoxpljQ1vyJAqQyv9aX
pkNSYOtNmxNmGcaufLoZGGtLFxFaaXFarpZ0epltnYYushRUxQjuyzwwIvT5ItFn15Qa5Uo7ZCN0
9eduCg/rZ2BzaGn9FeFxKOg28FgCQ4y1tFPz9cpGjdZzqIZ3tlExMHd9ME4FnhWTBj+aJug1qasH
x/XzbIx5EgCYHA82lAmxji0wcqGHNrMiOL4gX8dATHGlY+6O9jOVSCDB+B8DEZFKVtUqiZLc/lfj
8YAdN6btOOVFb8PKmKlwk9v80VZy9Mi1pq4bchbipi8N5goMz7tqMCQljrsI6xgiWwfHJg3BUi0/
NJ3Xka6NUd8m10IVk2S3He8rHVsdZX3e5P2c/SNMfPg3435W0CS+87YFNbDj6N6Fesx7TsFxxNzt
ztRGq//1TSSyX0ft2Y+a1kHt3FIUXSVCInn9bm1UYvj3RddyfZgjF1wEDCYAjSavGIDIVz7vOYom
EJa4C8DnrN6gyIoT/DFFdCHIi6hkqtoOphgopSdfRid+TMmNh6Tr/AP1s8qZG2RhZVLoybrA5GF/
nDK8/4BubzGS0Ma4Q0xu47TygjLW6p4mRlRToMDVgY00Hvj7y+6oKnrlaIOhEVRJ2C6tbZ8/oqJD
iAsSjKkIZYT4pJO5QFI8I9pp/LUHkAbnUhHg36vx1oE4+orpU0KRrp4AWkqSsrQ23bcX8NR70BAR
l63vLtzda+sJV4ADr5JwXj7kuVaTbx5uUxT7fw2vxDa/KHargNs5pz4VXbpQv8DVpPo0GILCJEZ5
dNf7i8F2Rb/jymLUyWEXo8+Pmy9p3tc83PsS7aGhceBFcx/2fN4965ZKVfM2D32DBqKYj96/tDRy
kARnat273FbnO0mtQydD4/Vl/Pomxe0T2+wYwXHFMOwUnjNzfTv2h7bT/j1pXL/l9RGjyVD1/DLa
D/iP+AlFe7RENMZqz8T3aRuzrzPP+le/km1FwMC6lKwMbKVzbi3HdXkrDyzt4x+/07fBFeM5LzG/
FtFkNP2HB0WXpHb+VvJGUmxASroAZFJBIrdR318KFUlG2+WYpbC64i9CVbeGptkRv7vXtN4aFnWw
fZtk/YBzlmlfWpeqFT1AK+QFLGysdCZXKloUd7TbVgjcWKg4IWZDSP57u6x3ZVZYwzGI5bwum5LL
a81fMJgVlndcZuzH/AA9IsHW+RDuKPqZTtrWMN7QxxoVXZaMnCGqTu9Ure2k5th6VW5yRPoNf7MB
XE3Zr7nPNa02DdoQPVHNwXSxybScfyXVlQkTnI4TcMnOfaOexvecu2+1SKGQVNO9RQqfumrL5qB/
uMu51JhYsATCUDRy8ivNUgZf/o2J5LPINd1vXce6bWKZfdfCIAVuDeh07l/+/8f+Eu1uDs/2KIwe
I3G0F51+hr2OJAMwt++i3cQf/wohfeQtkeqUeRUwrKB433dDto9P0oAIJt1a+r7Qcq8iS3ivqIh1
J51ebjNcv5VScLyF049fiJ9Aow9np94NEi67nsQ814gfWGlqrXDDiyf1tBSStmayJCUXjX/KGKhP
buH4v+anR1QcvasEvGWC9TKzVyAweRt3Px0u41qjKm+xfiunpdfNIcBCKopGuRvlJs/1aaQ6m+Bh
BJLhOEVRA46IlxcuTD+VBdY5slwcdug65e5IsN002BhIfCMkFlYHRdOPU130AfFjT44gX780ueK7
HmADUnSVeKkdIVE+aegN/kbCGhz8GbSsQoo0WTRy+NXvBnDOtgRStZ+6ug3gmVhkPWRnzWhWbrSv
TgwsJ2IZRvIFbJTx6JMznx8XDtkj/U0mw8qykV7N18akHM+sLJkSwhhmzfqmVxSEVYcBwsC5Pofo
l0LXOESTC1PRTFmzds4gdQ/zBLEQSPJ4CQ3inhdvtPshvp0U9zNrKsFF9N7h8crugAzg8tm67tWA
YwE5eI73qZhxHJSszCC7pEQtAxLlQkDeFERYoIDTNtyUTSpv1Fh1pS5nJPSejsmWB2fAXIYLJwrJ
xwI2j4qIlfi4awUuYPTGoHShs+V1u5jI9IOwRtBnpOJwJWIW4MM3HSmWRywIlTYLUMGm9DzIG1if
MLPwl/xMjtR84pMti911MRjFP4djmrKMYsBrocycQ8jMf88+c3ZIMBI0ZQhcKVroKpvTWCDxnF6F
uvcNbgDMJ+PGMFkR7mT+64LmwpMzT26ejNtkOlDXIIsvfL31+OCO/FLNsXCPOSfgXwhS2yB0f2QS
vovcF4ig+/mXi8IiHWA+tCWx3d6nUk4oM+gwyfEN/XbJ6ovihS12uhPwFowSuJ/4ieIyvUyl/SH9
vt+OOGOHV2/kA3Yjc95t6C7pWWVgqKBsBOaX6ppyIbQ2y2Np5Qw2Z2dxE10iSaLty9YhOjv6ypJj
lvGM4MQv9k1qiB66JXrQiQ56xicrdsZiB/lTpIVFnoEQ30/SPEuxDvBKSiozc0Q/DOUjnHa8hYm+
Rq7H0wMzjXK1rjyG+yzbhN+Qab94ASd+PyARitEwAvMTbxQK7SDPgr3rdN2MLY3LDJZLHUlYQyJr
vF7nHc16h9ydMEryIAvSmfdVZuwBPJOYBNYJp0xKfE6ivZmTZ6r5eCvTtNgjNM+3O+5QuEcNCvdE
M73FhbPQfhOmVxgWlXPBWTuM6D1uDGvewXSBzUUF7oOicz0grH7K9GFJ4mxkTn4YTWoHPTQ9ceN1
PFW22YaaZE3eaFRkIOIeUg5oBIjr4y+Z0DfLH2PiYm9K7udpTM64Pu0Dihbzy/mPc8SaBBMOGWp2
uzQj1aVITkPoVMCO6AY+aC/3bqu/1kUtzfsOWJhL0a1d1BUeROUxnLM/oB57xM6Bbk9ApAftdr8l
y7FWKfv1XeGbaJGY8rD7z/jRJ68VdTg4n4QlEYa32W0iKKm7QgaufpqspZpCAOFbHPhLsFUs2/sq
V3wpjpkT9ZqSWEcGqh2MvVoJyEG2fNWCrHx22abOHmFz+rptaak65ELaLB00nf8qKyY36g5xAqhC
qNqs/73TJmvvg8fuLdfjRAoPYYfq1P0wD8e8moc+WHdWGyOtr8g7/MBGqdMNmk18apsdquWYE1PO
zsLUXpehGJGFmjyDQTVS5W9t8Gy6W4QpeyhfDbp0gqCtWi4iEcKivSXMCHoORanwitz61PJNiI4y
pW0CVn+xM3vp31aFLjkm01VO0bsjWi2ANYmTm3pDoXDxbrIKsBs84uxAZXLPBUB1msa0nOMoOES0
Cl/k9Ka7XFt1yWaj5U8L0Yk4pK2wgiP4XukOpo1Ysr9FjtpHzdNcc0tmceRZQQD3LTJct12zdqUs
beIw/1R4lUXTIBEIzaZn1s49EWpyUuI1/2Ngo1Oau+PVziIOC4NsdxMWLS08Qv2Jd4hmwS0tWumC
IxDh40yj3CQd8F2txB4h4yClPSfovZYZz0YxTKym80vxH2a12ymzoZJawEFzfwFHxNkg84zomksU
dFoPwKn9SNaSVtwTXKkFSQKYW7TKtEVdDfwFw3cV4NWg1hYCIHNFZ12KRPU/LNCXaED9EEGHFRis
2IEhfukGlYwqJfAec0x3X+NG0HSbFDsdExEMzk0ZIaYMkkYpQnrnJP7T2Jl1y23+asO6Zfc9J31O
vzgjHgB5kaVWYWVBjHI18Obl6PM+JFFCIh6F8crbQiSO5o3DjkQqfliYlGMX6P0/3WEArUxmttOA
WyGLjDIQDVTl1YH4RXbrnobcjb5jvt1w7laiPQKpsmsda5gIvr+ntJXnEQyXMZkoDH+RblkPEO2v
3Y3ionxfiZNSC7FrMBgfGrjlwjg9G1r6QbgUepqLrp9hfecLEHW9l8lHULNj0vpDd08qxfM74Rk1
DM2yoUM0NNVPISx5djQas/tuW5VOdo8stJkeVwuhr98R9HtnJ7jPmGHyi5z2C+KY0z9H/laPTR8T
pEkUpsKU0tuD9VXlmZhTNrhPgdzmQBFC8kshP04ETuMmBJl2PkhQTH/EbGinU4mEEkNxdB03s8qA
pdbJLy7ho2ZHQfR9BSnkIeQi57MizqSN43QC7mkf0Ye6KeBjyZzBjelgSy9NECoSKwn/QqupqHCY
0N/zQv4W24bTPZTREm/tGDvTI33vOmSWr8+DJdrHWVYnwb1LkB2bhpDUC6y4B7JCTRc7vL4ytlTr
URzN4zaeOAlY5Mkh6eR7j3dlZtL2EXBek0ewG4wiA/T8XsnocGMgA6rcwGofqhyOrdzK5ztyxwlS
ihr8CProl/gvp5kdvKIvzsonehqUXVHd6n2kxZIAT0HGelcQXIDUrl3h/gdqn0zIHTtjLYqtBgdl
fDYLAVNR+Y2KkyC3c6kdstDW4OQ9L9P1LW3gSAaALGnA9NJ/v9gqHTP0H5n7OrEU8RrsHkCsgwy+
jVKcP/dVc3WOwyYs6hBCAgHZ++w8lHriVCXug1TOLTMb0TE4c2AVe5FMzch5InujjTTeSb5GDZGO
1hnn+AOzbwz/ZezRrazxdauIMsDIE2vn/154TPP8kEgDMQnuSbdemz0Ko6hfzYbt7vPUx2VwTLzz
6YMxQTnuSnWY70i8MZR5NlcB0EEPBZLXza7jTcCGLzj2dH+Sr111ZCAVA7TKswh0V4J8Ke0L7DaB
DSZ3N4NMf5SJiHLxEu+sVDslPhn9o9ItoXCouncqgWSPCq9EDhnyXlqRNWBgXQSgf2hnUV/C6poZ
tarStDFzFoTPXiJITckyD6k++5oAel53wAquEAsOVl5rshl/CRfJsdE4TMRVhhf7+r27tzYmLeFT
QwT3ZVhmZ3T4h8UVWlJwkk7L8LGXhaQXunqRKBpwy6TKZ2/i12G9S6iEkqFs58niGpxSeHsKGqtC
dTHQaRlG85yejhD42m+zdkExd0QHKDysa6MTodVy6oF5nXaww1ZYcH0UCvJ9pIsgySHy3wtOO6KY
BHlDM95yNArDXLR/wNlisXQCqAnB4j69EZQ8k389m+8GXqlX4XemaOwImQUKhI6GmU4KE8aRGNae
10K1WrMsqTSKg1VctGl1CDfCUL6Fy3f63jSKs5UCsB47yPBtCt8kez1u7WfEgzEMdJ53Fwmoim6Z
MKh0kZdMVpjxHRLeedVeBceHS5fEk1LASl90NNja84yTRiThf7dqfc0snzJe7SUT0Ar329Q93Gtc
vfVXYH60cDELrxNYvOc/+z3IpOQPObrXFIs5s3hfGWWYWpoNrjp2QEK7AdJbuV+CMRTSKQ82lG2K
0ESXw9D2mpTlUoaRe5Hh3/KTALRx6ul6cLuE1oMYf1ucse/hVRafAyV7Ferm37z8bFFhdLZFPO8F
p6Yq4oshwKqaXnR3bei2XM0bmTih1rPbuDKhKTX7t9m4WhNLxCiHLWp+ww8f0ly1O6ATNSEqU94V
8JnFD3jQl6OJRA9a0UJtNPHHnUS8CEL7wmzmgTAw4OxeTljSzD0203xISRiBP2HRYNMxGX+8CNoH
+C2z7p8V2obsvXsqPFVXUbGUPoBNQj2TTL9KBXE78jIZYPAEyPnkiJM56l0BxU+WzAFUhSafbmeo
S6irjt6aUirFmo7TcsUocIaAvSgFS/46fFq+okUA7zOzZxf+GH6QpFeJHWJvinTjY1vLCHbZlizG
clSfzKdsDInI/vW0Ti48CjFJM77YsjDkB7pvH4k2QapRV5c9xys5PpKmpTus6ZFqfeCrvpNX3skG
QopFzo7OzSWwwP4Qwc9uHVRVhgjTsBRpY0MqCH7isE2+h2AWOORx4MH9CoX5XSIw3GczvVqv2h4H
HRqW+u45TXib0+1KmGbdrJiBVaI1IBu96T9oWLqsqqDuZhcZIuwUjjrupRaW+NAH36fOwuKbkSyC
mAHhNywJ7Nq4mszAp4yPPCvs5LZgh4IqxwOaQonUXIMAoozuQHtqsgrbSMb9HbipZLKcQkR0LLTI
v61CK/KzLJR6GZvzFO2bHyzcG1Rx5L9mbDiJo0y8oSjxECUt/A9z9MYMysEL8JCp3V61VGAZ7M5V
TqzQfbC8HE2AWEwQHReexH4xnJzkxQfqWfKEcaxbyIQdjUa9UuaxRIXjA9YkkJNoNYwadqwLJQHg
Vx7JYaLZgLuTYOSk3JDHljeTB4DikdlU0Iqj9xAMU5Jg8x/Fy5aIafBNUOoC9xZGsyvSKbN1E7xU
FOCqNVXBfNSds+3t39jQ5ZYXx7Nf4vPFiku/MZBKGdoPg/P5SQZCFcotfhCHoV2f0ERgeDt0ePDX
xCUMdGhf/Zu+wE45kWmdHbDNGrz/KemT1Btv85amv5Zwkj4qbsAcmiH80P4fgilb5VWIoe4206pz
K6vxudytFV4ysK7hVHZEiUoq+s9Q8wrnw5eta2CsWTJ5Kjxl6q2WqIFoIpJvzAf1dBTympljftCU
JRPEGHvOq7WTZ0puj6vZEUIdmsZCrOvwIPjfXwkS7LhqUNulnHRRbbvnCY3Kr2M6bCYPUcb23sBK
DYxe3xrDtwiVJOyVpx/uolNXieduiuH0RuZxmfKT3imMeH4Vsbx7nkc6gKjsZDG2uiTCosNywab3
2jshI/huFiFcxO4pqwuaYMp1lXogH7Y5P+PLX3DXALuEabnhmrTH2YU2Ywtc70SIACUGJQN+FQO+
K87H9zDUyZxXeuhCJQULFGTeXVonhimdL+jwYfhazE7vjIMfe8GA3dQV/rwd8w9UC0WF8kDIjarz
1cNLa2AE5BIpQyzig78/lFhw04wjXZu4wy9x2EWquAtmEp5c3T8DjmVlUTB3th+lW2FsB02zUyje
x+YvD1RuYaOePIOhNX0xIlm+wGgm1zvUfdXjHMJKr2BuHnzre+EjINIe7OGLkb+z9rGK4frFwCVX
7BgDWJ+N3PeR9dgQxmfTVv2IzmwAs8trXH7cIIDaW28grkJoYh1S9n5nF6Sb/frRvPB8HAE+aP4p
QzCmQBZQbLWgusswno7fcoy9Ib6VclJL9FxtsSCDwYh7CD08FsITN0lKYlAWdhu1EM9xeLsCE+lQ
XImYhJVLltKZ31i8fJGAZRV0lp7Aj8ne2ewRb85IGyZk6mW0f6YyXFUwjZWIaJd9wsD6EwJHezo6
HK7sBavW7QjSiLKBqtPF77734immaebq86yrzUn4PiGz/+kaQH/MilDnYvJBK1ll36pNY34rVfM5
d+8YyfimPETq9LMapCr0nWO/781MQi6RZsjHTNQTgw6Zu2hmx0Y8ZfK04dB0XH9VH2i74guAXqAZ
0je6wvdHBWWDC/fXGdQ/yxCNUlHsdaNwrxSGW/7xjYc8cJrC1Kqk3R7KD9eRuJfwZJjzYb2zW3A0
EaymGOfvQJIsSuWGR6mk83XeteRmlQJG39bEw4eBT0xwLjivHyLusi/5IPVNdworMhIo8vi6Y9qH
CGW8M5UwKUDso1m1l8Qc53qUrfmtJbnd8C4PdBOcLu/VjNpy0Y+ikvQtXn3LwTHyPAUa/qvvukU+
9Oh6QHpkm3vbZy8TR8FOTZPhGFKXG7aIepTHY0dVlWXyipEY/Y6EEK42g0Ewv/DGS/qIu4Qz//W/
hJz+pBQKagxbDKBo4ILrTK3XbG4CKJCtdW69p5a22pLxK1wVKzvfB6cZ+OAzp7ySGq2fv4ZbevXz
NwBLXOCQvtFx95znlda9D9nuv2i2a3z+BOFrQlJKqMVWwrFFDdnVCILeS7L4l+5LWCaWIN+LEW6H
WmjmFOWKzkxoRaDnRJ7NvJlYNBdtDQNz6WbXHamoHnw3YsdQFtKixakAiugHUfl0kNfKI3R0WF6/
lgAn8pRP8L6V0myB/oJ5veE5Sje0ttcvkaeydXWheb23sS2SGGSMm/D6lPXGAX1i5MAwuYS9+Nvw
RC7kmqvZLd+4NVVzMZ/UBF2kJcG1/zVWaB+XVoWwHgSdFAVE806njmDi5GOzh8vkTXnq8KnbUfDJ
UETmixsCsm25Jdqa4UHLqNrCo/ANKs8hyLbgW5BlspCOsS5bkiPNVHapiZtNiLm1irPxJRjBO6E5
EsAewpW3ChTZ7kV18V+JT3MnvbWiLxWRKiAnyFeyaYYz2on7EakiDlT1m17gWelEOVUHOkFO2Bqe
wUq1bXJQPFFpCax7bormXEOFJAQfwejmyQUXHMCAdqqWti5nsOI6/qmKnWSy8J4CZ3AhYl6EJV6Q
NbwppGuJ9TbO/tRxdrJ0nlnA/vAcF+CudCZWe/YapDixA6W5zVU9lA3EE8hXkSzbOpJmmm39wBr9
S081ufTC8jDk/jPd6tXCeCTUcnHd5++QCH08BLHs630hMa5nmphEEOS/fWDA3H/CfDrT/0gae1ok
GwPJam3C9eqKlkprRd7Jz02ExzhEwVY32oFx+ug7Ik0ZPtOuGU0y5//EHg7nkhrR4plPRs0xqYJG
Ed3jJWPs7XE2fXiPui3KW8odX8d2Cp1ij7+AoQv8IAohZITJjC6c2V8u7pLh+aaVPTwmgbNpFJa0
skzUtmePrGIh7PShYMgXO8l84QgDmDqRW+mlh7gInECiOB8lK1HBwD9RrC8onktSzk8xIZgKjdzV
PRaM+dYR/1+9IllDa0ohwjyssGwdXdxqOcHf1fCi5Ksd4kea9OArdRQpbkc6vT6rXLAmmd5yt9sc
5SxJNkkqDdWipNfKL8sa8P2AtQKTttzBXvCEFVavW/MdqjmRjvkwybrRU9coCAaakuk7bZ2mWkok
SFTQdHPMLA1cD8PNS5ytBsf6QkBqtGS8cRQkyCPiUF1X/FzzgCqlorootjfxHlzrlIKvIAgubmoI
PbLgfs2PkT1z/a0sSp/wDmqyZTaKKARE7mYoH8VLBoZrzZpl+2DLIxmZGbubZofq03/zz6pyml3r
PL82IJJaVZ9JpeD3ZGtuTWQnroF6/yXPwmDntRKRaieTUlwrB3kbP7ZUUxTUB26KB8wQEdBydccG
MfmdjrPZF8T/IvI7CeAibdbd4xJ0oGhmvnGdrTvzx3rGJIJNS0SiaRl4A4UU/XOzij6cOHUJjQ7O
u0QGec4GhfSj26vL+EkwHokO7ZSULhW3Hyf80eN+DGyCDN2cZlPYlPygxcnyLWqK4Mckicsc8Dto
gFfBEfd0xBuePtfuy7i7PLKuL1CC7mLiKrDoEakFoY1S9DFsiPeXIV57Eo+5+MAdJbgNWaRsDprX
0R1mtrOZQoYYeJ0U+YRwB6+QR0AejsM41lBOpVSqp5X5dHyFAoUhgc5Dxm3CgqA/1Q6Axxd3FcXW
HiPUV65m87mRMLgWDDnGX+ablrBHaO2EoCpzEcERi/I/1tb2aJKW227T6D5X4tV5O8YM/LfEK6Ap
cFANE5AHcb8ACM+3o32adBOYkdm5g8Wgnr66BDYg6E/Jp9UzLCHrB2EyaRmojHa7/tlBrlThbOIp
i+xGAbalPRkWgr/baU4UxDjJg7jP5d5vxzDgs9vjFRluVqv2itC+sKTJKTZKxegXpkw7yTfmiJ6s
G5Y5rDuaAz462gvN9MMw7YW4smoCEExJLcZhNb4Zbkag9w0Y2p1v7wLyB/5ywbyxUANbZslnfWJR
jXvZgeKSRjF9Y42oOWvF5XIMeoQNEhJR7TbUyS8ba4YjtSWYDbqYADFNQdWZj8zUx8+joSpsLpaq
aiC9uodkEfCXdpcpy+hPbJng8AeatN0QxHjQGkDKBUiSfdfCYrlhJj2sKX6VIxoHiBfF1kb+flAb
SDTMbkEx08jYn05HfObWb4iPqZLWjEumYg36rtwoVs8dFiTvS0fd55A6rEGzVP+DioaAPf/2SQrG
l82yLthk7t01zjqXPkIObyVk7hfN6ywR052ZHyvQvZwNcN+C8ogYPPh26gihjztBWtrGZPToserK
V6t0un7J8oEeAAGju/+fD1h0xHCtTUmL0WEbfsrJ/H2PfZnQGqXJnsm5T+RtPp/tBhlZQBDTAxfD
RwhhhyZte1o4au+qLr4yTnQJdZAPGYkICi4P5iMiXyVD2o5CKOqZWUndyTGvaJTVkIQVuDpHLYZb
zVSwrleyozbBT7Se6BYXXsV4N2ud/1HG+MpJtQ2Y2KeMpGxg8ISkyJ14YyhaRSlyxmmnzNfRqUlD
wJWRMDjTqNBG3bBOb//9b+57UW+Wwp64UwXpATiirpWExwMJT6YtsA8jsT11U4n/5e0/N6xVDgBu
FEI5nbEevyKOPhhhUvfH8FQxiQQomJy0vafrIAPYUV7tncieQAbF4A8S+Do1aF+lpN+ZrLYEzeNg
0NGt7GmBAqv+KE5YLRzpLIAvES7xZWDqf0GCCiPBfAgLlQaaL6WRM1GgL2Q3oYZo7cee7DqzAm1V
T17mJ8vjpOq5wFP/TlfxfBYBCk9ZlGJOdkPRSQemXirbr4JNyMtiU69NH5I7n7WH3acmPIjDxwOO
7MeSHOVc8oA1q7sbjWRbj40OjYppB4hlKrrxaWRJHc0JbQHdfmZvqBDHWEOglAd5iL/wgVDtGAwW
K/IpxI5L9FkFRQf/GAvwZ1YSNk91rKScGD+p8vQP3cvKL4JrqbfveW/OIC/BYCwaIaIZbN1sznzs
cctkY7KCP9aYNbL9VIMuBoEBFuZi4pXRq/q3LpVIenpAhEaJZfkddPInhgAHdRE2R5WhVhRlA+lq
ev1K4t8OYW59b3y4SmvJrHyW/+Vb2wwAlx/ETihF2cUt0Rdp3NeB0E75AxwVluChDqwL3yOiVk3t
1agyePqOW/tlsslTrph7mNlh/P+EEXO+MWnxGfeVEbKxf+TN8ZV+1BHSjA1DEuizQd1J/HmwyLvM
vdSdFBdCFxui3V+K4ILnl3MWjzN8u+agL7uM57LuziK1O+PGeChDTKK76nsgvPVYhDm2CJipBh/k
x+pYa0bRFakiSNaHdhX742XuEOvtu0Xv/FYESWHERcP/es7nLqAwZSmvog14GxQBBML1m/QRYrkY
ACcfhlbvQnxQxre3EkKwbrxdJYRF+Rzq3g9a6/V5P8JuhkLheZVK8HEzGn6uTu/TyWwwxYMxVwVs
yl+nI+bOaeZ5mGy8zHz4+dE5JuP0oa0V/a///mloII9ccY0rRxyZIHgNOH+8sn0uW4WAK9Pj7z+0
UgfGzr+9syNbtDVCEY7jkxLunYIJ0EhKoT1wSRX4yPAGTkKDvP+P7PkA9LSPQq2CvgL8sYKqh+6R
jpYZvjiLi0Vvou44IZ0WSYlzltWtBwrirG/bRvzF6/VvfufCVKsOvvhIix0YSiVBUVjiUsaR07cT
tPSBbEhJSRCJ8XfbJrAn54E2s1pYWEbxDhg506cISICta5ddbgI2He2k0V99xTTA5LhBAUdy+6m1
EqxfNdV8Nmqab/ykXMqVz7iip3V+l8ALWs7iBlkwnoWGLJkz/j5RIScZcZMmwgy11Ai8ApnHvy0P
iPeG60pjkgbOTYdiHXAqdzUKyAHH+KMkuqCGOeNaiiZq0G4MCViAY31vv9DcsGBn+OtfdZDS6G+Y
X2EHr6IvCChTH46eG1IWdoYFBaUH7H0kuu4KM1UV87yaBWy1lYxfOauukn/eS7UrFgAixej7Z85S
qUpiw4KjWoNMNG42COy+tc/G7l3gtEYA8elvJArcJqTiA4tZnhnkDzyp3CNd2FgJ+nhY43uGruRg
URFgQsGfJwj5+k7sWEP8pdL/lHREctlZojwIOObBZUTDJgdcAxGB2h/dEV8uXhAwwsmaggDZkEPF
PcFHxlcMmfWWU9R8vgI1e36ch89Oyh2SYAPSSwP3QkstCevmiDG3+8zV6sS3WFVwVctfn5+ygEJ0
vIdDf7oZ1U1/XJTikmCXVLfb0PHsv3Xj6J1E2VQKmyiEzsGVrRW37OJOu49zHRGIRjoNIFDjZgr1
Qn5zfAsna2mjILqpg4rGFNBWEgPlht3zpS76qmjAJ6rl2PZIzoABuCEK43LBxTDUpCnl4ztBcqq4
DskfmHtWv2RzHZKFMduLnAjz+W6N1jJln3WipAE5lMbqYMJzRTJrJwYJcls8dskTiqdNq0GkwYbR
ONE0FT2DqwPJyaujJ3/98AQ+sVQgfOWOWenKqKXOYedKIzQHQ8ILmkPkCLH5AN3GgbNGxNyYsUER
PCquvi01uzKDRhpSZ4wIgpesWphKg2qz4aF4KTH1gL0W+2egshLto2hD7IcyS4g0PcKU8uvc2dfQ
szsJXO+9cjJJVDs3yI0CN6jxiXu9/EeeJ1OKJM+Qrt4ytvGmxjO+mIL46mAfcGexAF5X56a6QoQt
Yc6HRjQ8cWs+HAc+5Jb0iqFlzd9sqzyg/Y4IsyeBOzhkMsUiOWSWdN9l2zLHJnB+KuGl3wq0TmPj
ChuCTYeD183lbnmCUypcBIhmTbPDGkoUBoZAmkKP1jxdtVtsblz0F77cXuFkXDzsbv/0oxOMZkPQ
66ofSvsoxnkz9qLudCRuocRKn0dRtzpvJgIscCImz9IW793gHeLY8lk7i/7vxWqd0QfywTtDuwh2
mB56COQYqQd0yq4mLqO91PwST2nsE/1sEryxqFpaKDfuhHYGmQAtBcYnQQAjPX6juWNqcGhsq1wz
G3YEfHCIzNT9m2Su2IqFDPoOT/EGd/JIPIfQGqQIxKXFtgypgo0XUIWf/LXiYkqqC+RderHNO8le
wg49BEImqdACRWm2Je7MG0tapNA2DiWd0sOWIYn3ot4ZYY6wZNEHYoO2lRAHkuxa1FRdW30mXl/q
/xeNDRsGfHxyUruf5cGbuDCWW44zUIh4uqf5aQyUjhM2wFGAg/ouo7ocQHs0tcXHiGUr2DPwcni5
YwlBMlL8qOtRD9hBd+k2oaiQkkyv7C0jq/9Jv95SUQThJHwKlF+BNs47tvrnW/pTPNqH9eoUOpGp
STuHwb/mvVQyrbQ3thVQXuM+gtlOztfJsZaFkCzsYxDOeDTzNGbwaEi769dGmhvy1LBEnprKsfL1
55uBDiJ3LKIuQZsfZlMafED5QZ8JrS0IIg++segjSPkgQy+QFsWOiDgDSGzp7LTifOOPMS/7CLGb
BnJu+wrOUJ+agg3/CZPUn1NyImfMivRRi7htpE+HktMU093aA5NZPzTHXtl3qpT8ALltsCzd4loA
joylMbbaRG6vOhjs9Gc9oJvQ4cNwxMacvIdqh8q0gigT8ZRNujzJHIaIBBc8YIudAmHquLj2O98o
RSS4Bc9SIwuv4b0tLDaHGnchV6BHEXs77IcuTVn/6Fx7odd3sd0zDJ+KbSPDNWUafkC6+IhLf7vq
ZON20sJH4oQUw4y0xn0Eqjev0DRRghFdYuoOuofqn7oZbQtAzcUdmbvIAcNRofMbU67wi7Ds54YB
rmQPmrxV8WvCxWpzFQsJrGsi2w21sPad5ZmkyQrVF13DMnq2tNDf3jqf7I+2Cfa1sKszejuKG+Kp
AQvEC3CZ5NXQxYV68JGtj/zf9QB1anYjN/wQmazouFypZ39H//6sK5e/uDPPnvEPDgZcriqK7Pjd
jgYghPlRldxNwiOhiDxEoYDr0jOcc0owZR0+9MHt65/c0dyBYlWFbvnTnWhh7l/dAlr9Q43Kh1zl
c1QW65jIUyjZdfSapuKtXYkl0L3VAbmOj6s7uRkRE5znJVtYiRUjW99y7sM462+tnX4Xy0l3spGo
7beSGq0vb6EF7muaf1d30wPV1chXLhf/ml6+u6AU4GdEBKmc7L1g4rvly7lKJ8UvgiW0ZsUrSVSE
D8vzayFsxyudZrgEWUm4IrEGzesaOzsvOTXA1qvUTtVKP4e11SjpGYo+3MRZlwjL3x5BIo53GT+P
M2+3YiIC3UYJHY8HrW1F6IQDSONw1tm3pyKbb+3JBgwyPxA2ebmR6uqZ9e8YOymNOe+HLpfYti4K
TfPW9kybv3BAGzysa1zz5sSBWyzDpx3f220GQtNDmQr0p4TSqPmr1WDVaO8PQaYt0YnKxAjHZ0uD
fZ2EN9sjtpPu1X5GFmWlRvklRsw1pSSjOfsG2J2ADzHysLK71mOgkARf3VcmlOc1DMSZ1bB7gzdx
9DRxz0aoXsyUrvgvUcmoGef2z9tPhlQe7XOA5QbBKOrs0akjtngOB5A2KVblKbQguNaC2tQSjAfe
QDbRLtku4AWcH39YxbZsO6+X05Rny7GV+Eyrg2dRbagrsMsZ5E3W1lGwGMAYvQsHM6JBLajGbfQZ
kDm4T8eobh5G4MmKFvAkLeHkYH244tXWqLr+8Y9SqFLkQEsLNQcBSv//ZbHQegU0thVzAcK34ggc
dVgnuqdVJYhGXsCzV0cgHn0R4oMRs+ACbyjLXqCG8eb+ClvnEFzaxJRr53/zvgwyozAxt7aN5j6k
EaKECFIv5lhQ0LXryZEGVjNS9QxOMOliLNWdp80pwhlgbYh2fToxiMc+aIaMHii1sYLioX1seeEG
PpaQl+BiiIB4dxiXNo4RxURZPTAF9L9RsY6MgrRvmeSwvnsJY9YqtglDWm44GhHgPO54/w7J6x4s
91GcJqWruT1APQlPSLuEtqL5Nh53aR5GTmoxYqBFvvMfILVLH7yC/t6gw3yohamsoXM52YFuOiDo
fe0VVyhYSVfXWq2AavD0+9piNHt3uPNaZWX8IIIUOygKO0V+zZNnfCGfvotVx/5Mfix3M/GoBilt
zmKJZ5O2FRvPbC3OYyk+Opwg6Zqn6Grw+CR6SKc3NZJPUGap1+rec3XlvIBSZ34v9fIybeyNZ630
DkVEhJH7dmwWRNa9htmJiH/2NA3Kx8phZx+ZUzwqP8f9qeckoO81LsB3QX27tvs8pUgeLF449tcU
Aj2/vdIwTMQr9BF/OMjkyJarGvl3jqkh+QBihnkrghafQEEAToD0GD56EYz92QXrvZWhebbDeePE
wE1sV7LGX+vmCyABZ27JOlb/O5w9k9Lc/8VIW4ySSKBPAWH+32uBNIKc33UYIori6V7n5Vmrws9v
HS9vT00uu1myC7BoxIdXEYlftLMQLbOp+x2f/Iuknzp9NzgQx/pxXbbRQCigqkWj9E0pSHCLjAmI
mH3xj6huK2kglLdHVLCJ0qFeZjZ6X7KjCRQ2TkmdzPRHZLxxsvUnzgDuNC0ZZIKFP4eMz9JrxbiE
6/k5oZREPjx+wYbkZA6v55dJGOqbIsn6JYcq7RWPT5c94iCx9SrcjFxK5rnkVjzc15WI85t4SW6C
blpCF/CzBbZ3OY307EJyliAPyYZB8OWVgs9qjH/JHwXpoTtFDPnHdjOgj4qim/7xfVt10dQJySt9
GrQ1SfU6kXUPoWgABl4ujbtBRhYKOxHbH3VGf6tSZ9plFj9g5qVv+59UVPd3gyp2Rv7l7oKp0uV/
dCQ/ewVwVZOyzDjhP3GDM+MiySLboLU8IUsErUt66kmcErpblWvkemtMiopstz88fZIq07uSqOqz
bX2fVOvWwf3tKbeqjQ/4GWE0WhRfZY2h8FlIhhNaWMRUAbt4aDTTMlOOPkU+8cPQlAohRtFHNLWa
hcDOdcnmHNWP1QGcyT05blrWgRQKXHn6ZsMxo+5tQ5zlrN3Q39QEs5d/CELgeGoDitUx1SFndLop
g8x5gDBs3JnIJbK+oxpwdKZF+ZSEmNt3yr1CsBByHJQHSKrdQ/7ydFTRheayRo8gRtkkIZJL4/Or
c9HuZrykeeHKhtPPbGdguCPFnme5OaKpzPWIyWw8iUdsdltc6pBz2/KZFzb0ZMiouNoUUjvGVx+e
pN6U0BuS6LDuyk9SZPDXMUW2n3k/+lffTgkck60RTmUKw0mKwmuaGYdLcjZoG3xhuG3+N7TjAW55
ayO5Vb7U+FXGpAoXTn/JywUwEjO91KuwDiviR6cX8wtMAz5TZscyL6xnQ/+xGE3PNPhGcRN7TnJJ
AopqbGh4vv2mZTAGqM/GXupBsnKu/b1/6+ecqghvg9FFLNCaDoljkjwyKORXjhiYRoQ0COeHYIE+
FpippagyaRizynZExdJoL2uUZBs/UgWo0Iz9Ubo9x5tRC92dJgQ2/eTX9QXLOOGP32U0HZejRLyi
0w4YhjqCPa0gsCMw1gJkJgVh7hFLZz0E0mytvVEhgeA2u7quOBBy8gtujl7JuAoNt4kdSsut1b4z
h/dAgpg0neOL+oS9BAlEUsizG9jIKdBIWB3RxXNEMZ6Mx2TyOp76kOodH7ZOVFnZQhBBWFmD6SpI
+AxYbELoEpqmIhQlsGWWnkNzlCrdrrZx41GV5H84EAADPA2agEMkb2yKIXS7iOAbtJr+kSqkMaaj
8jzESKMCEtvNSDAERoeMyrKcIHSkQWM/fZyOIVeuPPB9VIGQYQqo2Dsu4rWHKLGqY6P8pN5fycGI
HLfE+66TQBXm8SZEn8YDHDMIvu8H3x6VdYyCn0IVL44BK14/HT/FX9V4z9BQADy8al4TcFID6KnP
fT5AV2hbnRw2UYdidlNwSIi0oWwjD+wX9I/CRQ68YQtpIkFCBhysk1amXZyMaUVltIqyinM4FHhd
KQYHIe7eFkBzMPulumTlh3I+73UxUIc3F1N5/JyRpg8OizcA2d+kAzDeVsGHqkUVH6vBhJ8ADOt+
YcgQq7SzgFy8zUbPxvBDEEpTjQEwSXR/kJZHW8h5r2a8j4Yaj8VrAi/eaKJ0YZneNAWrBaYXJBiE
A3lUGP7yCjh+LxeJNkgWiT+zHKcbaez/E2PnllevD853/9WsvtBKAmT1xGT9k1fE+gGgUTngy7wf
baMBjb0nE2WuGaFXhuSBQBLbCwHGNOHSn4QfPjrDUkOjob/Ws6L2CmJbGzuHcgpQUp5cjuDQgf6a
G24KVzxU6L3Ew2L2u5eS10E5N7AiE1/DuyiZIhJUaP8YyAMuJXYxgR9pWb5bnbsQ0pQM+XLXrYNw
KNFlCG/srdPtpF0acS5YqnahRb7XB9rze+QvpNpk66Y7bPb05vhg08p1mywyI9CM+p9NCLV4o8L/
C2XciTgESH8THJqR5IQmCiiy+CXZC6Ts/h39gb9QKF0W6gTCRVmdiHT/i4KZtI5TXjLZSUtut7s9
FAOc72qD28SRqScYeIihvMqnm7Yrv1fux0CyOM3HrszxVT4cvpZgCU1JAj5y7N3Omqd/bPrlbzdr
1j9AypABF8nn8BiolTv8VVWnS7IC4gdEGlOqgm1gbpadCbF5jRcsVc84fKfuXSyfUlb2YEuzwk11
ud7o4vpMrfrLxh0KzAoBg690f0rT2AO7L6MsQZwxEXd6J4gZZ5Km0aV/udOTKLGr17lqqOy8MQQc
EVcVhrEH6gBVAT3SGPvxPiyDd2CQFJvULdM4DfKMJFJVORtoGm2VGEAXgTa+KM9a7yauVpPMYXjJ
3FUFjFlwnQiWNOd6Abm5RmBHBtXYjXniTBjxh7GxCi3HwhM25bPH1s4YSSd5fDPelTo99UjWqE2k
7GPNEKmAYAAOdFcCXF56wW6i+0+LnUykX8U5jtT7T14jfzbJXEv4UyWLzltl9GNNpYUL7IHrPB0/
vjoatVXr/mKv2tl9I+whMK1s8+skAhmLomi7NLjY2wsCyri/CSlyinwL82D0+4bZj6ElpnBE8vjf
oLYVVy0zlBgYnvfZqSIScMPmMCD0jA3oBYFGrhzEiJSyE0GOOCy/8UN+aaj4TRw7NRYe+4m5JRga
/PvkZ1LcsYx8avBG612x418GpaeG5TjBO250go9gDmt04vtNLcSQ3ZXHbRvgnvMkGLhB+ujy1oi7
PYxzKuPvt6u667BqbL2LCZAXWBgiKGFhAGAz31hC/cyebdsNQ6MYXfTbG1HwZwGfsz7KuLxiJoOB
Gk7gqDHQJztD2pwEO2YPAC05s6WN5dADwjKubRM0TJpl/0MAnsFBgaoa5I5aikKvFUSsosq7a1g+
KNsT5C6t5oNrGmhYNVOIqMTpELBHfg+KsYy92ccEB7Pe6NF0bbWAVox2+GjFM9cnTgoBY7OkR5ww
c1av5lhYaFNwq0xjdMzPeH2kmIMn+gsFbb8cUvgTMHi8/9PuHIhWnzz8D2im8qS7hB8xiW690PJ2
JhIsCRDRV94Bw0gAE89OB4EV7T1dLWj2XRNEvK+kbgCfIcUwCcy7W/ESE64qsnKUlS6/OEPyxKAS
mTcZMVpiiF0HDbYtx5/7YUrVeWXwUazpvlLyLGkHjg8v0Kzm86XbcOoIE7grihZkpdeyUjUWFQKz
5CBRHGprRq28Z98vrHR36tAl7QyqK2ZiovL7r8z8Xd7TkI6fcZkIwxlK40CXVr5vB1p3IatDykND
ifaY3dcdQYC+YeMgUOwefuwq3S9XyceDYt3OtQlBIFcSTctJSOTmw+T7srU+7sOP9+zySo6CS9RQ
KUQl4yRJ0aF+1iLTR+qDK9ZbTO032loO9QaN423/uaskLIltGQyQm+J7r2qFb7nqMTlm0fxJSZKN
QDt1HbaWHiNLoRAvKyi+SwePck9uHbTCMSEzDxb6IQKvxdU1XUf2MIl/pElH5h/Ct7t1H2NxtXEK
vFoI3jdLfDKGIS+4gFMPnXFs04AnbQA/qG0fGzyAEvjbr2ATIcHN2UeGt6VRqHIlBTCEA1YYBFX+
shs0KprMIuEUqwqL8fkcTrDVz5bBhIWNZgzprCJNdTg6dktyK07fpb07WyKPtdH8sWCohZzkk/bW
RQqUWzCd7JUfErrTh09tEvV+77LcS02DdlVoV+EQ97CTDK7pMmO5vz5sqcbySBWmgq94NVafRR7R
kpdNYPpCJMzCV+xhTm9I7VjurEOunlGp4V1Fk2ntDPAnPJR7K8bJrzJD6HomoxniVNeAshn1/VA7
RwdGMC8kfown9B6XtnRSmS54n8iOur2EoN/lIr+NM4cE43c5PqZYtxDFpoeovMKeAxGO/k2qcC1T
76DU1JpARa9FVQ1LaE8Z0/w38dNwiDT6F8qdQ6f4fKAyzrppvFXdAAcvZG+e1yClUKyt+nB1aHV9
qLJWhfEEotAgT/7gQ4NwpDEFnt3XmyDUDvkrdWuEQX3TnmrSdtJlnupIi5ITky5R6NggnjJ5mFIF
Qqgp7PvrPrCVGBHjRuOBK0M0x3FmiBmwlfMXz50ERtSti3JQE/CVgzH5zCGQQJlwJB149gFsun07
Mwx5BR9MosDM1WHGngyUWPkTTrGXOGoSCuUxOmMHzMWssDX27xnDCWnrMA7SqU/qZz8zSpKsBRwh
yFQ0fW3NavdM7YpoeQkk28hlp32VHtKdUmLaPD9wMYXj5Av1p06r+nRX/51N5hz/4ZFareJ+lLA7
G0kBC14hYYXw8lPTe1bk9vYwRWIA5J2hVOzP6n6fwn3l4jdlgkRHnxxBoplpPu/ZAyK8hvVMwyd5
HoaFbTNa9m6Y9z/waYFKSgofqdS3eXueI2HdTA+3FNiRvPX5HASVM2uzOKe5C/PmVeFr0KV16eFb
IxLRfMqvTtbkS9bkuf9unYqE0anXtsMPFE2apzI+/h6jNEyKQhhYZbTzyO8OkvMODNxZaV4/IFnT
huQOGqYtxrlr3pVbLhrBu5JIoCq12IBtAc1lwYUq5Y4yiJSKg0JaPncWysvJojWDl3nEByzOUwi2
alXAa3TCozVOTNRr5+3r/18ezSfakcKFtUSZ694jsp8cJRr4WciRdJus/N+KKuojKQ/4HxmiUvea
lsi8nRdbsm9EhjEkHRCHXmM/iT5YxAmdwz3oVWq8VndLhzSNnW5XROCglpEMOBntlHzIvEuMK0G/
Sd5wLMtynn4t3ZDaGkH1R/EHrbAvKAHiwqtRsKX+HdLCkm4MjnKso2inkLmJ2/NL4GYIaoZppkPL
5OMwqUV98sV42yv4nwiaTVwAQGbTUVcyWaNDieYXo7dlknAZu+tiNIX0Z18fW3Qx3dHWUWu6fIWs
M6GSxPUmOt3YaGsEVj7ens+iDJSizS2IVL//5JDHsdhTbeOMtuEVdqecKvYYnBTsODGCmtoaSdG5
xRyuR9OYkxe/qUMBrniijEnQI/ooWMgPLJ0W57vmTxREHDYrT/0pY0Q/qwhr2TPvcjrFagJi0ew6
7DEmNeeSnembSJm8ZW/UpyHrUtcISnUxtHBY5J6rNbtl5sogfQt4AU48iePt6RVpKpmcyLLu4aVw
p4HomgfLfF1Tmf1HbN0+531kJzrUPGkfoW9vyLYsNVAkc8ct51GyDanUoS0Yg2AFSSPbu/c/Zl/8
iwKZBB/ag8RWFbhBitqX65eoExnrZs00erhqhdYK4DZhf7wfxL13uQ2qDKWRNpil0JYAgt8tsEmH
4fxPK/M2sIVYuzoyv1bq/TDpjO4vl+cnFYtN3V0CG18LYa8hfS464YmylnkfG8wtiDEr9iNl1STj
8inYZl0bhfIR4waHDnrwvx+GG8pngYmehugStlH/5uAd/+YlAzEJL8g4OFi7XXq9CCpHyq3N4vG7
tbt44ZASoON9bFypb7Fy4Swk+m+4pVi4jQkIZEF4x8hKNkFOQUdcXN+MwSTHE8TFO3r9eUQyCSAo
pIqYapoDrq20LQXb8KyIA1OKmTF5vqd2ZZsvioZkrwTW7QcBkwSjqXotZF0DwMXcRXbfwD835NSa
KkdEdhyGq+cf3xyRiqe2i42bIKwxMdUm1WPRW0cfUYBRvBWYn+AZpfRPdTKawx81/GsXUPv2XoZs
JW5BKdoW56MDeYOwe3Ef59bzs7BhPAqRYK/p+dT9OjyAAtB8uTDGck1i7o6reazIyMHd4GEDD2m6
8oUpDabvDqdrwJFID22QQCZNj9D112HiC2vA9M2NxM1Lvk8bBtBxmMX1uax1iwQk6QSHGi+Z2C3t
HNj9M/200EKm3xgC33ENUxnuHLW/hBlllpF2QANO+ZlUGXtIU1EGSzjxEtDL3wSlnV3V9KeDO0uv
S699eawEfsLIm4nWUdFEL2wDNwEbnnGtlR7fylMFUn4kbrhvx6WDLnKBYh+uj32KE0t5QdReLNsD
IYhvIF/KvTxnsT9t0RRX1KMncxvkVIED0dTy5yb2EkUbJBVYhJVrH08hulLwGKqKgGhgdvfuAMsT
nadYJvkOIg2zW91Ak86Bi14CSdqdTJWmbNuIUvLloAuinqybj1GKCBW0i/ovIp+xhzkrhINdYep3
SpgDt5wOUzcZ0bLgmzXtQHSqmZeGN2ySzpAuo8SK47sCwdPurb9/q7u6klUgcT31XRzlz3d25OrU
lJBe0soptTPxECApEF0rT8N8ndK3BRUrs/2GD4TLY5EMZ46vqr/a4hdJE7vWDPffEyyUuO0k8Xm3
WmOpl22cmIRNPsfHimtiIdLzZv+vK7nkqAiROAAaBSjoaPIuJUc57FffapxOHFP9oPgpOZrqCqbd
19si69SlFrzfHvXsj2cPbpJ+MwZnMYUjkkAzN0V3d3IkEuenZss8/16blN/wdmzIVSKxhsplIE8F
zjkhSJlTZV2CwstX9SARU7i37jN7D4qBkWy5Yporf5H43gl52XO11sVOyj9Ge407lTwXOY6nGwoC
22S/DAefljiRcxai2xiZDYh+zrgSRYlckOJfBQ2e99uMjSaVaVGObcewPfBug4Z3MtiJATy+9KAC
3xS4RxIuhvK1xm4phpw+MtEKVhEBzj+R7CUiUtFITKmE8hS4cqQG2ThYXakGinsSbBdaW/5bkpy8
l7AkZjzvvy37vRKWpKscfrC39F252qSZOvgoyDeJeuqRwhvDOA3FIllprle39tB6cwrpzvl4f4C1
R9HeQAm/xeSo/sokcV6UBB+SP/X+K1XgjlDa5x0nFdQvv3F+CfjzHWT6blxLhZNwoQo93s4DzkyM
8LtJjpv2Qz5d+M8qIgfzLqloJnh/Dvjr/f0vtxxLnnYaYLWaxqeJbJn9o0QjlJorvylZFwSl4VRU
ZsbeQRpzh153oilI3T+kLyxuPzOBUfW2drGBo1XtqdQRvgAK82ZHWjFm/45BznX3Hiy5aL0eLuXB
rK+62pFqHzop6PQwtAtwg/hgrT5vCBHgMi71yEkLuQI3ilZKDz+uWfAR5pknOfLd7VA8sJJq77DM
YDWpxPNTn5wkNc06eytou+wu4Vk8mKsypG1xh7WStUwCXsA2TrAjDbuOCAhjpVazBhPlLMk2zfOs
h+6eYXroVINgH3TzqtpMDbs6EzVnWgFEal+zNt5GfKUCLea3fXZpnR6Oqwj3jnytMTE+qZmzDawT
/fyxX70sADeGu/2QnkgCQFG+g3octElrQOP94xZR9Enu59INhHzK1pKnesV50G+5daBcHjFRZiWr
bU7RUjM79CytVULXiKOWLPkWfKZQi/DB9PRzc8JShMA5Kw9rrsZnMcy88HxSYSWZuvGM4skZlNWb
ChGtx7hlqE7aQksYIas2Nrt+1XcOcvuIg5zAohFnqU5TX4uS567i777gtQoONxMHZkmz/AC3oz5g
aOKw0nKEPoFtWm9tfzIT3hvtQ38LMarEZOFciVTTjw/RtBS02gxnyWVl1Naq3cz4dUV8tOKt8q7B
1wk7wwg98eWVVxLoLIwt8UjRVCKkxfZERI41KAze7gQadjUe1tsDJZ80J8XCbtD5YUz10HM13X7f
tBspQBbBlXP53HrDpEDnvPF5L/1Hl3uYBJ+9m8dWUkZM3EEbXA90L98JL3j7b6SCIWdT9C8v3TNy
N2Ompsmr/Z1P2E3kbJZPu4m0BIeJYRoG6OndPw/doyCt4dwD9ugo1fm/PkhfshoDWODMNumKiPZ4
lrZ/dS1AB2ZdSF6iA2bG9FBAUJIXqaxCZ1Jz/zE8q+rA/sN8q4Ews/UqqkYCeznSQml2Bx9O7zPY
QiLc0Zh1s37Xfw/WNAjjgSyVnzeQC4OF8kwAV6t7G5OjAlmdrrX6y6XevUmNpiEVf46522UgPGiS
IFp7JDKMjh61u6XPl5pc9w/G8TkfgTdtx12HUc5uHwbOhCFao/WNBfMwEnTM0sJwVP2N0mqMp0jY
wpqYxybbSi485NTmWtg+NHOKgXOQqlzq8Bhk3X9EamwJg88B/EWlIH5anPz/mSkJ9+xOBhQAqP3h
YCBTT40LOWv0BdeBfW9TclFPHHBo7nYd84K8Is7F3TtCjsr7rMlvxyXqI5L0gLqEFGAqyqDfib9r
xKcywB9FmFSnF0r0LyRuORNu+8wRcl6qPzQWEuOX7NPLM6lfHaRGRqqEGRQw99SffLPOZLG4DZvR
uzNcyPaQ28TRZ1wiF3MIyozYfvEKdJhvHYc1sYntSDhNRBDbH9gIQYcUppFSIXZwFgjN2Ayec4J6
grHdAl3+2C8kMQIdsu7p0lGPdqEnic3qDZwHTDxEdXDhZ77j0ymGNhWZzlQuEojJXOMq4oEjQ7kQ
oi1xZd1aQze/cP3jrKBlJdNoBsVdv05tu/NytZLdmXR1eHclmaKbVnV64vOHoS/1GJjJuQ4i1dYh
m3esTz6+x26lE7LqZ5UjiknagRdl4+b7tkGpIpxMnnvyg7qKiOCrtjbTODFkinfvm77RSBWPvj7i
6BWnIcwB09NcuPb0AUw2xNfafXQmOELMgzSHg3z3p6gn2WUXXjQYfjngz2rt5CVF9yQcdg9O8uME
yI3zNxricaxIGK33bB6DzY2LZUWltNk432p9DskINjHEXZdru1aUe33SB5SQH1iFUPQDAnIOHPXE
iL4f/ZkkIXnMlKfSaQY8Xh5l1ojOUrOkoYtKdvB1hoPjbfH0PEs7lGrFAazGLzZThJgFWdiGoUEF
7t3wj1oEr51uQ53jOJ5iH8JC3XmznBTIj04fX/EoHd8vjJCmRcCneTPTEppZPhSGb3D3lE9i3r3z
heddP6cwrboGIBsECn7/075jjRuMluZ1UAPPK8Py19Ath2NxrCz8T2fTX8QPT9ut69nfTQhlTkRF
SnuAP8q1JhnYepNILyTVfEJvOmYLZW7OkSqO64NXek1I1NaHJaR73R458mOeHhfMEn1vI5R85A8z
RtMJaINdCaWkhXUb2AyFxNupRAfSVPo2A7MiD6K56REljSH+PFatHvynU17eR92M8J/lAQMCMnA7
Gdr4NNMjRD6Ug2p+3mJZvBaPflNEPoqB65qa3gtpKB09tlqJ3aWue+punQP9DLGfIg1Rx4jkV4p0
+vpJvfVNiyet5yJJqOeOYWOGiU7lV717Oqlt02bacxWJfDcyZfAhN8qnJCILXGq3t4rBs0MRwoXz
yuo40+Yr1YATZ6qSnxU3Vt5s09SSJMucpMLLqWYIcHQ4q/RQ+Oak1/tELP9lCPvZ3zQBwm+MbGAq
ZnhH3GfzgaSKSAUBeLfLV0pc0dvcgeamoZ91SJY5W8CzhanR/mtM+/wrqREp3iumBYIGuyy2ArVB
rrcHPTULOA3T6/as1AGKNNh5ytqzLzqa3oxIkFEQY+KFDoBPztLyoEBvjo3lFFej/SEik8MAlq/Q
tHpdcVxti7hInLWeN9+c/SbPqBBYijYpIJgCyfH2lxW0jam9LTOO/FXGAiRNUYCLExtTiAIIqjZA
U26x/iQry+w9t1eBqmEafuWlWwGFMEm956z559yi6WqebTFioMf54AeTRp01ADmjOSq+H0uotY80
uD1yeMLQavVl3fq+nU+XSCdWKhL+J+DNnMgJRNLYsvsPhApDFMvSyQb3IQ6LBhTntNqvo/LexxPt
MkR8q4d3/8QgxcDJtbvgtE/WX9L3S7GgcG9wt+KzoIR2F9IT8jL5oEJElDxKOefsKUoPC/5IWTwH
0RAvFgBTA+JoLfFRfiVvgm5TUZxpeg9oG8uRHduEGKL+NW79IiNKXNh8zQ0nzuSQarO/j/GOZeMT
eEgU33V3UtnhVqATyNPcwqo5RzqPmutg/Y+mlEqjqVGUIcO62rrUI4opTB/zrqdL1Qii39/MT5kE
gA9N0jLqMc+wWgSE6uhUe59NBGvnLU4vopXh/VBCvgPvbygtjF8o/1jePS1Ed4gKhiYGVj0m3K4d
FXC7FJ+fj8M0UKJu5o9v8Ib+g5depaQjdsKyWXSGKabiPfQF7RrTXh0UxScU0Veuih3DtwUbtYHp
E+B6cffUQXZZ+xwaEexxZ1W2qu++iXKafudM3ZwDkaoOLNJj7q8Ym/JV2u4DH2nKmqBRakJsx1Lc
Wf7b0mZjxglZSCyKD5Z9z3araKfynsu9twQ1NMWxSFhIGw6CWJSvEH2WeBDotAjTNnDGy5vTSKLg
QIAjac84yPcz9C7w+JJ1YPfZF1sX52N7uJm0gK7ro2wmzCbY4vlSVKDYmpD+2ukbN8VZCBmBoaqA
3Q2eB+v57SLw3JZj0xnxFxpmKZ7g3oGI/wiJb2q/gt2pGMX6h+kSYJNeq2nXEwvF3RS8jAu4jTfX
eEzisK1cOVGh9qRMNhY0ED3hT5ctRCPlZa8R8iN4vWZ245BHDbLtkum+RcwUlv1h2jtcSJhOY8n5
F17hwcQ0IX2htG+h+1lc9WRN/x5VzyVedVAzEOJScJ4FcbDsXwikf8oDCW7GixVAsr9d4WfJUGFt
jMRgh+q6NOAzKpqmQFaGKRqs1ovVpM2fvxSNDgw/sczHNhOyzNnea7/Wqcsjl4FhFwXooaDJW/CS
iSBxzk0YttbwMTCCW5AfyuQkzEdP69EanqgKmg49MeKQfPIRTzcBeCQ96IE22OjV7eQ1SRJAdM1i
mZ6DrmITwPrRcAC1qw6k2AhavVVqevJhMcuNCaYjq3P8iPoQ2k8RvdoEAy/oHTXNslt72iDQhdTw
mrjH47kIoUgwbnMvLtgN+UbQFSl4/owe9AiBijb0xETCcllDW6cvGnVbwImcuG6znVPOdNQrj2oZ
A+i8Hnp/Us4+0NJqaXKIOWu3VeRB6CE+M10OvxDlFoEXolCYXVPTMvbxrIE94f3c7qkygtpxfK5e
OrMUOL3aKtEtqJlqtpl6qrB1jCb063fiM65MHeFYu4GRQSjJ3QBc/VAo7tA3RMDV+bM1Bf9SYXn9
tm0XsU0v86l5GmnmRySNY+8nc2CItzp5KVtqmk9XJtKrV17hatSQAH7zpOjcMvJo0Qr001tXDKql
9Mfi9XVRDXwwdP5Bn1jNUSSLh815E/sUJNzezQPK8t2Q5Z5cMiBetlGMbuC4xzUKzlzLHCVSeqgA
b2wgqtn/Yofc0IVNVSDfme8HGxcvvIoWST3vZkUd6l026SFH03zw06Tt2HKRoa5yKE7pjwJCXPwx
H8pHo3B2/tLdbSJAeMMxK6mjoYtC42t4gXNR9Id0dp7MASAxAauRSMAw+2wSgUeqbp4aqEoBlzsM
mF6qEWQk9SGs5/LN7iPGOSd8103/JjOdmcT8mDYRhl1j1AiWpk/qrJexQfh5C7Ja2dIXKrBlEMX+
jY8cENvY3Xul0TkRVhhKn2tD234lxMNevNcRruoUVv5UfO5wvuH1OKv2omT4X7eZI0KxNhKqJpDo
wLDRNITrfbnkhJgdY/3uB/xCpaKBIt1HRxvBChcNzXTR127lIPKuVM4Zig+++N59X5JWidhywuqs
q+qG8NNBPNVDxkjnlX3VwPl8SQ+RfAzZpgmdP/pWHcKPdchhTGAm26gKs2C5K6XxrgHCDUf57lk+
LAtKl2kHT0nMxNp1hmHItH8V0HePezE07ssX3bByN+/lZYV6Y68uv3NK6wSYzxozUsrKE5SuV8kJ
7ldT0/Pqhmze8yfT13eBSbkqNlxfkhGqowNqUF1xEm61NDRj9JHT7/dAstYiADsbV1IibCmVn1X2
P0sEkVKEvtUqSJIiXNhW3+bdHOCLcVVcAqNdHLccGTWuGb52RaHVct3vvsT8t8FCVGPsHVP4UBml
XZuzxl/Kl6bXu68V3WOBzFy0CMQbhZRsHAkQPL/mbf4KEAnUFALerLnAx8qYDzv0vMxWGWfyG9Zy
drLK8rcWm2GJBMz3MVBSvwXPw5XE+7k/HGeqVt1UpUm7tcN/XjVw8Rjj6QAjizbJWPC/XSnMoszE
M4louHjZIq24tApAGtAdVDaX3g90flOzjsqCXIjTunGv7smDf5W2Uj+A9axSZn9bge6Gzfi/IFoW
oB2aWJlEMmBE4mU6DUordG4/mx7zI8ltACelrgoetRr2zzHGbHDNmFJAHcmBfcxQB7zC2XAQFbC0
90C6swbfIgpVNanGt3Ldvr6HUuYEkO8UgkNRGph8t0cAhZ2Mtb+fkoE7c+hWKUALHvCg9DiYjI10
H5kMrUK/4ahP5UsdV7nL+Z86r/TE39NojP8Q8SXGDxr8nkWzUvWnF2zlzzDON5z+6Q48Je1aTsv1
s5o2xfgmyitaNSoJpnrVSpyEcsZtbGs9ca12RIy/edYWM3JZZopDf7X7pu7TEf4I82mygt2EnR7n
9gI1AyYMSVXqlW9rJPDsA8oj0d7gA8rRXk63VALRQKMntLwAQ0W4a5HbU/i5w9cVnELT3cXMIXLt
9fqhENDijywKyR78q6W4la52A6w8Y0zskZ/Irf2TgIiz94OVB5qwseMFoCxl0qV+0VrXpDYS8FJX
8aOJgvE+EhJZ9cbf7k3TJQW8ZxLO/XWgkDQ7JRsyfNtZ+Vu2LKmZzEPrwScszVc7gRhdONio0fcF
dm+rB1s38T10/mu2g1NsrrAzckjk3iDdhUqwYHnDZ3HEJGmHRgRY9De2wV7PAQ7NfC4H4irgOxV0
yShhWdy6mjpZPF6Pc/QZaBZh3LGdK9MYlUp20n9twh44Ul5UZk0F74iapmotwKqsQ/N+GMEscORt
uPRhrLisC1M91F6q6T4IbECmPPycWt2by2Fz4psBoFUr/unaHS72nKlbGFTO7PnafVYrLLeb8E1U
1ox1kTj1ofnyvNE1TxpIEIv1uxvXcbsIDV6awvEA5TqGwZ4wdRlq9Xxtx0+6EqNFTIEX1lhwEyUG
s27DlVaHPkYpHdptCVPsDByNQa+Dr/B9lcJ6bRJzcHxZCPP57YsftP6QH368EXY8ZNnxjbsbMOLD
Oby1JpHDmKKS/kupXtAPOYdBCgE1gQ5wbRlbSx00Tr+UFCD35vQ3YT3SWTIu3ax1H0uRD4Yv2OP5
YUHUWgKv2FRTLvSP3qAvYxDvZC2VJOZKU4AVAE8II3QjzFtR0L3gMaGO7AxnBunW2O2rZzdWHFA1
Y25nkWdGG6VSa6+4asF7Y5/GaEQOFMJiJJKgdqJgULENvVcwv53o8r85SFM0XUmwsTUsSXTg1DIK
DJb7VYW6rmfLsVLNs/UwUPp3sg0HQqD6ywnPq7bVu0L0gJZwF9BlFv15vFapSB0PSa6VAP0Voj8N
s/cERZIgaX4tM9Jw1oaXtuqVGQ2n8t3pkS2MCCsI1XRnxQT923+yKp45vcp0zKFiIKMwcN5wZ4rn
hN2ieYFbayifeJ21pvhQEDuse+Pcz9e4ChHW/6htDyPqtIh8jAucBsDfFdhMbvYHgf16g0raJ5Wg
GIhKlbnWFSAG4/DfJzTmDYP8ToHc1aHy/+EptoEwaTeFE3fF+b4XtX4vU6DmsD9shwOaNwVnJkfn
Dcg3rjROZ5GlmmFCIsAXJ0A0kJSRboo4iH3d2dYjxi81XyHBb2eH2NC8oyPitspqo8xCsAoM3i7J
cokqhe8wioX+oPX21hyKiFpqpHvc5Mitnh4IW8CU9v88Brq0x423LW6BCHEI0T9e6MfroHq8287Z
ftOOKPeIv/iHa2/RR+KRzSVcL/wlyJXwwmxZ8d7AHrHpKiphTKkxYS4qlyvtcAnJIpSUJC/AqcgV
NGbBm4NsoBitVQAFhW18ooi2cVg3Pv3n+Ak7yLfcqYFxUxfSqivUAbaKztmogXOt+6/GadCHVtiu
7bojPzyd7ZzZg2PGBOv94f0Na3VMRakg4xUHusx+CWI4RG8foO0lcB495qLdgwWxzv2yXwdVAsGt
p3n6pL+YKmrYFo0752flZgqwl0nlUd7iTIylF4KuzBXurE/KpwdEoTYgeuAhbWYzn8BOZUQDKyoi
UnNHXNa3hI6BNfO2jlFzYZtrYq165FfktHTDHnvROG5fEHI2ji+0/E01CKY5yfEdlEe6w3QVD+f/
aDPDTns9sKjPZoLqi33M6Q1wIGSJ/rjr3FquaESJBk5Aqj3HZaAIuoIyj/WKgUe0nuf9AtkIBIug
kwOz0nQMk+l2eASPOUMmbdoxnFwaGvxKYLrzusQjupozb970u1eacglYh2LGyLn/SKTEFZ8vquOo
RfVK4rkj+Ysf23zffsf20aCdEylmGrtZljUU2zkH/uw/3zwA8+0v81CdgI6rreQ0ZuMuckj2Stwz
f+vXagmkcKhFtcMiYnVziseqOCXkrIBBoeC1Upf7Y1dIVqroU0XnCzUavDW5mCAZ3to5lnRmLLYP
FHyOXZxK6jpP3Jjbjtlx4oXzXhguzHWKTxez+BDIrfqE3dHLZQGT0notFzkWDIredw9ybmnNjMOE
sdqvBH1Wd24ym35zAm9JU+0PM6bDAa+gITcvg69T/8jMn//dQEmh75dHcWqr5zBmhljtj4uaNbA7
lYMGYn6whREdyt/9G1tDOtRY5fx1ed5BSO3bNuXeNBSjRT7R/31tSHI7XgUiD5+9hSeZfRxFWVOk
seQkS5mvN3k9lO+g4EPcNx4EPw7tov/u1tr0D7oD96OmDa3hAsps5rGDju0ldC+3ya9dykA+tD9x
0iJ1qjFbc3u9TEn2aOvDf1n3F79b/zj84zggYc1vorSuxbVKpSzkfjv94MlEybEvBi05k7X2frLg
t2zYTC/qYMUmVWruX/MPq/Ug5V6IFKxNRWbcqjhWD5hdNm4Q7/8VhFHeXkcSQRKaIg4qE5tImz5s
s6DXg5WEhZF2tcY/E8xz/vb2A0cc33qwOGkaMzVJHirovpRWhCKkOCSPNQng+k9i0haj44fbJ/OT
qDOT8ILBFN6cpVfZP5F0DRnxa7FcAISnIJzJPaso7wP9t9ac1viSHxBAvjttoaLW3j7DQneaq/93
3dekuOf3es2EmKM3A40oSc+7N7glD7vd2yEC75RVJMUGRY2zX1/oHtUTnEl+vgTTFlbmAm9WZmL7
RDlYGNgr3RP04w9TgPJrfD/G9+uwcvj9T3dnBBTSq45Q/mSrHNUy6NlQeB8Y0a180pj0j8YQ2h8d
7ASsMPCfFQ35u9blvEhJ8tvlXDha3V/8gO6L8QIoeegZjyGVzU3JTw7OCzNp/+KE3RzDjBcRWuGQ
eHy4yyJ894PHlD0zTVqeLgkkMomg0+LOQz/Iqc0nzvo9d8NzS3fblrsDA9klOGG4ns65i7L646Eh
BaDk4VVaWSm3FsGIUJ/HnrlS01RY9cV37+w9x285Jk3KG2aFKj6mVXYc9kttfqHfPRWt16bzFNIB
5M62dtbWy1W7ObGQvuO6U+OPV12RvVS3apyT8x3IyeFuf0r9EOKDUwkuNUOJ86D5bDMTWCtzfXQg
/CLbeKIWZL+/2y4K90/gMZ/sbDOafZqip/6MtcPEGczSiJUpcmYx6pB2jq8kcyPwrQ1AoiuqtxH2
p/pmLR4dSn6FpI/kFRnVPdHWAbuCQmyfa+QaQzQL87aQljLkVMaqFmWcpQEFVD5hsutz5FHnT6iP
GN0BdEzTbi2Jtsr+H4T9iWBO35pIKqJiEpO+4lcXUeftAO079GA1pt2SXz5USTTM67WXUZCpaMAq
tGiU5oqTEugTy1v49hC0bgfF0qgJ2sBnmc9yP2KK9oCSwy0VmvgQn1dKszX4yD9+1vVaZMXTFRE7
5tqBkquYneH6vfa+RZzJCCSx4G9xwk35irat78YyEM1476MkrZYoU+gnmJslGOvfkoDmeZ3toc/D
/jOnjLNynOuBhCHG6ka20EGADLbd8YjP2wu0bDH37U/G8B+YOKNGgkEOB6rHSpEHNxl1J6yT0KKu
zkpT7KFY2XjrBFc5+FkPFTlGzbmeRjOHyFgEFEvaV06XrWeBMi2pGjFLrniDEekA2yBVuJRLaUYK
KTHyKhg2s/RscHLei7ZaDmOD7kcQ5d0QqLWhKZU02NWElKLYtOrv8QQGz+iQM4KZZPw36cc0BdiV
Daz8eReqdHGcTykIzBdFxbbPYKr9VYnR/K8DZE4PUA6Og3S1C6AcCjF9A8zNMfxWSOx4Uk/N1T9p
wapgcTBEQuwHYTaX19dnH9Kh4M90jNmlbs5uXDh8WW6jbwEgbQoS/KH2grWMagPXmR0kDS5tJJyR
DmmV/dteX9ZYlZp/EX2QrKvTX+aY+1meZLEY/YKK/3KE1HqgQ0atHEOPgcBlQl9IafPrZu+sk+BD
lsiAczLnS1SgGeSk0mYWqhm1ozCMNTdZPol6a49hX5atMQdA7KxGGVKjluQZAEYK3eDHKHDDyTJm
FIxqU+XjjR2ijytmVEGnwZvTYmc3PXo4/1kLKxkKz+MabOz2EbaTNbyRuTh/F8jFjxHpw43Be+QX
9A0Z5BqqWvTMXGexbU0bDL0L+OJNIuX8G8rRo6l2XU/haG14ETkIhSTG/H5urVlzKDQq5sL5/F6o
CAuJVS9QPgJvPLKf2edd7LeH0hetyWV92LL/UDSVojCC7yQDIhJHbGhYCrD4+xMCCenOia9jz0M7
utRoaZo5hel6tKSYuQ96YhUvwg40ybolisQJCwHkuv/50jFO+ogEYoywiOZctjV5jX5IeIuLC7UK
rTVSceVY+yjzS0z37rJ8F+2uecobE9GzwiVfF88YPWs/0NsGpwqK4hx7kSkTHtT8N2hLb7DOIyhq
qRtnkcwck6GHes7ZVAStPMPa3UZTkdzH/LExXxeQC4nSqqIagIUw80MQdDJGwpN0XnJ3+SebLE5/
AponPQinJEBSkR3gc6WJCPlRbP0KcuuHsiTrq9L9mSqRs188vMTsbuoooy/2N//5c9YurKlE5ers
KCF+WtnMOYmFEebuuhqKxTdLaQ9PE64grdYxFeVgltRFvJyHZYMz39vjQpfD7wD6eP2R4ekWxn8I
+Mn/sN/n+AOElcS4EYrBV+4eQA8uwsX+yHKcXdbS948YmwBusYyJKLf0hJt6eMgQJGGRkH38Zb4H
/vhLAWugXVvv5tg8lDO/QG76nnwiOrZonyF0SBg4xuLTmIAgF46tmhmMH4M7diPnny+QzqaxkQgI
cDpwVC9Cvqvgjfd/nN1QsBbx/BL1RN4ubmvQ9GKR8u9UOR1KFqK1GOinT0GeiIhNpNrO5OGqnvXU
9yiMTPdnGD+2eaGC0BF3iD32dFqoIKrl9VdYsbbE0Nwi4qXTAWGH9SAENkIeeeF0PBPHH+xckt1P
6xAtrp+Ovo9BJBlTQHURGvG6KS/aIaebFG+qZGvknaz/aWGIwKVoNMrI3RUYGOu2uRecayrbK0fz
B2ALpHBHpFHZsheqYCLV+1c+ZcNbWco7Lm4hFL5F5IQm3MCelcnVKBJl3eMQFWiKIZgED4to6PEm
I+PROgp82Z2q4ERUTHdJLqlwpSgZpq/mv9MZX6wcF4UheBdhiuTv2DWHqyGHioHgYrb+ikj3KhZz
fe87wzkUe4z2SXn4iLDHNNkFeKTbqQYuvG1w8k0aHsRCK2afSqt12l2+UoGbCng02/upObKlLVlG
fv9cW6jQDcELG5pTxslCa0X1Hp42XjmiWTV8hitfI4Z7HatQ5xj7pw8RutCIUBmQgAZjDJeoa54H
u7dAtGZ5Y4b3FG/hkpA8nkFTZEYxiSy6yMvrYA+7MJ1UO4WLJqCg24HZpVAPfMrs4dvUhoA5DOg8
okMbVHq3BQB9iKQmlfcCFmqNfBt8BMHe+cjx+Su/MwxAkDJmQzoC4JDdUaZHUAva2h7MVpjlVi0N
BTNV3boTQbkcu2POlURgj1YE+1gOOCHniaKsuyLso0oUyE/n4ohS73md4gUg1H8sa/TOYsbSB/qE
vjaRrdoTf5+wFGqhzzPBCdp7NDtu0l8bPkjAHx2kpqa20+snJ1spPxacgOyMCcc7AHxuTEsDK5D4
TxEhLyyplaKIWeN7zjh/MEFQGjF9hRq69RnhtD9x8ypiHqXfL834oTIXpIYTq/riEEKUoSnHUJeT
lqJjzeOS7W7yKwLP46KiHm9LEa0BwfjTGPidGlePSM7CF1eiQv5Ns82pGWZtmeJj5+gulcAYDoCJ
XuEfD8z61/m7BV9LihVyAXuX2N5gkoL2ZlbhXKWeBQA+tIZc6csmO2hyPKUG+pBJU1r3qtF8diPB
koUbWMjQAoCd2PlWo8kiBTWA0WndsdIAvN8SDXyJ//xzX8SGvICHpCxuyln6U+0uI7wA+Yl0Uq16
yCfvkbtaBxUOiRmWH5hlFJlX/0h68vFq4p1tKIQH6zNU6N1Uti7UV41jOeo8yMqa34kfcvdmpW+r
b7TEty1L2zXZNv5QFiFP+jhefc2iHNMi+x9uzYSP2r37PXEUksWgdUcboB2+uvAN1htb315WuBYt
lAqjzL7g+Jz76etlHYtumV57N87QZa5d6cvCbnnzDnpk/o3a4HAQ54K0PRM0tHOcChoKrXgLkuMd
hAv22v53fXeqHRVSA8ECKI/K+sCRevPHFzo+z6Vvd7tzqeYe6ksTnx8RsD/BMjAMoyFklNNw0I2A
9bBhXyBmFkF1M+mpahoRdODtbWbq7EFBkaLfDRfx2iG91trFuB805lRiRdyOgXGlOM1o3JGtr5/q
9icQRqV6iqQwBF2l8R1YnhLK0le+iM7bikhz/muOrTtWr3LM6e1ExfnNp1bK1J+Dm1n3xyk2RJT2
oTjm/myRWXkNJVbrEBy5SfqbYul0exYhWZ1tG0hxF1KuouDpAOy+mS423SpP9bUrGgL7oHJJkNva
e1elGZxSKXVxDzY3isHXuKaKL9s2pryi/pneYcjJCz4MrxjTNkpxHy2ConUNlbc4evs7CU2HH8e3
gy1rp2iUVG3U5FIs/LAIbTB8rhGM9bzxhZlNhsrC1hnIoUphszXni79jhrfOHmM+YNOXFin4NlFT
6oCQe960ngWOIJpPlb5i9V+FuVyrZX1kQkSVa2rSDLlxJhgslh782VgQe83GYfjXkBUNduEYuoy1
uiyB7qS8ZJPcNbPXZKDWOzgxu2YyM2uxJ3UltknC7hCLiRxWVdqfwuMkqyng+UYYpiRZ5IREBgoG
LL8e8zpxVcrUq3Ln8xlY/8tk6T+63XdrqMtSBW+pcTPgRwG/VZOKnR2IUraPnR485TrvGn92Nf3K
ojpPXINJXc9eXZbLL6yX5IXM3oMdjVqRS/eIcyuSW81t4tK8gMxrniKubaCzqCGgeKMH/WgWCCbJ
iVQJsokr19VbfG5TbCT3DZlwkYYwgUCa2Qq8DEIYWgoUnbPo42nL0uFdsQi1gA0DYGTeQJ+K3Y8S
JefNh16YlRVnrFMTYqGVTwgX8M2pav03XmfjXQ8tVVoufVhN5TNegD8zXbA4o+RiyjMUE49LyelD
d2wfjpZyUXMXrgN3PO6sHpHR3QTkp+KxwfIW/4g/F/m16cBUkMO42Sf9tFBNAUM4ZAIx+LpjmAXR
Ev8QsuLH4tZyOoDyEEBsHueV0WsdbSmF2ICaZB4pjC91oa3Nl4tLB6xbTToERgnH3czGvIFQY7PH
u/OnNCeYwDjIbWur+Vbua0+Zpv2ur2lXTOPCGAa1RGlDq34InCSJLCcsGNNittHcpqx1jZ102L2a
5Y1l5rQMw+D/8bcPMhP3psxHe3z4AgCDPTrmcwbXb9KGtKmrEjroDlPgrbWQ66YC0vHytAW118yy
GJyXqPbW+VsTEU5VcluDTa83WP9B0qykInsN6wcnXSIEGfA3YYCKmcIMZ/bnZ6dmm7/UTObnFieT
B1IuPsEEvzK8SF9JRbXjs/hNawZA8jWYZvOv5GMIqt2BkH9uF0ffHfdSCE/+A3PVAXOg/iBlCeRi
copS17HOQIvtjOz2gOK69O9bSjkdG3I5eOvsHu8WKZQ+VgMOtF8WgTe/MvbwsnMNckvEK0Qjru5/
TqSwpks3WDImT9KQF4q9zkQ1q7BeXnxgoy+sBIh51iU/eO3W7EzG6QkD6feEWA5PfUBGDBdRe5wg
iiX9ghHe1EBiS50bXklfQF2ocrTnc43ml7o26Rr8qYOruFR8YPaC+NIidXKJOkbNYt+v43Qjgrq9
fColVozfoKYTJO9a0L92Toa7RTwB4ZWVF5EQ7m9ds6oiqhqo18+YIMYzP1N2YvRogOMWZHG4tfwj
1/NNbZ2XGgQMOCz8hresOtNe+IEMePDub+NO3dTThq05Y7h2ghTC+3P69dHBj2tFWBuYty2xPjec
jp8NxCVI4rZQzmTSEvYpp43qwhi4f7yASX9EfObHgKnRfGTUgX4yxpFMYGNUcrTwbOvc9PXucpZZ
Gci1HT3m4eD6a9uknFb7vm3D3ZK/j5pXKzsEq2cNrQwfJ/Ar6aa4d/aK9XDY8H5MX2SGzuPYvwU/
ymekcWXB2/GOy/B1xQVfQoWqM3Osm0FrGobJSnO4Zhs7HaFJsjF6kfXiGqeNjHSuasANF64MXMjW
4wUUB700rIVOr7og6Gy4saN1G/jboO9JGq5Xgohb8eiXWAL0Kpw9XhlOLDuJvJfDheeOKysQlL1O
kd6trI2g9hD+NeOI5H/VsEZ9bMPJdfwcJg1TqEqcckAHCRbCE46vdAMESauBBh7QMvquXJZ72pDb
6HlvZRd+p6OHYnNZ77pWeJkKpZGcHYylZFD32CjeXI+LQREZLopvqXZzFmRUWDUZV4fabCx6m6K7
CyYSaibWgDeZ9kyo8sgiRKlOfkg/6qsbeJBVDf93eJ1TaU/sYBU9NcjX3WSoAkoWn9FbuGKaMI7N
BKbTQgEUjjkm+9qXfN+TheLjNxkUurXXSDiCrnemPzTOylVdUDwSuRJ8qG6on1JaX4k3OdST8nnJ
CoqQPQf5sOc5JDVTuzEnOjeE4sHcfolt90Qq5XNWd6ub8Jx8ODtgScEHuFFzX+c5mLOCUoYaRlxq
+vlf/TZiCnQhc3DpzlG9k6HuuULdMgamifx5EkfJk7jXBVglJhAa29Lz/PSG96DIPwhBn6NSIrN2
gFeloExAu9npClYo2/t3FmktNULsd4d+6aUPpEsQrgvdWjgJ60mIywRX5b7uxaSBMK06ZJKQVcTV
J08o8EEKh4SO7ybqtmcpLNzWwcjMfSFPSlOWnbeSSoLoAHLJgTS74VhanAkD0bA7Ma/rD91wyJ5p
P1enD79ScjuhvcyHAGDK0sssmPW1sNr3liB40Os0GlXNJtQ73tIpiEkBzMsooFHbrkmjUaIV2d/i
UmbxeDj0/3zFAru+vOnmXPah0Or++i1UFvYD3Pyvamg7aKhqeXHsSIf1iI/+CyiEiZWx3zM1mZEU
CBe1BLCPdn9zsNkK3BOotiJ83hORc/Cb66Tbn0hDNwgmp1ur24kuK5cgASCEfPSBPx5AAoHpqZVR
MHMNeJuwEnOhkOc16YtSGtSsZRgsxmbTlzXCJdncCiawu03urIN0glNMLiqWarEDWxElySrN3ioq
WHOJCYI/DzIKh/1gRvVdK33AXAL7W/XrvUaTf+Lo/rx+osjuAEylMALFQEK4eSsgxMlD3ErkBNZr
nuxLu/hSBoKLRVcAwJB3HVL6963N8enIy+Nxx4aCcQk9skdX+05AKz+D2qLCssNC6aQ60nAW//0/
5YCo6PikS5a7BmA7AoDNMQWRH6IYi1EBDuuq0ZzUJgonnLpqFiKPiREEC4OzKlAQGDKY6K16XMl5
5kr5C5sWcj8UxsVhfV1QWmiToidKqsMXi0FORw1cIACwLY0h3OzFwIfUd5Vl5qqgdylYZMOdJzH6
hGol3q76wp3Ls2YecWkf3Ng3kj6MKUxaJcGa3pQg12zSiC8NH3GiDiIhOWdNhyuRtk4ix4FX0YWD
3YryyhSQC+2brWnEFXcFNlPiY7kpF/DoEMXw+qnL9res8w6sYjpYjzWMY6uIwH1MLBRlimcmZtwK
MD5cxEJQISV7v//7auvnE5aQL2ry2L5+Qm6DPQ7OaoYb6G7gW6rpA33pUm+HKJCoh8Ky8eWecErv
kVoY4Sz3sOnrCKkv2xaWowUsjaC4s58kApLXHBwQO1gXOtB6NkY346bt51EJmFlUFlsukcvOp+v1
WRrg/3njXD3s1C0pN98SoaeIs3O8cTfpV+wtAEB6YBi+gWLtT/k4hZxn1+sTQgcMN4SXCIHnHcLN
3Qi3xrNwF9jFfJAhZ9hhr+4yNRP6MhPsG16mnZ+gbrDWMkYez/hFbb3FJK+sZcodB5jG6h5fv6es
O1BZUsW/XFak38uS7BLRo5SrJU1g3hyJe9SJVd7ia3eSVihY/0jUpnf0RMooJn2Ay0AQmXlTvhvj
3aCMMGaPjlhVz8wtW1rZswzeNnzauJpD7kumXnqE1yuSuvkWtfg5DpInfK4ko/SCVl2fH9dFEpiA
MvEoMQ2saLTQz4wMgK96ppQMAMqus3VGjWl6MrkMTgV1N+K+7e4uBAZSQT8nCXydW0aTKAnhEmnW
zbE9YpTQy9Ff7TDs9NeEX6usgxCyKJaSNM1Q0GB1L2M86TSNgYJ6WiJKfyhQWBPg6YSdNpOE3CT9
62QMFjVlCPCWFiCQRjY+oRWMx5fIUpytvPvovWjHMq1VBQNOkvQ7O3ISS5al5GIqKOnG6FeL43cs
OZhteoH19AfAThefrxneB2VtxhCVqHY7ZtcJdqjcar9oSQxXeOCz1PWr4jd3VjuUfX7wE8MoJd8s
nXJ2armZejzw88+Hu1lHspBPNLmXOWFAPZJjoLP3qnksnz1oONk51sd72AXcPqsDQwgqzZWo6Cl+
AnFlMHc9V2PLM5NCrpVIvsxMCrL16YvppV9hgVQFZSWWHVdU4vyyBGvgaUv8cgHJ7zlksR0T2CVc
XwFY012uQWzf7en+sM+0Y2sQ49qfZc0qfDvOGvPOGxNF/JSirkC+IB35oG5YIoLvqq5GFLlJaTzp
YY7DtsQXzWqqeA6uACE/AZAQtEIUusICu1rZHbvDBOYgjWEgXWZkXV7XO7MQUv3y+8joGEpPKBkj
CNtIm6/5qCQEHoxYLUCQlePyFWDyzKm2m49l8ahR9EOoErxZs5THJ1jjFAUc3lYPnjRfOJ8HRamV
ELN0bAYV1ad2pAU8ixd1bzCtY/HrtUmA0AYDwOAnGUhJuFYprc5ZsKOAtXkFudw/+TS2fWYb1boE
z/hFuyuNnANc1ZM+Vi+wKwVLvDp8yyU+MiCPbABh1ON1DC6ccwbZzUneq3gOgwRTmMRdmGrlc3XC
2NvqkgddBnd9PbucbcXThQp9Mic9/1B70Ur2/HfGdffQyZ6qq5UEW70BmvJ7+99M+3XzAudFLmqh
E6oecdHXWClku72sOeXCxd4jwp9xVJPOoJ3EBmklX4CP7a3w2deIhe5T458+Ek91eWPZS/0ST6yz
6pGUs/3vadF9GWq/hNfoXIXoEF5RUk9SLRVw3Ni8bkMSgvjlhqDr8jqbHmuLYb/fnx8MxrQlXYqo
yOusGfIP98bMr3TXeI7fKHcK22k8n6JiPT5AZlpHlMn1V8gOWYv89ZwVHjImeEskWGNvgByErEhS
IiDTWeqzg7Y1Y7g/xSnWQcdDk735YotiR6BSHN0a1GPs+Pocw+Gg6Yr291mZAQIe3kRMMszmjdHL
kL3nE+BGKBxz29BY3yZwBWO73JioD623oqe4OvnjfkG/mOc2L1cZSWkpbb23TXuTHstdaGI1xtyH
4BpH5tPRg4EgfAoV1qsQYhKr2I02HTnJumBQRkaR0BsH7nVwzJ8xcdPcRR+hzAkpk0GPO/Kdtzyu
ZbWHhIZlLnNmMTEl5iaOcrcqDLcyjntO3YT7zWyMUQMz5Am6gFht5/+YrDTloqPkIJzZ/MLWcT64
SGLQ7u2gWyoK/caktnrs0w83WkfWiRjsQqrBlbsmJ5NjlKQ1gJlvqEDQi9x/6bif4jeZlv0f6bkb
PC2J+EC5kxoRmzGSRHimJQL3CjZYwJtXr958ck/2flQrI6Fxq+VyRf27oEoC5BOSkoH+4YxiLd8f
TB2fcR0n6jL5ya3DrhZPqHmYBHJIsCV68cjyXPpNh1nQoJdNKNib7sX2H7xjo6W9nxIxSNTV2zGA
0I77qeVV783r2tuyVgK+M2ZPpnjiJFe5FR6nNR+uYKJQnQPbyF4naIoeYW1UsgQGdIhJ5nF03R33
bwtfV/RUfYfnIUrP4YXi8zaZzSpf5W0CB6w3tx8nLxT9XdBp2ZsL6cUK/hLf43ezZjHOvLnqlItN
N32QEy/mFcJQS6rLvtVwu0+e+zwVsBmkujWkQaCAWzD70v/TL09oDj+UF5f0TrlX/1eCRGlwz69q
4TJzOb3WquPMmtsGpjCJtIjb3cF25ENCQw51I6PEHXENMAnNlCqm4VnWG3tbnPPQrAZ04t9k+AEj
pBTRVQa1/e5axktcdnEbIujs3s8ttXgHbXRM248gZo+BrI8si2n4HPU834G+gMEHHaDXVAlFmNT/
fZSNEQwnuCDT0ePFlLfc5nypX5LFzJGzxkSy0XxpjJgkmyee4B/hUm5KUbWmsY7+334Y7DGrCRDg
TvuX+V/Jeicu7EOughJQ0Hwb6t0HuYHvymfu1/wlBP3/YRbbG+N9JPqvDDTpCh5ZnMPkIhyRjcab
jBOajOUc1sW2LVm1c6yoejOuOasNaiTurJH5RdJHQozcOq1HIJ+OG4o19GjWaJ5vjriLHYxIUaXo
Kcmw6PxL/dpSiedhAKl5eVm+SP+fY1xpql1+EwH5S5US5nM56Vc21hgDxZe9kEMfOeO8PF5kBg8q
inGlkUIkfWOq45RvUBR4FMJ5pJ4APNDdroQoIldAIiYMuBnzi1DTUd/gOOm2skrjOvsOnQO7TcOG
4DD/BVod8GvfI62J3jYnveI5bowpl87IHxX+9qtvkazNVc/geKAZKSPYdu7twuQzRI+GErlV7mD6
lc6z40WGNX2if5spsw9iyV5q4BmMnnsMw49/G9+AADaKk68baXlIc9iJBMTLWOczqFlwAjAQy6R5
Tkm1zF9UhtE13G1NME/PvNEzkPbRDRPskBGbLT1Os1Q0f96A9iN3cIpaiTTmD5vLTqEUNOhevxhg
Y/lI+g9W2J1qHrHq5AZJs+szaa+n88Bi39KqUesEm9gv4dxuKGw/PSBKamJQDdF7RPxcRzrWhMnL
r/gc1de34qZC1TxSCMz7ByEwJx06R0qjqeFC7V2vGfsk7qei8eH2M0GZHRiuEeS/6EuC8Dyz59hG
JK8WK7GXJjlCHng6SbrG7JVFXruh4woBCI0ojvTXbD8MQVm9kl5zE1+VWHiUQKRUdGy4t/qX+7vK
BBArs75GPHIrr5eaYJEGvwx66oROETuMXVTYIeoD/oKHMwdkThaYBzMC2F3kfPlynikoKMhlrQt1
13BW0fAwz5i/0vSMNHo8labHzbb7kEr9zQvPhvnWuQxGEwQMisR6+VHqZrAOivhAzNY/hjoiT73U
lKcdpG5f6QeVainyI2E7JBmvRddF7ioWp0HKO3INnHpPWuL6OxiQJSJn6leqyN9QQ+QDlkhCQthI
71Huwe0+YDOlt09SnnmWxGPExMsbtEgtLjAXtiMl5VKAT3EsPuqhd37McQM6R2sViueFtpD9oIM3
31vBZsj0Z7xIqEI7urian/koHdwkA5I+9RxcB0ierOXUjOn5W3b/7YuWs1WkUP/IV+r1UvTPoZdW
LXrEDTU9CcjSQ0EqJCoZ566Vwpdz+2YbHv/294lBr9C4sY5I8jYmQr/KzC92M0mkuBXTfao7NlW7
ExXqRUhaWP2H4aNk0a83mCcOvSV4Nt700Yxu/oFFwxg3goxByBpczlkfNOgAeDcald5UrZ4CXxY5
MOdO+XYrawV3DYuot8A5gNi5kKmQiA84NFUPlDPTuVk4LkNyUXhBHXi9FzvZIaE5hAa3moRJLIFH
p/nPHc0PzoBuisZIhezLGiJdcFa7C9SoXWhXgbAngTb/dKFbzg1W8CPMYzQUGwQRPwUeqm0LfVN/
e+jKMqw2CXvFPpLPhXDIWt3UKegmCi/XWMD0NIu5cPsd924eG2bd5Mnu4NrlaaDd2cJn8g3nIt5r
xSkVFwpRbKHiPs67Vv1szWn54pZqoMZwVhqpJZHgSV/WXkT45GS2JJWGcPvDXM7jjfSoWtSIAGYF
CZNJkNdnJSijYVO6dF+Yk2xYRROlG8cQEsNVRDPWHLPaTHPGPLp/HeioedqwQ55sgjNb2T90zK9P
KqnCPcuCgMfeLGwxXxa+0SWUubUkgSRDS6YaX1aXyX+7s9dZnQixDRhZHycEyuKAXIsArvS/zHqD
SZNRYOx+a2JtdGF0JD5EFuRLO12kOBBDHhU6W+CuLffALY2KsHzI9KUvOl+3wVHkbwg08tGns7vv
F+0OxMzmLXZweaqsRAPmiCP++LqRrPdpJP7Jg1ILLdze0AATqu2rMCnib6JYduYFKYnfsAqkrvg8
XRCSC4W77hYfNJFsO4et++It54iCUo7w+2V8s/irOE5wtZktUgg5gwKUAY3verZJQGfKQXPw7xqO
WHP/rEIkqmpVs9ZjvdedTwJyXwpyg6mexTP5vKEwU0FKGiQnXox52o4VaJi6V3tVozypR55cF78y
GqFWfIz0yzFDLZ59mKEJlb4c7S5aCJ+B0Vp4DVFLzLEhJHKkTB8PcpSqRvHwf48H51PE7D366ZLb
w3Ua2H3GdVNSO7fZ3DFyWFMX03u0+YcWTxd0wZNELfyjAmnZXLJ1A5MpEbhKUwN0GaBgMAcTdu/f
fm1+Hrb5xeHatedwf6glIgg+26mNKrWOyPfUct6CkItMus2lkbg+sU8EpeyMlUh18ApsMXzhyiCl
cizQK+9h2oCWysMWvCMnmOYfniyNNoUuDI4QF2T5vrf87oqg6cOK7iuAE1MRCyqY2CnoJslne3w+
/ezyuODwdNhsus6TgQno2abEYxpm/vsFvioJLQ879Tr44B2wS1rRpeY5jWEX7SrYbEfNs5tvFMJn
qXC3pfmZ70WPwWLtGvhsY9HpEQrOg1KHwJ7Ngi0GgG+SOx6sU06o0QX+90mtsmDUtb9LQqru1zxb
jsRjZHLABkkHifGk5fq2i5FvL8L7S63sqko9+xqTGJC/OFnpd8rRpO7W17oCf705vU1J5KeCv2hm
YFP5cAG/gZW6YXNDaG/VKb76Y+Pfzht0Ddmm8R9cFxNisaY8tL73HObf+ZOHJI/scOGUy3irzBLF
/AnfsKqNY0KN+95AtcpIiOsp/5t+OBEE8WogtYyUxPHZxuXHZCr6yK03C0SI0n8zaDY3MJAnIFGV
ua5cC6T4uAHTVK1yELsPrm+BuhPm+l5U4mPvGz5EwGavAV6i4/C5L35YZMkrEVTETWotnJYckJN9
QSDJEYQ6t3e1OJSoMbtQtKWMtUsSFNS3lgmDW5xKj/gYKUqwk/h7u8hl5mIF0PyuOFd/cujbZAJD
NVEkjpOZUE1AfrQoJ1Shy9ImDW6LdY0ryDKM918MXV5slglYcjFcjr8sAUW+kbptj6vW++CNhrKG
nuBKT95wezkNviYdqY3qxd2ute//YT7sGYqf+Jue+QOUTWrH7L9y5duDFWVNUV38/RNnJoRDprjx
w+FX2GLxG+L6/g0OpozXlHkYjP9MXdCN06fy6mGvgBemc5n64ammwLtLMrFwZADkkmsyiLX6n2jQ
GBamZpy6LEYGpkTIyJRuXsoE+1SWph8hxnh7n/w7TK4vmTzSscJQ4LWxNMbx+fe1RqWYkuzMaLyi
jrWRxvmEpjNE1HbdII455pGWBLnd19mdfSsrucJdtyy/K0+nNPGp0KIJm3Xd1Ez9+DwXHhQKtzVP
ArXEbaeqEMG2/4E21JAeqO0jyM4hjt1hhg3OQfBYbnVK1KiJ4uGc6YYlh9MT7d9/jJeKVjBWQ+Tx
UEZXZKNtlqt7RDs+zZY4FxlSA0uPQBs/b/apIbe0aoBedpSEHacJv6QpCIU0vMDoNhyK60loffUY
TQUWy6tqYI0+TZ7EPz9CvERtpCKXgbBZetURXIBFQMp6rgs52w4uYrFRp7IgcSOAo2y+1DK5yKOO
yOWhj+8x8CIyl+31H4hAOZ07xr94f0iXPlwYZfse/6aE7XvGMwCTzygJQq33MHnVfeK2zl8SMkHE
I+B5RZMPNrHLgBF9NqANKa/RKHqJowbORGZlLq98+G9g5xFSnszfp8Z4euK9U9bxwpAsCc0mcm3r
c0+SpogPfqdsbMNy050OQzYhXrDGnqJqnbRhcTVp9bJMhQpGPNVFck9eLvXv/ukubmdZtVsoVCqT
BkndHV9m9DtCS48YDWi3q6hx5w6fzSStGsRd+gm8sL/CNX2W+49Ttl9e2+qvB4RELkftI0P0mW6E
AuhU655yAR3R7Fowc6kcxWusrLo2eTHzENm44NQKrfI9z/frhuAfa1fG6q3BcDA5r0SebdPLvPDh
g2UvCNVK4twX2oc5Nx5YC0MNcCCQ0r+Y3bnro9XJ+XIkCWIvymj3zMsUU9eRBEMCJhzDIFIs+tfM
XAytQ0gOmuHRvA9K55zvCHHvcG7Boqzct7zBWy0RRAHP2mqGpVpu3arU2p9a9E3P2rzgIzCmxwdM
VoU/Af2FvcYEwzQPwvIx5IJvA9fByTwlB338fmns/D2qsbwBcP5hJqyLs8VZ+LHGd1UWKMX8VtEb
tTDqv1d0Y3Q13uxJEXAv2OB32cdGs6H5Ak2yhqlGPYegYEn/blCin6EKgHSmhs+ng+E7um0OzbTI
mEum/THQ05ak43g3Ogm6JqPQjSrfKVMdG02Q4tsxMvejWz8fnUKDFLO/mgQaUElRNWn7Pw1Q4Zyk
8BZYghh3wV2u2wM/+2e54pQMVKSNJpouHWLPuti/8dv0gyzBIB3yKNwW2UfIixne/CaXx6UkKlqT
yoAuBm0QI1tA+VdLpPTujy5+ihbvye74sW7ELk+XiG9Sz/2BC2aLu+RflwTRLPo3VpXwDhUaA+5k
gbaTfiMcEHy3xMVwsefsVF+V+ljk7hdBQC6S0/bdt3N29DRbTGsVoE9Jg+MumT+Qb/+lMExBqbaR
DUlLpIGAOVykYvmnQT+BL/mX7EAVdcbWUVYAKEf4zQswhN5N3bgsSH9MYNuecXUhxFgQZlQ29Dos
LHykpAmAUnT6P7t9ipl2q92WEPesXu13MCmQFZfJ9EuO7OpVPk9DkM/MFpmsR7VVu6aMn2bRXAeW
n4ksni3JiEjjAYMToKSgVQiTWwt+nJ0OEWDcUTVv3YlXyaoy0yzA+Mk14QvIYPS+CVcKjXmymNIm
Oxgtr0VjCdP9Xi22r/R/MM7WKN9dknbiDp3p9rMyiqfJAmJR9c7FRfz8snWzBqMJyGrM3UVV1BJ+
DT+3AGMUpWzUQYTD/WLqWdzktzIxgd3VGtHwmNRNE1SHcJS/fhDmbaJmnzr8yihrsDm/ikgsXm8l
BrmBKnFo7vxoIHGeLb9hkKne8mrXN6H+VznUWg+DjOltgNc8TUB1xhlhBQjMfsE8+2kIw9Abg7tK
XIXEySrjnpKfbAt80Fja0NBkJP3vEATfIkNLvx8K03RSAiw7O6/RdvGEOTHt4BTm5Kqrlg7QNL/B
+9m0GDAyDtGuFsd8p1rMVdkj31htlD4xfAGbUaojws2HCBp+s6BlP2aL1HgoaOGgJ7dZeFydUmVT
UbpLdmNcR6OHaLmDVy2nE77uHOhwZmZKuW8xrPaqMRQ9sT5FsIJJd7p0+JNXlbEl3fwuO4cJuS2H
KdRMy6qo+6ervcLUOZplEPobFPnva6v6Eu46jucQ9c2PNr+EgdZI0jGsq/y1X5bna/T/9h5ypxjI
3dopCjt3dbOxz3ARgYlj+IRgKDSu/LjUL5FDvU9nkkzPhNuOyy9GBoedY8dYtTTMffinq5X4wBWQ
FQzSE4NPd82FP/MBTxrd/V7RC8yqsgV+kGNOvqFHSfZ0BrjXPFd2xeqJwgMAcgrejVSYeR5Hmkle
z0SQjsntkroVX0OJFMPRPCepcIkCtm00T8zQAV38ISZIMjShEFc5wHHXHrrb8gkvm0aPEnXQB7IY
e4gMZOll0k5u8os0DLjOEAGbmp8gmraA5a2fuAWBwOqHjaYvXKSfiFJMQMjVs7I2jwB1KkAHM44Y
W5NozP/7aWz6lDKYTTNn+H09qiP6yeVmX32cem8MZiRvQK2TWf2Srk1fT8ol0NYD07IIJkqZNnAz
WADlg7PXSSPCp2qFDwn09ZVGAOUo7EKRGvpQEHD3sfESWuHAPN44dIH6Ipt/JHIrsWwm1XA8slST
X/8YSezaGz/nNchNVQEIcDGsCXhnVsP0YkElEXKxLDLd2GS1Y9QDxF05PruO0CRnHGAM3nu5yg3I
XPxL6o1jql8XTKpO+jmA46hlFKWacieuKk7hePYLwzCVJ1b4DpkHSW7EIGkp1GdM1mHSSc0ooon/
hVg1PRx0a1x0mK1BA1DrNX3Ts5KBnxN5goamwBA8w27OGiphKwSvXuqQ0WEBBx2TkWYecT4nnTYz
m1zrskMRpnfrBkH/unM/sBKARU38tpMe96KTTHJ7d93S9IGOSYx8pu7Q7G81vw7njRBoH4RSyC9J
twNG6elWYR8FpJ3zDi2aaf3TclL67xf+jP1j/pTJDT20tC/3ac33PgmqMjVL5av0hRWUJEw6sg9m
RCajxWRenw1gWiiz4ChKD7p5r9WfdX1nnkJuA0Zwkd/oVVgz69ZcFTyKXbF1/4dc8L8SYSGvG3/D
B8lo5W3QdVW+BS2EO6DlpuAOeh1NEjyLvpD2+x6H3kIhrXuEHQNuoKbdcP+fGc+KPFSExvgSNgsB
5p9EV9n8LeJHWzcBhY/7GR6TR4i8gjw+F7qOyjPCmFwSzwTQ9mq0QMsoSgwjBMvU0GIaEpnntnnv
SYImsEch1c1PVM4dRGwUcN52v42ImGN1I8bjDs076BIgBAeiPvzMZ2zVvBon449R1NvrDhzu+1yA
BxhN6UouCFJEKNOE3iKMtZ55VOF5n7NMUqqCaM4vIEx5zUaU/bgQPq299w41KKtQwwcmvk3STRHI
7tpY2jFHu1FSJiGpyijg+4Tt2rKg8D0kv9LscjbLdhCYOOJRwFCD7qU2Rmrn+DOUCHh48Bn/ZRis
Jxe6+5dz0G/swN000m4ZWCryfub6AuWo/11+/Cnm4tcIxZf4yinHBS1EIP5Mv1vp2+td1JiURyuE
3CYExuOXnVD2K9FXbRotpkW/8iTzV+T07ETwmZcSz4iAuaLrJckXB204IW/uw1gayFtbmPP85Kmm
EbNi38Jy2Kr4L5wTOg6bJD3zLmSLiydDpta1HGKXm/Ku25yNONkXySSpV8IXEkWtb+7/aAtHfRKc
gxr7yKjviqjTwSoUCZ6hJ1NTZXi2wS1ELV6BWBtk70HnVSmHQ9p7Q383NjrydWRBQ5Lr3WVxhblK
scwVhs7kLhkEdsmQZn0aeOco9dtaiIVqvPCTSioWSE3BISDS8dFST5JID1f1utjJEIXNpaFgIYQs
PU0FhAeZyXMFZ9NZJTz8aoYeQNSJgJcCPsxbcSpLTXlBvqT8JRyzEZujK5Ddy9cb2YTGRnd/oKeq
D6ol0e298mXRL8UwcGYXW8W7HT9IpnvIh9H/qjXq15yA8j7Coyg+wqJ6/R5Jw9WbtDyId+W0wQRj
4M8FsmjYxnOuxh5dZU7CLj+AGHCCeybImK10KorsNULJ4N46bsmOzORqtaOZBhYGuxL+aCkP0mUY
FGx/tnI3Oj2oaeMFiEtyNN4HvnSLGNMwksm22OS07G2fssp/rpQYReput5CmO4OskRbpH+DL3LGk
97tx1ogRBX1XtqZ77StCiVwsvlfKRL/TOHv2kayz9BzqjxME/8OxaXTgtIATBICYLBYxZtEjzDKA
GvovstvmYEtxPj5ui2F+W3Ahvc9zGy3Q63D3iOHqOcWqzveoI5FXLbZ+L3AMk6Z+0mIR7npkBqaI
kNaney5gOqh7ZvR2LULz3/aPEHLXJHbmY+gYzNKMzIJbQUwzmwDKf8D10FOCK68YeXB50iLVFNv+
QLTs9BsbC0IURSDPX9kFBa7beb3uFYw4wcfNMhmCyxaQRVasLwDCWrSRDxf/bW3ed//k50adVmR6
eSWq4AM6Q8OJL7GZybw+y7QeSf3QBS43M4xpY0aPK8VamMfhkhxJuNl447gFeND8Mc6SFmGYGIkg
G8NL48vkYlqgXFeEDDRP0lGjxAMvO3iH6Nl1zxjtbQZjkSHUJiLZcT4Fg+db9TrV6aB1CVZ/QNC2
W69yJBTMrnzlTZ0WSaYvHUxxijhzbMW1I0CBFSTboRm2tF14j8K1Qj2JolKPqhZHYLBs91q2y/JD
EukDT6LlR11VbdaZ6PPK5GccETXf0kRZTGo+YEq58YjV42OqsxbCPEm1wRCZxz2Rm9Oq0GAFhn+P
h7JnkjC2OIafpAp7gScB+JWNe+GOhPAwAPJuRzQrzbVX46hfoD3bzjns/GEr19PuUf+OQjDmaeoJ
2zjhBoMFCazB/nVDYNQ9mtQe8D5M02MopMcoB8+DYfvorELWsMtiX5of+e82cx5vV1GyWN6bRsJx
J5lsZnt1/34n3G2Z+h2MUls0dQuyTwkOL/ubtjzamAbaZrtqfW17mKmQKEGe/6Mpsr1nMXoGp5KW
e40+Hdf+zDKHgBuHuCjYREfkX9r4QqpDBXBQLob8R5Pq3Yd9zbNNsZmQigyrGFAVnZz7LSlN8DgY
q0ONL5kRwpVIDVB21Qu7fje5idggCkzlRur7RPfTn6+QMCWsWlWfcsy2GAFpm/4BM2THGbbAiGEf
U0fRmxNMSI+NdmcrtKEGB4Ui+N46O598Kq0qn5ZSliC+FjUWd3s1538YCBrvoVAhiiM/LZ/ErUbT
qO0YLjUvdZdwUcn9eRr+7oJrjE5NSLMT4RUjN50n+rSAXlvBUh+iCeGaegayZpSCTDUF2XxMoOFr
+GHFpZBNLk+KQuQaAfAcoOjp6H9l7KXlHcCGDYtystlTdz1nCM8Ci1UTJ3FeYSrEDc5x8L8XkWD2
fvOz13Fy6N6BjHiBGtPy0R5HJ0z2VtyJ+jze8lMLHHw9T9BL5mhacda0NKvN5Lp43F7LaA40CARF
RNz/U9kQ93YIDDSb8d1XOsF0HGFHEzwSji1+wwZ2gVfeLZfA3o1jtYXst/aoO/W728UZHy5X27Xn
Dzty7MzPQX4SYkt+sJ23IynFwyZ3Ww72e3efgECWibJNRCxLSCMjddfXS2tmYDxPyJsG8a04OvS6
6OWV1XyTJraBa8LtntDIO+RYDkAeSP94aj+kgLmTxVcXBv/VESt8+hlRPVRMnMZeeDskZDkOWQZp
5s97NpZ0CETc2DgZHcYh2m1ho0P5FuC4VbPYq2gQOJydB5FZLe2UqYUDPCQS5WXMkWYMiGIQFIFz
zDI/WYvxS4Jx2OcVvLvOWZ2uBEcQn9gaC05lECSYTYI+vaOg/MBt9t+cdTbciMua3xWazeWa8gMS
oTaYEsm4t1r0Upfu1HaEZ6hCX76h1KML3I8G87x58mIXwh9GauVRnT6CA5U6KEe8y4fh1v0mu1P0
5XHzLrMwe3Ahozw49HvLWDy7fhv1kky2QtTX6v7enrdwM3Sst7wzg4NlcvRET1rqr9u6TkqupZwA
zTGqsU/wSSsXag/ZN0ZSA/PxEdP1YO8l1ULFdTg5SL+ydq6GPERQjv2FVjK1nrROFgOxsfi+KXoP
RUbYu9btTA4/QXAC/Eau1P7tjXyY3yRz1mj6CUK2JCu1Ramswt0RKHhvkUHC2uXc7yrhvpWexvRG
+X/BOHuzGVTkiYye9Zt57Wewh5P/9WaEnSJdzLtJw7kGiH0vXNs2gV289ublE9pLpKQbiGB6rrkR
OJDXUmy1lz0Pxglz9yTm2v4hoY3mh4bXp2zud30cAfkDXCsJ6i+pkdpH3J5P1YwzQ62SMJ1ec747
YUFSoHYttssjtDw+FwAKo92Gaa1/ticIYKTEsH1bd4USHq/wbcyeCuG8PMry0zv74YAoSKnuaoVY
zFai+jr5WT++dOZIjWCeI+vBUtCHP1RCtMEC1romGZvD+ZEQTvdxE57JcARDGxslTSBDP0FCEAQz
1V5JW3mPrvAXEIAgrV2zkK48breZbPB4h8qojB+F2PLHYJDAnFo5CbB6SvNcRHzVdeM5lRyd62Yq
evKvDrDYDLGNG2usVWRgzCJVmr+UG7/rPNVF+IYgKrGEZd35FCKZUtLIPDkXSjC24yy6XhUaKcj4
thtHRyrzXWTcBA/MSvkOhHDD/EfqikQrXgfQE4ReW5zZBD0GvrCqEfNGkRVsVqZwOsYv8Z5Oyp/u
su3zJbZlOt9JU07TQLe/XapoB4iuzmXV5GslJi8TGtvGrzE9uknB0kBFZYDcrXCrqvdY0dEzZB9+
qdqv/clojdMXDEt2addmF3f3f7+FrbSb+RYqE4bOfBX8pQbXhbGR276NxXHrju2WMeWDORB1Coo6
lDdKi4AaarrMdH/Ds8G2krQjhn/aox/V4ou2xoAKJ1BYf9iTq8AdLQe+Mq50eMVRkxxBjYb28kUq
gIbEVl3wm9m/jpGHNXP8oVPWeR1JJ9pHFNCdaOox27huwOtBwew4JwpsLGE9DGoij2+VBwv0vDBt
DaLTOXZwEwvuwtO2J89uuf6AXgau7jBaVET7ciUZHblIPHbQ9WNl9TFxwjmEFZa4HYu9EnGk+Unu
baZhUrDLqmpdiCitEyzDR5x7FjqVlSqFAwbh5KzP0CNCpl19BRmvbniFP2LL4PwqYEwR3trEQjgK
/By53zrL8Cu0+OCdEsgzE6mUMUZ053H5Oz5TgpYSpAKX6gBU2l/CQgF9ietcTKUyZWbIYxcCSuGR
JPU2PYP3thqpi5oXDDE87uJ6ot2xAOUjEm7o+P2vH9psGDNcTKCrR/0QycRuS249AnSdxEhCTyeP
vg0UFbiDwctzlAiuAVeOIgA/sg9ej3t30BCsadYpmTgBl6U9Hl4xHOVyD9P917dY+Cm1Sq+4fEqY
TYh0N+8JRRjaC4TKWCPn28rZ/Yv+wXWqaVyUTk+1iEnEWkoLTSCV+nnkrGhFQewotLa9zAh0ZXA3
ktfV5pQpTWJi/Kefw7ufkfOqHrvQfrPv6gIfal/C3oUVkr2OW9bmy4NatrzZluyOLolnp7/idfYe
mLebsk5tFGQll1crJzpwSfXIlsx46ULErqb9H0Km4AIDc6X2Wt6R8Z1paDt7Q9IFBx64ZpO9Hfq9
kwZyEC+CxcpmJd5fuRKjn6umDsCxiuwuKlmdREEvKbD2TkMJ811gbCldB7A9ai2oMAFRTrhPUKHT
YfToExwtMKPjwAWw+ziTGx8ZISrvn2Dha9zM9eHEVNYYB9DonlARue60KEQfAlhKjL3zLt7KRFe6
H9JS4SZZ80C/saPBV7bgB7dC18DiZ1stu6UiXEfnkERM9IbOoTjirwlY7A2v22bgnAn5MMtJzoqi
95GyzsWsvSAxjZntjEeBbMs3qHfqjBKenxoV9imNpcw5j295PWqgJ9Rkc/VdHEfahv4g9ZreCeDQ
/3MhVLfXS0ZvGeNnTZXMp90xOvRpRzo+fcEXyMgX+JYkWWgkxSDVpCPJ369lxZSd7cx8thCwLKyU
nPnyapRQPyFWshbbB4EG306BHbWdIBviqw8Bc2wLD66xh6k8HFjMF9NJxswAmwz4DKo4Qqizq2W8
Dl34TgVtShpdpSs4B1AmQovSyNgP6YgmmcZliA2ppF6ruOd011yyBRGzaThDgMHqkUS5DmHSQcsV
jLhsN7poI0HejhCgNdwbXq/oLJTmrzKUC6VkYIQ3BLRNclcuAT2I0KEpnHZZxdvyJ2NjuV3MAMLz
X9eUhY0Z6tVUGIe41iQoNgFEXscc7gbudsmo7mOhMQPOPEMtZfxlbfK+HG/+tsfh008QqoHTqeI9
BkCWEvDVRrymsdXCmKF2tO/mwr7F8Nndkt2J2TynN3snCaS8JaNChcahaZX4Vs7MhUvFgkQ6Yk0q
xH1nXwFDyGtTo05MCoqb9jmSTs5PLY8/7NJXm6ljoxAc/pcY/EBaPdsTph/cuDoqTRgSALT3s1U0
I9OrRzOThLLRVGyAqckVwtKazvHKq3JjYbhIT5JSNNnQ5kTC5SsbrX8yQ1N5lWE0F5mz92lrLuUz
KHhLyRIH2aCfcYg4hsqO364qxZpRigV1fbHzYhcjsVPrd7e5RWGAFjVwtcan9FFx1GE7waRL8eqH
zeh5wRJ6JLCsCqsvIJEe7Ar//nBYQXk1bmN7qam+BTwP9r5c69zsPxo/lDT8XNCGLfw3RQP2Uor8
T1l375Z9L8JSm/yc/SAvAGRem9MaKkotnvh9IvScf8B8V9hP1M+xy0z7Ay8EJKZqYvqBmrR4fnqu
jUtCeIAI/GzZWZZs6VULGG2xAvbOo7P8RzeRb+ti22/hbZRwVh2pSZ8/TaTafmEBaEIMA4hdUPVu
Cq5q81ETWGHQRoupKj3fE0+24RUf90hux1SFPQBFpAdwLL6rqlAZ1CSWDWbdKszr5fhzEMHRW8kG
5lFb23oo5FfR+GRm5JpBjEzU5oWvPpw5W2ba8aDGVX0XCYArpDRe4RGvxXBpki0z6qviG0Fukaok
fpJ/H1xBR4EatmEH2sMLkC/z7kUzLn5b1ssu2YapY5JIFEUlMnsrpIsASuBNowucHtl6eMox49Tw
9HCaRrENPCrXY3eAhsWzrrQAAv86PNS1G+4Zh/uoviJv5TxSxe6h/IiDQxyC0erCtef1npHW3zEi
xjznMqrrl9FuxmxDrsG0nxZbgz4o6e3+0Rswv0100tMR6SL2lHFU0sS2/dAZWgWqbgfetRaD3F8v
1vqIlnJjFxk9XlhnTAqraXU6mOp6jHv6zbUfYOWWCBpxbylKI2/mHHxbCDH2VgQ079xfRdt5+q9w
kY0XN6fD/6RtLpnIyOnvEWpHLGW0diJr1Aq1EJvOJNMxUR1MxtozQVAdAhrhzjEvmxPz6M4GxgLW
vrIxncZWZWlf0LHKOYAz+hIxULemKHkmrJv1FpQmiHNPcCl1/WiCwS56CTk64zkmyPX4VWjUwaUB
8y28wcgB/acoYUyH2v3hFLNXojioB1azYzd7/DcDca60W1Cpf7n8EBj1yrqh/N1bYTVy4GlKUrF6
WHjrvC+eKPSMXGvD06lZBMUknb5P7qHLWdr3JmX61nOH2MLztivPfUju0X0VSjqftH9+cJd08fPE
MTpSKysNPyT7Sgu6TqIyUNJ3RsiCE0zBI9fyZIG/YJsmpvpgwBJ/UFi0urATyZNbdd7ffJo9KX6q
Yxx+/BlU6A3oDYRXAiWUTM91ML5AwL+D3hJjDUVG+ktqYaHP6JzykZQLWBbeIPR6kiCjpCa+GWHw
weGJNWj/uNCPri7ytOLg5dsYMITQuHfq3iZI29JAS+m396N2lnzUZyVXbr8skG5nYwLMGUh95afe
7sNNT9uQtccCYDYSC3OMbvTvCCw9mlhNS9a1JiHUIUIv6LXm3yaOM5XRI3xBBuqC/iS8gmP8SowJ
pBlv+aSYrxiSQZSsbFtCHDYifLenGn0fHx+OYmyPHhGBGnfSXYpZJWMzaWWM+PVT/nRM7ln3ecly
YrcvEV0eKKUG24KeE+rzvv0wWla8CTxvELmos+Y+0f69NzdW3/uAN6eFIY5+fUbQlkHA4nF6s/2M
Kr2+uDkdcBIXraZ/qS+FgoCyzSyi/7R9IkxM34EsGvWvzeKHdZASMVS0X8A8+8Xu7WEgRhFA21Xq
y9hl9LDiEZnzTGZ/NxZBl1pe/0AjAGjfTNVYwjzvffXRjnIuuDbPpVbpBRRYacgZWrZ08pfIK6yt
7NrBPtyMyltMi/MeE+aht6dPdxNKDGfbN2kpFIxUAq5sL3kUq50d8/FmoCQzI8xt/fsT9ghIv5d9
Nbh8Rgno+NQW6T4E9K7QItUS4CdLdmljdLkuUkjoaUfi8UIYnDXUJ25FBE3jHloW7dpsnfLio2kk
J68yLSmlnfrjVvZ6/96qgk8BAXFov6zYASobjklbGEdT584R8QmDMZT7BFPHDphOHZPvE4y7ZkH4
ut1XojBZ00QlmrtRjpUI40jDN90vm8WvkV2VM9+rJC+fgANERb5wuYNAY4TBidzJKe4WTjVvdy5H
ItmrpLVSEELEJpIM/ghcRLbAw+cWDEXf0kySMbFl0f4EQqKkPaEABad+a5T+jgGPKIGkfMhEKbh8
6zhEUDS0j3Y5gcfBlP74ode/qr9y7TxTyiDZpeiDtE6oEdySr5sbVY284lOaaGzigiJhQohW8ph4
MJ8mzy7mOktk/7Z8OXM7zBxOX+9E3wNepb5YE6XxAAjXGMZXmAXi+5GWBmJQ7JcgBXPB2pSkt0gs
iorfxydwGv7bUWs4R+A+RnKGpXC5ivX1Uoe9BrZzdOCQPyyy6UZRt92WD5Caw2QF/vQOZICohndv
vqjJrq9baIdwJSDkKNu9u034BkpfHcRrC6aYjNPNbX95GwgdafNiSEcvjUqVy6ESmzILkyCHAQyj
F+mKwRI/xKRtLJOnKnTadHJhxCXszy1NfzgzqpwU0Hi7dUvaWzvLTuuL0yc0oMUlTjPrLELG71pK
eWeXX7ir4AgMhKfIr5ebomV7kbwqy5x3+/i1Am1f6di9ygR1/bdCS4dVN3kR9z5KK6gZNKxYoAST
BlQ0NAik2SXwfBEJ4nvwYUGmREHCCVxzpPHAU6ammAO2VnbsX5+Kxw15Vw7a/72omDAwKtUpnjkS
sBqTeDJKhVUWXfX4t6vkBa7Jsg6WGdeNs2BROSaRQwv6WcI0A6EFvxgjgsGkg1ff10CgLYiBeHea
OLM0M1NXuqUHHPgxRIeYi1Y9uJ05xUm3FpTZEyopm3J9jIg+awiI5Ue6l9JsxyszRpeq1pgSvoyu
I8JoMf1nCXXMbZ6khzoGsCbOocEbnuyjnEXuGyTr3sRQR+6yJaHisdoZyaHkCUWFzl/NFqawhGeo
ClzQ5RM6AkvB5BbQbga+X4XmeeXScq/M4Q4wjXdBh8BOz2sHG7tVCI06InIwhobykRb8xlsi8A7x
FIU2KTjZfMZpsSlQmDbki/E8ZD4UIOK5hmQsmbCC74XmyjaHcK61oadO1gdfWdRdopKUQbDl76Wx
6OCMSEsTyJ/7eBCLG+xfExi2/CSb46XExKs7hn/kgVlBDbXhIP1FucZ1WRKSTiSOgBo5jilyrNAA
ea09t8/1JxQkulF3xqn36iC/hheDoYLe1o/Uj6dz5mAOoEdA8k3TEMDWs/aIzAMxqK8JaXsZkgP0
5KIFXgveigj/eRpoRRlkCrq3HNS0XUyMqtIllKiBcQnlfNaf0LzdwuH0/p3sgzQkgiw2de6AijLU
1I9bbX+Kugyhy6MPE89QBoyf0C6KUVvUUxlpRtqBRdfuXqwCV8UId6kK7x3YkT3eeBFrpOm2vLKe
alwMANoyxjbFmkfUPV9EGMXIHRdC2j+JlUg2YeLSQfL6iOXJguQGH4ZwCy/Y5kr35qOlvSXcxjhx
mJAHjrAF+Bo1EroglIT/Mq7wN6ccyRBRM2VdBoc/agxBGG9/sH8Zvm1mNkzZB51dT6muljpblXmg
jRq0G7+IiWNi44sFmf/2iTH/K/1aFLfHnIU1QIEmBhffI0gi0TfnTz+ilWHjweRtswk2GBh3R16Q
oIWf2/t1v0CErEbHbwqDnkXET4+gfxSqoXVHZdazemr5sgMEknb3RCKfR15j10GfeWwfMxKDksG1
2uRjGpx/RTYoSkdzUJI/HazrfaxqNCTif9HlfbiqaIhXkQAmtK2rvVeSPySuD8fAm6FOZgeGcihx
yPeC4x9Czu0wATC4ptnjZzGuJoZs8Whu9tbDSdnXnSoKmkV1y+HqSo8GZOSaK59AeS7tTyvdQvFg
0XcozJoP12jayRTbocqn6YGI6rGDQrWCFDxwZHhy42OiB6T54pmZtiL5q4cdYewW/NNkp758ognl
aUNHOu+/cCqo9US0Vmllcn6Mf55SrKKJcoGvcpzEplJny4HO6AMUI58BNoZPzx/xg5x4la6Mkh2u
FWI0DfF59UFOKzBXky1gT5JeVotG4iGi2idhSdPTYC2t9zh2JBaE4eUvroxR5Gn8x8QBf2hvoLHz
04ikscxk1bnqEwdhGhrsJNXElNIzgGBQVJvFgx+Jo0XZ4rQR47clm4yzDcOW/oLBI7OGRW8iMl/I
PT0g0Z8ZztSD2lCqtxI42UAJPusiD7OdtCs9Co1kdCBM7sGaOn4xuAi8EKhbpr3z3mwsq47IaTyw
Nh6gSjNj7QMhzd0vzAvWAvDCjvAhg/+S5R8Xwxq6yjRzUFbsX2Kd6AvKjz0yz8PW2hlxuTOJSB+N
xsAZ0gLjFJL9IPdh0JiitDjoNRT0DvQPOKVX5efjt3L4ARyVlFTtZsN3eQQ3VYcKPEShTbsnIfjE
j/dprE6Ea25QnUQbGukj096+/kx687hfFvVV3tAdc815nXLLNzaIbLBBgn9RBG2Yjd/f6azZa4VP
iJXfCOq/BqZUOuB3pHXyQ8d2sD/y/nLXggymMmbIpjPhCjLO8MnR2zGQ8RwbyGOMVcFqtOkavq34
74jLLQ7Wavzn1llHTsOGg7jKwoOVYwQuW+NqkaHYigv7dxV49y78rgM4JskbwVB09pbLT4HDdxLO
UriDuI/g5Ehrvxq4Po8rXex976QkOk52rZLIBXz0TWDV8s7HnO4xEMIXZF+ARFU0jyJlpicik1YN
iBfbZ2uJfr2NIpx2+tK/VriZGORg6EMkPyblz6wAuwSnFwdFqQt1QPT2BUFSsG9kDZZih/PEt7nr
NR9NEd1fPVKO0Pa24n4Wqtl3wAjHeXv/IildNlK5GVtyc1WF+tY4FuRb15IkjOIzxyHlmgBuLH9F
7o+6tdQ5BQZ5P8SzlZymF7dxSsEjhLA5diKvHqPMllVSWg3zU0nJFtioF+rX/YPZBLWBJDY9DPtI
KCnuTTEl7AwnmVEm98VBn2+5coMgPuaHYlyOTZbhitnnCtFulXXJ9h2OD1AcVO8Pnso5xP9oQvPf
iV5iyISr99ui5stszBsODL6qx7Ji37iXhY3Qm9IuWamimVA1oAMlvdp44pXmqfP43xHcBRto7GkU
SADUZ68s7wlpuFkI6kKaVlZP7TTHV3Xjg4FdNLOjVfmvOR9kXXD2rTJNCDMDOZSiy0DgW112IOIx
Pw8Ktk+lrTniMVWyoJHm/NBChhuY6BTomUwcPLwN37a15eSTf2yR+n5sbE/MkE71LC2OBnmvYkAG
MP0SRmuDygJt00f+NjPK1r41eevCG1kA36VGGB92ZHcPrmGRHUS4Qi98ctVhf9NWIHE/x8Rnjc5a
7EPQGWWYhjUTCZc6XeV2KmIpN7z6+xyPePTo4oEN4YUl7OBwdvP238csFq5PAF/E6lc4vAuOZuoc
Tc6DbsSimsJp1jJTO2HJjUyvrLW8W8nPs+QEGzd8SRMo259QjdYMyBbg40fEDpTSb+fHGL1YNFyU
83iPzFlyYpXq7lifPeMXT1PvBqW8H3w43CGkqROovnhBn4ZLfNdW/tYI8JOgkzhuYuAu6yIxGx1a
MdbZvBtjJ+Rjn9mdIPpKUFliX+Rpwzk4qGMKWknll0FnpI0K7qsnd3npb1NpmuiVA2xkgE0frUsj
MPaSRZn4YUEfq8j0C9fzh1vF6k0uhw/H0mkAtWpEpOjAYWk26w7iq8+BmJL8L1e7h8e0iUkf8UYF
J5PWOM2tcy+mfNysGrlRhl3BXv8xbBLujW4SlcPe+AfjVYcrb3r04kiwtNc/BWM0hLnAqtG4uj6W
kqAOzUFH/I7rKeeek4D6/QeBbEFm1zJtqztreVpC1GSxnsFrThIdFSAJWd/fwdM+bGdVytRg0aKz
aZDFg5Fn2eKAdx47t7Hpl7wjhdYJZqL+FOC0N9V7Cp5PTY5zfKt9aweZSBbSn1czNGc2421ZNPPe
teyvpIOqTvyyoPQnDqEWKA3R9iVk7d5/8pmc6rymabb35kosK3cZLB249Alh26OgZyfSnXoLVn5l
OsgzlAFTEK6DSLvZ4jkv8L4Zs9Z6uyZiV/oUjcEkpHoiyMcXj18ZDbyX5yg6DJCT02WMd17vjXGP
9SPQh9x8j5/vIs3GGnjqVRnnHaCw4CsFt81+dllDwGf0eYVdaTM/+tsogyjG9kXrsSRQKqTzg293
wDx646wXgY00uPlWrvMzSyKn7Bjd2N1+ZpUpD1btI//RTgIy0VehyjI7DOyuiZ7/OIwHboR7pzaW
MVRIys67YL9zufZqUhTNW5YmQQh9GZN6ITDqyBBIUqZqpx+4kWXfBnRUQbqB9vB6fK/QRGY3YQY7
08MPJ55vJPhTNxtem+92i9EvVKee2jTuDuITfVnoLspLO3wEQiVkaL/ZDkze2i9dRLLtRYO1SAiO
7e/myxOP3VedonMRjBzW0NWJTmg8lsethfNfzHU+1Zuv31mqeHQIWRa8XQ2nXIx46PbWlK3kwT99
DazQeKfChvewLwiCRbZuhd8UL3Kc+Qd7UAhtRPURgsIyqweN8UK4+QxvIzUT1DRjSXFyNZBjNprt
5Dd3YJ+UpBuecv79z4YVHoc3Xq5uaM5z8TNZ6yVpooo8IOE4H0lZKGZ/9K50oqPsFieTzH7rl8UQ
BjnZZxn8KdLvyxVc91ChfwUFiESO3RfHgbMcaAIGMX4KkYFUlH//PM2hq9bT3SkIA7ciBYzSguLA
vuVR4NzQOqztU1kQfWMQOd7rMkUJtc/tK0w3PeziyIgnY0qycmUGDeb7Yg7m6v0R6EUO0fuh/CyG
Pyf02YEb8EoK+BBnKf6uq7fCfu2JJcikVoC+2Ew95QL/YUdY2iyA43/zNQI475jdci8/sd3yHik8
I3tBIYFKjgMb1gceF6aWSnMAQZuiPrxbD9+ZCQrJmiIkX4Jafe1LczzIEZN+8bU/qGv8ctvkZWPn
WBLKFjhGzSF/nN1aTke08w4KK+4ymCL+R/N2trNNgJzC5mPIH40fuZaGlpdvuvZr960MXjWSK9tK
QpGoG9CwPQiH9epEfQsCH/1BrthCCFH+zlAEakMKBopa/yRfGkDKKmBApaB9+X8n0R+7Po/kk20e
8QbMN7XtR3t1WkcnGpZgbR8EYSGOzWrWDckw0mZVnPxkeK/O6lODElViZCokXvzq0bSkjZ7kZV5Z
RYKkW9POQ4wnk0wzbGIuLHQVvoJpFiBdylj+4B1qVZ9my0J9crCrA4bQwV4SvbOwRo6csj6yxLW4
uXktTSugZcT2gh4xwqtM/J8JBMX2dQfSebenyj92YTst1nmH0rMDIWn8O8j4kzyjS9djZ22MIOHc
MBtsPY49SO5ccBTzqC049aIKacmBymYN/G6U/bG/Xet1ctuT9fL3PEohjLM0owhnxB7l2qXJeqDp
pgD/bRnpy6v+dqf8Qg9+RbqA+DHJFFNP2xFkiht0rTvaloZrT8LYwbXnDkMRHJhGUx174ASGhW/k
aOHye/gRp4xGQGdSy9EqxPStngkNsflLOr486SSC1MyMp6Aeqybpww8gZh0L7Xmpsn/vnU8UpW+P
cZxEZl+2crNzym/l6yF6283P0+ad2zxDtHfVWR+KkyxrD8zaEcibKde4b+W/wQBwInpYjlBUf/wq
M6TLnBm2E24qQl0b59aYNYVt9g0kQL0h3Ub0G3+IP9K0J24nE9gcJHp7BSie8e0wVIzkrlzaj30e
dk0PZc/MzoeCDYUlqxJ2N/XYy31YLgwLgEg3WxJCHbQDhwV9PgPXU0lp8z1q8ngTT8RL+J/qWOJG
bpUqhiVpPbX6/SsRdh4/lyCLgvR1c/ARW18/6HD601Fjk4jV/lYVHIttxXsaKYGOQrUo3Xb9Xse5
k2c1/u8vf/ZJCYauiNEbIp7FBhafDHBUnSSey/YUG8FpRAT/4+hd/70hhsFoly1vlz299W6SyZrx
9uqQzORGpn7nLt1NrsOzqBxQU0ZtOslGHnuQ1a4zAP+0gcNzPvFYbeKsgs5pZQ+h6X0LYqaKDgF5
7Pe8TKsj1XI4uLl6B32CO5wtU7OaHAnG8uvxDCszueC5a4/GET12nrc/KZOVdhhQ3XRqX3P+W1Ue
EjEbsf8SubPLL3V5Pse4ATtE6PtnRoMCJNj7w7KLBY6YUd84GTjx8AQmgJxvpMlnlGilfUmumuEx
UHdOUAISB9yqwbi/3wON9VTVNQC/O/Jzj99/SQGtWTP4RYspMEnxJ7pJrcQ+rBRAx6Fk1ed0b49w
/XpB7eF73p/wJ6Xqum7/QHppvQdDrpNzN68PTj+XvQJePRiPlHtGVsYzB0+adDsDwVPz5yS7DNlL
ImR0JAmVsUi1X+eKHChy6vz31ItI4Ve/QbRKv/8Eg/2MbrDfWpXhXGZKQJEJeBSoIvCm2QbmuNbp
FD3CpudyM8FrUxay3MqriYsA8gcMB/htK4Tw/bwUb4tfL/k0V02MFXlTrT+BU/Sijm+oFJP21A2O
YHMDwngpIoblbm/+ecb6583wU/R+8NIF6dtJQH9lknSBfznoNpcCkbH+1Eb+dgvDMb7gikjv9EQB
hE0xU9UxVhIsrA/rrqiKIhtFt2NrC7293S2Fyo+8GnXesppCyqrp7wXibC21uVY8dRSs96Y1kxPO
YcITUL1HsVndkuWoC+D7b/CLS7UQdulftCPXyhoyHKUl4X/PxbyR19XWUjkcozkTgNtj+bvvlOZY
nVZiAahPHa4ClYB4ePAVIw1FhmafDRSvbBMwpb6L9+tQxs+/LovwHKPfa4tYLsQbho6HCIKCl5tD
G311M1eYbATthwc6EjQq4tJxoKJHwL4BzwwUMBluHGEgNxYPHzRjtd2eZblhskTslscOsNoBA0Hu
xlssW7xpBfvko6Xnaq8ges+ORFa4k4EYGs5IU8M2WxP+VjlJk/NN2O2DtyTmOyYHUVZu8rMIqiqA
YYMVjOJBSFA9QJtaQZ4n4BZOsgA+GcPT1J00bBAUCYXqsFgGSurzXNcT+45DB+7t1gtRie8lx0dX
KslVxLbwLSrMk1dtQLiB8fFPbFKvkp0KEofYMfTuUbFvWXpJDhBxjAAwQ3x51QDv88GkLIxgV1Vh
BG/7NqVrOuEemfVgsWG5nbMk9GMNBKTVJ2Fgw/Jse2D/kRCXk8OgZKIf5Iq17z4IfPxTqZQrh5yr
P1RPQJLBdnjzAOTUu420FC/BORGpogOxbSE9TXs8pGJSFfa1MD/+ZPEQQCgGisp/iteFe7ihSIQY
LHlxw54KyvE28U8boPtvQtxRda4AH9gv73c3Ksxsh4RMZBH9x5laQQTLxdgJVtE4cdeIs5oyCS8V
WYzTZQ7rbfaap5vufo9QgIg6PXqiGNaigx8SEddeBd02Flp2u5YdAmlz8QyWtcjxt0e6ZkfXDmH+
W66jXoSj7VmcGomiwsvkpPP5+tcy4M95u2J/nVVaycOMXgv3c4wwoiYOIgrYicKzGh10skdo9o2i
FHzguXpVTPdHCibT0UlGfxyyTAi97BfRG9xo4Bdy36qKcfiG/7D3rlgWR9LmPFqzAfqA8yULTzvW
mZ8VVb0q0Ija1GJvtM/JR0piEBWr9Pu+3fo6/SnMvXGevODty6Pl0M0wLKRxQuRVPVqziqCTJWHN
t2PJtx0+YEDwNI0Hb2Ca2GeWZwXyJM5zUKVW3lgAuffHWOPPy+JB0hzD42AFjbh+5qukWNJd2lxA
9cojsR/eITu1vtbAbE1dBWy729nSIlC0uwvLURFjywefWHA6uo6BJSVeUDZAlfuielkI8MUFXxZh
Ss1SjZGhFnblXxBTxF6baTBgWvEQcG2LceUO+fhbPt8RuvQJJi0cXFLa2O9UmPs22lvSdwZLzm/D
WAi71lVLnKn1XoytpPYKpo1UOhrSrDg97smpPNewfpDsLJAMXTPuoa0sYCwLC4Z0HtiLHn1HZP74
51XVd5/sQ7ZWw72RGksl5f7fuhEkbdfhZmm8+iwZQwZ+XyxsnKUBaaub1BrZ+sLMbgsG4x0BXZeq
2SYE/gbMvWg7Iu8HL5scbCMPnWeISAWMM9k0XBhHdwhQqIcJP9uGPwOc7N4kjASOB7yfRpPR3qLU
EyvzF8fxHzKyTZrlQtJI4PuCAEEY1ZyMkPRV0lkbDTgUbgBwGDvdvoUmxHGnAtglsuwOEONY+reU
YGX/18S+eOdoW1rKyjclaYL2ZsDrpqBK2vmIjgOj1FFhjIZ58FdvT5SWSN6b9usC01tQ30JslBih
2M/Aydi7RhhKC6tvJadaWWwV2brM3dR772JAOScW0PC4TOHOCFk9t9bdwwtRj0yS7ZFmH3qFjWoQ
bnnOjYM5Gx+/iiDDGYZJvCnJuPGVWoXVGjM127G5OfFX64sKRz2xPHn8WAWz2C/HwTbsmg4wZdju
873SJAWRbd4/GNnp0TIpuMUUAbaj2wgoqzT2NDhaW5B+QgkyEMBy6wmfzlppjH3+6c3ZAKBjVirN
T13tlcu7GeIvD1Dv4UpU8BhlezAmSYlVmC22ci93pH25rI9nSww9hv/A1/aYkzWxOKdftgwrYtMD
lpwyP5wrv1pV/zdPNt8dhegcCajsLj0mbbH0oL4uiU9ovGn9Q9xdE9svD1Dq4B0S8A8gJnK9Y7/1
clS3GJhVDfyL43AjaIp1S507tvsRCvmf1tt9/KZqM2RU1X64oUxrH6h9NwTDbpZgT1ZNYWFKgAEu
oJB7ZmK+9Vcsh/JhblHB0PgyyGB1BL6V0e8JT2+2Ts0txEdY08Do4/UFx2AEaVAllbD7zIljCiD0
pkzzSem7hPTrCFPJgP82Hyx2vOSVgFas3OpyidiAseVH/lYhvE1CyXeW/3g2ImxbSziOH91Li3vh
yfBt9yhQp1baKl+KXMX1Ch7pxr3AnGVhnjgwnsudHmGPdzND3kXe17B+s1w0Lvt2ezYdE/xdCf+6
O3DcZh2eE6Ze0rlIJ01xxZBIGEg4Vs/HGAsuGyNJ8YI13DBLu50OVXWrldAoS09pQy36EcezA9Zq
JprseS9gP5CiC7/vCcmquyt4nrfLsQRgOzXbEH7uFGqqPISdqFKeJQLxfPFUqkHL6zUY9YNV8bOF
VZbPLZZURkuv6+ti/Tba4fYH0bc/3zSfUVCi+RK5Txn4gynpEJhuE5xubedqAAC17NpWSLrCfw1g
wb5FdwInialjAvRgIMtYQb3BRI1OhriNKD1yBK8jM8uKa5XwYSKOBw8x6rRbGC+Wv8+sUgCGIhSF
vD03f988WaV4frTZsNJiMwbxJ1EawiWVgJ+5euP+8Lg5fL5tnMqKrIH+dWtNdCR5+nyholUYbGl3
0xejLRoZ34N0KyasRIKCPYXRN4q8Vf/4Yqqj7wB2wJxqh2eESJ14EFKCJs6rd3MSFU47LlhMH0sH
PUFSsntIcsy/1YENNpOar9VrpcBQLhZYL/xX84ZX6whuGLgp99Uibum/5LW7un7zhljJs9W1Vx4L
HOM/DSRgMyMllCSrRUxUY0Niv/Plx2LnpDgfW2/T1LZFECa8P34OIv+LFguK4r3sddr5J+NVBHWD
WO+Wyq714PdnRdklCQj1gVtPGhT4atwXodntQL1hXgvZwoO2BE8aLhzs6Wy/fJ9u/1cDyDPVE61o
bz4vRM0XNWfXbPKTmo+t4njDeQvJD+WsIqK03Gf6SJMT0hBvi4Fy0BgDwzI800ZQWjzg4ustzaoQ
+FsGpJ6hdqMrMjJKXjh1kubXRllvm/uHpF5wudo4QQq8o4L4b5rCK8Vr5d1ft4ooCHLAKhnN1jTd
MIyeVi/dSDNFYSE7hfbtNtPV5sq9TXqtjv11aGg7kiZc/N5VV77A5SD1sxSjIoLUMpyMl17g8HOG
U1cX8wsiqFzsc3ryAZUzZtBhUvNB30c+l7Ij/9M0AYT1ys8clrAt31DVzkAbAyLBSKTVtO39VlHS
zBNxihyzR+7V+8Hvepk/0O+rUfDd56VUc/6grCO1R0JvvzwY9VisiC5JLn59tckx4ORXTGu9PGx4
u30hodjdhmSmfOq8vKTsj7ki3OWXO/6GKHMJBr56w+rhQIxMVRHE9qhv57axBur26u5Aj+56E41K
yxuwM85G0oF5MUMblGVgh9rIYXxoiDVHnzAUjc7EdR7RbuJThNaDBQRXSeRROnKFCxloiWdjk2OO
RkL6ZUfSQLrub5zZ877bNVzL9pJDsvNg4ua1wMj18J8e+WTeTUkiSZsamskKvwv4YieTdYlqGDnC
IesLoFOSEDGSHPUuqvwAWouhlKNC08N2CRwr+C+r9JkIJoI0dnQrqDrgVTvCrLJL2SUnZ43iwhyr
rYZRVasC6CNBDYOfa+PomqdJxqgcYR6O2pKIIcLB6ObaCwONPhMyB23x8otFM8glWWkO8iMzpLKf
eRYDOs/a0krktpJEiMJ8zTRV2gWpo2TA52pJk6EVtBai5LfAK4xL3EzsGYWCAP455S+OQw1oNFD9
GzarXFgiJtgFlPmabFBogOAMoHeLF9tQO9GnIHjRcWFHaD86MVPrfEUW2gzzxoNqjpQkb9g4UeJ1
A/t8Tcwbh2OmER6A4qvu/zoTEDmDGysytH6aZbKjVtv+KY8dd+nrp4jVnS6kA1gd0YKxKiL5e5nP
SKsdgSwF0JK2ZRn3BwBhjDCWxlV+qOdNzOT4V7kCKimhqxUQ84TL+6VzcSgYYODwgQanGa63K6K4
vEB+24s58sTrxJR8Jf94JIrYlt3EoICyvGX4Q8QVL8F/a670u6Ni3b3ztqApSKacRRxNi9z+0csw
fXF67eYF0g5YrDzpuLFNe/RrZzBsjfDg1mPdBudiEtQBP3s0focmb+t2tEwZ1kda89miOUVbyokE
5bQXnU3ta3zwRymUGqv/zTlwzrmTyO9ovZlOQJb7yISnaq5sZHb7x825kpd3LEl3VshBNNYwTiaP
Sh1uRW5VCYZ/owSVWDil0/8bB7Hhz/xlPPWj6z2IVwrmo29QjnkUJC1kFyUFbkNu9VLlu8iFt4Ao
jlIvgNOxn9nVnBwra2I50jK5pfc8oyOvWpsTPiQrhy1E0HLMvM/SEMeQfD/eriF1VetRgJGoQf5U
qf6K2zR7PSE5dINLORlpzrvYrEH2P36wzOWVEIL/oROS9DuwHjNrMvA3VeNlLzrfBX70fu5DF+jh
AKi5TM0EzLE8f+HP6ylLCfZWhuvUpUxb8SAhY5d9wsvqYeobJnb6hTizNIu3IXgkewVJVkNq9nCM
rawD8FddPPlpMU6ihYFDPrLj0GGDsftC+IpvccRu3YsZejFtP0hLLnUfTsU4ImF6LKq3HVp6rrid
y88/aHh1+qafnvov8WvjoCcMGXKpopMpEYDRZ0ySDvcdE01N02cKnavOzajYRkDE5Eb7zwpSf4OD
MCSX2a3Ef7xXxFpiMzQdJ0VYOxt8r6hUN3YoxrWh3UyKqsgB2vjcbTCAS/AIl9TjLboTwmdCkzyQ
T+eQtwsfRbXqOChcoQRFH203bfKSI2hMTg3gCosNeNef0IYGVgPK4UqeQV4j2ommlNcGua4zwMZ+
46ZXbVclRAYDUgZu4AJRTPyLg8Z221MO2oGZuOvXN9lDudJWysy+ngnjXX2Cp3CRJy8a5KBAmghZ
+1bYgnN5N40h/WF7W3p8mavmmAn8DvNvP0gfHP3QSGPmAwQMYuzwr0STAL1C6Iqt+ZKZpUBmtJMU
Sz3umzIGWBIK0QjWnyGNBwoL7dnFmRpIj+6/FhHnXXUAS6uvKzB26rX5SGweTaedlEKbSLdH3LLk
D0ALVUbkHcGOkumsyktLgkqWUSaK4J/tKThOpwXu1yVlwxCV77z4mvuSYWCxt8Uvm9KP4FhFnl+i
xVeoozjdPyGts+pIvZACZUjQrBXIZj5MAoG2CalzB5rIG0Nkq08qrucJpEh6OeID12UN2jv5WS0d
imDuZdhm8maKz953jK+69eZpZg9y4kUjf+f7AT94XfY1p35i5GqbiPUJgqOgWzzVryk0altYilO8
kPIZF0Z7lhss2Mfa4Q54y7xEVf+NyGpyXneAnhaGhvahMG0J80KzYUID76Y1rVmJCoC2oKjY2mPI
dxKAStIo14bPx7g7iaBJQIpfhDTriM9yANnn8VQYaz09wJNep7Wd67kk0y1FgaskuNtUPtyEBVma
MIRev4YR0I+LDlFAaRlatsA6TSQMf7ohDDwJ7cPDEz/mmQhkj347t55XtfG1+0+dSmEgUjNLxdEY
XIFEhU8a8Hr7xul7LZz3cmq4L7FlKOUXJwZmbVNPUCixk+Fy5IRoRBOm2dncPXGDZeRikwlyiu7K
sxliDRgSRGHRBXYrLHTAKasHINpSYqi85oz3iEjHgPohTdZBReojkb3e1Vy77KSE5MvtXat/toTD
HWA1axHEQhsegtC4Xd06Twn9XYKdIxx4q+4wccbu8NearRXlaMVmNxEQ+GAZ0ahKnX8Qi42sY2ha
mkTzzmkeXPSqt2zZaDpQAwlKIumAGQJZFaOndeIeHWR9wJvWUfxTZ8fB2SBI/DY94uo8lAgRID1g
g2TOQ+vzfb9odkmO93IbiAoOjQGQu7nolP3fBCz0Px1JV67780/b/V+F5YVesGANU0OXyw4xdY/A
c8FzOr/+WW6Q1DyaMcjpPfIT0y57IBszWhc14oqSItQ2mXmJl8BEBg5/zU25VCUlEceiiocfuhQ0
l+llnVJWSii9g+wXmiZqKZ65oSGY6KGxPM5FtJBof805zWb6vP06E6xTdv/t+bpGTclXirtC1nJU
EsqjZTr/Bq2ltGBCajMcZh4quCUj179mMI80JObBSg8uBUiA8Uk2aOgFzjZNuSe5O79iFNbZnRHZ
kKBOFjCU+rBtwDl1VtGbP8j3OycD5+W1/hkEcAoenn9LhkfFZJPLGpHVHp3Zmu5wZy27X4+zy8TK
v49MJnSMNjeiHcBdqfFW37qq12z5ye+X3XNKxC5L3W4DKQ2tNVTf+o23VANSngh6LQdpYv4E1YzI
3EZF+OofAZ/aKUzD4VBqDpnMbqrHYi1HRzje/XSuTrDArJ90PQA9vMpb8H0+pmSF9L3FkpbK0+qr
j8nJQkzVdIxdkxUen5bl6xgF8ui9mC5qOLzsPIuU288yR/fDoCWXybqMJJecF3JtvMi87COqmJt2
hVbZEs3BRSxH/yWaX4nyUeL4ndw/i9hkAji/w6JcEEF/QmfisRFgJxQHS+g9xpYE1xqGrNBhJRQy
GkT8V0fPY7DqwGjuPjEM2mZ+V7KHNCI1VISEswiiJRqmVzkCtpx4ztv0/RlYu/G/jcxvvicpJb5O
yzmjuWGqQBM/cy/N6/w83nRV0v4EE6ejaYSz1LayijhMyrBuhXGomugppwcpTShTiVoNPl2C1nho
LiiWddBMmw0UxjN/eNnDAQrxLacv/Gm/6aj3xA51GOA/yVJY+c+gxdaMXpvCqdtQm/TYi0ko39/U
0WaNUWjzmHUlJnyyMAWcR5qGOg17exKum87bI0TpWAQDRN9Ga428429MegABP39UsCzLgHnBqoyO
I+WGJQlmaojIlYwMvGPH1dJPxsGa7hKsHNylfFQKXcNI2y46FTd5QsWSZaayS7ukNVT0IgSX7HGQ
dcAIxKiJ8INv7VyMlEn0IJJVr/3VodIspG1pCbO587Lw9QJJvODA4kWO44xBGXQBQM7bvw97+x3e
+ANc5LYTUfFS3N/8Qv43rm2r60IkCgBg0XkrjiFxEAGekFw2426A42E+9mOh9rqN7kRMvyhY4HXV
JeHAz8V7lyJMSp2dreGamRyksZwH2EfOw0hDIquFCMTwlY4iqqhR6qjhtcWrJk0qHFHVvaGpER68
OdEg4HrI/3YDSyaxm1D0u+jbyLaNq7OwIfiX50lMUWM8PaPL8TD8b/jcROyUpsLx8GYGlpP8OcIW
3O462/TJTspneXfCTm3zfQaHysUoI4c2IHUw01E/kfSLi8yUOqcWhSoRVksgxtP23FKpBVhkrfOR
ewnXsrAJqyUQZOh2sqd1XWhDg+MevK5C706xCGqbTWzak+2UHKkWW4HlIYqVrlBOM0USXRygu6+t
xjrSnX2tAWvVAjZTfSWIX1+F8dV5KugZ9stTqTPt8db1w5cTnhEAjojtKIhTBpJZl0K5yD4rJg2n
vfnlntwVH0yECECtYDdfX4o2NqOaB9wE+YocYRrLJN4nYOq4wC99pj/AfigpElUUG2PXc19ZZvK4
RpCtvEmr2wb/iu0RyzfhEQMiEQ95RlnYmUdLR2+JF6hZWzFfEnOcNuObGX92Fp1ZrzNE3GauAVvq
DJ4iXZfFc5rzhsfkf0s1/fRhRv7lCLpJbl5Kb606u/yUVB2qrV07/S7/qJnWOHZRw0CwZJrwCKS9
Sl2t4DNjme2naRlKMDO/AMmsRRmq1ruSXyxzMcbVV9E40Ly8HgMxDUt1Dlgo5owcyZUYsdXka1mZ
b8hEpzjkRs8AoPgTZ39QJ+TotaIJuuANTPArR4Ua9A2ATajJsrJsSI0sRQd7t0YA7Rqb+W5A9XU/
vsPYbighlorA1qAWTtgUnASMJZgz4xvY4qgYM7Ic2n8Sovg4/zMxpDljA0HYJsf01VlfZQuEJj5V
nyCq9djU2r8MQP74bQRIcTZnSsBneuG7LGDWo54k5bOQKIEA5SvLIvLPJ2dBBy4wNLpKO1r/7OgU
TILh5irYUWhXT5kZdOgbisamtVj3dCR4yvzVBipijhWje4d0cUbJOsak/8521eTbbkkyJFHJOYoe
LSHByDd1+N2eTAmCCfTD2jlNZzOaMB9oK/ujw38JO1e0mIJdDjpure9RD5H0ucO03s2xt09/uZLk
NKPTH2eB2LWyO64lc24RYqj1VhMtOr5ilfqq4KFY3h/SxXPZEWsOR9f/I4jJ2a64vI+fdLWAs7aW
udnvHAF/gThpZzrUbiWrjK8tig8zJLBYk0HBRR9DpjcoX19n6jsDnu2Kyx/YmVuFQy4lIu+Wec9r
FBP9/nU4zC7mOuDwCKqYWiBay+wHNGCAWNXs2MrHSSpfF443cyVh45XLTkk1v/3eLR5kWmoWe745
9tuL93Jn34almtGtsKnkLASJq+NjbdgyoAqi21GxeBdFxiX2Ut33Jv4I0emnj4jubfVwTfkxXSJa
N7gW+ArpJk2CVZLj5iOrLSJq7Ouwpi4H6WXpdsTE9fBQEerwkb50jHqZw90kADilZb+epIiV7As3
pklWSWlHqopPtaJhWwY2wefZB6J3b6aMYQ7Iq/ui4W6sVLP9tXhNiPzkJXm6OXnLhu59gPocT9lu
vV4N9gg7VgaB7DF3iaxINvhTT0gjyvseR7HX6HXjU4hdmhihg92BJAqaVuuJ1AKSzIOn2u4knAe2
wr8zhwzXq4pqZXLuW/7edwFCLYKxecSTyEM6NUrrDXjIzRM5lMpgYNRflocoygDZjTAWIitrLMjK
NQFUyBkT5S7yQ0dc5ft/kcNjV3VqO+fah+84WyRZi0wqiVDSsk5Eh8lOWmRCLYd0/5Om1bRK3MIK
b8p3N7REjTrH4v5cpVBl5s/hbWvMalnBmyHStFq3bKeowPfvXnZ0ntT2LuQlgIgUsnscjETBYKYM
zPnkb4Prj5qvb5sNxAdJTdhE09mdSLV9vv0KzdZc1vwpBYGvDr6LeNFn534Y0ptxFoFp/LlhRLAS
ktTsB8cmeKQlhWOETzOEy6mCu9OhtLdLCOL4KpE/m45hC3/lvKXTsBEzfAhY55kbVmjFr46YBewY
BI0sVDOWctrycwSab3gAQ/jgSzb0Zh6kynzqpba6q83jVAAuwU7kGCEID2I2xHODFNQjoX0V3j6W
/bJxyRVwGI0h/izxO/s8ljkGbtWzjzTlZo+JVBSQM0Zv9uPqHEbYmdRY4ATPbaF2Zpt7Thy1EnXz
csD3j3kczoiWtNJhoYQGSAfgYCKHTDVDDQkvbI1tt86Da+oKioWGGpBdRtzXUf+Re/ttlxmSldj4
Lb4oX25ndDpZ0GhRpx5Sv68cj/mQDcIaWy6GadggdlthFc1TkGM5HmztsDpGQQbmL+w5RAEKS1Jy
3vngt6spj7s75Omr9MPoXehaxMuAqnTAOzuhApBdh5yeSOtPbi+ZPDTAllvjNE9eux/gL45Kavkw
lqrrnmrR7BC39XytFlgCzY3GkXFh6iuYI9Omd08rcU5P23Br8Q1UmfLLshGVDPNYwKU6wNHV9rYx
ogFuyKj4RYEKue1ImZAAw8XRTy+u1BkPwV7dP4V9MKLyIv1nS37Fe67pQmOnlYUJEi1anf5Kn0pC
2aAPyYIL0TZisEc6UuZ4VToODAYO2TllItZUml9N5azjOaYc8FEXZo6Raw3KbyagBs6yBoOl7QZt
s8o3+kqg9A0WSNfZBye347oBmQralsx9cIpv0+62AythuLLQEgbJpdHdPc/DAuzT5Rgo/Z3aVTt9
IoHuniOSBsBoXWG1lOi9ASkkphXadq2dnu8ImDAVM2f7Jr/ctR+LL79VLc47Kh79H8XhMX7fycWF
iwrBxpIxQw/frt3apT3gG3EdVgm5VmXHSVaC9gz03IWlkJrGWn79toKC/xk2Z2GT+uHI1CrH3gGo
NfGqNhLhVpUDLgIsIM2iG7RLL6O3tD7F+COSZ85xQVtpEq3i84Ih1cxuPPmLynEZ35/DAjXruFwY
BuI5TSkELX0zyALcXxv5KHkEXAcivXYDIKTQfbZD0X/RJ9XUW2UbRX3W8SNjeMmgjYIYjqi7k8Jo
KZ9xMIod6BNr2FU3hBV3e3+5XLb7RYfta2PKcNDT/XVr4uv5ERK/4o5m8XXu2gFqam0QtnDTEsbS
OYQvUlEuVihgf3nMyfjHMPYQUGjlqeyHEsVxAFYVQ2NamCmVK6Ri7r3GrDz5w2X7x+5nktyrZcni
DlmcdnBzSP0rc8B2x/W+ugoCotseZIct0pN7ihU/qOVLehhA/GK10xJDw5j2Qz/QUEY2hXGyMh3U
9z4HQzj+DgFLVS9gfRteSeRDV9VdBE4/iybJrfpt8yoy4+BPfwp1hj7Xhb27ZtQHB0/z4KXqircV
59rLPb4pelSX38NhxTE5vZs6dtAnzNXy1G+tMXUmXjSxXufls+h9Gi+gNPb2WKdMtP/VGXX3bk3Y
afF5jb6cH1RyTZiKpq75FUEzc4RRHFSEkHs1v4H3lHgn5csnh9ZBhJTIud5EtiZILwxO47Rzu2ub
p8KWQUuEqb533/7EapbFw0oG5CYpKTApAiLeH4DGncnminvVrUf9btG0lZdnrX/Gdn4Qb6mkeFAz
YRwG16ByDlabk5IZmJfFU6UpluZ9Qop9hnUWXxj/hGU7ekY9NGtJGJPerHzO0hu+oWTUy6tO+YY3
Ajs7Fki6pU2nD4OhdieV6X3AbNr/DszaC85X3Ksh6E9nJB0GXsrvqA3zdlHlhP2/JF2hywkw0Wh2
7wi/rHbToboWzqNNfsfPJ1/C63UABhdQbh3bC3JN1/99MUehXtJLbtUQP0Kzk7lQKCHIE6Qd/bi0
MK+XGDT6ajAOo6hGgxiVNNdGbv/o0lrAdLiybEYhSZkg2o8YBYVj0smd70dREloiJi7RpWCwPN7M
jA81G5W9ZxNirecs7b7Uaai6D8ZPgC6iPnm9uD3PPliJEDUtEr+pzvIxdDenRJ9wygSR4CbbJigb
a/tWJb/Yle6r/q8TEYsxZKbk1Zs7q5tm85O1ByaiZu6wN+nykWkFU7A4vJQuGqA2r2FL5/ZVpmw4
J/gbsQIrvRuocXI2ozArs8jgihSKZI9rKoINtqiz+B5MiQ6l97NC3wRE8D5q8UnxwFdLZC5tqMWp
t/w+TyERM+2VTQKbjj8DlRrl09BF+CevLEIS8llMDekw4HB4oz25v/Kybj1fEEtyhC/O0XTcvzRq
KE7lXpw5iUjBNdBujSfZf2QnrMQG+JgTtjZ/DJXaqyfbysO+6A/UDh24Y8T4h5pSFRgnbt17M7HL
uaxiv4JWh8JJWVuaDCZIKT01Q06094gbQaVwmzHa2vqNMBaqvVWh+tYkucmlGL5Hr9J71Sxr+ltb
bw1PrtQP2DXpkToZ4PvxGKDDVUjM7cxYRrHi1xIop3mgXcFys6JU0NEROG2jfSlYq2A7ova/wteb
zDG3Ijx3hjFoa21UamzuTWnyjzpRm9Jvz0wqdZv64nmzQiWa0WZ0sCKWBSk3mJT3rwqbadkVrUbG
eKj10YLxQFOs6UrDgFcU3v9XNOk6aQR3PBnDRfHnD03WIxtcg8FSfbYDaAqFsYpZP0sjytsxVoa2
j/I5wsemKq8qd4zb9sMUPDmFvDJLCM/FL52+o7tbcFbKAbGFSQp7mwX5prbKsenmXTea5I6e/36d
oQOezPjGUaA+sE8R5nhNfogjHC7zO7Ik9k0eeSXoNF8/1+TOisO07MgNhbNmk1Pxhe8JUNgrc1Ij
btGU0vrUS+WDdhfCtyZwlR1wlM5nJRqeY0z9o26io3PLZoyIwvxVUDFB1qZzm4V4Ci95hMUTGh2e
Fn54UqHQjxuA6mZHlbkoQcyFrdjaGILPbSRZEnRtI1gnrdT/MgqtCvqqyL1fKdsLqdGKlRm+VmH6
EGXZk36CE0LstCTNahS1dzYgLSo2WqFaFzfIy5GfOWVzd+8ARP+L3bdhN+eDP6IVCU7oZB+SuwY2
UamIR6oN6oJXYDESCIikX43LI9l+9XYM9+radBp3B48L81/o7TT1cAtIz3Dunc2wxSU9ASiFSnKk
HAU9aPSD7wrWhuLtVlM3k1k4YthlHM64yL260W1CNNykQfZ5mSIj7JniCtP+eaTQdHm9xHpPwMFk
DxR3U+Su1UgCu0StF4i9g4st0Xru6kPvIcTZw1z4Sb/1d/IM0so756G6gunrv566ORhYg2eETlXN
jnUlQvJB8wpRwx2iZshR1xIknVdJksa7PmcR8Ohl9/clHpNdaBOHcONwasibxM2UrvF/fgagXej3
VFZLpgn/BSlmiGo4oD35W11v+dQwPgX0AF9oU7QP89Cdvg85xsFB9uh8Xhn3Fx6q0LnqVrn94j8k
F6UZVhtEKfW9qpVng63NXDqs6TJwqHcYFCYkmlEup9FS3FNZLYyoAalJXRm+/z7RiYD6tkJOrVJN
uat8p2c5N0D28q+ZLGzWDY53hCrxHm5ShDTvAgWWy8qbQpyquLH89+b9ohZTLIiRTfxRu2shtMUe
zTXaAHBBsRPLgxkXQlWhjH5L7M7U/3qgEGT2q3VBCQm4D4dbk6Te5qLt0jTRCG3nU+1cl7PO4bEI
JsZEmT0jIYhqkBvakSoNinUmgCQlaVf6tILriyWAH9ll/Jd9+3zRuIJpf/8YB+P+ueMcBaIfSO+s
EfnHVH64ZOcZiPQCMtWlNWhCTuePHXb0Jkqwdr/p2KBkYbXxvdkE5iBTRpNxoGPT3iZPQLferL+m
FYS/mdGmqXn4kUAgNpuahVFQ8AVyla/MMWlye1itwp7q79sIpO9acSqCvLZDENMt2Yd7vRqFoe0p
BMOuJCInhEdLvZ48HSaOTyh2W5tEPrdjzUGvr+7P+JhXYT/BoWChaqGM7XSmUmc4Wv+BjSATsdL/
GRjVm9eqsW8A3mIfI4bY4IVw5J+ZMfp+ZqPR4k/FH0XMnRkArpg5/vpYCZK/8Kqv/zbxz4SmU0Bp
0EC2u0HKKzf7XNLX1LPM/q9mDtH3S6WOAuoCp/4EWWg57WJLbxQhaIRt6Qk9iWRNE6/OMWXLnJpV
taVAM4Dbg4quR3jvdZ0aADMLS2MjVklNh0iGGGXfrf7sFHusMeQte3bLtPgrPYnFmTsuut0CfcGt
G1XlP0V+YObc11NAsNZilv/nMeSs8MjmL+kdb8G/OMHE1UichDpYvLP9OGNzybRhJjBOJH0cW63/
gqbvmlaT6yNehIqbaTlqcYtlsEJB874H4g+yUl94fi07caNiUoLZcbsqZaMmJy8QJIpO6rSsGMLZ
PM2ncBKn3K8c5iUtkeA6UO/EnEuyXClek7zhH//1jP+G/Z/j4hXrcpQG7aayQEqDYfPjjI8pgJ+H
ys44tROUnpWJqV+jFMj/Ya6mvGwkl5uPcYnbbw/9VgMOxqfOcX7hjF+8NW5Bezy/tXlDGgmA+HCq
PWGeKQDDyiZbjs49QiJ0VTbMIPVuesTJvtM2+AQ62uEmsW4xWl4S/pc7Wknc1hYoanGWYTNAF5cC
VstdvYUZ8WsOFxa61Ut3VhQPsomQOxZEXkJ2bUA4l81GZAk+tSMvfIA305m6kXD+geKtJKK32D+e
uV5cILXSjNINBnAn6/2BWNnsrhUgMi1q/GiJq62n1UwnbvMxDYpjdKJ1D31hreH9wxM825Xjgeok
JbTheuHWcnVWqbEEeomWZ8XgrQWUO2cO+QMnhUfmb2siJZj8WzPjFJHxikei0LIgxfZdpp9SuzOP
kb7beCkq6uHYwG+cO0JjfHyeQLItnjPh69oWoFvApyWZLfD7jgugiTbU0iv+Tx3q6yaCQzHEKbTf
8CdILah/yjkwSsetOiXb83g2PdTkuYilHcMp0V0LOnM/sU3c4M6sIdVakURwUNMRDFSzDUuD7BJY
Vi6oNvckhvWY8aczsAuoCSDsFJaUDYKPt8vDDEB9VAsvqO7Y7oPTAFcubi12DAi3x9ls0I34Mph5
DosNBQkCwP7JRTdd4FcYO4KDAN9rp2KPoI7fG9BnstUA2vcuv87LiWYg8ij66tf2SFOQwsoePZ8G
6mGlsJI0iib2R1yqiNdMyS/WmsLc+UxfAcq2df1F1sYuLVsewHfUCmxxgogsSGrweKxTIpHoXwn+
JTAZkyiEb8kVmBMfs9DtItzk6iv8gSWHMtPz/SqZwBgd6edmrzVLZXM/Xt4KDoKcF6BtXNzrr2EG
QA5mz8g4OhMxmeuBmIyNwjAMZn4rcjSzoZVRqlZRKehOz8PiWGCY93q/3YRM1QS3mgQQrRXP5kTf
iu2FM9kQxtgRMkZ+IMcIwdAIcOWmSyQ/o67PghkCmUTsgcUQ6qxsCy9t2zroOJ1Y8Byp8JN/eQKC
/gRwF9gFb/y50Y4VdDO+pVp0AlE3eG76m7RF3H08kX4ETQJSTYx6fhPUp1TdvsLLlMZjiAjCQaa1
S5ARJDnIX34Ot2GaAqWLdboS0Qf5HZsv7Q8gPwi+/O87x79sZlky9SZ1jZG8zT5nF8ZHuhn9T1jD
4paXIZxOWpUD1aSmBxmLE9wSGBWI386NOOHgqJtPBwfH0oqcGUpfxVOvBbtWSV5XeeCY/sIz9vZR
+lnvor1XarZxZBd9Jn5OQSu1LmhfDgqcbwhjVh2IBWsyhgi0ugOl71CiM0m4xRC72egOVTOrnACR
5fDp+C3e2sB6f4Ugu8buow4FF9EM8GoHdFn1j8lkk29hv4PryuVHQwyNd5cTRyVr4ienzOdmWyVn
ybDyfgfcoA4U9lPJL0s+EJ7vzx8mBfvBZ9AwXDXfdDkaMSCGRKuxlhtuX2a6rh07J0abBFXOTVJU
pfeVrkEMh2Y9VVu2alaMFEOYFjYXzfBKoF7zfR7KiRYr8OmtbeGxRAbDTBYeyRxiESxljgQSh6Xf
clMV9OuYAz981fTrXuYsahOzamP/GZB8W04h+DoO8g7SkLoV/FzNt3z8fx8QDZ9M+MwgER+GNN4d
QZvYk5uIwcl5lPz57WHzQABG9Vj8qHdcd5vXjcvq1BopqmbKzT662Y6utCHKpCcn6EOCVmKni7kN
Q9qzNb3AqF1d6NK1rmCbokDT5ealcYxoIWAjfqz0nYsq9xVlXvzcqMzBURQzfFYR74DoCP0fvw7A
0+3m2eqXwK9IAAvGLKKs4Xy55z0ChZiGn5hpgvJcbr64cwQ+tFkjZUCjOqzbHIatYUW0PJuvC59K
DcJAHx9COCL0giNh3r2OnJe6fb1ji/eS1i67ErTn7lv+kq7kpIgIbLV1rHzx7Ff4+d1PDghpOKbU
+UgBYxaDCwT94m+V68/eksZ+YB4Pb1cOXCMZuH0s2H0SmWA6S/DSnmdnRW27PA2cAdyQe1IEFFmo
9Djil2gZsJ2ABWsHkPMGXrKSGmBWI2nbJyZDZ2bbcNT0fMndzeqt2EGFQEQK/MMeMiI3dmNnyh4K
sfz8V59SpTR6Bq0ZEtUbg5ZbyeCRrsTFammSequeRPoX2Aw1wfEteNqfPEAGfikhv7kZ13DgTWuc
qWwAOaFfXX7dfSfkb8NWwZMA4YCKRD6fKIfJV/Xnyd6yfzPAWK4v5wYgg1yZVTW+Y0wTVqwnM1XA
ho8uVgsxmKeBblAkrsnwGeqITCyR2lSPe4Et4sAex7QBE0C3OsZfnWoM2J0jGl0t+/YMB+ujtiON
iHEQ2tMaXmVYf7GFr9PPJ9bidd9p+uPgS4QUu1MneIFgHxUziXBxtFRDZrr+qviWCAcEY2I+suKH
FvfosafOSCbe1ziDtgqZnF1KdUDnP+60QJQkK6MP5lL4dRlVULe2Mci9zqlms5pUenFyUCYX+G7k
p1GJOmxjIcREvNErVleg2jP9I4UE+Fpd3fuZoircBnqNUBxzrPKGipdkM1PqpzfbS5J6x2EVCmx8
5RpWUPYUZipCGoWuOkS7/cKhgfKDddbycUMWUSIv8+QfN+hRgV1g7cMlyYhgnWMniMgiTIuJ62cm
A0qYy8LI/M4EQjT/6HHH2m/RINXUCHR6bqIsO3D0f1X2bPmHjFSaR58kxehi471QX8dwCLg2xJfh
g2gBo1M2f5CCKIVSl4XRQkDx0mR74bMRbiBuwD5orcQr2gUBbG+k2PpMjfEB0qhMpwSi4JMSH78N
8aXSuMF7JawLdTTvjzO6nSCsDGYyVMRLB13Ho9mv0h8c5AWRY+JcgDrV/D6qIK59IjqXxho7M++B
13nXoIRXYNN7o0eoGn06JgDEs6caMPSbzjNSrP5eRgfdQWFWTqyBES1uRVH7LVenghk9pX1aII3z
FJOxF+u2F9EdZAE5hnqvaR7kPqAWQViKx2wgVuU49+KKtqj3vRhB/zj4u4REls0hgJgkmuAbfeu0
GTWG/cAc1gNeyn82Y2TtBQtrlaK0zXuPgPg5Rm1qCbe/FX6vjILKYtJ18Nq81M5yZ/Cn7ktJXjAg
e6Q/SRFygSy6ljOCjCuGtrk0gQMaB954q5j5xY4f8SydK493vUjJpAi2EDmyG7F3F2n6hwscfH09
gh8NdOobDFj0skcpqIwtBVuV01OfUV29Ydf5Vz/AaXYcYlnbDQPoHq4vevYthuGriYznB+NfFNOP
VzlezLwyFRfH9dJQhHD1ODWUhRYIW5DXPP0FKHyNzGH5xi2RIjYgLBl/6ETS4zEwdKE6VTVf4H9C
hLgsH1vduVpW0L+IYGrbetNM27STXNSjYBIk0EeyD9f88EE8T5OceA2CouF9IpZoZ+P/0JNpb+GL
pKy9fGNm5xc1rxDlAWi6wLRNno+9WCn65JqxFK6sx9J4TWmhfiuvAhryIFlkCnOqyJ5eMY/oAwtK
kQNT3fR3eibIagLjxSihQRANHPmYE5jV0y0A21M1bFfUPhDXyP3GPAgHMtWaOY05G7rTGM4GW62w
e2X+O59D8b19sV9Z941axutJGpfbRlbpjqL/yaVkkpabRwcG90qZtGhxztfeROs6vg1eqyBNXwj0
ISMtFE4tuWmoTdRcGT4EtXIJWoEm5ieEhmmcThCYNDTs5dXZoWboJJ6AT7VS/KD9QtcyolqL6g41
b7xuEgOWm96iurin5X5/pUQHYb0RBxomkjh8bYa59Iqnd+TJo1KRKW1IZ0RNb2FnoRFWLLXshoCV
arngTYhC3A4iqrQT4GHeUkoRw7C752P8K9+CPSOJbhWURVT8pOvVfo3P1yrEhgLZTGemU9N+Y2jV
uHKlbMdytKHU0saATbflXpVvYzWjXwMJGau/MVRyEg8uDDNjtKL/uELAcoU42/G4dGtSXaghRKON
XExraEE7F3QiiMbnWOgcnfucxILZ3cGiZmWU5vJjsWXIwIbircSewh0OokHtv0evtNz5q6N1qnJi
cWlhkyqYG7IuLR5O/l+ITAVvU+OrwZOXOze0zi/4fby/L8fhgiiSnQAf+6RxnOZMg0h5el3i8KOr
lYkXG2SP7yuDjoW8VOgN+cTZVfFwTcVLtkvas/88kPid4jKvbU6dTIjpYPePHvXxlYimP4e5xUfU
yNdk8D8HvCOp3gy975Rb0Q8qltYyedwr485/9kCr038EJM7raofRNOmZ7PEZ1q+vnkhTYLEg9+hH
qtWFMH4vBnY/bpyOfslS4AQJpo7l+jfOV3q2kMUHvIFePWSWe2G7pZkpyck8x+JMR1N9P6eky2qo
eOkfvaim1OgFxLiL6yrorTIqhos7EAJ0LkGtA6/Eq5NJ9K4pStF1HcD1zqonJ6fJYPwRjOq/fzA5
EVZ07JoI4gG8R5I2PKONGQxuInqfm3sS8G8XgKn4u4EmKYXcRrRLss8aBNdWN1Wa+cH7WhlpKU3D
VVdCjd7hGZvqaUEpA4tW/G4/du0CnOFgNegb4ptPYMJ7DdanXenybWikJZGDRsQsQO8nmbUhPiHO
xZkdwCf9+O7gDIQFUjId+NuKnfZNWRkIdT5zqfrAowXdyHjvtsyNQaKikgTQw0ZyCU5QVdRNq1j5
mNlOb3HgyOx3O00ediza8KM5u4vgjeAfRo0qN6sSIUzn1q96jIBxQhRDCeC/HbVO8QyL7ZGe0VLQ
QY9gwDOiBaCsTW73albNzaKbaWY6KuLGa8bC+5poJcBm05QcL+VceYmURmSUdgc2cWS2WSUg8qyw
VskJL8jOSYGlUyTjjSjFKj2/pC357jSy3pwg8/7U/oxgRYHdtXNZOaIikh7hmP8SQjYmQ8FE/Pug
eC8CidtvrvIDqAfUP2Arm6HdkardJnqY3gE6Pp7mmffGrsNjZYEi5h75AYqpLxdpg8K3LjJTylpA
dbxavFMvbiluskyel1Mlh85vrZfUu0WJi1ecq0b5Z9xK8WvxbxWQ4W6Pnb2Ya2iqI5Yk0HAG7kgE
6fNahgflvVZvQ3iAqmmgof2B6tE9H6w/ruyVjgkbZIJhIzhJ33inA9wpw+EmEkucmAIysEIQi+H4
bkZKUVcgf1mDTPvM3YwUyMzKPAGIERZj0/DP5VpkCzqDx2XZticwxT6gZAZ4GZ/90Oh97ADGo1dp
TiRGcbG8vkAyhUyplLazn1lyZWXDRMWQaFQNhFf/mObZA4hSM1l0CM3ETQBF0X8dh2sn2QxpIxdO
E+bJ2TPEj4eR2HrMvQ8Fv2PcfZ8XSlW+jXC7pILd21eiI6+S0gej4A8LwyZizOYPEDel5mgKvjuc
DW+m2MxO7KzkxMj1Taycuq8zdOTF5cnbpwCSP0+Ntg0jSbDwakiJMCknZ2iLQexVscmJuyrmcy48
gQWKcyyMzPHPV/ikuQ0Tdm8h2JTDrFtUFhcnZTK464VQEkNeO4oJrGiUECXMolh69j3sk+NEpg2J
wu8E57q8lb9eYRSFP86LIv2gJycRXIjxCc1eedGoVYU8AtDAyqLb8baa3EqFO5bESxbOBj6WzYCP
T0pZw+PP+yswCsELe6I6SvTjk0g6cUSU9ahD3SSgiBkeCRPh60iNenum/N+qtZ6naUkY+rWDyNUA
klc2oWXdbuz6rXpbRAMdd24zyDLZc0xUjycyAL0MsB4jtCRMeWPlGRxxb5QvpiKx3b9lUfOqgS/A
KqzgwYNdkRMpXgpEFIydqomlKraUJ7MoxealwlLo2euuqOeEI2WJdmYZqkg5KJMNKm8+fNO7dYko
t91A+8kS+VcYYJxOBLJUJQrpH6QItJpFE5ccjKa9HD/gIHpigmBF8YAhDUC+UwyAfXrhb/v4Qz41
J3Mb9QTzFZFt5QDDI5YyuxpK7SX7djWKtppBYveqmo46Nv6C22PSJSqDPib6rM7XMWVrvLEp1X/d
X/Rqp4d6KN+O3qW0jMOvusOvWx16HCJPGecFcnxIcwP5gjdk8wOPc4n6tWgMbDNkETkssRi2uWbR
rLD7N7RGwG9w8LTVFixdLpJdR9aiY6s8YF5o5RrN/sxLylB6tqS8O9GLIzYzs39sXzuamX3i+JQj
L7EWGZFZMD0/TjdIWrERwvOueakrF6ANu0OikuxCEKAVk+At8ESgruZ7W0lirg8vfuKZEBcEiR2z
+OXdH1zCHLGKqA1OtFy0F2soDtidofZcjp8fADds8IbfWMAiuKkqjMD1WiUh//h2k/2yatF7fWRD
4Np8I3XA1zE6hwbDtRjST+2cc0/3k61MjqIvsuc8L8sY8+ScNQJSEYpYjGPJ0lfZaEsDhehSpBCZ
1EuagOpIe2WaeXTrEBwV7+u+rykU3xVKvVR7NMxTWmJnwF8HJLkrElUTpWrAtPtl4Lmjc8oT+g7F
Dw7l6LR1P/uJxRgR30+JK981RwXQ+m5yu+Y9vxjA0DMMy/uomXHpYCua8w6g8csMO9IZkA0S/f9A
pFa7Rlc8e+ICV+ha1OYn4PN3j3JqIGcZWsMSqioCREkYMFI7RMHxj41hZb6gJeYT94154Og9H4lV
DZSuqBa5GU9WR6y865Nkvwg221kIqjw5mJlsONSbLOXkTjpLTtuwrGko0EtWpZmkzuIkZS8JK56d
Ciujiist/tNwkNgYG4NAB0uIww9fK8eOX4iwBSdDrCN0B5cgiFPgrp+hNf1NNGtGeeTJ6uwl3cKB
UpaIb+XI3sHkd0logWtxAASw68TiC5o6ntNslVrovhLqlXJpSyO5AyM3acen1BzMNZctQ+PyL7GL
y4wd4PBeC81KEu7SHD88ToPJIL2cO0rVVn9gRpgh80GViHy8Atvua8WGm0vQUaiiaxT3KfKa41LJ
r6QZ7i2dWi1NiAqeaIawQdJJxEWMHwGjjH9Zw9NE2kcA23sMEw/wZiAPFPblSh2bNCTOupQRWEFF
SlBBCCprAxgW/0DfuxIx9dyNslJ/Fxgq4UbE4Y7swg/NvoTmBfevfK3/NPfYnjQUy4AeqQ7iPGab
uPeQBhEZG6RpqkINHnWhoUifynrHKBiHfi5yYHD8tLWzK/uyG4HttKzY+C9QI/19WoAPbSTFT0k2
51rqbNIKLntNr8bXQV6i34H647SHRx8hRgsQnt+Ebk2Z4wFHjDley/BDib4UYg6toQg5SqvBS5DO
ebwp1ek1kb1hBGBm0DPqptI7pxuKk+svdXoD5+BDbQ4q173wjyv6UM4/3fGLBRn6SLWs25pp40yG
grGW2MHv7D+jkw2LZ/GBLgsBGrGb3WB6zPLlabOzNZTbBSxTz0Gl557aRIy+cEaHlH4gStxWm2Y5
Rms4sUgvDPdA2bm4aieSUgLfAdJnhD2IRZ30Bc0WgrNUTvBsYC/wq1OMalnLoeXrK0gfrgwI4kdY
GxI4jmQuAHJytxU0OJ50zZkY/O9V/G5i55w/oXrn0F4sN0oN0c3DbiacRVirM3zEbHeH8g9VGrbx
nxp1fR/BeXxeRIQPAeGLnfSdp1DK8BZ88hXeNXZIVkQBHIyACbvndlR0E8Tp8Klr3BSCMSrhpA7E
hdZ8eqPyCJBehnKRuNVhGVmNcqp63BmSh/2jIRtTyZ2EdpNy8Qsv2oGJXoRr+suHY+GkSrMuRFtw
VsaWhUQCNNBi9/GHigMSpF/9e7Woi89aIjh+U4hgf2Mjyw7D/pdKjh/u1pHj6TVLl3pEXXiTzkFi
H+h+q22kWoBazvKwrFyuat93d/1UJ5cpMrFVn4DyVm2PvvZt/rln/y2QZZdgTBBGz3BCNyd3pvdU
r4yvGxEGIehSkT/M/9ctuLYiesvomYvNxOu6ZFUamL0BS1mb28IG/Nl45dzu6ofthYN5tWkQeqvR
9lJD5hwNOqJFra8aFCtRnQGDUPARsPiBkjCiJDEgAB8ehRXfcnG8/J+2o0d79PFrn7lxnhLCTxB8
ZcvoOMwCPmd7lUV1zFXaiDejwsL98qKPRVL7dPz0m1KSCMcVCh57STt2M4D+3ntrXDkz+Fn8RWER
f4ZOeUl1kSfpbUW6i2qK4ZK7eDt7zEVBPVlur/LnuKWCkap3CD3FBhSUMR4ZmMBYc0bbDhUQO6HA
c8xyO7ErtznxUGLuRXHcXy+MmgliSCfqSIQBR7FThVtofRpwjnrPlv99qrEZKlGT/C83kBedvM+Q
Lc2DkH14DjxAaM8DZ8qQpUo35Kcic8ZdoYeQmWD+SkrF9xXTV2meqGcggcRTZ4//DF3kZejluvqG
TKpadsQckR6UTxsFwAJDqCZ3gugPeqmNikaadc9VPrEWlxsrRfDVoQkJacTEBgSsDtJg1SYpEFS4
3yGrlgO7qfwrozascURZYmQABJKEvjKrjflKpVfonvfoKxmJt3pc5OwGgO1hpJPJTV0BwNfXtt/s
8O+1FvZx65+2GqdbOyUoDRdc4reCu/RukA7Q3tb+kN7XLbn1si8qedjBtEzO+FnR3Tbpwqqgw+Vt
UoaBBfXh0WrmNy3bWjGIbZ6QF/a4MovH8+zsDEVMnNUWaEifqIYjiYJ3VwGAA/7NlPQsZlo6LGZr
TMZGTLA8qUg53GRfXDViG+smOOK+LeH/fTDzC+a0k1AaJiXjF7yHA711NUTo249agN8vwkj+wq4o
IE72Sd6P+Le6zDclEqfUiE7Xwuo45I9QIzZ1hX9AMS2Ez2t2bBaZrj0cMOMbRZM87Y5x4My6tsG9
D7xIwY6MwylQhdQDsdSiVc4XP3eErBM48DQvPv75fQbJe8pC2oeYl4esKv4QriM2cXB3DlCjdAAw
WALG0EOtC3/Vn40BN1D0lj8eNw7whuo2BfW1oVmEUFr1ApYFKFtMtypkdwhMvkPBC9Q2HztmGxho
9NoZDdmiTbS9RntaDYpKZ1HTYo9Awy8jjK/uMhG6+acVwAc7D7pxdGnVmK8c/iVbBDlybrZAwree
mJKmBT/LfJEtnUYOMoD6JrJCUgiSA0z8YxZYFGS/tBfCUwhswZYIqcVsqIcAxCFBof7CC0Q2T8Fd
Uo59NC5VSn2a2XXRn+5/5Aj5Sk0pxNt9Q3z+ZlY+YP19BgVCd+qEcaXbXmXD/KJBg3xoTwAJxCFO
mYouQc/KYRlvObAtA3dgb7leosgRCNh34Bpr1AkQCG03C4n6/FMi7Uoa8OxykQucfdSam8ORFUim
3297Bdm8wSUxRCVV+ChiTnXMi5NqrOybMua9IQ8AvlVeg+Al92K5RfDbTXVqIqmYRvJpbEMtiPqu
dxj3F+HFqGGXg21TVWeJcXp2NW5qnrI4BgCQoQlN+5p1Tp7RBzyz2NHwA5vdGxlolX0i8qT0UHtb
hiavuF5gukAWZ3tCMyEQI42DrVnIAAJPRxKz8TTBafNdz6pqxaJiZfmYDtjIOl35q30toQzpfppM
4DtZ/Ytpbmx3W5gdlzbrO7qJbegmcO8Rlbw3QZn+0CsvY/KZ3N0J+jC/1+ZT9wKpz2IFy9ewEjfD
JHHzjzEUeSIhw9Hgy9QlFIpYTC0UmjBto8r/xoPdt8nBwm34clbp+bB6DDTBrHnadZSxpYD3tzJZ
+NRVvObWVGKV/n6wQ7W5QxZXiiyWRaq7PC6GXkWVn5jpefDrAjKLJaH4zXpcZcRcaVivIVsxb5oE
JDWhJCtzbUSRYQZrW4AU48ouhwaVsdsLpLRumtQiO4jR0J2qTqa8606UFAH1A2djx/6vQEXoH77n
YKpU/19tQZ7ya5TtqZ3lHF8qJsLO3b7pfKa4tWT0uFZ9lWXK642d8DTnZNxsZU2B2xR1yCoQMYBA
oPi+viiEfjG8VmimjdVo4REkogfCf/kIBoJPk6vw60668GYeUDp1YCOA790bBjYS/VtsQ1tx65ni
jIDtuzRgQPuVNOK/AcIhRuFjaTvsh9FiQntT1xS9N6pij2h5IQpJe0IO3EqHuN4C0NFf6RSz96yV
2WHiYRF52cvBYH5KyBC/cMmfQz6tHofEPY7309apXpegYEY7pq9+K2h0MVwje2ESyke28clfi+1u
QY0eGvNVvSAn2xDp7P1wNife0t/Ui+c8t6qNtMTOfD3kmD9sfCc7clTlPZm4wWmslhtnPKy7Y9CR
dnaCTDOkuQD8ZZRdJjRErjpJwmw1hWAagfJXC+Pw/FWF6m2ut+sNys6FfLQ+OsJPrOmvySvm4BU1
nD/VPUM8zGMMwu4C7zeWRKGl97aKLYqJtw1Murf9LUW56GTFfPRbF32j7Y25c05JNfI0MZbACmiX
erxG58o5AcRa9zNCsD9hP9lhW04q0HkgbHmJ0oatMErDJ+Qwq9rvEw7FT9nd/VzMX5O7RrecOPWX
rI3G6V0HHwbQcbEURPAU2c1UEQ33KgoTYraU4nYkzcFrVT2L7s19m2rFgKl3klVdhyBZEQjTabTc
jpLNty3Ooc1qjD3gxKWwcx2kQMKZs2kE/4d/7GCHQ1yFXSUuHP+ZfxkulZUVO9fJpvBWyTXiImwG
7Z6culRsRGo5E6iOMpl0XeM3dJi2jPvK6ekerB3mMDs5CZ1WtHVLgQrWNYM9nxhIfMnZX/tMPZUE
vXaaQkXmkE4z2x8xZajNWQU4YCeK9vkXOQzGXAk26lC1nxtmNgrf1ooWwDdInPVHbvL38KbDBGLX
nQ2bjofGfQzPlTNAAXx6WoXdlzkcT8L4hFbmkcaEujDw66dO/5W+0+9j0fQRYhPsBaN5VmxMyjkH
MYz7p2LsvgjYH2IFYNWb4nfM/aZGY6C6dn73CtulUmGzOTysVr7RIAdcKKXlyjoxoxf/KEnBTcfy
j9ZFsBowqa+N2BHnONTccTXbZ1FdqljYgVntu74eaiEbB7aehxoqsJfqJFvAylNW0W4Pd14CCKo1
9oztg6FxovSZn/weUgFdIKPg2zgq9YBhkj04CPEJfV2MSCftQSr6EGHKKhrloqD1mX3I0ZrrxFvi
Sl8y0APUEBTY9TT99n+zW09WvqCdAqQ+/cD+oLDIdyFFLgqtY8MrtR+K87Mf1NKdKFGtBz22q7MO
V7fP1ocmK7IQhwo497mapNo/wg6EawsGwxUPS4nEGRqOp9nDu93VJlYfBOjxTvBSaKt+DGdfy/MO
Fm1cl42DXYUQVPPkCvmLp3TfacZz50eUHLKGySJ6XuUg9Uwwglq1DGDdjSiOuRJF2VuCY/vyEigS
kPp+mykQuKwb5fHo6C04bv8ijemOGzRClpcWrQRIN20BzpnQMkE6JLVKhWxcA/eNHIZ3afqZq4mQ
7R/EkcwAChLFyB9rqszFVQOjVQCGwPfkd9CAOxBICQTP8rhPcfWjFjTzKPkq3A5jtHMqe9cm9DJP
FFyfujH6xAdMTvAvoggzVXtqwNpvsTr4jPwV7WaN+x1WD44rcK5RqwVZF4qaO0muWbiyB1sKrUXv
veckby16m7kvuy8xIenxsBWSKtHNoxhO7OH6ntsVIWm2zSSb3q9BuEk5GSptGfd9H8IaNc9Phb+6
GhROYET2T/zEmXzG827kOUaS936vGXEaDt30qBge9yEckcWHNwPtJepRZATw912nVW3QMBYthcd3
cosG9v+poGaCnVQClmjbaHSAcEbznb4fI70tRB3I7XMVtknO2zgf5A+nvdSUBauJTBH+xQ5LIHij
9hfYwLcTSF2uxKyDF6O8zdMUpS0zHibfRvEKQUS2sc4Ohs6T30C2h3ZbkjGEfk501wU5CvEd/nJw
7OA7vQGB7fF3vcTMgjNBP+8O0zMCdV2Y9pBiPf454QAaJ5nA+ghipRucqRrhlaQaDtUPxPKrD/rB
csmoMX/lp3AVmH8KAFBjuH5w/nPvkT8zXHltrUEc2DDfQlHRT/dt8Url4TjGHz1aq6o7t+MYDBi0
xQTZz3jxvPvVBdeNiimvd7sp9u6machZk2UULzwjg7kAQshl51VrbnENAjF6OLqZpi//YGXR+wKc
j8DFkOUO8z43uprJZcj6zamvMUcZd72CdmfPHx5AlgkCEMJmmE+iT4iWFvRiAvdPAoYNfX3IRk8k
ghbf9oro44YLmCzN7NvBH3X0zXW0rQfnM8zvVk/vIVYD5UwuwePrQb8lxBgk+eMtEE8KZHR4nnzz
lKo9ksKhEaBM/3r7LghKV/yOwymW/c28B4LcpPCinapbqJHSPbHGKzqD4UhbxJKFywcxxuke4ZIU
OHuUmCg/CW40VuU3THHjGklbtGFOsDE7M2/NWE0f7RoD1RUk9fE98YN1o88gL9En3zZrG3qFRgE+
fnx69YmBSO7a7E6/g4sg0oXMesOCckipix3x1NHE2fJ+XiQkng4Hh2tK3Y6fH0qETb+C1aLhl2VJ
0SHa+/qV3rVySeXhmymBleM4ZKMoh2lpHIAOY865mgH/4Awr2aUHBNZOO/6qdxShPmpW+dxXXOag
3RKX2UuH2pg8n+ys5sw6QfRjRmVB601Op2F9Ex0TYEQaHakQwyB1r1u4Pso/gqrULO+AemXvqKvG
GDLS3qM9dbVPNZdiVLMKIrs5+D3UY6aGRnawJ8FhmcqitcLIWe+0NPcNVYlNcHP1oEOlPzO/SuP9
yGh1/39y4yvmhfv7XUmT2Pr6sJ/ZPt/N07pnn2m/i6tgbvnJKSA90p/75nIZWc3gvStcYUMehu4g
IDVduv9uFYv1Izh7OFM2Gy2PnI+s1x49MCedqrOfaPR34ro0OZ88zU+sSFXG7/r8NXu562QT7dQm
P2Rt/atNZ82SCfG/kYrhE4eAbKzQXgeacYmHkWs6YQxftaj2BT8UrwP4KD82exNjvUAA7TnEQcx/
cvo18AclaJ8Ly73SMPI3tZzIiZ+sVS/GKyvDK7Fqs6p59KlbpR5b0/fQQN6avKWxfhNfo62bqvOB
7Dl1heeJxEn+oNhB1UowlaxaR2bnCCYBiVnMAztjNqRbXKOc6SMiGZdB/FRP6ffsW3JOyMiYB/ms
0hjPHYvrhQMHfTrl4AKEfoPUCSD3/dGbQLFEmG+RWnnHlIjwc1yqhz/04fXElp6K0krUiEioTYeZ
cSRMjqbcCQaCeWOUuK5PWiHNlaf9FwciggVuA5wqf7vW7jD9m3+6Vv/9kpxx6xC3VqcqXt7N8Gbt
kf6A7/hHcR42i+rpQi95MCModqbawuwD09j+2VIHYfuJhuUzzV6Z2yUixQ1CD2z4AXV+of8m1LAr
r1jPZBfyVHPBaMGvt8n0CtgbGLpuhdV5xq3WgGlyjyxlIibwxmVaOR8Ozvyro8z+wm4On5dkqJRf
ATIOSmpaE4FKhfDX2cVaorWrznUEmlYnRr6yCvgumCnYL2ZLbfyYI4uDaNfIlzaBjR/atBq8D+i6
/LgjxPguxhTvgG9FkJuYhRlZ2uoqDaestHD8AMYSuqe6ur5wZTciLOlaBHlzdzycC3k7RCvNrI6s
280A05m9ztee7LMIFP/Ve7+i6od8A1IcjuALdTJkw92k5vkZ++COO5icLUpX7iAu9pIqZuAp4R8S
ZofGmWCL1MHGEcV1mf0/mz5YKu9i+PeHfUjGGtMVcV31ExzDshRQvbsYv7q62KT0gl+UT+juvpxi
VYVr9gk1bziF/vM0KSs34rWZxKi6ozfOSYA9Ae6Ery0Q2ga1kBTVLP+5EP0UxiAtl4NOI5bjJa+e
C673WxKpUyoI9v9Zp/U2XG0fZv4aX44kZdDelf0CpzDJnGx0FPDIksHeE5F/Y+opiUvDpKJISG5q
tZ6U/tO/8a8v4K487v5+mEUEi/r/EP/voVr3aILiYMLuoGcaS6FLVnJkMCVQSrNki5Jd9hWLJ3au
ILNdsrLDWzqfuKgUCVEdXTWrzZ6Lh1R6WnQP6egm56aI7f148dL6UuTT0I3Bl7W31QBiacghP//j
WGV/XycUDTBRNIAdhS6XVC3qgjzDeMLEm8zakwFvwPozs6ZeEJGtpF6ZtNEsXICAdSaQIEefCmSC
MUIkf4KaZ4O0xxRo2xhwmh8iy0Hv51W1GYmtpwdACURU448mXJEQoaE6c1laivLpH87urWVX5p+9
HmczVzTowuFxJ5f8A+640Fy9q2KRtLybtoEZSh+DTSPkvsnCFayokm+Llf6QzjWf6tAwnukntXiT
QoORFIqcR+2/OJ8CXJU2MBJ+LNXqZFfevlXEX87y7JacEDBdw0eenrExscO1JiBAKpMj4xIQ7Qnh
ND4ftks3WE68pVQ9yNDQVwBgNFPipAodXKfjRq340FxFZKz1j5pOZBzFRIoTaDPP824R5AmlNpBG
JcyOkTkSoNN1n3iurYuxQ/d/dzhSPlkiCD+6QQ3KFlxm6etnn7Xvn+NgidDw1Xr2BnvIxycegMuk
ltUFDVxHjh2Ry8Ti4n2IMQJ4mLzR0EiKrnaLxM6WKd8YnbJYPqhtUsi1Ek9E1m6UYPAM6s6/wvwI
tQoYXkFaTG7B9/Yui9S2KNjhbpZJzqc84Xj9sVNYxwtF/EOnde8ykxxkmMRD9ZoG6DYA6gw1Wm44
bd60PG6bp/bzc6qZKaCNhPFwhY7SxC+LIhuqsqEnbbT/M7BFVQgze7knbKgwnZaeLqHuPuCDRjJm
SBzUDm/lpf7g6NOi5z5WnWJphzM4lDt73DC4rQ63W0KIB31z4ZgvVUxdqY6AIeVNCxv8ecByQhBl
+2egNsl/7Xi1dhy7NFUUrPkcpzFJ9BvsAnxCDKB3eGCJC2xX5MY3fKkhf2gnDi3L14H442qQ9L2+
IdlykaCACXvtw/AJ4MUUvwzZYOCXkP/nU6E7K0UGyhXtTjI9x0WkMp+ilolo2qp+SqwOE9YH9tsl
OaLvjRUgqocAd54iQV9GbQnlqzWPorD4BO6tf9Xj9ntxVnYqMUeAk9Jo++CpXILuZV9zYzVQb7Nv
yiSu/ZlAjTYekGDI2U+6y/T7Us51EnvEHIHi2EyjHQSTPADONgfUgAJ3oa4Qrre8dczAKk1+0YTc
+xiPILLcemcgBrYvvQsfEidRNQzSm/SCLzG6Lay8qXEg60RhD2GO+SzB3T0Kgr6mn6mDnNUqCbT7
tg32tang6929keDXlEQWEXrsu72DMsb/PCYNTDJlk4o08O3htOkxWcRbHsokBdIgiON3rSSw7v8P
xWrp/4ZSCLJncsEVGd+SBFakvnH8HreERt+QKuvpa8cv5Xb8cQmUU1k5k6GYGjFDbnJAsWjBDF8E
fgzP9BqdGqIuuELQcrhMwkpGMUoX/ESp8hh1Lp2bDcPtRMdONTl4fsQFqT/te415OmlZQjzpdw0s
pHPhN3WXf75j6fhWs9io9aVXhuECOfGo4EfGd2XJRouGG/EMT+9qKQHLkTTDLsMF5rJFXOb5mLz0
o/xgUYGG9wa+6YNsML0jLMGdgPp4Gl2KlexqQ+rjqIxg9gYKOn9zDtmC6c2Ed96RnT139pOr2wtX
1+tFMI4lDshzxYe41uuFDBERHIuXSxPdafx2NwY6l5mjx6yKnOkhzL2BcZ3B0QYqw6Uy3YA8zGWb
++pfvuqeryZXr7WNssfWUtGpQBZmZF2lxwejcL4YegS9XlGNtHYldDo3zk+X/Z/XaDMsPF5nVS3L
BYbpO7b+zO3Uq1rcCgi3FlUQM6kY86hBryEKxbjtHqcc8C/n4VzYEn/BNS+ZcYFT4owrzlfYk0nD
VFi06s3mSsi50Bz/vjv7znGgVJ+L88DZ8xSzjk5EX4e/XrWTRA4c/I3f/7UAp/LZMLbWG+NMfQZc
jvMtuvAESFRoxxirI5qa3Dj/OPixHP/0gksYdTO8c4D2gC7njT7/lPyQQaGipBggzpIaE+KCcYFP
I1R2Py23IyIYflprxl8oB5t1oiDn/KglQnt1NTo/zEg31ffWsrYuQthIqbIjJiT/6Xf5QFWaSa05
g0rCHCPQzvjRfQoVbcN9TB+/VMzZFVrLXw8iKoM3JDudsEQwsvH0Ibxbt4tt+Mh8CnWKiBCpDUYP
gWnHMsdZ8MPjTlp7SMbOtvEAlIgoi/iIkVQaCqw6cL2sUEtR9xB+7xF6Dlj+uC6yR45cJ4lT0Lbm
q4Bdofo+E+xyBZWeEzLPcqZ2Wkoy9Z9lH60QK21AbcZ5XK04ARf3morNVpS3mBIPQqTx5uGcrd8y
/4TuWY08LQGNiKsVfq7XvX/KxTEv8BYDawCFYw5DigZ4FoBSza5jJwBdRBq3QdX7xkPOrWa1jDZC
HDxrZig7+CN5WyfJ1+gC3IiA+m/mp0RANblGekD7Dl1JYmJHKiTE4cnRR++OCCJj4/+2FVtB7Huk
EOjf4v6Sw6P8GwEkwng1jfI88tk8ldyRx/KA/nOp9RZddcaF1cHEsmqwQitrQdwcFKXIxDjF59og
0tV7IkMQ/9Gc8qBwOFoSIFtX/eNedKpPLCnzg3WHpMqo/pwbODeUdZpB6xps0cRrcXVhpKc8lRaU
WgarPDoq2t9TLLoBAtkWQeWbY+kKZemrZM8ifyD9zSYWiJ2ssbToX2O05oPLQ2fFggRKKWTxXRbW
SuygGBCcwO7fBWh3VdO8S8giNM2TZEQsinkrgy3lt0/3EZdY433hjBhbeynkR/03SHg8m+8DGcG/
Q8gJCgaP6iJV1Px5FDqAVehz+QG76ffoZavoUyc8hfHzajW7P1jRfvc8LBAWQ5zBvQUOcAUYMOmH
5IyU44WE+UELVgK1QND4lUjWe8bMMmwFvkZvPdcqwjePfmr/LKQhwvxcRvmC0RF+FvtZZS2cyvAH
E0Ne9yImCmeiKwfvG6+pzMpMCRlcOcuWwo0mmMSV6BhAU5krVWi1trzMouY1e/AqKszqqggTCGXC
EpHP/70CZtuki/94cCyZsvrfAnDNykDp1stB0yIeX0LzEOr+VxMvSm5vAlmIIY8OHXb3kqhdR1mp
QHfSuwsBt/OdsZQqt3R6c1+obQRjjaECDseqlYhAa1hrqg78o2eIZoqVRXksY6iuKXvm6xxmPuPG
Wrb4kDkMW7DYmP0VwjVPFHmiPfugAhWF/rMROF9fGdf2B8FYTutIkMwNkq0TPxWQHQpqqrRr18Hj
RAPwckezyfYrTxUGhYKtk6PtzuPJAlcNnqVeHEhGXzi8A8s+RnN/R2AZjPcZnR710JK1BO3pBba/
HVql8P6UDavCnwg1LEIHFb5aODAYaBEaZ/baMdfFfn/090C/bLGj8wnXzevAabFb4AOTL1PtWHY0
IGrROfG/u6QAWn1bUdC1r/Wb9NIFUW6GJaaE5Z7pcQF1oyOzxAntnkh7fKjyAm7UNUjEqoGcPutb
rdmvYtmdAXt7digDF8AvXg1p5Z895PjMk5uxXV0XePal6QlpLPx7zTctJdsh/7jnpN+KZvaf5Qdy
rrykpZFuUJWYJaTQG9iCjGEAq/HXhKgAktIrypqqWov67qcqvvXKaYdZxzzWA19zUJ0RnSsoAERz
9qKskotqzoglg//VOq8lR9JnZbAYpPQZVx2N2y0aa2sVzNqVQThmlgygVDj3MgJup0QIc5d616or
l1/dF1B6cioWgKokGD05OjDSzxkg9jdBhh/34C2LuYnS211Jkgsnyvp9AsFA+WSCgxANMeNrtqIJ
dM0G84hb/qIrbOn6AGi08ps4LOv6xvFjU9ZFJ4hiF+AanK0YaJlZmyJB5JgokTNJwp+i3ZsztRue
9rP9TMoESqfqp3GWgHzRNswfu1HEKuf8QhyHLlutR2XtR31+slw0CMzpgyDTl+9Me/SWOiblWiKi
i/uhYg+tyFOWTUZmXt8//z+VUi/D3h50QFY3LY0BMfGB2ydylMcIVJN86r4wNmfgRUFy1p78LfBQ
IZ0PcP9FupXyqscWjq9PWuI3TSWUO3mr0EYQjhFTvCATeJNPeI8vwsI/treXGxyGaYlfBQsjG/5V
W58FUUc/LxR61v5iqpJGG4Z/myiPextWJbgGcE7gONC1ZjtbjnbL0yp6exsN6KqMzy9DW671AwJA
I8xPfg5mQNHX3Kw8ggigYANg+/U+fLjN7BFgX+NWerzDvT+kaFLFxI+dlia9Ihwbjrdz7dmSMHSH
5/FHUSkrKanLJUFwV9hcbXmHvhByxZCundjhXvxbXPA7cFHGNNduxe9vNjremvYNkZu43/UbLaqf
E2kOYcMsF++99HxvYZX9VMF9k73sbSLYB2BahPbxO3p1CuBORUlWik8p6SYkipt3v4Q5vM+nA2US
5iyvk2P91h1l0BgKa7p0YAeej7NHoHCl0glmRWPyOWGWcMrzO/zbH0/Geoc11gT2/QKRbGg4QdiQ
6oIgTHeCqiseyZEZKO/SwZfN4h44e6CwbEmr7pEetn9o/8XH9lZp0NTYrfOrVVlzC56Qe5M3yBwy
2Terr0Ei1Ck84tDdRP6M5AWtAMjxh+qhTSp/3CVGn056ztQk033R5SHecOMiO6tDZWYuU4HFsW4Z
2yiBV4ctrgvVK/UvQwtWU7588mnxGc59ncUsuTyThfkOMJ17z+6ThMxeV79umcAqJlva/8NLI8/x
RWdZCddTWL/EulMi6WzH0McvW4jwTp/sOW/Re/HvdmBv7Hqg8/r8h4T2aUUsOn/GvtA0gG+/jX6C
zAFFzHY+/UgqhfUspZUxFJTtXshHi/2WGjAFzKtDWwCtIy656NRG2TMHswpPOarJTReYtCvDUokh
Ee8pNWRQ1xFlU/5mnAg8iVIezXwaAcMrCFSKdwExkPXndWh1JRR1OaA1kgu4NoXgT+Mf0mCru57q
6jMnMkJo22jT82fQ/eayyjQwmA+uyEpPKbD6mAbcy3VjCCJ2pEd53lST7ioXlF6dIAQoo7G4JCGl
Bvc0hCnRXF6PFFZCqvO/GraNRT1bpyn3Y2Yo6hC/W8wBbrfYwzZ/iaCWq5flZRJ4pQyjwLYVfEsA
LNNE29r92UYbsjCyYu6tURj2tcRzZn+ENreZGA9w6zhEQgnbyOovn2Oynvmc1hx884YjgZw7nyz6
sAx7wcut+L1fPVfEqx+6EGqVU15D0JDhEPvjVSIVWiqKvrVfqf62qmNfR/+hNOtTo2+5/91MiA/+
x1smNcakdFoch7OvksQew6+E22RGPJmpRdCm9aVrniVh9go3L1XSTqjAaeXOBfg7klAKNDU2mnUP
4tkRWd9m16hJkKjJu8ygMTYD8rodGbsOPK0lWvc9ul+ORqruhlGn8pYU0+DrcJgF6VHi79h7bWjs
jsSujDeFMx+DgW4dbJFRZ+UXEHewJX+ixc+zXXVPqI3PyAPG9qF/pbrdwSPlioenGU6vxDXum0xe
rZuqT0hAvgQbOuTEAqAjO2qPKqJlMCTJCgoC/ZsoO2mcDw3fHc+Svuw43ZgeA6UhGJ1nF1cHTNH9
P6rkKgDdyYZMIu9BAxCUN+lG8gn7PA/MN45cUJnFClP4YSTNlqJhp2PhgPH5FFfcYKM7EGA+cBQm
W1D1rRBifopiBfIm3r9Sefd6gE+NfJ+dGxgAn5AefyVarf4Gm5ZH3qRXP6iTvs2aSMSHr9pGNHdU
cq12Q2zb1FcZi109eqIxFtrIYUc1MfrNq626NuDoDHlQSqudBl7dAWyY9Wtjf0ZVG/Lg5CsVO5Xt
l6EgYDsM6Il2Bbce7DRXRmikbZQVWNM1aCoxna3BkUuDGz5DhsjlldU2J76mK/NeEKciz+76zXcH
HLMZC1nIKzvx8+hG/NlF1RpNINAgxamCm/wmc1LZi9HNVmpARxr3A1wT0J4+gWIdg6pXgivelbaw
GP1+symTtQ9uPn2jNNQM5DnBb47rN8PWHrKaWgoox+zpxM0zb3hMTdVHCovyvELstTNgjp4LdK8y
ktl8wdY91xD4CuDNofaYnFVnCuozgIaGJKksEipjWVeUgAy4FbME4Okk7dwF6bKdi2Fls+mWaQwl
s6qS84GmInj7Zf2/bFoB/p+t7fTXV26f9bBSYkqxPo5uO71Jw2cixoPuSPV5UH8cr386E109f5Ss
l3tKY7fqrYMGbMek3Dvd7PBRUqYVT1l7qkqeEXJ4b05Kud44yDvwoCB4iYVrvm69/EJB760XFDc5
DUOVx+U9yD0ClS81zw3x1/KQekpMtzJ6WLoja/Ca8vSN/dwBvb7LqavqzvkpvSoQwC18NXWfn279
1xdTy+yRWvey9QDKGe68H8qoMkMYBugB38puyKjNDP7q32s0XoYU3eYN9qk6w7mPqkxZVmSYGeBm
DxQabM2tqW6WsF9qliAiHyx6khjNwqBaAD9+M/t1tyo0BGnkjhwOkibcLv68Hz0R/wlCIzASWgyD
KrA0OW54/Mn/NtG+BcYGO0BeNHMzm/sMU34HVc8XPgcLjN70SpupQjbAPQhiIDKK1IKavHhLAdHi
yuanLa7RWB90DWN0nn6VQvcDg/W2hco/Vgx3T3UMmcY9K301efAJSHr8OMCApqc9mWe9BeW2yJIz
OzgKHTh/jI0NCYRD9r47+avFafVvbQeS+iA4BZuQsY34TA23CaOvMr2ft2lIzPQkO/yLfmOWz9Rw
EMrU9U7D592wu8Hs+01MvfHc01gtjCFK/fnB2BChJ83MxFzZ2TWG5+13c/BzIQhsGQY456Ze8HXp
P6fnCzgw/StJKKFuSOMnmhwO2b2NJ95r72gJbha1W2i4N3d/L3SVRHlGtXMCqO0i2rNNXG7HOzMg
VD3MdqPm4AhW5j5OsTRwWGVvBjqfyD81Z4OUiqY1aQwxC/QqNWKMtFzsTq4n4dWWQ9K4FxYOgc7F
1aqsZAyGBF/Xr/hRp6m5OLu/+TYtuG8LrUuhptxK8Go/oS2qctjs/XZ7YaK9dvwz9YANAYVSrQVj
UDDsek9FQgeHtwFNm94hp8pydiHPD7TpFDb7TNJ5YF+KyMze44TKwv/qGQS4WoS4XpMQ5wiUbbbx
tsroKVAledhVi436Lr9g57IX2KC17dsV5IFb3pdLw1zUoFzUGI83O6efMnQBlDJSm0SEukuno55t
G9OBduWvD3i9q7+1VC1kKULIzyox4EduFaWc00U6f+yVzgGqKR+wBsyq7Cw5dEFyqfvCLjGKK6R5
T11lUuLEG/aEVC1bs/EoFw1/qRKiFtG/hU8SB/B4ACMMeUmWQqfwHtSEPRSXZn2CGYkg1feeIm8J
gJwkbDwDX6EZ8mka14FLIdyILLnFky59FPPe0coiuPaXZ+izsKiLT+Rp+1SWmqPm+Pma838u/qml
0gIK993aI9wj2ieWEIZ8SD9VmAywrJNc/CiKUtxxR/2JGYutJ+4A679Vl0f3q6W3wxmB4+dB7MVy
OpFfzqMDtdkAkzXEMX0JY2HfyTwgm7LcObvolWMPPXJc2YNN/y5tGz23UBYOFr3VoUeNhCFUUC0K
tK84fEHdzew8Foo/OFrzEaD+UfkMvSWXFl+SPfb/j3yKpzwZXvSpolcPBlqrPTOWmCjvsOXja3Eq
MQJ9r+XTpOfTBBKeIxxFhEhm1nVyaGbSIC8ApIoDKWzg5C1pTY1HphFCXffmU4/y3qzLI3XRRqUj
YIYaUplxXxBo3QrdCD3Zf96Az8qUbICQThhdyePtu9QatYK7x0OHkvdhcgvqJdvv9d7uPMNuU/QX
Ye6Z3+HtmIOQqWH0/b2bWaB4/c9nTx5jHaVIuyedeppSpmHKw/6Dn3p3vFRLXt2KbxCEwejpNIfT
kfX7EGE+0i3hFNcBoL3hHhbXLyrPA/v4L6qkuRB7ocjTLby2siRg/Nju9YGsknPetj5pQTUUMcTv
rPi4WORPovxYjKwH4wQ+RAgCGRAw9pNO81Zyg+/xvI/0XEI43jWueLtZNJVnkDsVfTCpezhZR7Aa
UQBmb+Snu4Z65dtazRRY0MCluRr7VAUC+4q8C7ScRasxC7hcWLIVc1VKmwHnlikikuPNfu2gx/N7
BB54WbpjthjcvTeuDiqCAZK9zsiSVzaNVP1sJxmTixOUHkJEwXoWKk59IuRUVZJh+8Co6QKBts3u
A3B9z4WOr3hcgXld4tpIYvV82Gn7wYUVvA2hOx42qiwoSnwXIhWaYUyfEgjhPA0VdySbO+VXLTWp
XCBc6bZHKPwtX2e5WVD7QViMeBZLlJ7XIsqCIohsS/mQudUbNrrB8DPxuemC/Ifvn9Ff0DZsWz7h
NITygVmK10XLu8/sioDAmxrq3ExCEYWu3o6cNkP6sRk6RZQgl5pYbu5+UWquetFJDDfSp+lFTNWs
9XGEGuukZUTIt5qD8N90YDJ9rltviCPXy9nAbUpDYlN3QytopSAayIbHhBmv50PkTdBuzWflzl+3
4LAVCcaBxA1hYOXr8PDg91pyrfCMNkYjlwSfgVsDvuQOHDq214YGcosjZBlbowtZt94Clzu6Bqd2
FI6JvjGvzQNLnu4veCCoDljw4bch0j0NMXbzesAa8EByXEpHbUD0EXunYNil5YWwrnPUwb95TqIL
ZW33xVK3Xmb4xHKhvoeq9LYyzo0vWgB150hBrmwHFAdnXg0rYcWRiZR3nwuHqjP1da3L1RdsXfCt
GQYKnGrVH7LeyBtOqbIhQ7h+hl8uu7a2JPJXxoyMULdIte4OdrFQs5qTFp9g5idYKH9laUmK25q/
QVJVTPvVXti08mKy8ALnbJoKpI5GBb8eS1ahb7uD/HpaT+QphmWAxdvGs9DgXeLsZfUVqLWGSPb6
XTjX+uk0Trr9Th3WvNb4gGFf2VNSXGFYfBZhJwKJBLnxVQ5xhNSx3HNo0LLhODjZeg2pkw5V9XF/
iFDXxtA4mqENp5U+bPu+tSlYaycBcVG4K6omcWw/fA7wsVLK/gXOApAQ7NxEiYYYTEA6KGL2UO+d
AIh4vIdB8JV/4N6MYvUCINSPJnnkiI2DtzmOPVuWOdoX+u4EIjuZNB87nFCMxusktkm0ytXcL9dD
8S1OESOzA2Zffb5eEPzboxuK4m9CkxERJCeFHlwbL7OYymiXgaGubm0OQ0eqz81mo9DXhqYJSan9
+PdYYGpwa7fhzGWgpS5IBflYCU1BedDRteVwlIXh8R1oA+Ip+A+D5N79Yj1l7FjZG0KYpy3QBRTO
V7EkYKTxczHqgcLNV1j1sEZHQN3j6aOyGWrXnWZElTYVP6qs6wTpUmb9pWbKjnEoQm+nmVuYUJ0n
Zreh41AU6yMmrJl+yRxB5yy1gZZ27+oNRPzJ6p6IwIMabtESqcrMcHMihq05HmZGTQiYGl2+Xyo8
est3gUzM1Fyyl20QTfzVp1XDHbjKcWNqhRrA1eJ6fMTLLhE/FQ/X3mnBoRlkVKJGnXoCLtr5d8gv
RF3nEbr+UZ9HdvbIqxJwcXIb2XaqnIZqZ3sNvRydXYA2+nualfP2V6q6H+lmeyT77BJPZiv0Oh/q
3cPPVkWGBWMcx8LXNKvDSJr8yGFf5Oh8XEqgKEEJHhumLWCQFa84h6gnl1zgL5fQ4orKBLLwePT+
3jUUnoFEDNdkU0hLsc2d0OPsAKBoe0DE4hVbbWStnq4FdiIaqoUZOlSIbyBRrqFRPM5YcUdvwX8i
jpYTqkIibAERz4lKLG3E7yPIXbMB7/kqsaCE0pT+zQimWf7SGn9e/82r1cm6L1XWRLms5hXDcnsc
ZgNLveEZJJowx1vS4BNGrpN1QBBiRCY22OBcsXonE/TPZubusdJm0ggI5JsmE6grDET47C78HWBU
6tpqWDIj31ayueqT+nDlDTeYPJ9XLxcNcXPjTlnlTD9sjSeysg8hJXB9XRYVlxdR6chGixpLADNi
raUJCfClXtxnU5K6v8ekN6muhQmhVH/w6QzD7orkCTCSho53o1gzbmHwYYECcEipoUxX01XHBalt
1bTiC+KKITln9wReeyWQmUs9464IUKKn7LzmvyqTsm9RqmLncKfWt6Bw6jmA5Z42o/OY2yv34x9b
LkZ3gTMfVJ70xsuDkO0D1sdoFTM6anWnqviOM7esg5u3ufJgoN4rj1eYeMbHyN+FR0X+6xqJ2/rq
xY6JpDcwrwuqoJdaGZM0sf3ULwPVO8RbGJxqO8PSjKxu6b3q8XZ/JXTJEPHfYQb+YXNPOrjjIN4c
ci/MKJOewiB5oADdi9gu58TjO5YePWwhDkkWpsmDkIpUm+kV8Z4bem4JsC/G0gYWekxD5snFA7QD
glxoE2PJv9co1HvDzJeHOATv9ocVMQdeJi+ZnFK6qpJFl+tUgdrv2cnl8vbST+8tMeSpj4pr2JJo
61ciOQdMnGEYLjODlZjpYRYFJ4yq67g2VY4VFmhB3wwY6jBi4WCHSGiZuYJ5TAVpFHcRf2dn6c0Y
cwWVW32AS30QPCVqPEFcDSjT58ADDR+oVW3sY9PV/953WQ4zXbDdIHZcpY184O7481VfCqgxDJX5
EJe5/ERsVTSoCZPic6TLx4XrOIaXI1MCuHzpiAQOTa5yMgGg77hB2Tkbs5gH0JrUhNSNAiD2JDwF
37xL6x5Rj4kxAzVe3VPGT0t1xUYpzljLQPVlSBSBW2is0tmSj+uNLHq9xNqNveDyTBdo5QN/xWK+
czWE2Xv7RyfoneeoxQQKP6hUNtGFXz/uvazBbozqaKVjJxy5ovVSS5VxQpgvT+BGJoUxBmhNsJdY
GzKAevp8ZoTjFFSEP04PRE2QwRVFOumjWpsCIP42XAkeMogpUTHaYNL0e+8knHtbSnga1gQHj+FM
L8MabWpA6hyWvGEK4dgWYUW3AnuoO7b/+cNpI7Pb/SSX6948Tw6T+v7SRQLOJq9zIzaEpC+PX7TT
EPXFugStGNgXsDhAYxKx8c2Bly62pUM398+Hya+5T7/AjgCLlR0mgPHLp6kvF9dQSB77qX3hY6Xh
u6PICl+Ki5bV6WPk8sRqosPLTSLkYuTgbW8xEsrUvsB7y6kbS4ABExmlhAAXyujJL7tKrImAwtID
OMtuadrCrCuBwQfvG+23yCI6KP5U2FlopggDJRVTwTHJvuKE3N1cR68CE3Wtr+GjuzOBxHlc4wev
JZ/6vzoBPLmUdDoRtoYSSRRfA2FGdZjDw0dMMq6Lz+XRa61AIcmap6hMDn4neXvCW+T9epGzE0Yl
aEFbALFsx/gsOQHKUJ+2wFmx9XTKscDkfem4MB9fuRUqApgCxAFGw6zlAlRWCK+TrRTSyee+1oVB
Wc0N2lObFug9JrBTRhwhW4OJw/bVGmGO5tlUIlY0D7LNPLU5R6S2SmzvdMZ/vj3rVAKBmDiHSWm3
/t0+6ijBqqx/grfCWr8B30Se7/Ksi1Qzqs6l7FzjoJXFcBRw0WBGJK/EGV1UhvOZziidoRlnFhDR
f/L0wKKooEgW4I72iz7aJdbN/uLOI4swigdwj6a49mRE+ux5NhGQ3UEDXnQkZTVSQEJUCi5E2BON
77vYZZ5eiHbaTjauToxQDBIrHUMuce4TXRjz+tby+BD0rVge/HdGb/DVECbVqJaNc+R+MBQ+MKPG
uryJZSN2SaVdZKGNcOI9fVgngdEVW7wz6xIw1u8rONakFZYqOPMJHAJF4zFXTpSM/CiZvPcHqmdX
qrDnxx/cROamCEuYlYs5J1sZzVFH/MPHtYiB2dK+1+qf6jAKwC/y72ljtquisWiESfsyRQgPPcht
kvIYeqDZLCqyRO3AmMjEd1d9nvuJykxp3UeEBUReKku+97HnWNY7JVgzvtRBUFsvZ6U96y/2KijZ
lg2DrOxUqMwqjnCCvvXx12qd/v+iBmEdfPD+Fr9Wq5Gm0rz0noxjqd+Mj2N1A6K2hzSIL3LvT01i
9he+Sz/3ZZx3XML5j4/fTa64aYEm7V78OQ1q3Du4oRtBzJJ0t7qDFHgQE9K/5jaFAHCoWb3IZ7PY
LJN1ns/wxuuqh/YQFysv+ZCNbktMvG2a47MEDdXyDIo05QJQB/2fZJdN9XXxnJaqf0K2049W6xy3
zHqfKJNfzWHih30/n65rDkHiV24arge6bMS2DeZNBS7jBpmSGPPSU/2WZ7OI6MapHvXZUSVs9JLH
+AHnAeeXU47Q1XLMd8pMYN1JlWuo2mFjefL9JQkYw5pSQb9XFw7ZP4zt++PPmJHQNLRSQRJS43e8
vFhXIFAjJwLkJG+ZgMGI6trtmdU3pmAlzuwH/hDWFHk+2jvPJ2lG2VgoxGu1PKfOculKwZs0QBio
EscKep2Q5HPyEg6hA823dYOtJ3EUc+RjauIRsyZTHJzYVPpyP+WXrAnfc98lZiokBRjqcooFt3/7
q9tTIlXPI6afypwi3k+7TTNq36IzTq9CXI4Fza1o4j7a5O5cmGKn/TsjvdErkgDXTQNSGY+3vsvk
Xljdb+hMzMXlHV9Jkkf4aJDtLAIyqxYvzuXfUZKh/RurBz0T3RshXGpdqoOfCy0CxYDC0CHq2A+y
5sMWtpfMr9SrlyRSmmjNtEkyg89Nqot39w4KojuhzYDoQsen1YCawPKF04b+BiTxDKw8cUmtgkvT
C4bgrtMa0AumBV5A1uklZNRiLR7j+w0rT45C46IY0ynYIfIOmpLRWvjHqrqIuqZJmNZu9NxpaYkm
f5g7piexlRWYrSWlQPgMlBMnW+6e5ICvhWFwZay1bZsdmqRu7AbimdG28203AAVj/lOqtbDaC1oY
Wu9SM0FlL1VJYehVSYmaxNkU0r4tvfRWLIvCQ4/Hj1QXESFLB6BreqkGvGyKQOtJWm0TMqgyWzNI
PmIPTe4MnUdWxxcxNR+NEtyV4rxMYIiVzRwvmEYPvCO2liYcLX5EVMZxkwVW72ql4pREEdB1BY9s
i+03fn3379vi+hhTQ7BQZMbvwG1kNphWVh3Jq5+CuLzH3OH3kLn2rLxPn5VevQyURfy2Wj8tJYw/
HoSfNbaKz8Ps/HTShc8Bhp6rRrwB+KX7do5Het3PTzAiVb2wKwMGgWK1b6KefTFqEQqgzlS0WsMQ
I0uGjmN3ok10wtkOyFNJautQQWoTGwteDmCbuz2QgSsfbtw8uTZKBqVl06F/r34iv28PkxqHbU/N
qjxuR3XK5TkG4vuDTcv4pvbil/AmNUVAYVd5pEit1Q4x/h3DBnjT2Gir0Yw3lW7XIuWc2/LzfjX5
RNE3x4t1Y1IQfuRSHf51EDB9nC5Re/Jg4M2LBXmOrJcJ8omVnIT9t4SQyValrVfg/HXCoAeV18JD
BQhDH6Hq+ch+L90OwcN+Jq6gV6TMcw77s97mMZsraJOE16XiTzPVsquHb3VYFutDRKf2X3zAaZIO
9aq5LWFpW0ltKgwKFvPzJBZqS7TS6GY8Drx8VH2/rg1YxwKy8DTDOhEuM5oN3v1S+om29XxH0vut
4XyYHt4vjjX3ijMMlKDvlj/dNBrd1IWlURk75A3UQrIFBboguhCd9nXcTyn5BLJms3gfzrMvH0ra
qKEIPuzKIJA+/FTpUav90vX6Jamf3bTna4DjwhxE2NbcfXtXbs6lcNptYISafX/2Zzk8O5SvTrbG
yFODUGYpAYE9BP/hIPB0LhGTANKCGI8MYkS6fAvKAhM3D+bz76feTLN9T2LlY0ImJacohBBFA5QL
BG31Wge/elRA13y0SxpIVvoLBxP8yMcSikYmQ0RrQBT7TJsPExYdjYHB1accceqDaVMMEN9UcMeK
uF2OidPxhATyWp8IDqyg9XUFMZ6fVlBn6vlNYX7TJtjmKsrADfNV7xzdM/gLqNHRlelV5FNxFion
BntyfNjJGyGwAcQSuH9IMZGlA7yeG8vZtT9DaLceFylnqCp30YL0ItRemN3WGbvROOd1qfdpxEGT
7mbrcaqHeBjcnp2QJ+DHvy6TsvjIMD2nWldRspXbdW8ZM5WjRLM2fqvZChi2LW8dg95tqx5o6XX1
1JMF3drV7OiR6my1/zYVEZ1zk24h+SnbWHaSYQnrUcX8IuKfmnibQRhuoJD5OnOd7HVEM4jnYj2/
AXhMEkrCy+rw6OwG6oS25GrPGRiACklMEn9/h6kaqX2gomFlFXIU8wyeZerQWNITvxobYU/25Gbx
5nGrMBds5K4PfhGYl8WJtDY+j5l6Sury8FoaCHFYTHiQCXgaQFRqeNhD7ykwe2vtxr6Rx1S/fATQ
Pj6gHfZqhJXQBCNG1Aw58lW16NZRATrTDwhYkIWlYEscQLMDsctXrGu1frJrNatSklV7hNRcr/+Z
LkoTHYA/7GO+9C4NbMZhouaburL1gB+JbodyOd+P9LnQvxN7lSCqhDtejfCXvqCE3RxGBbWvZJYN
fKvajthjU6aYE/0AeQcHybD5a4QpGnSTrfhnj4wD/wmtgiQYksTCSrWs0uGki2Y03adecdPjpI7y
oN+8gpLf1naqsBxFkW6kgm9pTZQf2GtQLwCXHZUFMplYsgii44pocvD0G6lno4ruDlGiqDd7za+w
qYFlJRMdpVuVWsQdoRtpfG7JlP2KJl7Yu+4A9p9YkAjgfO3XQuGy4PcweK8KPSw7rKZVdvHgDTIV
JqWtCqO6CQ7SnD3Exb6Z0yTITENpir7yOCku7v8F3dBmMOYBDAqZw8H51Sp0WJ5D5WmU0AVOk/z4
Gt3LPX1ihcV0x2Ma81EuNNzY06z7xhcuGRZSFqa44k7Z5/KZdQbwfngT+FHpuBzLRigLRBchH2+X
GLvH0KWM3j4ndBRxSp/X/wklZf6IX7HvbY9o4tD4BQlVNfrMerQhWsL7hsKw8A+478aIZr6p0Asa
Tw8kAQ7W7Z1X8SYJFEFy/uhhOS5CLpAu1UUj7Z6F0wGLyaXJvgpvkLoxUSJieOVBP3KLIGrYxNuF
sLWmwv/DcYvi7LOQIyLC9NmFn5ZnsWRBe1Uw8+JG0nUNbcc8iXHZO5olK8puNSNYqA145dUlC/5z
E7jXhTIb6uU9CcQDUboplHadSCrVppKvpSG7lUiwW2IDsjq7WziAiw31JVb6fTSsgKq05rU/yXhl
nDUtc4QFOk5X39Bsr9N3fGSiASmq2r+CTHN+0rpQUVauV0zEmBckb655Mq3EVQsg3xX4MaWtVcmF
9kE4hpDfu5hjO3iABKIh7hHjR3U6AUHa2nMGHWwJWuwSbgZSDuVqEa56JlSZO8V+L47/KSgJeCnI
kukRbDFPtSaop/9Bd3im+ZPIrR3T30ZKOjClVWD1yCb3iD8CPJiwMXx2fgSvNVPm/Vw/QoejOFFO
u7zZFI8dkx0RDhY+mp1uoqrwSF4eiaujLxkYt2jCXGUm4veKq81suQqUQXicGDHLy4ZNLXqKc8SC
DA8ugJZ5TOxrASZzX3Lh5J/1NVPZTnwx0eDvD1/y7MdoMursWVgDhy8xYhi3LAxqxbUQ5jdHAZOT
WhP39Ry7F1KWQezc9cwWrK4V9BXK/lV8Z0QOLK6Oc+lnO+OED+0bdsGdXPeKYZZdmg5jb0w+tI7c
RuHDsZUbz+FOAanREm4zl/j14bmiT1Rl/iIED1O38ehhpoR6VUfjPE32/UShwCVEZuupRFrDh0CF
Suj+7waRzyfqO2bDT1NpmqHVnDDXMbWYnwZNTEypK7x43KZwCctfqlcwADP6+SGCzpnxgPvyaHwF
qbuqxy2PaDeGSyjW3Ot99ZhYEUns1O4w5U5EA1/aj71W+sd+ir6/erM1z0rHHEdFnNOquoXZbQqF
RcXLLNNd1/bopolbvuPOt71UWuR8oYLNhYAxdlAaBc0ovP8NltlHUbx2crvzSeKq9I1zOA18DhUl
o1HaG/x3ot7fherzX1zkyJAOyJ7PkF9j5GdOV2LL9XGV0e+4lW2B58cwtPLMMklDLH1QmeklUgBF
f6bgnQTJl4g69P8b/rih0D5ugWX9OcZGv+CryjkkasjDApyn7W2RLShwqOr6xX/6wB0DjSIsRvWE
+JPa//jxyanCfbmZNdHIKaniNViOKwZZjejNpjzGYFfaSJRu1oZGcK0jnsrLFiUJ/GGFqINXTLr3
Kck16yaFN4691hqaZyjxonjzulN/nIPBT0CRDS27fTEJb4ZF5qbI9c5zcXJiU6bI54f5mwu3RFxe
6+T1RXmG0FJKiuSRZWCtlpUWe/sxoApPQv4OjvenMwxsGvLLhMu0Kd8lLaxudeabGm5h5umKZe+5
oZY4DLdnIM1IV5mCzWOq7QlvkXLymKs0vwHnzMGlrirRsSb+NbRk1RFCwDEy9pFLbFBwZ6XnhMti
mew2vI/nB0H+eI7TWOdjnxCS7x8uru8fEfuczKo3yiB9+Shyi2WT42/FEHK5bD3HZPfQt3Uw6J5Y
nN58Vx80ll9E78KnGkwB3WMb5+NELZO2V7BRE9W7WWRMy00jMR6CM/1Q1LFTycNN8yg1XO1JN45d
Ylbb9JsDXWJ0kSRQKme4M0dm0vPXlg31LY/t1Z95eynSNi0vN9IGyhek7KvQTsIpqPKLsRgvEYlw
5dYw1vmGL2EkAESvhV8WXfKmDZA6+T25E5g3UCLFQ+w063jm1BCa9rIsO/4qxZ3ya2rdqq0euMHM
xn5eKdTbWEf3V/NYRou/S6BwVE5VVV2Xg9MSd/TOoQXbBubzP5H1oy+z4sa8ES3JdLWvERvZXhzN
3y+ZvEinCy3Rq70hWflHyREw7WuWE+ffCflNHFvz1XhHBz2/fozykhTG5sHpQXnH64PGxvjFeW9C
ntv1AebpUcw+q0o/ROT2xe19BF32S0sdBJA6EWAvIHuFcAkswUTVkxpZiHgUgGaIM+I81JAoabW5
59602hGmaWlSsfVScXBkxUwYD4e2nEu51zHu44COGm5XZ/WyUAlYRt/xO2qzEd6pXb9pQPBH572h
TE/tcA+bJcH5cgesPc7W91qt+keci/gA1BVTRHuD7ow4eEZI4ogBeAqg6nPGD1t0DAq4KraopGzS
6TLQIFLE5S/T88Ad9LrVhA6IX8/czZf4y6+erzbEECpKmwkTPL5jfw0QB8tEgWMcU7/7fyt4SHn9
/ZMLKQlAIu48C6bQEbbC3tS+jAGQej92mXElSLaeDwVmfaAFT/oCjXSWSim7BnFkJ3EjzRSSKU8v
8d3+Kjym3S9/i/Ecki5dvN9FWoxERB579E/WDZin8OMbIG68s++bih+XkRaHDGgYhNKnaL7SI6HW
6v52AkKcT/p80bf270RsYkKbHFU2JQsYKHptyTpK/NgrXisa17CA3G/4obv+CrmKoW8X4ml9cJmR
Njz7aRlj2xKwsIyVY2bLO/w/kNVY/mYTqNgDy/KJTfvRAMymdXN60Sei3rfPThmKxALJhU2j9usu
WJi7/kAapaNAMPyQyg6USBGM9vZLpImZOSFvm2QFAbfSDW/fe6feVmnO99mj/NpuvuEoF6THGmDO
IBIUY/U2nwglQDjdotSuRKc0JCiPHPHGutxjGzI4/hGupQCL/4mh1QPsH6hzn6jLgF1mv4+vN+Xt
Cgij3+25h6E7PL1EQO0KPVE7mEJvVDsnJvzqQxeiC3mVGNJw+sOOnDPRKL0vlf/59Nv1l1tKOwyc
9pqG5wW9Mxpnvj0C2hq/mumVmjqfgti/BL964IDQIqyDckVFUlCscWx7tRih2yKiU0M3qmmfIw6u
mM0vChu3BnihrZjFOJyNvnIg+6wQQ++BPrNNECtwGgBmyHULkvwnfIM+vg7E/UilHNkwN+cUrTKE
AtANDooDCt7ZHDWUAzpbETfEvJtJefhrZeyUWv3CKyuFWOniUODrUHK4tokJ4t2zWr5/LDMLvFal
S1ZnoPViIyYx75qW/44Tn+Jif0U5rdPVSOYVsw9VsouSDnhKqxqmcTP+E4us+k2eZVPmQbUlGLUw
jxGz74N4BaPQsSQFhpBOBeSUHbXPa907Ps85G5j+PrJ1kfksd/bJ+LcYnaP7YTqcTYAoitPRYzbP
O4wPEIpR4FxVspbRLqajmb3aqrgTz3y0dSgLgvhKkt30eYupeLa1jai43pFCFj8tsmV1MzxHh3O4
l6X8JkmgdtkxVNvwqHqAyD/f8GmXeUjyvTbxlz74fTypFAEsxc48VHF4xUgZICu6i2mScDlMzDnD
nI5c3TknOwJxLCDS8xgk1YbwPeU6R79BdP0cprNlDtv1gMgsXFXi6MoxmnczTYeiUawymTmfgM+R
YoN5r1a3APj2/Iz0nBEJ5hUB7Q3psOBK89899pjpR6ISUiN9ESd0D5EQz+OErR1APr8/x2dSLjZs
HTT99fNkq3LzGbV0v8MJ8QdeOiFA445K0c3zwWTLiDMgk4nB5TemUWrndqP9IA06ap3H95kF/GQf
i9UsSzqn0bur8EY2w8Dzs5sv9uDxt+LZ63R4ajdvyXwsd532FaNMMyY+ZLEuJL6nkeRMAGK6P2Sk
hBDery3Uhm2kQDVFo4/uoY4aDmhUxFl5SCiJpydTbfHy46jk87ByLHqeqVg6gXlesInpwyPpnn0E
4IEioRtRQ2rbbsFEh5hni4f6AwF9IXw00SZO+8mpdhkb8rO06b6s3tAhPv5/QP7piUtR871gN2cD
z4W4lPdnN+mtfyfp4J2ssl77Vws7LZkJjWmTcg9Nez1XQp3c1tRASWBK245P+g96swL6L39OPrTG
w9O2+aKHorgv1Frl6i7SMNVh5IwCSanLq9W/hw/HnSbeLe9Z/h0JI/2YWPihgaqs/zhwV5DaEDLq
OXBB0Qa5O720jooecBcq7kz9kdjE8mZ9q2fXQb7MuReE+PqYALLXKHdZyc6wFMvC/mFQy57eYo4R
2ThEsAdDZumsNHjO5lzqL67K1q+P8x53Jtbb2+uoU1gQQieMw+vmcj7MuYSN5Gc7yBEvs18vR0jG
9MQZXXp8WJC5q5BwktWQn1hVsaSsjHDG8Yb/8sFGEZ7ojTWU6OmFAmK4W6ynho/mcQikiV32wAaG
l3xYIhKH7/NAmpfTHgwIswzhXY4eHmzZlDi3Rdkff1wt1S0CaEouN85j0dTfrlYQ/w2J5KxptnP2
H6020g9IOEs7/wSWODSfPQFT12JBEhDj1JQ/FOWYecgl427VbPL4/2NjljpctFunYtP3rVjeRMFC
QBFdCOMSxWXOffPSnqojpQuwG566+awKYAfVqnPkBSLy+Kza2M9vgeRbnYfeSiSXTj30Glf8xGMA
+2oiHXf3/m/N/G9I665D93pdCtgXtLRqQFPxcei7povxpwCcobSHGTIIDF2MmOzqaDQMpVve17gj
nSRKQW4/lzh7we1idEH22dWyzGwHtZLUp1EDDtrTqUnCZh7PGmdMQlX66woFP5mtx78I5w49gkjO
ODEub8ditZdEb312nh/+aklTWsaZFOBd1ZGfVP0J4tJ+c5g5qQ92Oyy4pXBELnj9g/zxzPOqZgt6
ObL8O9vPVRz+rtfN6RRC5P7FdYgNHzI1xULe7f7Ow5Vq9xTbJx+zujHrxfvUL7vBdc9Bx3TMFRE7
0hsizmf54+nupqysmoojEqBMv4QOw4mJab9Y4+zV1SqhOCxTwtCdvnnaLiax2axOQRO4pUq3t1VE
b7FS0CCAGOiuQxAotx+nbNV++9sEE+kzPgmoF3wKP7DAlPlNHK+F/aWsOBi2jQ2unjvizRIhRxaq
xRRG/CZKZQHxh/o6PUVPUfi8s0FXpBchh5YGK825BKWUoKdPoy4mtC9aplVpBlse5CNA/62jyloG
AvACWjgSor2Ctovhrqlw0Z27oTiWg6F9DsDQKj2Ddnulg3fqEu07IbKuoifWClTbO/78NagU91Fs
amlFJIgPGqFDesnr0w0+NfQ6PCH3cgcsJ15aBqUCfSR9hqVoG4zD8qIXGJO63y/H5/o3/vzKgFex
gfuISuFVoS8Afk4WpP4Kgn8PrfgrtYUcOm2qmOi6gtb0r50wMijT0dufs3VBfkaoJaTODOauXoW8
tHaOVbeu0J2UAuhgTnU5nkT+jCZyq7dSNYmiCMu9B2ntdX/E+i9VuKipuTHA/VxbZA+QayRVzINO
nVd3qjOjPJud7deKcd/ULKu47q0xYvA8a1wrxon1ZVA4pFWVIt8TmBkzJvUZ09Mbd6mRlNvf0VT8
0SZcORrUKf+lUKEk9MWc299hnyJDtaJzXlAGi78+OXCdj07gmCzc2KpVbMDByayE6LvlUZ1rKdyQ
H+jHIMXfQHvB6eaWe5PC7VjirV/qPe1Ri4epI18SRkJkSiGebFSP9mTh7md5PVS2pKuxYahI7cvH
mM5ffndKQ+k5BK/tMncdoMap+MY37zlYD80AH3XgaY7Myy9YXSTaLpGD7FGKIrPFZM/jWaK9JfGE
Q4ral6lzSOcd9sv879oUEYG21JqV7XnVoaJwFPFXHon9/Ee8qRoc8eT52wPc3LHfX1xDebsRf5rm
n6oG17y/+YQXveyAveQboI9hbhCHEKIhhjTZTX6vQGh2FI9KTX4ScwFwpLhBpBCAPkDRX8saCi6A
tqTM4yNpJVRWbS1v5nOm+2ScGk7OnVstuqAsPXsrgPcWXnl2D54wORhijX2sCG5r8SzGrD1qr57p
jRh/i5KUUpGPzzoa/WYGpNCdc8QNPF1h+lILiVKd04lB2q+ohujfZL5scRUggf8j6SuxGz4klP4B
Ax0ETCGa6fLthRWVWABCu4XKvecFMdto5CmW2ljQbdndC7tpytmjtxegAjedJRbVki2s1ClA6WUw
/MM/eoANVxzeZ9WYuxbgS8XlWgtYKPyRXHCrjSJmlQOZHtPZ5FHHLuRl2LgNBWWR1AEUKz1kgPGn
m/51tAukdzpHcGOCuvlMRTZ+q5TEcr4TxtWbM0DmgwMrwYN5bS20R/XViWVYLRuZH5+HatDvAZV5
eNaimjc5k4soqZnEm/8YNjXpMzuKn7AIgPfUUROdlJ/F06Bq8lMXXoSwP0lzieAKOGxXySwuNK32
Fsc8Udd8xHqUPxkBUfmbbSxEjwG27CJl4syRMJ1pyLQaOw7vjozHxDuDaequvWAHS2oDX19rcB9C
LkRnaKkGAr1kpDqitIz7b1OghjwKGB5ZF/KJiVpvQDs+UVS4BxJmbDNVNQlLS5jiJYAofvAB2Kjn
BVqWQ0z4JcMvcKEjXQp5OPqvQQPMQL4D67++bl8FnbzKmHh2ACvtW8yWkhwv0itBAQnXpMjze82Y
JQ8rSCfxfOQLQVQe6N1Qssz/9Lz121BCkYn6lOei5WhiKfvd1Xqf/1Z+7pZKQK2XIWRet6fSeT/j
3cz453JDCrS8Ti8h0EjU/sBOnBT1AfxRTdQaAdPKcM4lexqC7qfZA7PKvyM1RTCBGQ8DlW5xkNT1
LBj2v5aVD8491ZgQTOroGrz+XAESIixoT6yCTAVn/9UKo0PoEugic+4dx/Zm8BeIh8bz1jt6MXDE
9Yg3gRhRQgOSzShJSF6fPtghapygukfbAvo0slLu2tH/D0CzgvN8QPaxq/58yGhoVD2dyn9+/ku5
VA8Ai8NaWgphfb6s1zpf3PdSi4u8OeZvG9CphXuK9gOWP1VKDuClvOgrZvyqhgAM9N5vysiISRPi
Wv4MMm8s+u9SWJ1lLiq/+T7xRo3XgV6x4wqGm7OhRpo3QyBsZcVUmTu9KydqOWJd8wl/VLiDr0eO
PmT2NJ94oO8RVupAm49lElSbDu+dDkaGfFmY590TR5QGkYvLtUz+TscD0ZTDV1vwxlKoLbZ8G+W7
VbD59Hf3+r2hIF2Gvk5PuR4b+FSUlGb/5gNWFGS8lvWh05idftfM2ZyxwzCI608dma2V0lsQFPS0
I/p8Mur0JMNtkpY6FIPevnbco/TzC9nQthwlAwt4HNREj2Yd8iqZY/bHR6d3w8yRkLCc9f4cm5oE
CZkB0hyhR2zcW5/ee7SmNHDw12XIXwNbL+DObEaX+cLqn68DPHJ7ID6hXonVbj7ACaA88ZrGfi6e
1Kh2iLNq2XQ+EozNwvbaxjs4wWh8M3+k/6W5XoD3fTv/ygdvf/BoZPlT+kjq191hrcF7OSX3h0g1
KgTClVM7Wc9peE3imGxrT8ehJz3RZOeDoCpdiV9x19AJXiraRdekMQ+tt8upAXxOaFWhkIKbjgTs
B6qJUxe6gqWMYF6v5ymUqO8Rdql/8suiD7593Yxb6PLNKh9Inr40Qa5BdSXo3+IrkRugH/OxKA2a
tC5VeEOkJ+nEU00mjmqK3gkcq0OiJ+t6gGqe6C21daSFBxeHRPQ4UD0a3+qJJI7F3wBVRWNYSait
PjVOXyD78cImVtrPM1La21LDX+JEKKmpS7Kl/akni6XtS21Ut20Ndx3SoifnhiiJH3lgRRoMP5VB
6eN3g+JF4S350dimVMUuTleHtKOhgC9OoOcjEa0jZ6J/bN2zw7iVmLxo/ZUtiuu3liBG+rsPKldn
6JnbOcKiGi2WUHvz2A5tUmYk/niwr4wdus29N0PWueJK2TNSo2RaoOKTbjMHoHL3mz5ryOwwMIgm
Q0f3KqmPm2am7/ZIOuh/RhJnuD2P8MvP2JoOsFdMebcahNrd2qBvpo8wmLHsPYqdWUqXA9PKExBy
aC5Ag3Az950frJVFRhxRXL8dJS9auPHrXWhuY1uu0/ZPJBU5AD0dCOGLSSJcyehcDPUxYUOoWreu
e3916OOwIKoQJqSFdxtoRT5AkvkoGtpTxKE/VEhrLMieSyLHnFTVAGOCGvRtVny0qAvUMQAkybMU
uTChVzop4fLceR6CsckBLGHy6+5sdtH1Hyo/YlvcQJgpkkEJnj75JB8EwHpzLsUZn+yQbkPsLK2w
ZKksfruwClyAkGkcUq1rGDMKrfarPD2QhxWE+zxB5Z0E/V2WSxyQMc3OVEejFBTH2xODVEop1h0z
8qMf8f+nR5Z3CvLmkGGRVR0/2NeH+Km/2LTKhhskXsRfWWj2rfKlrZB9oqcOyKeCQmoNg3Nw3Kq2
5YaQKxnwJ+VfZUFoXqB//zTgcNG3d/c+plQCUxm+dKb6Vy8D65l+2HCR5ClGWGjo79MF8W44k63t
iAPMrBU6Ay07GnJdii12Cdh4I6F+8jc7ziVYTtXTVOpc5G7GE0kzqj/QE9SdoH6KhLWshVsab67R
7qNU1uJFPWKM7e29WJ2XPBq59bDQO7ScA4yx4dr/aWgxl1mBzxNMu1PfBFd6blONh0BtdHL+BZ7M
QDbYNOzpUL3f9R9lxKhTSykzgW1yomVikjVrClToUwyJp7uUZ3FCVV+y6yhn+2zrNVIjRAySo4rZ
sAB/6/FFlsDuj2xDs+AIV/MrhmyB4MfkmPTGPD8fg7nmuXlyvO/hcx5ZkYYm+bp89BEdG4PCI8d1
Z127yWhpY5dmsaDvTIpZhJcDLcfRviFjmUjgxLFrFTm5Qcb/FjR5aWEloWEJtb1AeYoOg0ML1T0S
ofp0n52FHiW46kLz9ueZWcUs4Mt9cikOh2dAtECHco8dCzuZK3nNP8b34Gm8IhCC9KmqdV0xQPUo
5zJC1s02yzh4auhSKJR8WKdEhqb1h6Fy23UM4iRaJiVD8XWyEIBwPBkROe6rHQxXDfhXsvUEkSmq
agseBr367tgcJ0j2gAcn6J22O8bfnV0S0lsBRjxbWET6UFywnsdfg+SQXQ8hwX0GkjRi+q81W1ZY
rQYS6zgNDZFvWb8qDk67RNRWl/iquZZsI05Fvktaw8ss1oEiNy/3Wd3ltlzWsWtznKw3x2FANaSU
Ef5vJX3r9JAi5gAiLF5bxsIT1G+9wVfc4gmBXa+S02O/5yt8kCHFdgVuKQ+z1nm6V45HDLwgXXem
KXupRTuY91v8M7zb3BKtVTnghTpFd0BcFTU+GBHSMSMeXagYegRiywjuN6lAqMwLO3ASlyzoIvhF
DqEJnGJn6Wifet2Ok7r133cCAmptS/kdaTSXxJnzZfF1HKv5ZSrH7Bj8NOvHwhUdlqIS1Sfsqjn3
IxuRaq4qj4Mm4z5MMLt/5vcPmfSobcz1p6sxM2yfjvIraBWtDeBIsLjODJ6QhRWj2cvrP8Y7CaqO
U+I7LeiiZzpAUI5zA1fOJSmPs1EjuHb3H2VpPE4/qzUhZzO8v41Y+GvxUm5op35AAiWhX6mslAux
pq7SzmHMpKByjnNMitjLyPPOSPcg+p1GKwL3RoP6GactTe7VPK73Jq8fa/rGVH86ADDkqjHhay+M
mwXrkWlnE/PgZfNmuSE06MtJeQ2hIa3pz7Ts18P6xRt2Gs6hLMbG5DJIh92IVU/ddDgp0uIw+ieK
oxDq+Ty4BOqvawduEdVW/FVvFcifo0KJdPwEEjHTcDc6XkB4J17YzUI1FHKa0RRGQWahhaA1wG/6
HJwGcJD2W3IXW4iOPmvUxPXTkP36Ftu59TP4qqbC9vVKFPRt/kQgwsXeTEHipHUm70hrTXM2Jq89
rwOwkRCMYNM/B40+kve08MgOl/14EV/9uhfa3d9GSBQbiLTzK9rWnYCLQkKCItNscOmzJY7Rj4H3
TEL244kJWpWpqSgpfOm/euTTyyXgfQosRTSGROjCZMBEuHnEOmRzK6e3Fsm27sFvtZTRKiMKZ8uN
sIMqdpfuwTt7f9N9P4527c8OJYln6usCfqsflRG/+6ZGM5nw/ZRCAKHGJn5TPQbSUOvJX3MYh60O
/L8EuDxIf53R4OjPCrCKGLBc+SnD6y9B+BmwhDz5J2G1e+95FbdnfrnywunTJWjav7eVAkiZkv7g
+c0QMqRlj/5SmXJtGfhYA/K+aTvEh2KaEckim+rY7zlG725JK63jAUrCjTtbKAaTU7GL+6U2LHub
/jUkiTi5ixNvzRzkoKzuQz9tMadKAg2WVYXTZIt4T9D+h9i6wNL5Bj5LOW6o1ySevVZDp2msR0r8
F6OTp8NrdYQhtyCpKLx+6sH0CrKn8HQt2AdBSUfdocICTbAZ2PcyexirPWuEuttWZi19MIOQD92t
GGxSEKxzKHoGpoc23iyqIhlSsg/puPHa8OENB2Rt56JM1H48HqPWdJxcrx3m3vC38ehlKwLFF0qm
9N71R4pkynKUH+pYNenTw50IFN2llkND9GACR8CJou+XRZZ9pLt2S0ciDqF5/8GDK6QL+GRGsXNS
exHSRMbRM4NFzecSgrancSREB2eVG79mGf0XDhmu2KSmcZZ0/kR3hyacCdiBuLTebSC3B0Lkl9ZU
NDSD0/yt8cXnZp7rjfTEbAAJbmwE9UKm8L9AX0niOEjhELeknOtt/COk5hY1iXYRi9UOKDcbyfU+
BMTs1MZmfm73xfrbed4Q8P49eRfxIwFa8s6y2dHA/uyK+BPjNm/O28WE5UzxF7i4qalsqqyqrmpp
i8qStVpGnytDNb7bZgWK7Te+WPoqI55ZrvaQkp4jBU62MfddU0i6MFFN4GA9mP4WOGSNbpeXMs+G
roO0DMyt6Yy9+rV9QDlf75mnfw6faZKr/elDr/41nRTG9JLQ68oUSOpF/HocdtgBoYb2k6+zpjXI
xYNsMvLv7Mwtrhqq4lLyhKl8Ztm5tNY6cvafBqyl/5JZiVK1qjEorkJD8eQaUeXvIofmygeqPdzf
/eORjW8WbBw8CNdzskUUPkT4+WvsfdgH5+rDMN9m8Nlev5SME4zXpNH587BdBU+eh013MCcjyhss
xoVqG00fhSxmt6PAE9jAm3angppkPZ7UOYQ/tovZAnLF0yyGLsHFFM8e6KdEKh2BH5T2e+Hakq5t
y+Wu5hjN4fKmLqGEKtRNqqMKDj3qn4ArkrLbtEaZ0maiXQsota2mDKtXX00wgqv6DiNnZCJcRcwe
BCdutK97sSYxwQqTk+d4IrJA+h2H2ldc/N1zqKzm1AMkhFvx2Ui+MOo+lI4dkapYbFEFvfOHUzKj
qtcQzvxb9FkxyYRsApxw2pcT04us387rGuu8rdUnP+FD8Z80Pf5jPpnbAfYp02L+9Yuu3BJlRGMD
o3k+fjamK3DbKmjnxvrSRksyrwXha5l4XO5ZzF5oN+WvdUX9pr7DXYwxStWFAKDWJnE25xsXYu1q
nA9MrPnuRQiOJHo8dZ6v8JVKvdy0ycTFM86Cobr29FxjEeBfx0JgID+ojb+pI2Fc3xo8j58e4+Op
drAWCl9r55kgNsrH2Iwj8iho+nnRiVC9MME3ZC80b0M4/h6zru0Y9WJ4Xdq6mSeAHF2yH1zS7lCy
t4f11vkwxYxomRXz1kb1R4EcuuQhi8SZsb6IYFozky4d9wyjiLwUV2UlstT2fyy+Wb1dzuO4NyJU
i/Dvt8wta9LOoVDWIysIe7/8NuzdorMTFsd7AiqXj3opEy1F2p4SQ2YaEcKwqPz1kuIAVQcc1Ygt
gm1bZuHkyexkSak7YtBxM372+utAi/1SiSp3dazDTCNc+0SIYeoSEQkAH9hS1WgeYKb2beImcAj2
HahGjdCjTEbhsPPY2SbB93tiUlytvDgyxj4++LkevqDvPyFiASwGi3fMYGgSx/VJ7KHyW8lwvwSh
VYTBVVLVcMNfI0+H8Ma7VcoE97uC/dYgSEsIDvw//f4RjhKgV4hg0nKqtBMfO/KEpJMSMpd4wl5/
rBr9U4yS8V4v7ktGwChAgDk6NXpS61kN3fNvnztAnsUTFjmu/Qr1V3KAfs6WRdmRTXkhLO6JHH/j
ib4CPC45rAw3FvyPyc2OmV23qU+4DWNoxBKQEom+728Z3FJTuizay6nvgqCAC+h6kJITxyFjD4n+
Et6830USXqSzbVOsNnZfx54+IOQ6PF5JoClcR7VyTAVCROqjwU0bEtSUKtj1lCHNUsl5KfhQ6A2m
pItmAffkA9DOpzz3YXqSj0r+gHJibmMBvW+jJSXFMYCuLcNf3GsleGFciYAwQVfFUhXvovxzFgmT
isBSmf83Veud3sa/obpAcqnr7kosZ+T+bHIr/hFqfzMZoPDqwhQ36enNSxBGw6y9xHuPyMRMkbEP
j5EmjPomyjoaKpsAXwDMHBOjSB+sGtUH2KPsOvYz2JgrrSUysRepbReDJX43Vm1g5beemdgFR99C
o0LYrQ2WC2mPoZN+usuw0jqVCZyGMwmdX2oXL9bd+RD9lA08+HPgly9iPoiN3crG9i7Y3hkqRMcK
k+VdO2Gv29wNohq9NZjOslbA4hu5Ruzp4+5dQSQetTC8yOCImh7HDl2JTQFXSyf+mMBSjfcAaf84
xDwTAiq1Dd8QeINT1I7Yi0+pN3sY7Y2DyzExrePJIspT3c7XxQLmxqRQljVyO324O0flc0JqxCpB
VTpaOU89gEpPuQco2faGkOfwJELArTDOE3jo6GuKwvX3ILPAPVF0RAD4JO5APKsrdK5XEbV7ma6s
pdNxBS2m9tWmj2F5NUUOW/KSENp2fGu52g4pqke6gt5dcGC0kd3DZ3wPyffY9nFI5XPuMmsurOqC
IciNhlpeteGPS6uVRSfwSahItTTRz0qnnjmFfkAEdgV+y+5Wlx6mR03EB/7K/x/kXGSSqvqOFWz1
ZLRFX28bbXDPx3Q6LT9kERr+03jRakrHn+Vc8oBHOx+JFwnFGlellqxMCKzWRQKoxGIAF5KM5iER
jfV++nXNlSuDkkR3GIRjMD0skfXgCneKA1Qs8SuO0iFxDnTotD5rzJfPCsOQ+bC8YgiHnX8Is/I5
Z5kzQMGNumLoeXGteLj0bkb9LZYxgSbdJcE0GrlCOjHiKNc5bAb9D0UQUyk6x2qzoxlCV0lXUB3D
CPQuzGecCO6ORSC7ufWj9Q2i8V7WoctCFj9G3EXhnNxUXkhn9+27Z/TBpm20iDZHbhVyAmoZ+rxW
0S7MFJ+xJwJ0XeZlD8MaD1R54B51gI1IF7n3RVQlVkvzFsv/cwRYncQpPs3WG7U0boDJTnsB7nvu
9bKYRHHghb582v4myNPdzww7bdZ0+oaRAmWbBnTh6EiSyZzZrwUREiUQOaAaLS0UPw0e8zR8TMW2
BF7J7sVyOL/d9A0dHej45Fmqr2cgLnuJmvvWOhTCyxdIIEvv1IosYB46NNSZMyXdgD96IjCUZ0qK
sg+9Tbi87pLyyvYLYafRn0Fr5Vra5ChzL65X9gnkAjn9TvXJB7JRXtqX9m+LL/WWfv1YXyvpF0NE
9lUMsm3aH4YyBDiLwqj0WjCigQX8WJgweORgO1yxnDAwE/l82+mXPqYoKoaqWxkcjhL1t1K5B6Ki
fsKIyXmbhe+BZ61m3l+8IoeWWVQRZWYlUbKKJJuuPbk+17OKzpnu3TUi81XnBwVBKmnFzAfs7nkc
Y5LPkYgXPjg6v2752ZLECllTcwdfETiDtR879thbXOtb33UqJfddzhpeFVHk4wqrZmVcIIYTrHKr
DWNNvxq45CnO4PeJ9SPrAgtPd3EssIfB9lRDgJZ2X92dsQZNtzK4LkLkJK/+gNs0jfJVu1A4hBZb
nBVwnR3OqzuveNazgPgxcsQzWgjJm76QKZzo2uhVknluu2BDC0dArPni6mOq9SId8El2p69TzBnu
Q0CpjvqSBtD+Kx3fNZ2UQwQ+9By6UsO2HbcoIxpsvkSjo24Sc8ZM142Vg7wRS2J7VbTf80RkB/Z6
WYRsmnEjpD0qdrN9fZXAGZJ+qHL9+KLjN0l1jfELJ25doAZs5gJeHthmzRbNGTJzRLnC3hbz8XDf
omyhZPwH6X8ZSsXm+zDOkFqa7ClxUHOs/MIN+uLCcdQCugOYfsJt9vqYg1vCc5PhJjDKxRlUh9m1
AzB4XoYrjmW60YK+TvSPj+BZdU4s4Mmh4z+WIyxq42VYgTNQuGlin8AVNaaSeXgaayggq/hoVphT
FfgZ5ssdwrSfSI7xMwc9qSBKZepDwJyBd0EXGMcuCGqsT1KpQud2OMumpgp0JDn6jUrkoXoTTPd7
fiwYnSJ6maTdphxhViB+rzJFQpLgoTG+JG69N9TclbjIvkBww4DciGTgwLkiNFU7fEAN4lJsjvGR
QT3Wt5viFJGMp3dON93Lry/Zdxl0r39Do7a3Nem0ZWvdbezFnI+6D6hwjPKZwrzEemug1qcDoq8Q
EyCPim/3n6VqXbVPE/aZnsWTAylzH1bZuuPgMvO+j5EcFmxnp8Q9JtKqiAPbEcRWtVUfr5T+5yXm
nL0TCfSem+kUemBn0S+SJfqz9xrMV47VZ1o/i6UYb6jVXxSJ0ImLqj9T9TLd+cI471UgMx3fDzN+
5/Tnzn6y7bYfwmw1N8aF5ci4TszJgVoUOpwPbc+J74UHMh11bKSnSIrDEQMLt3/UFeQMbPaEHzcy
sTpjw/HNK7ETsdwj7TUMVKErvEB6hjqQP8+uo0u9gQuDzP+pAW2xtCUjeWSGpo+F/b4vNLY7dv7w
kRWkQRZkPXq67gQ0EQO93/JY6sF0rvkeU9Q9dSY8olkZuU5/Q1tnVxbjQAs/qzm5HtSMU5itJork
fAr2Gi62RLlPjZ1gAnkzg0DWmVwVauOwsCY4WeN29z+zAmTlwXqrU3inNwhC4PvdYl4wEyuzkMe+
3p6FLQpfC7stn6YHyUEFAG+yYuq/vC+QxbouXJ08UEd0bW94m/bPdtGk1fDxv+09I7ZQVIBlV/WW
qpmg9O3pYV9L3eFcbApzdqH8gfSsTIES6oFwj2wR/Z6dky83LMB9Z+brYMnGdONdknYoNS7il2F5
H41FbMc0Lt8FSqmkQ4Em9A2iWO1Q8TBXBuS0Iqh/r5HwL11nbmWiZ1uAClYLjWdLVTOhKIdmQPC3
Zug6AeWBCHhSX3uXPIcvz5uMZ9wkXQt+96SdJOKaYNx+rc0LfNvsSMlQ55gCMZG3i1D2S6Q+aU3w
m5Ra4L+cVUgl9Ydc0AEjBqgIfl7KIAQSQfZYMsBoOFEpA56zoE6DrfXohRRj3kIYXUzrqx2ng3bK
bUgdmY0EMG+uE7J05JLqDp85kUdus62Tmw7QN27KOGNayPOuCX/BbF29qwL5jxQP4wwTJXjQJ2PO
I1ChZgeTCq+CHG58OtFZ0WEe+bG1Yq3KxOC5C27e23EayYycAmT7VK/tPooObtmuyh0IFLsciuIC
1eOw5wLQyFGrMb+t8hXLE12YP7osXaAiu3OB5RW0+IudR+U/XcaSh3YS8YgSTET7ZY14ZjChGR5n
R8V5HMoMG6yIQZ02UNcmKexcjKnRuWy2/TQqVdnX1prLM3QTxhqhYixHj5zgQLBucirhPxdL7aDP
HGntUE+i+uqTUAnxgdUSbSNMJiMXk35dYJunB4tiyOQb4VIq4TcU3fG6lMpsmzGk8I4+MlAtra1e
OFCP5RqvhdODgEkFl4gr/zCSAF7WtblGlWTedksW6CJ2ofmBnWdQRfUmujDuNh1uHFPjuowcqg+8
vJn4bUgSQTVM5cD0j4mwIYXVwLy/ceApv9GvW7pmvpVKgo6vewHh3dElOfw8Dt2QDBRtuWarB2tR
nnda2XwV/D/uKovB561eNv2E2nOohPvUecwk6QtfqPi/Ic2qnqiooyTvOd/rcb+oeYSzmhoczJUu
0dQeic0tka3unu1kh9f6h+E9VPqdlMC713O5nvWBpEShobvP0xX1sVo+oOFoA72IpNt6HsjBIEdP
Eg3EsOhhpgXjnMBlcRyGqOc/JSHXI+eiyzf0a1Cwxenxpt/yqMlR6tCh5sQZ7RPXuPevLaHqecL4
o1EXw4iDipUK/EOdR8cw4+a8PcqWMYVOJE//HNtNU2sNnB3QlTtuK64sM7/iA8hAGSNEBtJeGjl9
Y0CALfSoXJa0DLSkcCYqMkukDNMyM4jmR8x7E6cno//KcUMa+nkHSSss5RzxLMnHwF+mFbjV7oEx
LYpN+32q3NHwtQPYBcoE1rw2STfIvacZIwCdUZBhslYdh23qn4T5ONQ6VC40P531fFryzutiHV5n
0ASLqDxPj4GbHrHDptfNIjf9JfRL36T/Gpgf8vD7w6BtGqyiysbQhUZS+Wfw6ixxBzFhUeg+iYEf
Z5u5O4Drp1yvRGFmroajUnc9TDKDTpbGE5Oho47GMOn1UByjzbc000Dvw+ZeU6q1/Z1JX5toibYp
9yz1MoNmiwv3zV5QCcwyhZojbr3yRhWqPqKdvg/sYBa8ich4mnCOfhaVlpbGiTsrDx5nUbGwqC+1
krMSMh03iASyx3HmJ+wpVGVtt1nOEQDf90ZIjh05N4jUdTFUPMmlAqr37L+0+GVW/HY9bU1Tc/Ew
otjupJTSpmReIKwaT4MsXIuG2Po0YYeFY5TpGMNLrD5IxcAdZf/6wz9bTIJCCvdfMG6sgtRpWsJK
rvB8EdcfHYcDNIAeKFFhvNcXkGjCWHQFkIGfZTr+6xFBXZLbIsUkRyVp6CBRXY+CvkOhziQJGOvO
ZXJSyYdDya0eGjipDTCe3qFXyUqKdQg8lojOCUEOWySAEmD1Ghw36l39Mw4FmHIDMhvBsxkiYdFh
dc/V1FWPNrZO70yu2VX+ZZpYFdKA+J5profNq0rgCltb9gmEN/Zw4KTinpT55ab5HdktiVbPWu+6
/b0V8Jbg0YM/UACEALM8E9DSEuCAEGzu9QOTY8eiP/twTdDYHny1oaOTNaDUx2HdbOStmfF036b+
AyPVHL0uXpuFmRECPfopZXUbuwsYMXhwL/TTHWxL5cOnKIIt2ZzdB6qW/PM6TnX5kNj3mNREQzF5
AXYFbdocxJyEQOnXHsRGdi2t//bougn9Oohf80FArIyZt+2riCKbPatWOYMCWbpMgitoDaaBSAOy
8bk713m03SVXowxpHPSDzw5IrO7203nAyxXbx4RAmKrim29PDEEXk8V3YbAu32b3bHkF2dNv5Q4T
3nDDlOLgT2rwtd4Ygw+mS8wl+m5S0Z5FrULedFhp5S1LKLjxc+7NbaI+khwdgx+JwSTlQ+f2Ww9v
S/a73jCLkh3ZjBWB5YAIMLjfCaUPPtBMwjcko3+x3YxBeWPSk7PLMTlcZ0mjRLuicz/kmlIHokuH
+oUS3R65RcQyZy1V2m4bAwfunVhr0eB2WULXX6t7TCdSPfd0xHAhiOMJ1elWq/q5v6Xr+8kVW4jj
viBG0FswpYxIlAovluMLdiiBaZqVvQ0q9r0ZR+xWKuzBqhpldKCKS5JK0ZpIzm7fFoOkEqKH49UD
pLrTvEEhqowCatMqq/KhDZn4aznTCxQM3f1XAjF4ct/+BBkVdLy8eV/xtwkXq1kHJGb5J8ognfq9
TmrYuPSARDE9PMbn451g9sjEpQRPSpAeuJXs2zOFgoSfkjVhPqvmGAAHeCmN/QPVg+nR3zxHNLl7
addKf0+wmqUYQC11yDsm/Q20SSJxazkTqVJdnVRK3H7I/jlC2yMlx4quoFjFeY78tUQ4mPN+J3t5
r+d+yc9F6weYogrA9/qx1xt+Mw6OCQy7qufvSPRhJOqywIrMBcOek60ObCUUZDfZxBFTYOJN6+cA
8IR40coKHTCtiUnrfUOqg7BFRl+abVT83SUo4rmjahhbBcpdEWRrip1WXQSJgBcUmNLs6eyEr+3G
SUcLsglspmKPHMqp0nWWi2nr72I85Fp9/uo1pObH6RhRyYroVNF6gtrKvNgcddSEbeyzL05H0BPH
dIG5zoRBlDwIIfWG+XcZSfGhyEXijSq+NfV+fqjxgsF5ARq3SsxLIwnpw71o1JGRFUrZKMht9vA5
dPT3fK0Z1sg94czv1dp9TLFy+XOCoSOCOqlIEwEazoshL2/nXpxbiDjoe+V+9XfptpO0CWCq3/7W
MG+Hx8JwSLdR2b4laTb8jyz1EN1lqZxNSRHCQYW3VNg8nD6Mng8aLHijVOBzDLmpZE/CPNqs7HY0
wXaJuacXFmbZWXaRRoZip1hT6UyEogNgXA1OrumWJBNZX01eLx8QMwl8TzbRbJFPr4cX841/mdJF
UnERxW0DU5/3BWvUjItUN9MeQxJOE5B/uNFj50pkLaTNU6DaRzF7ewRwcqMhyDUmkYzNngZQiWmi
L5ySWuGc2fyrJSRwNvraosjr5ZH2bW/Z/LZqea2Uo9Cz6SBlsLmUKNRx/YXIicR97VPlhCwk+gmY
WkGonFdl9j0oVCgAVg+EKeCdJMLBeFxEEaXGh+EECAeKGzw+AMueBWDP+JewKRYcybl17MKfznoM
4JstyvkHlI1QCLbydbmB5CZOwLCk7q1evcE0joVhzID8xJiqKJOiCKFkq4OdIAnkbGNSmclNwtZ6
nu88ZaHqhd60HXzYQhL1/dzElFjeFIFkjTUDc4jsgVMoaqd3VyNcUs4QPZ/48rcp8VkUQyEhwTeH
6SRG7zs0vYIldnhhZ/BP7gbUjj7X5bumOTfAjSNeyMVhw91TwoObY12ePzyHQ2dCv55R+s4EXsev
xcZX6o6zDP+Y0SKB9Dtoj3MFZfLn0Dn0mYhJ1JV96OYDXtHwcGalJ8DlYh4u8J5GArwTUVuMgdlO
PVq6WVMFAtUqm83+dR+Xjo+DkIIGdQ7emJf3pKFIkD4Vn3rnTbCGAZGdjF5H/rl5SswdZIFtO4s7
brURmg6Tln7FnRyVX0cm4iTp5yEjq5pWxfxeBmNLV6A4cY95CMw/CpDXacIwQdXC1MwFin+0/y9d
tWyjQqdrYKxI7BEmCX/bGRZVRBUX7q4tKSX0V/YIXBDZ/gt0LIK4ec4h/PSFB3A6Lx7FwHVro52b
Ay35RO35XY9Ga9MjcV0IP1uwdv2hUvVVCbWWBB4uw7LFBddukYwJwquar2ZsQePC3sTdTk079Ij0
/CmDJuBZ/69FxIIqEjgJrZiie3urRyQUN0/lHqGwDUjPzKbqFKN6Uc/8eGdqm1hWpa6/rF6mfZGp
eKyL+Ec5Wiqg5sdg9aVbFCLUxOYTZbny7DVs6T5BGXbVGeuZ1nDXODC5L/Lf+BXbmQ1WGX/C0bws
c5UbQH7CFThhRE+Dizcz3z8WgNAnNzRlEzOCCOd6F+KoYEZDPPMG0CPtJh/PBCZ1aCSybHhClLD3
TkXi+lwqozHJAaWN9sE6+RTusNZyPr/1jG0Ms5cUhgi46gLUmO5c1bxm32Nk7+qg3qyzThp6pGdp
fc7VTbyMqHSCeznWuHtOqu43+houQ2USwXTe4XYFSihzosVISZr0lBAas+33bXhyfl5+ZgQobbGE
Y1nazLbbLb10v5f80aiqQ3m8A2LXBEWdP74q2/pUF9QEsaiG/fthnZGiKNC584lBc0y64DEk6pmb
90+Aeebcdr2kFFgzUxyD/Lh9PqT6a/Nyhx1Bd08pCwsw5oMCFVKbMJAaXRS9hADReblPaEPs45JQ
/BzkYowc2k0wyUihI81CtPcm4qOLF8FqHaufEeHvYAlQ67rTZGjMX/YED2yYQzDJ9hGfH/NJk3wv
CEw7Avdq1gxKAl8WkMhnGYhciKlsitK4WPV2STMBRoKgcTUYtV1DDWyztO4KtF/z5svnh3uPq4ty
HKbLZNwPRlNAiQZEJw90l35md8NiEGQc5rPWk8xtFT16YNXo0FDFV1CwMMkaIdJMwXX2NESQkHtJ
7aLyThVj7GHfJgFNJG1iD7aAupqD7nqcMGjYi/dXCR6ZihYDEpHwz64nRRpR7xLrNHM6C9/1Qgr6
kY3nsUo//+RJBzXMpNNhNuO8bYcGfiWC0Jofn4YL/PHkQ+AtWNVwxizNMVJiDvN9P9qglB4cqrX8
n4zl9m8ZOd0HnQehax62dKwawlqRiWCRItfIIQLr5V8egYXAV9BMu6x1ylNrCATwawYfUPYH6R1F
1kL/nJ/1+vdKnHoel7C6MZnVIikzlucgjEvm5sIE0czs/Y/XFrBbIgWJSJxgvfObHNi5IUeP6gXY
RSzrA+14qs8AITzfOr76cDCdx0sgbA8WTq1LukeXs67pDpV7csFTJMHLSsNT3X4I9rk4i8SgfEkf
9KI422OrNw6NZuOaMH27ORvz5+wTfIpymOW2vqBYtAGWNiT4t2FrMv1zwKVcLr/QKYMACOoUnfSc
HzeAGUY5WXMEsu3mzfWEJpcuvffYQvzN7RZPa9W/nCRlY5I3Lyh7wMG4FJZrw2F7QeFmPxGWM2f3
M//VZ7yFUJjPWqDVlHPhGgASO+A2wpEfCwhGMoYtanQCJJQo/vaucFpnQdhK5u9LzDG8xILBLlFe
7NlClRenNTaN1zI58W5TVwPBys6PoFNuvBBL4aZ52YtRFLALBMmHP2HdZT5P5yaUyMup/dzGh6xz
v5gl1gLa5yXh2canIhBSwZmtmuVGv0qPG2f6iswjLoYso/ETwxjQWP66O5lXIUEzgTorgPEjHqHr
amHMYtqN6bhRhmDdp+FV+4fbVxJLgkvYEezaegQHtFlUfwhkugsAo4YaZztxV4IPOvh7Uptq/DA7
/BjUZGTM+xOMse73d1VoR3aTvYSglMkCUV8QKAUq7J+Y5GHe+o+TXgZM5J81O8XXDbRo22V4uZAx
you8aqfeSnJI3wdq8tHAV0MUy6cUWmihk+slmvFfncvxLU7hle/ADCiSUDczaBV/bNU4k/Jyd/2D
T9TXD8013WYP/Zz4DjiNn+GO/emcuHvWMm9b1+7DBM6lduaXDmTpkWBk1jltnCAUOOCus9TyIjDl
cKTJcdCCnbLE4RbDzEXFORzVrd58PRqAleiMmpkWYpLsjAgQVclPznUiCTMfCsz3u5kpHfPfANvO
2MSMFX0aV/BMBdExpvR6pBL8kAHlMH9zGj5ugjzOwXe5VlpzHX0OzVYqcmMY2t+BnPCgibhNNXXf
36CxrugRYH87OGvgpcOMRDPSPusI6+MvOPESRLBuLAWuqmC/J/I7OuUVywrb6DN7gcS1Xhr65H2w
F9GGVfJxYGBtHIi4D+3L8+Bx42hXpqMInGFmaZF68uK6auOI21KBPxE1enLsg+3Fxlrb9NH/uMNa
n8EEX0PLTFU3FPiYO9FCl8uqylgE0BYh9It95ZDoqg7YooKUKPSTKfE2vMAQrT6YFFoFlCuxeDpR
H9WS2Guno4vAxs9cfcm0zyfoQmFuTCwC6QJ3gwu9R4Musfhpy8p4UEtblx3+RLzkJWMBRZMCLmoW
wipLU75KZCKVe1G3E2lO6e/DOfvT5q2vWpNxz4mRukQFIYnBdOaXRgMx7CsdPDrol67Y1xaFPW/Y
UEsii+h96sdGHpO0D5LOurvYMZ1tVptdFx1tRE3fYu6ddEnlBKjik4HNrQ2lTw0tmzUbQqWcX/2W
HPwLEGQ/5pkXcLB7RwCLFXAWqy/Hsk+Mf9E6cEBnTfM6ihkb7kH7jbXuLVq+3SAgjVRtLbdnMdaE
Wt2JWgd6lPSZkXSCw1U8oEWT+kFyqVXiRNNAmwTjxXiiAXyXFSEZcmBAEuCSnxk0QQCQzy7kqN4H
QDCLlQ3Eyrs3AcwChqGpqpEjUPlav4gJr4gxizxUNgjlWyMMZ1xPeeyAjhxG5IGWe3hRz6um+e6Y
lUtNM3yuA68J+BnnKp2NJ1uKb4LR5wBiirBC43Lxsi6VMee/WscOFmFui5LtRiE9XkRmXEHeWVmh
GjMl1+KqDf+Cept8sxfbCy2MZBUf/ekvOcpEJ6ye1eCa9zHNDbypJSdnTHkHKmd8J/SabAVExuOm
EWvR8BM+eiedh+kVrE+iQ26Es/IhieNHGWv2MTzXBC2sMi5/JM8fDGRN5AdM4kCB1s6n3uJqVE4u
TmRfC/FfXHrQ71fxoWiy27A7owqlQIJ9WIWugCpq+0SfFPLDGbXha6hGcmNtaxQj2vsE5B+cN2JZ
+cRbT+g66gcXDZYJIVSrzATiigKSw15ofqfkENFO8KfjZV3XJvEHFaoPuIMo5v8dRd7mPFibTdzy
jQBGfc5t9+B2JcF8KaMyEzhu/hc8C8R0D5MNHrPoPpTez29fUxSjOT4fS1BvRv6Lkydd5k2rXHLP
CFBnvMAoK4QYn0jfGtvCDsz/+boc7n07qa6sqQt2qpv3QxJBIzkLpHkh9pcNIjDgKIDUat3orHwQ
SKKTVLhNH/V5Uufam+rXLolw6luyw514zIX2ojSpleHZN6p7XUH/Pqt1K+CD9DwjWB10HjPm+MMm
45JgIAxNeowTbAe9YfhdzxCstfNd+ehGUzxoadODHr7KxE74XH7E2NrzII7uHcO9AFsCM+2cjEcH
4W6MY61Z6lqzCSfKf6n3bU6Mr0Sx4si7/gwsw2JAGwKjWENAPvB6cOtse+PqoVVFoD0fFz2Oo+JZ
/jM/Am2u/+9CnTdUuV+yQCg1Y91XUX8wvdOdu2CiybARLRZp27OuxIcWDgi2dUerqStkq8cKuh+O
I+VfZbT3vt01evHeQo4RQK/CX6N4Pqpdq+Kef0VmVAckmLO0Ff/bwZhEbWx9e5glxtMegnesdpRx
iq6eATW9/aFuYCd0f0JIwA1Nb7ZcWlVgymocTXRHZ8Htwc53ReSA73Q4U76ORRPK/BRWhaCCev2G
RQDBR+35rMrbY3Mvnn2BBOo80JLkBSFpmAGA/6aeoj06UxRB+ZLA2CJwbYxfLyFo7pGI3G9HCR9V
R2OO1asUlDX6VeiNp5N4sU/3zucesYYogzYOqcIjkbgwncrXorpYNXJIXXOQtm7B7t2c7d6X7Rm5
1G7ZBI9KBmJhy4GH9L4KOS7a//L95siXqN7MVvQTVP0UOYYZ0MRhGDrvHPsssR+5bkLKtyB9OdpT
NP1Y7W+qyyO0LQdEGtxehT+IXaNnh/JfsObbKcNxGDoYF5sZbfGAyKgPCPUMw/WcBW8s/4z4Z87B
mNAV/i1hMvPGHx3Jvh6c9jhf6oJA1AQh3OwxMP0qQwz2Ghk+h0yl3iFZGReiwv4MtgY/aW/gDu1W
ArNJnQwKW/2qaxEds7FsPJpJ10BwCb/KTTdv6ajUlDSycgeQFj4mNkmVneRvaKyEa9WfdyKp6r0p
G57gH440v4sVYTnFx5l0lryNhnd295DUIDWvBriqQd4P1FnAIm1HMcZT79HtsNwU2/ZzvbVq+B2Q
wCAaRxk5dV8FloCz9oFoi571JP8JsdCfRxqWayTbPi4kuPOjaNt0N2fnO5ZVKz6qG3ijRpCGSBVb
5YC5elIc5ANl8hqLzGBWBUn1jAOZni/YqBGS6sBRti0Ljfle8xlUkaVTVemqsw8SMzh4fVpo4bIX
DUrbNsGKuX42+Y/wRDdOHpPkxAYxRrym5O+pP6Wxki35GV3FR4rEA2+owC0jDxnNvIvSZk1KzeaT
hhaTgJoPTMR6NC/9KcqCCm6yugbeZv9Ua54u6Is1KNURaOUg3q/t/Ff/DtppDYQlbLB54IN0qCFL
CKbO+TwrAYtUzMjfxvX4e8+IRC24FSDQsG9fErf3V0kuZLNYHuF3acLpGjoxZ6Forgx9WrVhZm0m
KFZazX5Y56jlmnxd8SsFmk4B3yHjyHISx9+/ubAvLmObs3X6w+iAlcivVO7tBQ+ie0duRWse1Yny
zS7As+YTfb1yZMkioxfa3z4pZrb7K+Tq9MpdHmD4V2wKu6Orn3esNGFMmrhXW/V9RedFu14Lrpw6
V7g0FG5zCGhNuvYKnS4R/h8OXzXcjYZRcDs5HeCLNg0wMFdj/HORh3ibvJFqa8bgRqpmDeTXou2L
/A4M6wW8UM9AXh5737068OSIB9UyhR/WBSWbnbSlQ2S688eerjaiI8DjRrmockT5nG2rUqEkISfT
d0kGSSlss6pWz4BbrYGrSAWbgTJ/wUh/oXXfPRslruqDxxrXnPxrM7MLVmhxhdmWyXH7rw8FVtFh
1CNzRQpJoUiiGJ2EyduZ2JSqdVEahfFUqIvcjUEle7sEYjokh5PAwQYE4xArVDFGLp4Uo9lhWNYR
/amcQYVZT+PxQnUnfXn3NR4QI5bsidrl8/ihwfz1Ph/G5tKO8vcHaHOjXF5gnoHamulqbSGcLE1Y
rUf9+R6ceRh+uGGKW89UCRwd/JrnSmVh/TO5GLgiJZK1txARAV7xk68uh1cZh+b56LWt11qjVVXE
/vpkbcrvcFkPBO/WzrCGT1WndajSr633aPVVFLiyo0dBMixiwSO9RmUYz1kp1S5C8ryjX1cnmX0H
Heoc81rlOCd/VGoV4eNy+arp2aOljhkMFe0JdvnDz3g2DLeO7gvKOCpfuqq7EDBWrj6qYQ2cZo4E
DEZ8HkcSloMCYAAxjlUosOwMg6wOgYwKGsXbVtofu9e22EUl+XsvdP7xszk++3N0mixbLvrlShMZ
nH0PR+BUw2AthqBMBHyaC8J6mofxwu2wc5+6h/2RwTYLuAdjKDUPOqesZbARJj9A0AhglXgi6wdG
4dcQhy4AqpRnIVBY6iV42qFPGSKbhmaCemii3HZzJT+BiS7BY2iqyGcMoSNITZJ/gwYIAUUYC6Jb
kUew1gx6sLpn5lMA+gUa1iUSrfpiRc9+XaOm9tFbkL6iMNWJyLsDIiAmJSqG1RLF5H04K3ESYeTT
kVwsDtoBIk2nYlcohbpG6GOGkZBrIgCQE4deoeUsZsejLqyLBd+odBr++nusYHozJtjv4YGxs/X5
V4R1b40SWMr2tZHLjeJBZIfyZqwxzkZ+3odFEwRYp+xXEgwA42DtFcNULxJhdja+PjskKTYG27eP
Y5tW+9Int3mOiGHhKYk8cBVseMN2X6VxZ4iBN5lvVbDtg9mfykxPVcgZCMUyyrhgY5BxkcCC5wxy
DuhGkhbNrCuaB7ADBK/LsdY2lWdHs012Sul/lfw2mLd0MPVsTkEABDBQmOdbjR1FebkH8/83xJTI
dm3TO3XwoNBQu032v7A5h0tmLd6BdoZ06VHxuF4nUzw/5pexn4hP+4h2wNkIRBDqwAqALbqJRtYj
ot9Ae1pkLmH9/CODoNT20ixJC/mtdguXG/cu3xl107VqFUI/BJYC2uPosLDo+gNiQmzG+O5z8NHS
Pw25BWX6D6UzJgRsElLqeQmeNoB/KpQPe5/3vLvinOKLDGrl3NWmboxRUvYSkqP1G9+Z7v05q4SJ
oRjaf2Xw5BSeImQvHYiUw+y+O2CdoJfgMt1bic0OeevaXLy2GBhLg5EFNu9rYMUcOZ73O8Iie+zd
/FT7PjR2IIGYocSWwxlUvaPDJ83IJEMqllQp4rpuphjj8MlJEVRhRz3x+cn1vpplemdm1cKR/3kV
E1Qvww+N3oGN9WbHDcvEdpykLmgaJRhZeTp3Z5ee5kISdA2p+MNb0HRx48i7Tr1Rl0a9evOjOCBo
6UELEf5RjJLJnRaPR0zXFST9O1F+u8VY4y1Ntk67QExxbRSeCzH3/PqbrU0dRvD0Y0QHH5JSNC7n
/Hwl3YMsSdkEoBlnmc5yPts3tqKWse+BvcBu7xJrS2LmZHoE/idH6WA2WqsDvTPyVA+f+B+flDvk
21hFMGFYKv8mPVF6jWBf7mBKLWXPaTwToIrVMU53lF5+7Y0WdNGr9wnhA5V0VZ/fQxAKsFrxNuCM
8iknsW0ItDQtAjVBFYyG+AD1uYmk6LvZMJr2prvDUm50Fg9MuYZo3FS+qXOryrmB0hRayI8yvp1C
0V2R9Y/bPRY8wVtwa3n2qElLFAos7vxogqVnxT7LvLF61pbJ3Qq1pn5jJb31UVPknh5wh1MSKK9L
3d8A4x/XQ28jtezNxH+jU9+ZFmFHtS4R4j8v6acY08VVFDKqFuDfBHcdYSfIrhlMMMIjSvs/WZl5
4uGRBV0RBXg2sjnP4WbsUIJmadMXoCBPz9U4Pka66cq6X2LnMVjSSF+rJKgOv2uP84Kij3r/wafe
AamP6/U+RwA6d+S7fzuDK8nn0E/rjaiqv//mgYfW/KBzP1mdZ1qlvUPKCXv6A9af1fkAyv5kcjaI
YjOCq5lhfwpqTk05vpsrvAn72Vc7fNUOH8AD977GNa81HCx9xxnBWdg1dbcre910rwiUKPB47yYM
LE11fU6dFwjnrxRtrTUSMbx/s/3Wyhtkb/bfWDeDgbxF8623aluGY6ER87mXLDIk2k2hfJ8sZWS9
uRvYZrI1AjdMnUO5tEd/Ar3HwsLLEH8NjFY3VAWmb+TArYdGjOjq487R6c4yDgdg/slfh5IN4i5U
Qhv2YhPC0Ja8mon2uNRwsD1LJEbBN9QcJ4xzKVzsyY7UzlXNHa4mzzCZuNmxYwJMddUKtZULXWtH
vxEuTZev3Fd0GFe13wMQr/0F8mP3S+YEbukSS4Ryg1AezCuiKFUW8G93vNqNevCdo/e4tUUPp0mk
KWd+qAOUT6/Rgzhf4lDbmXd2XCntDdboGj1wTMwDhjL9EhGw3sRpnbrWZJ6r3Jo9poGdIGhPZLXu
hfC5Rff+wGZ2EMM5GqABFh4ODbuP/L+inr+Ky9rT7rJhr68areJB1BK1BEiYEJIZ9qXUcgeaIAZY
QTd0yLdjJWZEjnqZ53Dntb3YpXAaGPPIZnY2GMacQyD9jEICzah+eKj6wy7KQKkFYBzubnBzl6tV
uF7oTA8mG6k+FnKoF1V+madB9ajCNcXzKN3qMZsakLKlr/ly/VIrafdnU8kW2T7dum2Ev9MhcqmO
2MsEx+0JxS/y0fgu8nWuh5Kqb1PzW37hgQ2N9fBhrvEBPujSO/6qt2tCclF3BF/2MJ5LFHcCxXql
LsHak/tZsU0JxyD57MKIeyBI9aNXne6kspfFh59ijEyo1OdVSkQvSVloDhJw9jS2AdjyZMN+6tsE
jC0WJMYmrPy0gVmxalNTz7Bwlz/OdLgTQ0n1VkMFbJ2lQ1+mpNhmQdrXmglC/YNfkJ8iDyUNPvXw
ezWaaRZfqB559pma5ZnGuOpwWJqx2iHcNo5vJdhVQ81fdpKx8GtjOx3DxX2vQXEZfz67FZd0VNnO
lFYGWHbg2Y4CiOtn3IxyWddlA7zUY3Qhh6Eh28cbIseFJIiFlTr0+EVVYIvbEYSfvVTlxQAPLSxx
TMjpjNR1RGl1LOHyA2eyhSJ1HlYT8bRBsm1N96YMiwwe9MwLMlXpJ/s3ZWiKutRz/dUVrG1H3/ye
QG8C/sLlkm3k8IxzQrYkaw/GObSnus4qInEZSjNMMtbmcX2BCpaWEdcc7HguR2DoNKfW0MkNQnMI
W/3LQE1l7DQdsDPICs6bq+D3xCV3Dh57h9i/nogo5z+Wa3vXXsuuZRJinVBhLgLcXb/+vClcYgUE
fkunymDbHCbg0B8qfdq1YjbL+rfMrU9r3zpb6q9c69ddJEangRIH9gl5EwwPeFI1OCjYYhrPQMR7
y2uhfhoXzeF6ZA1u3zac7buII4ZtPEIn3mregxPEyYLL+qEJl9LNzJJcQndH2z1iymT2dK4cx/5A
DpgeLHuF5zzWlm6W51ABQqg5zdU5JLUlmGfOtg94nxBypBf2ydWWIYfWtdL9wLNbmb8Pmo7A9xzu
Zayor/Yiq9uGvXKl7kh4l1jTITaxg8xC7KESQ2N4gtJwLqEVILx3Bxx5lAhh2p/e2atqj19RsLK5
w7nyjOrNSipQ1g6rijA9TZONVajN46DCTLQZsSSJ/nwzPZaz8KPxhBmGJGINPA6OkHYll8rucpRL
eAEEOrQW5wIF0naYVqCHJl5gUGgB9pkFZmG0Vse5m3Ip9TUfoXw6ZnnnGl3IJLBVHJFRZoKl23LJ
GLLijNTwNCq43HIwR6Bw4lo82zY1tiTXpcSYIz7KfRG196vyjSwZDWT4SRmFTm8dfy6P4eispfkh
dPxWirCgrAY++iMHKoAdTtkRuDPITBH+4S10c5ZKdcF/GsVi75lv0P/j+EOw8fT8URcDJ2oy+aNy
GuL3vHdRbLw+F+UvFeJW/0L3aHuYvKLrMrQIMa4ziLERARjS1R3L1bHXRNfmUMVcYY1hhp8DLiGh
MYV/vsV9SFdtlTAal/F2P69UifArOpJMGiy3YAG7a8kGJGA2Xh932lnPmN/9JCubdy+RWvtxKEdy
oPGSnxMo0gdzaZgdK2YlARhJjoclV3XTrwzFgdmVzplanwwjX6l3tq1COBpnXcQiPvzNtfubaQMD
qc3VURUUvm97Sn38bqxDQ2yaEHoeGwcenrjM6oM0wHPslE6HpU4h82in5aF/PhFW4rXgzRIg7Yn2
pDG1+azWXOPcGxpUIeilJux+3r5NJuY59LpAB8RbvieU1cQ7hUYSPZqnM4VcOsAlL5SfNNLpKCvi
QlX7+nbv6eeZQd/OXKagIg4m09yy8DAsNg0TbqYKM6ujRxxstPJ/kR6ui+FWho5PIlOhlIvaIdaq
xR/S37PUiTt7yMWP61N6GGMtjpPJmi3OUibHrHJt7dob1rzBApOSzOk2ltIhiYABr4nl/yMHwxuY
z42X4c+gCY92Aqc+GfTTlJQLIKZ8qRo5V3yO/JRQ9+tpZQeH1TeedsKhffypcHqtzsvqsm+PWBe0
YPrfNpEhuB9zzk93jEat9YC7DNYFwT0/A4b1HLszqmKyGG/OksHxHaa24TxFOhBjI7gKAo3mpJJw
LC/uTZo+C3hFksBXL1py48rLTLErQfpPUSe8/QakXBG/K80hbUFK8gjEhLEEiRYo0A3yYQi3r78q
wezlOt6YB26NSKpgdXVXhIetpNkw0VSruF7ZLOhNEmmdU0jSwme/MSTPYC68nE1840UsXHJU8Yo2
+Xcn5FmowAoAhM8YnM2FsaannePN5hHdamM+o5s7JAOB6/nqCFwGLSBfLF70kQnNWkQ4oXHWYtSZ
zVQa3dqk7Gq+t9QBN9EreYGW0ccJatPQAlygen9LWOg11ofJKsjsjw35ed2RJYLDQJsFu0LMz0qM
FgOhQXpyX9bSOU2dGIMxr0WQUmeee1BSsHmvwQZGsrnr5TToK8qRLKuPSMKMv02pvLgRV+GV4cmX
oRedU7TjypbK9dCnmdV9heVjMGZ2Q3PbToAJEqCs70gqgIet7l9VC3NcM0vSs903ddxON9xgk79v
bCAJ17yYaH+7GY63UBOSbA7CcFo7arhZeIwvE3pf8iX25op/h6sYl41ZeSxAdgFtrQ6C/2HuKH1b
i1PIAV4jAoWNhIdSG0LC2TV2+gVPfo/LbimQFRGvXZEILW1sN232JgjMVSt8zh1GSvrwuxjHzLfk
5F0RVi2zQSwiYlp7WI5uTzyNPvxQdrOB0uqsBEKsg3LdClOn5brRMvV3pxnpgPl10NGTrHSqeb9l
h/Oa4C6XwbEj/xCsVLShQFjcOQL3khViFbd7RpFWlmuTmR6ZvEOm6pErk5dvHNvJgXAm+u/8fi71
aw7dxU8PFzgP33/nzV8KWmowp/NL/ct++IG+O4QbHSf51s8OZJE2Cfn8V+iIdBZDX04CmWU7Ej4E
lfCICyb+N1fhe/sgzn9VIywGr18jr5aFEFNuHOCL4TVJml0sgvQgNi8oJLPrluVqvIVQgNoGsEgF
R1jnm8HtqImD9Y6db/tf7qyqpg2R/Su0+Djfsv1Z4QUsS9Vwbf8spid3a4Ez5T21CaGGdPoGAedi
K4qnH/kaO3t1VvGE1W7qyde3Qd1JFUIvQHKOZebk9JEL71enqHMYgpXANHcwv/5N1gpSop7g1Eu1
H12+mfDVF6deCGqWNTa7NbDjt68UKR/qkysLX3EK7xoUm+ZNmwVCJUjc2WOJr1h4Cp+Z26eo8Lwu
UaWydXtOTfNB07OTB+fNsc21e12xu/vOGyiu3tX4ysINoDYu6lMd1lwrnBQUnVbJUO2JpXGnvxQN
/1I4sC9Bnjpwu/VQeBWwTwUh2zXl94mpXe6pDKE/7RqQE76vLLe+uxDy9YpkdX7vd4PjvbsWjd0G
OOcdxhGH/b2JO9JQ6Y6nwMH7TbyTVNU6dpI7tDnFn4vOfMKkfMP9NP+kukoHAwtQBYJes1p3ZNcO
ywSSvAA2xZurTC06vPzoXemijMsvc+oDMqKeeUZJH4LmPQset+otJb07NYetO2Tl6ShfmPHq+4/9
5J3Gtxo6jBfanTU86xzEN8fHv315qFr8Iq8Ssobgoq7c877USX5T29ia2BpbGCyTnbaaODbH2Z2w
CTV5qwOhOGzE3YeZbyujVrLEI2HPEqIkFGGYVOkqrlpjBiMj+Mzm/E0RjjeVX2ydRmsUgIEa52rd
8gDW1TWyCw1DGr7+WbzNvLaC2+x4nCW/Rq89bSyKhSjEx9n5YMcFxserdxYAUP+XxH2VCRoxfu8p
dR2uBOLpPA+0R07BAVGORdBUtD6/0BX3MSyhNWmaEYJGdx2iljznekL1qXg43uIwOQ6a0KyhOy9R
RgWiWlIaXCwKmzAAbTY7pIook4i6n4MAhzctOelGQd0RUH7lC8vefSe5KEbpVvvnPOf0ZJphVtG1
cbfbzbT1gw5379RvW3Cb8UnR+O1+u0/hCfK/8wYl7hRqiIL13RGRJ2SqZxDG7pZzlV1TYFB639cs
1teDTPKCW7rL+U8YZdqf8v9zm6/pxIAhJjSo7K69+yEo5fbAWLjNraqmJYL4qA9VG3H4gkMahVTz
PwGZf5ZBvEE0VwDs5kVuZXxOzbMHBsLEBswaE6yHQ7S+YGqjX1sdADkGPZ69kTLNk8gNrkFzc5RV
KItFvMK6ZG7q03kNFWFucgQwJeWaxHWYrxu3RHwl7deA2cOYVPOmchjDK8o52lSaicaWsuUw0o22
OcSvlk0cwFA3ShdOK1ZoXIGSmowaY5fhreTrDOWEoWb8CI+CpRhbEyGzFHxG8RW8a6ptV64OJxht
NlrIzVxKEyLw8KHqEH7qH3ANvpg8OYhrOHCmzp3/KZfmQRd9W5fipbrdwndygS78xy0Eyp3qzHl9
sN1MSxURhDLRSk0v24fS4y2rULez950p0ticiHERwUnawzTBX63IG3ysrv+nGlKFOtf7BOVMVlzh
A51sT91y9qJCFARf+aljXhBWFr/GHMTfmnEGNfWCG1mMmRV2QTv2qPHa5Xuce/skGoD4GAEn6Mhg
dxXqqz8st+SnAdJCADMmJVtPj4TJS+2Cpy4nhpQXhYUdhkr2XngafVy+EapA/n0xMRO3SoLfP92T
pV4sw1HDhRez4QyP8dVmU6d3pPeiAl0/WWZDxXcQKUgIXHwMnYmmdm6+e9uFmHZymgixM99BItwb
OCrYqnpSxvi6hdIJNj2Z3CdiZvgqYBNC3nDshXz06cn6Pkwm+BN4KBDWPIZt5xMd9jvH54aQUICh
3FECj11uKEj5aYLQ0MkTlJ9CA/dlQykp2FOUIBs+xNEXqo+oB4szFjUCzNfP440QEdoaFOnh6g/8
Lk6QI9q/jSiBOyGqjf25ncCZJaR+bZRGUoVFjaKj9NvCRwtPKCzFpFTWwaVUbbyBHxC0IYNXyxST
Q2VrDx3Meidq6EqitE5sEtCuBZVamE4DToJCvSD07aKD1hb341c39X3r9Mcde1ZIGoL5Cr7Q5d3Y
0AImG4XJsuGhGzsPPIxzr88U5/I+TSxmGhEqawoil2J9bNhKl8QXMtmAo6NuD/zklbnkgRrJN/6r
bEqKGtN4c7s14iXQqDBSMmk96GMzZj1RYMPvL774doHqsOwZJSU3/wJL0/EmYNO6D7iFBSVTYTii
CzKcFgpQf1Y44ZHuOMU6y2ZKy3oOiValnBaj+UHzIP4leAEJ8fP0wzwK2IDGEGqCY2249uUXNW95
MSr2e0mBZVutIYoqZ/o16R3feSxPaqLVLochjsgO7c9k2Lu/BVYOIeljBHX+Xl89U7kMYlUnZHsY
2Ww2I18Vr8MnOhM6LipHjCQyN+7i2G7tpd/JvoNGm0l7SEXFlkctIlCXGkm2AspvT3md1q2eP5VU
/1TZkKm3Pyx/AfyA/J9ZyinvXk4Ct1HJ/R9b4wnElevbVqK0lNl853fSaEe/jHB/g1iCPsB8bW5Y
ocKaefkXN7RdT0LXZDpJ9jk0ImEVxb+FaTAFts8ssujiQxjYN89W8GzRDTjdgye0vpc8jpRCriU2
DcobU4KTf0i63W8wh80uQlRSlvOv81SHlFW/hh5fw60XAwfQmCNukIeObqEdZHKwQjdbd28V3BJt
865hfXgPkdJ3paz3m3MHurqb5ff69GKuLp7HTMMa1TVy3YBrp4NRVJ5diCqPlbZEw41243Aqdguw
fckt1ZYvp5l9USaTzoPrdN09AoUQb/tkm+ovlhWn6N3McKgrPxWtoetOACKZynoi5NWmp+2gnR5+
LlX0Pb6xMkiiMu4JzQOHlTaV9SOahAJEg/AHiJBWVDX5949HX+JEpo0qvbsuTKj0M2uhJCby3jz/
AbLfI3H4sO940XjtBZh0RusoMSa+mkAhYiZFK55yy1RbsT9KU2/fbEG3p4QR7Wan74VzjcwqeBCb
h+TadaSAsIJDFNfwoih0j4oY6shZ1ye1pcC7Sbe2DShMrX3N40mmEyYPHGxYCRKXUVaLsdRCCB/g
YZoCCBLWLW8a2hdR9vAFcpkc4/KW3U3+MpAvpR7+E02soDLlnSXY000eONy+K9St89igKxIQUgkn
lswbPGWDaD4hrtjKrFhsljRXHwjhE4e9SNnjaY2O2o69pyF6IloH+ilPuELLG20bP6a1hhM4Ff/a
ECz6SHuI/AAkU4C+QakcJpVwndfs/RKUvJEkxTllFzqAcj5qlzc/uNI/XLOXNKc6GhQ3y1zdL8Rn
hoZOCYRzbnyy51B7Idc8/FmI+kefHo4H+nS1Rgj7Ftnsz4tUSCpZVObU4tEBhsAXcZ9AluVfIFWW
2nwwd5DLFcpNrYNhUSVzFLyql0K471z3vPELx+qR8gHX7MUcJonOqdUl++PUXfFaLZtZEZmUEwnV
mBOXJjVdifrUucxn77fcBgEYSE77U3IRCPitltxC5bZ554ZRAVy/zkYN/WDthztCrj41kT9q3U/Y
hh1IX9pQTAzDg4J8uOcIlvNJz7yBFudgPEJ5G6o3nV/SyIIJY+4Lbbj84y4b2m9rDSegypFX07+t
A8AuPMf/XtBJU7+KNpqCBv8O6UUuBh1t3NEia1avaxsU5tWXWc+jvDMDpc7IYyCOGpdcaJT4AGt2
iBGDhi6mA/HGH+N1ZFxqyvin8TzB5lwEmzACb+2fppTE8/8ZpANMY4R+VMj4/Fc2VOAD2O4aBDUB
/aE3zQOxrfEwTsw7gqLn1LUZ505ASLkQ4LDSrD+U10h0i+QkhSJYyfnnv+Dk/uGwpEyqNvNidb+r
8hr7zZ2U9k5YyiLm42InevhoI12RQ7zDpTMcYWmFyKQNfeH6yYkVS8l8xnjRFRyqkEBV6Yud4PtS
+nfN5hCnJK7YQqaiBkuZv1dpuC5j7mz2sHRBIhZmn4z0sumjAiSyATrzwGgCu9h1bQ9y51F0YgtI
neu+9QuKSvTEH2gnuuXC8b2tsmr4q4tiejyhLe1qStN9xCftlge+RVWKJycAvQfwALtWjyJqyhmz
+ttVTt3+7sajyxbHV/8fUgySQU4agEOIg8kIK5ERcLF5Ogj0J3SxldzcqbeNLs4dAZuzyTXkp61/
pq13PAfYWueKf3tnp+aTaHNCZOLhDh6cM7d/LR0nLMlJYC7T6kPdSLm+cghlca8DjFUtLWgrVChw
DHcIxlxNM1u3R9yjvx/xUn2OpBrj0FoUEi1cPdKVl/8ETuN0KwXVWHevsSqq69brQC/K9ydEcjn3
s/U3EWAqGUQIAMt2K/aZkad8pHRX82S6rXq2yKRkVHm8EvJk/R7E/kTfQqDk71UkPGeeTLkViDao
itKNESKR2YBzOfkdDwR61hLwAeZBze0SXSMKN4+roktDsN+zT+5thW5hBDkGqRbRlXbeJIi14RiJ
OjKhYjv7rSrzUFQyJVOkXeHhntwZSiB0+ZhUrFCOI9zKQbzPD1cxoAFIA3iy8Bbh8xVHiHCXvS9N
XGqJjxAIRKbThB2kUy09u7KdzSXNnXb5V9NaoC1OtbUPZuaBok58N+Z3/aIZlSa9oPtAJvB0/ig8
SVXxqj1IRdngwH2VUIYQtmER+QWO+jIpwg3FISWfDzdcLv/GO05iLWj224tbS/WdtQtp/kfa+Ah4
fmuMHYp4s6J76NrZhPrH+WM2e6Q2qAKgup0YuxJBkQ/WxYvPXDKlwPUAb21A6XcfaN6MR8Wzf8hO
DXtHLCwOAIlKCqMVpHfhy4uutu4JRCDbhumVaKrcbhgRZ+Ju93aRfxpJY/GN+s0vryFQVv1VOZ/g
3QOyxf0TRzf09TSjOhl+22Ug4K+irX7aXa72QDF9mT4dJRn8xm8WCp/524ggnGRMUUlMWqxO+p3d
QKFYv7la6pCIf50TzwTUFaoFm2tF2loQAkzA3wxIEcmg6BIlnA0pXF1rphMQjs5JHcmcXNi8gSqL
KC74cXobCUXmAQvvVXrS0PCoIDCbKgNjp4G0wREOMcrTN+4nP9FKEBKHbDt8m2ff6EH8xvFNSuLz
lsJoJdjaPBIRVfpw2X8y7sMFADPlz1fCsIPNONlZjfUKdEK2TgLgQ7OR1QBaMiaa1FYAGvd+whIz
C3l/CMNrK8wZ+Nla/wpXMfZHL5iLj0b/F9o81fnpm/9pPhKyQUygtplzo0LnH1qg17FIjE1K36ee
cchHbt1GrY2cRPUN24ftNMtT8b5Kwutps/nFkBFt6Bfj2aVgumyq0LmKeI1oQgrcn7PpWUBXZGh9
2IP31h0avCA6CaLFrxRY3l/LdA8tNkNtf85LOj86gC12stKgeSSLXSR8zwh5oAeRghCbKuAvAC1T
0bftZ3s5OjtPu3S1Ice5Z/A4adg38XTUSVH8YpyyvRsW/4wv/2edxru6Q8GhBAcJ3MX1BRNWe1ZR
pPIc0VxfCs9MzSIl8TDOBxwY4tzTobxbYc1DGAFLJt9bqKNaTv3fzZ9v36Q5WIBvjW1KEdp6Rq+Q
k1jKZwKN+OyQ1CQ48BONBaUw/AvIlgzcuPyZh3my5Y/3tM6wNh5iL1PlHq+CL42IlB+y3hymNl4B
idybW6oUCqZ7+937r4Bmx7Wj91GD0iLHSuPwro8cIBJvg3gkhgLEzruJELOUoiBoru6wjQE+Sgy0
zGn5ZFQU/MTSV0ja3uiVh8SI1Dmi1Q6ZciPM4AfNYYN9Ht/guTLmbJKJpkRV+5UeQKICJyPlunCR
Xq0o1F8hGSU0triyn18tQ1V+R39rmqeQOm3t1bLaMqr2moY8NFfJL9Y2UqtnorwfMeAT7B6snFnG
2cQTXoDTE1d5gqzShlW1OYfZmeFz3E0NTKttGMapKiXnxDioJEjDiy12ePXi5BpXTh290j7nuDeS
/dyknLOW3qAIjFj09IL5DtAqNEEPQ2HnArxR65TmtS7iYetukxrjozQ/pSn13SS1qr+TSPnAHMNM
LMKmZQbF2rOhfqyrzBma0hZniR49Q0WNt0Icr+/VfAVIAR0wmwcTmUidPxI8NdGM6ikwKWdmAuL4
civw2tY5erdqabp7q9o7IaEk4f7HH+C0RYsqFH0cco7d+jBHaFbcjWhfO4SDLGzH0YqEnM58tucD
AQpXidpB7aTm0cetJhySbjQmW7YGtqQAOAUYQ2bx7iHPsaxDBxjlOp66qMklkd88IcvkmHOdnLxn
af45q0P8VICoaHlAKnkhes4bJtPcJ41KSGr0F2RKzGtdX4sxjkdXh/1EIDJ7vNunsJhGN5b/QB7v
zbeZmmxRRk2eYjQOglFMihO8VkOTNvubCn0WUtUoEkQF825WkP/Ccv+nkM9kFl+2Cc7VhRPEtHJM
RvTdN8IrtxGJKRga6/OzeD+jdRB3PluFjp0G9X0CmW6Z5twEaHeIItJ2GDuKT/sUw7yFq2TvgIK1
h8ano4mmLhy2gkTbYkuV+9lLxp4px4yaQlyHC3qBs1phEPjI4DAxQU/3hLB8YEF7BfIBSjtTIzj6
KV0SVsVCVxxJtkpF/+f0n+Pv98X/RPjTwImVo+H28wIxxjJa//tau6oWgjhXQg+PQVQTIurUaB9f
2FhMPB8u7LhejFrEKc8YWp6V3tDOcYX7v0sLaMOjMurl8JXwvrprRabcVlyHMabOR5kvcXZz7AAU
AA+9XfaZ1KEWaO10QYtUfVFdaGCTK1cyN7Vzox652vFSKPPhejv9O+/eF5JzEr766T+7/uDyJBUd
U87EyWfy05b1+ICuxDstR3cRmCNC9qRq/CpqaLdH/oXU0TPPHHfAshjL/4UDnDswrG/mwOjXWNF1
fw3ni68gKtwoPLMSCi6NAs0RT4ts4n0PTuCz9l3jN+JglTBppOkZRHoyFJ8yhF0nI53DjKGlbOwx
qq7lOJZ1f97T3CfZTYdklG1K5wl5RxC4FnM73te3Nr9uO2q/cHfDzUqgyUcrCBC0BcvkTC4YcPPH
F+YhMSe99YHo47LxnYKMUlyg+pnp8sG+K9l9//Vuz5Ls4lOHAxXq+6Js8zzSIMZLOH9x3tVX271K
E8bsfLDL+oTKsnYHk5LKMuMD2UslQm2uoeIAV9OBYHVHlaUrGbsYmOYG5PZ6FsTpoNTOvVoRKLbA
meoK14XWqYdLs75+kcNlOJv/pk/4fGZZ22WNxQt7Z6CaMzs+tbfR585Nd5lYdYxwnxU82Kb4r5Mp
C0FgMYZIHMBfjWlAhKIG+nc0UtehggqvASgOxlmiRHWtOBscoQInOwuFVeolrTkvacoKMZLHgcJr
mfWBt3vTyFBQuCEWbWno1kfvJY3xf/fqDkFa2Qam0p+ByCo7EqaKe6AX7LHaN8mbj9uyeVJdB1L/
h4e/kUz2SFPUytQCqU8LLdtq/6doiDZiVefy7lLFfyZucju9wNkRdYMxT2+DuR4ea9PZHjrarGY4
B3KcmbINGMeRb6AiPuCWz/8D2niTyqQXr4jYloAdszbpwDbBN6YFww6SXffVpGvWNqsgj0MwlqR8
XxZcYf0TsfCwmnlZJmQiDVdOXgeS7STkUmvfRZgYgOKm1TKsAvLaQztJNjwTiLkoWqYhFjDKbGQA
j2fXs9ILfA4cijdW/Nt0s8p526iuYYeDmj19tVfQeyr6CgNyG22mfw70Hv+gR9FEUQy3C7g96z/2
nNj5AjwA/oK9nD4W+P1ZFd3dRYPRdZNcFpoCVIgfDdbSNH/dcdsaRpIA6M9nuUkTxt0hOCPAfI0v
GPrwLDOJJdLSMsTngO2G3Pfl4cEqUaXw+kGGSgtr6sOj1tZyqlIA8jZYxD2wQz71wFfIYP9vnbKL
BXuPABKVNRtXBXJhKoJYudVtW3FhLBcPPQ41nEx/MsYIsQY1P1NzQUewyr+yIU1Jn/SxSKzhgxxD
wixvKRrCQXpyZJ9CQZmJcO0ZXRqSnIuDjCMdyMmpigKB9yJaum1E1KbCRnZEuKHvwef325i5nlNr
6cxs3D9fuOpqW6F39G+DTgiaO1HgNQHQ9xKBnksE8XpdrnQlO1ay3N8L7ioWVvc2NZ3PO/G6VZ5V
sR+oanewpsvMWvt2F/rMyiv2xUdvRtq492rSO7iFNofTIE+tDuxxr+2qjzvwjMB4Oabd/NBlc064
LVlMKi1/NJq0lyBA4nd75GoZqa0j6hGFmfvf1vVaaC2NKPSg1pobQtsEmbiMrAvtvhLxepyFmJbv
yeyah3UUhlc7ZqSlr4PibiLIt5fi6MDvEQs2DzNVgkM0ZeyqRLEdGhRzfPBR8JlQBamshEe2GKgq
P7KTWS6oG5kP9PE7UIu4HDa5cIziqZMQhVUk9MSlNuxwzyw3CJS0f50LYG3PWtiBFid7yzo8pqwB
TMgLv97sB23+qrPqxfBkHLv8+mK1Ruy6BVist14CXvJcmHH/o1waeNMqq5Q1vA/lJdWxmKvaDquv
Ki7rbOmF8KwFdnuGCp03P2otQNiFTVkcGvFvuHBro8ucxvxqfzn33y9cgoWCaVx+SsIyaIgIKkyR
vq1y5vKPazwj4NHMippHdZffjY4o3fgJkeeH8IJgcbcvmHyCmyXdX7/LwSaAYC7QssU3Xy+Z4X+p
V7AINO9rXJDTeb7APgx7UdvSP+dtW3jZbZCpTQGezaMcURA2+NPn+SA59FcnCj51YEiSwopjyFb3
QFfrtnaTyryURcx1y1PopZ/7mKi225I44tKVjNo0F2LdwHsPWyUbMHV4i9LQL4zJUPMcer3yqq/e
Lf08l+XN0kW5k5X2hanCpNXWAJSlk49hUpPwP/oNdCn2kMeI0E/GdqLGGW9/brsv/K34GC37Z+tf
37vdi26s2u5NQOEpDQ0eFO2QV0nAsegPHdZJmL43KqYzYhFBKbBtQYcmPA1/RHfhd6b5uCdAapor
fwCrzSemyYGv5aGB5qKLItG/KH06vRfOG/cWtmDm8000MTCTYDrrCWGSmM7hjHAZ3nc9RzWJUq8z
4Ty2i3+iZollN/ka7AV36LcT+n8kBRS5vVC3I2dcHUafmM9qT3Sxm/TaqvMUTvJbJ9PlvTl/L+Yk
6fJUguYTowmpLR+a6hH/G8aM2KoWX0vLschyDg19llcPCjncDmzywlyEUcpINF+Me5wHyCRyb2QD
pZxpFGtWSdmm/qvz89OW2uFTR2WuQP4D+J89y1zfJ2a6gCMsz4PqoiNUolQs8xS+tI1XPQd/z6+5
68Vla7uUECPIyMpJ6cUizVN3LHgDcAOhxHtizCFELKj3IfimHiRGw+uvxpZHE03aFRo1ZI2qL6u7
SHdKOpb4kzXtTBIN3zwGOYq5AXUZFBndKR1n+L1Y1azds6OWh0gCMoA53hyHCjTw61v77IgshWbK
Nxe9UqtUblqWNEVxg2GXD5nl/JSraHjCdSSwU1WlIzzPhN8/vim/lni5dRj8GGQ0pQNsuW5Qoxno
kf6CYTmEqpBtFtI5dnF5ViAKbVMAPq5fyjan5f0Hh93gFm8l15JNIPOGoxu0Nl0xPLQCcoUrja5Z
it+XlrSrm/6QG73iqhRXGtSH5Mytd9Ya4uAzRpaW8NGY8m6e2BO9dCL7VLFZzNUYWJBjQfF4ifBL
f0/c4aeTPWae4nIYfhEpxRaGItG8DP+qxidzMVkqAyGwT8l1Ln69fTpHP+wynVi/tTgLDVM5ortz
gYgms0q/ETFD7Uq1fWK9Y/yn9kPrbWEOumA0Hbc9Bva2qPSMLBOQU+tzH+Et3zS4rOX2+t+322SQ
DI2H6Js9qPrhgGxhNrKnsKS7rzqy5lirnz+tSyQJAzZRduRqezFN+D+JBR3L9UVfBEU60bhR3mxp
dnvYNrE+Kv98NGA0aNcvVj0bNcSqQasUgowu5HR/zr++Mw8bINtnVL8sZq743K9ws2Y8xtDaRHQZ
wrD+6VebkQn0LB3IzyAIQHhCHCVMekRrELesYQwjTcDwZs3DFOp3OlScPv/eiIhxOPBWDrPh1uc6
N6HaM2TpsVeD4PBOHlAyug3yLdMzd1dPumiAZyPxqEBhH2JvX3bG1riG9i1ZkqAroDHfzcf3A9FO
0Fe8BOm3z7wXKlv/tEhOkex5nq+ubwqRAVOsmPwCejlBPiwqnBQzs4xiYFgSGhYqXGOEGMxtsWZB
BX9HnmsnpnMQLDSyyMElydlO6u0SWOu15kemMW+0FUdJrJOPp6z+yzZcfWR2cLcXbYuYLL+LLaN/
RE4+m1QKi9MS4QLtu6AcfkL9UGXE1nuntZ688FzZ92HQ02McfNHjraWlA45QR8ElOT95906ALO5f
CDAEuntXul5Ls/jD1VHmAA9GijBUcrDK8hR/6FTtqjFHARClPzgKOFyqkNXXWdHulCLP7DY1WqI8
vRn9PtHNc7OaVTYFOzHdgtFn2Wj+hBI1dYBD7AYqp441VYwf1du8c33C+ikUTiQXrdSntVBsf1Za
IC+0k+dnRAAqrkXgndgCCOWFLkFaflRFvZfrd8+fb4024ULbG7L/ro3/zLUAD84P7HohCtbejK/K
uw3mxP5kXbKWB3uXkD8W1pfAs/hYyQKzv4BUds7y2gaXeCSHYiTb0aXxUGU6WFPB0rKp0Vjf1WQE
W0r2fDXaTIipLktkZboPyt9JT6Jia7/lA/8KGsvce/+tjFbxZHPYvZ/6+TdKWjfw9o/VNMCltbQG
ERKRm6ej3tI8xeeCHlB8vZrPAAixemhkkOT7ujbNgfuXLTTEe+d62dv8jR3rtyI4GqPlRgHhedq+
enLiBysyR5kfyF3FY7cKbJHA6fMYIE2PR0Y2cj5e3M3n3O9gQXuoD1HXYQQS06fJg/3Myyehuyi+
5g818xTnDS0UprTnsIzKafqnA+/B5o6kf9HCeRPUREjDsQG4NmltHSb2x50w73uNKiqvyrvmI1K4
sjM5KKJuoM8vr17VGEmy+Rv4awC4e7kNb9cJmN4rpDzQmjP8oBvag85XxUUnsZL4PWoWOd9uFabc
B4OM0YWHZ2vBGGv00KcyjvnOvu2duOTdnBNiZ1g+afejQC7qpx6J3Dw7VwFTXE6SVDmmAtjn38pA
dE193mTFGCenGPxiFYkhPt+MbB5ZqlMrls4aFYuJGRjTCpQoZqpzQux4UGsZYA8xICYMHTOLEQmo
7vTuCjjQ53yBbTDiWL//WzNd38FGVua7iOaPyIQXVTvW2IPWRckg+d3vPYMjEwY6EX2rSej6Zzaw
LeDRTech5MwZ8l6DO/WMdXzd2yWg5DPZDElIAYEYFSuQ+R4MkR1Kn78j+4wbTI8kNwiLsv9jy7qf
czmK8XVlQDxM/s+fwnDWI0w2QRcJul5WDXLf1WGAjFHrU45IlVAlzg10znWG8oV68sNtdLFXcDM7
KzrswbHlUVOLeFC3tjmMwQr7TFgVaP1uz70u2auHyx9Uc5tllDlaZjYlpR7oZTcYZMoOeOhLzXO4
wXNjm8crHxY4OooVITFDXEvhEuQ1yJVOJ8v5qr5IJFPkZz7LkyDZh6fRUamT8mkzTXwkCMZUtzjz
HJroWmvLd1A5hOjXJ89h3kSpXG19ztqw0gm1uTv1fAbtU6rENy5rUcW1MzefPiUn/wblrEZwbBCl
1g6DebnCKYjcV3Q3masaoA/NVVbc5SE0VTCEO+1spbKbEAdZN1kD3vew1kNxBg0qIsifBVFeG8x4
0ldRfPyMmCqubHd05UIe3vIMb6eynH79YjGPIflbo7TznCGZXXwTlMyeQ/mH+vMZKsjZqCYQZ5ce
/JheRFlZ1VrhaarTVhnLvJbJrd55EVB8of3iO6Ilt4pcsM5vZNlJlswgjidnGQ0hSep2MS2hackl
ulW541Iip60yLGahTxmnSLIIzh2Z8DQAN8yA64XkJPNmTPjbngYroigBrMZSV9Xx/Wy6X6ahlfr8
Go1UGqbFVe1FRviKO87gxBMzToQOUPtKVVGLO+3lJkR+H7k4Rn7NCwYorU1bsZDV6zvxeNdfQ14J
ArtlDvMpeFuZB0fVDpq8HS9yGBa4L9/wgtsEubGQ7lmlAjJMoC64cGS57iUUAYigo5McTBl02boB
4SA39q1Hld1xqzUCaAHBu3fQs3jNmpHkairV+kUcZmD+mfLqRCF1Qk9LTjmDawqQ+acnYQ9Gtqci
vDYH7XxkHhHa6173r4+XK6/Nux5SJPcorjfkm7IBy2NT2FMc4Po8f4JutXAhNdQ27UbjQMVjz3cJ
qyJr+dhYxzj/yYMiXmKAtJhOk0vlMQ5bZsmd0Y6CEdJfStkVrKhuEfak8Hw+mYNyJRVBoHheWFLC
4jp4VQDv3wpix0Ayy9PsljblENFHvuJRK3MXUUG16DCT8E05K7A+XFJLJKHe+io+yemXtXt94JUR
JVDe3YoWxv9aDMbbDoPmUXfsZvH5caOm2TTQnrTIw8yye4/vxscaRB0afWlLTtkojMoUQRFbRdo8
bSAF1PDC5PeWbxCi1vCc2k4s7w0ePiPTWWOthn84N429hbOm6TTr7FJgcGS89kLUHjpJp14Ke/Ll
U2ZqZzrOBwgZwpBYtC3lGXZ2zzpgWleK06jSr+fVeOiOiAFAPc0vKbOXawwIB3To7QFvPgEDZJSL
H2os39Ri4ObgScmSwqW5HOm8c1uL0NnstTqPxyvpo/pr4NJse3Q3aYQujVyIRnz41Q2RlJEq3YNN
/Y2Pt4ZtpqkzH5SPkW+/azKHwrIw1zukk504nNH8uiy6ovdEjKvqZqkCVzZisp7I3oVbZO1mJeb9
xXiPioSkPm+p4HC/75KDKCOL6xHjxN0IMi1KLb2bzLcKezq8ITrgJX1pcXVEpxKSbabCd+vOtG+w
CctrxpIbHXb1K7b5ZUE8N4Xw2n/fcgm3Rwg8jk+UTMb5NNTiRipe+dYzCTueHjSsu+sUL1UpJ3VG
fL+pYi54V50leu1gezUQ43ilEvOCSS22P26FWPhjKHO6LVgXXVAugGY8MX9qt4jR6aRnaiHB1tcd
tlHG+HzrKEVd+by30pQ0XcwV1Or+fzSmAEVVQo01GvhuB6Bf7nNVU/9FFlwMjVfeG0YT5bP6OzTo
VOAx8zwJbFEwp3HwNWS+ahfuWaR7yIP3GD7c2v5TIW2YrB/vzzNoiB1YJca74nzh5SosiN999K1W
91DgPdhCKVmAp0S1TZ1LEBX7rkOt3KXu/vhK4ZT7krPesb6nYUuFzpjRdg7YPoXt4yaDtQW0b7M5
s/dh/X3bVSeOR6KxIy0eVZFyDLhtqV/7Mqu4bTRHBVcFzL4SNP4+rPkckAJ1b/w3XdDmLbxgeFey
FedzKurhbCx9QMsizU9M1bXxdvwqGukSowmK15k+jFC6dMbW+XiExwfpXynO+NFvJMENJxzlLomB
zQM2cI+cXHyfGuvM2SjFObW9CTBxQnVUiP6RmaM7S+Btvgc4lczhBRzr/sI9CYUlwsnE9JXS5Efk
a7j9rvJAzNittsqd+GW7QGyoubiwPSqh4iJtYgynDNVto9piVExBWS1fmbbq6nj2ZWoo5GiH98wP
MLbv/jckF57XXP3AMDifQ4IWH9SFRaR8+MENikMUkfpQkf8nPag2HDbh+57ON7PmFnI/MG7pDjdZ
4iBcptK54pqmtRbsFGG9vM2gvKq0NKsXHk26WvpV5lcAchGQk2I86m8siSXnH1/kJ29jEgZ+JOyo
FZ2OUuEKfiipDCoJqkC9v9Nf4SSJteJrsFaYAasf8KKmTpbH1VzO6BzkbCkrGgnyOysXppzUinH8
jakVO8HmW/DDUAWirVSDgwswA2nsG/J3LdGou4KO98rZDPa/kVXvavB+qPf9YPyqKSQRKmNff+4c
CEStRBhkwwdmK9ElkkqFTyBYVD0N4rJ8iE1hmXfKXiake149wYZXfre8lisUPWFlDxWKprQpGUdS
mvtgm0BxJxQxGLs43vVDzZ82jjHuJdloybfkqVyjNZFbvDWpRprKmNg+zIOMrIF9iiuxPixwq+NK
sIfnY3ABtdZJoY9LhvZbAUocpBKbRSk4mJixX28eBexuyl6VIkNsc3KtoyWKy3Sk+WOpnPLQPjyu
eBsOVoScrTUKnDxi7TvnoYLb4oYz3IY3dfxiyEIVQB61HF6byTIhuva2mvw7FGwG+RpBblrkShe2
ey1r0YnDenZJWsVOXvRihlU8/z6YsvZur/vB05x4CBVhLKM5Z2BLRFc14fGjjcCcHPPOgyV/Iu85
qHpS56S2XAMJGfQPMxxg1UbofLIsenzz2lyyH2z7U1M2xLX8QTJTEGQ3gSdGnS+cP1jnqYll+24J
yyIAss+YRGP5WAURzStfqMFw5wfRK7KentyZFIV+4BerkRapXc5t5v0iBNaDkRhDK84mgbbKJn58
o2cwMSvoJkSwQlnBmUzGwY9Rlw0bkXwb8FDhtPpsQEvHNsCpuRc/G+4LlT6KU+cQMbzx91XxoEfY
LeqsakXRFP+ryZ7skXcYdnjNXSUvAm1dtuO3BNX9Ke/apjeSeF0RCyVfbR4YcOZabrWbG3ccZAUF
kFW1+t4l6UY3+o/Cdl9p/AlPnt/8RQC6gvfwHmr5T9NUegUUUZe+f3EzNHPuzwPuufxjyzfC5s4R
O1NvfNUk0jcQl9YesX6Qh9XMLnKVdOo+9KATMCAbqguJztiVYljSOx6cnFMHOEH0RXZE49MQKuqw
ayYRv7MkcMkTDb82H/UGIX0/4KekmUu6XJJqRlGMJbE8rBgwgVcMLjKnHHsOlpqaCFJo0oikuIVe
I18fxN7YqV9/lXO8BBwsR5Wc3xG6GU3gcYXH5Skq41HfnprbNtci/+8m0fk0T7rTh3/Zw8snVrz5
y5hIgmpQj2KX4TAVwrrAk0t16zWGWPHCvET1Hy7wUwBiA0fe+clYcJTD4V0SKOIlUMNvH16j08eL
8XI+/n1SRseSFQ4fqLQm8Ag2uwiBK4kKAZXqMe/X5Ee5wyRxRiaCYLN/ThY7Oa0o2uo13dHcKMCd
iB0XDfUs7/fJJyXB9gCoU7KK2pMMWxj1sDuM3ORrZf8WBSHHzTEM+e9MCJ4P005MSn9KFPVLuW8e
1lKP6JVI4nKVSR48n/ddyVRsmO4erdplnSXKKqzGBPrpcZEwK9HrblKwVjyMxJrlgaf8i/kVJ4Vh
ywlrYH7XlYK0D0Tg1OVZ7jqLgLZYVLWLeant5l1Nn/wfXAxXs53InilxXZFVzMGEo+hDwSwCmapU
57f64sTunqcNyGDUrjrmt4kDQjcb6X3ftvu+2EV/EbtuPZrcLlJo5dVtOTh1qdoAjhX4Xc7LLtaK
vibCPPm8yIgCgyPL+/sk21Mue1kxcYSn7A7ogPnkwWAFxCn8iXkheOn87sv8lT4YyRJdrW5ii9jI
1dYY3HaDsqkMIttOqURNftqV68ZSFUlx0zPHjMQ6OGopQLRTv3rpG0lGoi/aLROpfFf2XF6JN3aa
GM3oVwvXOa+kBlAF/+D7ymttdJgA5DgCXuWVkaEsVr5eL276yz1Rkf9vexXZd0kiTBYv1Zre2eCv
jK9Dqw1/7LrKCpWOwhU0b7AfY0h0hv1bMhOiGMFAk+Q6hZIz4ZNoWgsMpoXHR2y3Lm9+pyM8EQYc
8KhEE3fQzQH2Kja5y6NAaMwt0Wx10dTbasOpDQWlSts36q+GbQ9BmqS/jYuo+MB1v2r4G8XMWPxl
AzsODcd4Dy3NbXpFMtNAyr0ZSA/HVZnS+tdv8I+kFOtoJGa4OjnhxgOyzboCmPiNpxrNkzqECM2j
xhE533ioYQQ9gj2kiBmtOUP4291gVgWBNpL1+crTFb8j0gAb0amdpZ+0ppk5iQm2ndN22ochUP9S
dkQFW5Wo7BQnpB4BDM9kKS8d1BQ2IEV2YRKnP2O0lGCLc1lWrAunOhjq/l3pDtDPAbUCqlefDoK/
LJT3Y7M0Y8a3gOWIFzdvtkgGT0rsYSpAIC7HOFSVbmR8qA7XzN2vr3BCdv+8Fo+7opsY1z++BDKX
f5D4uetKetS7nGk0x/VRmHZYvZ8FkZSFd7BZ+z9bFO9GpdNUAPmwDZnB/hhr4TneQ2TKeH1oU0zr
bRvYxw5wqj/8+2yGFyMg4dM3FwBzroHPBrWCLQ3su3dWbZHgOLwf0qjD/1OO9RVbilW/2Z3K+QlG
Ez1TcJPwxKxGFbrdLsst21NQnHMdE98KkP4SVcRdGKCnwryuW8CguPwWbNk7OPaV8JpRGAf/k0ib
0cnTm8bMvD3CTD7z+Gbd6Y+zq5Fvcl1d5vhOmvzjiglGDpZMUNjmZFjb0R2/KQBR3Ssu0+XUnt5N
XmK4gmB6ouZNjKH5qShmTZxHU80bPpeZN4zrwOo18/oyt5jKtpwWNS6PpecqeQ7XM1QW3SY+AphQ
/PjnJrS9lP0yaz7T2JYTKws+BqyaQKmQPG/OdVBLv73zPTnOnBUpz9qZAWdNd1n6u3OzwV7OAUS9
Hrsfy6verZsUriNK5Lq8Kr0ZrqVEDeSLdKA3uhYFb25jcnzo5SPpS59AandO4yhoX4xzD+UIIFF6
bokEfKHMv7Rn5nDkCCcKWobOLejLoNq8ynrMoHLXtir85xWCjIABCD4ubp/F1Oz6BYA4Bbf1fWNZ
J0M0LCLRwVD852zlsY8ffC4fWNsvobbmyyKXbpKIQhit48vRjMwrFJZhM5GlRlD4XeR0w13qFZjg
Tm/ZvJXvX2J2k3X+OUw10Hs/AQvHk/oDvJGPhL/nZe95WYqo4VzLYHAp+fW8mHw/UVoT+lw2yn+u
PuNLHSxH+Wf3Ib+5KM3xpjd3pnTVw0SU4jWNZ2ZNKKLGFJyBvFhXG3N912wbuMLlGzKw79t3++FU
Sdz29Tznki8uhzhmuwNnh1T69PScqYk4RWx47AaYe2C0/NF/j8zYiUsas6bfURWm1ZwGfFDH+upQ
kk32h3CiDBb9/DR7x6oI8C7RDBGUrjbhgNovMTEYrBfs++ISf9tKx1uyksylFQkVWmRmCJjfRZiC
Ro2b+0J3lgAsb9rXHv7Ktb9T9SHweKt6NeckXCYphV5FRxdL5W1CZrjvlps8oU9qIQFlbztGC3Om
D84K7/JYww3y49QACLE7/Qf2/xGihV2l0+gnooLy9XpwwxxWiRdjKZ6tMaRqByGUz+kJB8LJrkvf
V65iBtzFAPBDWyrKqcLUONrILnUVmlJIqci2VFhDV5avNWNlzlyBwwI//rjxGEm7jks/5hEn92h8
ACo8W+VBrswMARGWQr8BjNZq0RxLB6emQkqMEJ7lqQUN1qiVYCOoLufQagbcgZH+Vdo2mgP+DIDT
3OJCfZ7hEnB12OcnHx+ydw4hrU9MxqqF/qQ/1w3jfysAXOOX/PQiPV6m3bpbLaTIn1kbJR2kgcuA
QDHxJVYi4TQS9funOGeeZB1HSLt63TbnghlPgwOdy1YzRur5k6b5UfCOBN2I67kXL0/2MeRjF1Ez
R4S6UPK7GeOwCpjxu9yidgtaxH+p58BkGCxfUhvfHra3lyDUk5Rs8RpvZd44JnEhMdm9wfPFeXVy
b5uzcn3i7b+pFCk2wJVB29EfK7xVJaLoeVXjJyz6KP1LUyQ7t/ZQZUIXx4BJuU4+qj9nX1f7Se5P
c6hbfeHbfAT2hSohzsm9D6eeuhDTfmeyQLrzAfUDfGGBbVM86oiZGy4mBNcagf2atJXwzcCihg/t
iStfmn2ozKxXGLfh8ufSj/lvLtD1rk+FXNi0Q3bZSz+mK6r6qZRzgOmoAgggM9FO7SBHVfPACwQv
UFoeSVvYlhwhmjfNBQzdiDGN+WwMoGIPlbc1R+tKrMGe9MY0js7F0RIqhTlL/XIl2tPY5w4epVPW
wrG6JGrQqzWG/pGPodseF15tInik8iCPhitURK+7KloSJ06S6TazSW1qLYajk6vwx9NZTN6ghW0S
dD+BXuJIeakDjjkcsy5MjkGLldhFFi1p0zS/9wfXFRYpiFnOhQXLh9KvonCJU40+O/2tm5XELy3Q
7Mftwdtqq4NzIPKybyf2R5wf3SweiTQPRlAW/x9InwDbBH5kRHhSx2s8O3UD+dXmfPULe9ccKFad
to/bi8Mvs3KaAGNGwaZojOWKpChH1JlA1pv6MaZdEDDI3ThHpHgLObFpU6pdm0AxV5924tz/aIs/
nrmDXvzRfvo5EdpnRt8mN8hU4Z2Ji9k/Sx48fF1+Ily+01wU7usl+lQVo1sNEYEpDQRX79n/w9Gw
zob4sGIOIEsgRw1cjEp/QK2XB/fy+3twRVljxbX9/H84CeErhXIGz2NyQRyBfRjPQgMjAiWaTAdR
ImoXs2ac6tOeBgYjDxTvPUtbiFXcyk5+rSevrf6ns0pKO7VYFosVmTdkTTTd3z8Ciy9jGSFzMpw6
vsKGIccZy7euuDcS2IZUGQ3f1JBiDvyMOMwCijfTnvYvVNWkWRoKMekV1WL7/tPJsOzi4iBz7OW9
DrTwe2anFXLC4Nb7OaWgQaXe4LlLrtIMvXGY7dKsLL7ZZdlxmR5/Ck315u6CEK88y6Av0WYjsoFT
r0e3AuDjWr2g9z8AmGZKNDx16hiIku7O2xKrj45U1m/zGOCtXGTjnJqKSX80wg+opVsjjIBxGk0Y
z3fMlmJWDspPfCs9AZlhlWBcjlnT6RoeFQBjqJEPU2fH9gLuRlwNrIMT26Sym2A4urXCLYEEV0/Z
b9ac6BR4BG6xr9tF0b/UdtlWqVLbNF4Qbsg3MRTzQPunftEkFmImbicjGFAvcktRLWeyyh26qhcG
nj7bP8qv9QEZBhmGySNAXFUi4D4XmS8b/aaTQiB9Ws+UGLoWc/TalKQNwnylUouMN+3cG0uNrEKa
++gu7313oGetCqVrgKEeimnQjc6bEGVq0+kOqlZvoHgIACkKWL3dLBCPTxv87S/L18OXjOatHKZU
W+HHPuJJBRMGE82LAmBjQWR+cPWw5JqBujaR73GrSV1/n97PTAVcTUMj+3dT093X8mWV+Z9YI8L1
/Mn4r4ufC/MbLgnDAh0QJEkjbIxZ3VIDzuinwFI57zVUBYH2FyZzpvFwsId5g80IltXJAUJsoC97
K3IlVMjRs9woqgSLuBuGgVAqSn0QpZUpg/L/wkCiTao3ZXUSmGgeKuJSTj9lhGH410oOgUVnE55A
QbejfjLkQRi4YuW4XrWmH1oFR5YN6/t5xwErSJ8kwgGRFHgRz53W4g/AGP/tq/kQu244wWxj78ak
kK5iEd6QZ1kMhPEmxo2GQwStmE5Q+8Cex/UjoqMBpoblko+dIM4nvXsFwnBomrUbhC6q0PgC+f+d
0QJ/m+uffot8fy0t8Kgs3TCR0Mb2mhwW5FOcKVVfdUZAd9PtHgHNbKUDR/Sz4oovF2v1/7IXawZJ
En/52e582Z8mRAyNNDvBN+kWaRwIN1wg9nJId0DB5aanG5nbjimpVfcMxxyOkBU4rO7TH4tL/NuP
cG6DSidr3HfD90C0IKaqjbyFOHSvZP5jRC307wXtwzqsp8L7Fi2oCy0f76I5MotKFJ1Fxf34OdDM
5UvDHEvjoCbcnzfLRCVzY47vAugW6dos9DhDLmLMwIPn7v+5i5RyIA9mJQl2EtpKtrRVsv2E7knR
U98k8eTQbYPe3FGoQ1NFmjISCFGZ38N0cZiQVGn8g3HHJi/NQkhE3i7qzfRA5aIuFDHXCcaextvD
mD2NVlkCWCwFyEdw7dfVcPnCmZRyubC1sZkHoAU2NgptWkDrtnbPZrmc5sH9/FMT194svYMGtoIQ
vkZTY3inr0ADB2NGCafimRdtKoelWvrWJRLYW3Myb9T4dWFMjGAt3S48F1YeMG7p5DcZepliADm1
y9Jmat93lEz6MNKGdGp71ljmM8FKjJW8rXVW8AOXkx2cFEmukI+yRXPw00DX8zA2UWjrx55Dh4iT
YNWEBelIT35HZTodbEqhw8uNWkb41ii6M+vPqrSmeVDYuv9/JO9Vc7oZrK6rHd50QGGlbqdHQ+K1
0Cbzit7tfqy6e43C5GMSbJjMTfZrTZnJ/oyAAddfUBR3cEfKEcko4y7WTvosdN9Zh0ns3V/JTbOV
WjzSNtsLii0E2JgqL+puJhWMMG5h4FJbpENVct2AvmlfbMZiE+V+e/Qy6+B4hxehUGuDmRveiHwF
1w0keU23qLBAM3cIwObrt217LU/mWvXlmkXn/zekRrxiGpZFbZTs6VBDm79xG2FFUQUuGBRM5G1X
x/TQV7hvSorX316gI6Tcudolde6YF7VZXV/SEEK/BK9Y8u51p6iinFhe+A/C9nrB3AOKAMIwNZlR
tr/iNWrZ9PO3zhxoFFO7bz+nLUxEPP9G6gZ4r6rOEfhq9UxY3LxZMiWh/Esu+fxOrgyEYCxoalmA
tZ0eL/lO1X9dATK7Jz5PyaB/tUVC0kwX4O8jHKR/yZAprLB8j1du8oTdMKMC+5xsiHty8GTkS918
ZW6cxfn4AXHxMuPAqKQjoJDdE0wS1XwAGXhWQtACVJBkv+/ic94ob7a6J+8RBR08uIHZhBPKFsW3
fDnAOEhxMIXpOYRdHyRByGGwTl6YdZ1+mZ6kDIowg0KLWEc/ClvONE2vCn21TbkvbXI+qDrGVoKA
/CyzX1eRSxeE6ewQ4S1YPxhsHYsN4zlcqMHR6eKfnpvdgJt8T/d+WKBBaDgRyrw2zLUn8EZ3jUvr
NRAq/tlHWs8m3cKeqU6OjJVtLj77HtUgE1xjUus9eSFVJUiku0wR3QQ6I/f3knNreWttVB5hCPqP
04VyvCzIcGAnjBoj1k8oI/7h6RD5bnkbD1IR3wtz44s9vZjgJMTus/zNrgbuxqunEvJUHqN5LZCS
j+MisQ2iI9MqQtz0GY7mkqnIIX+oXTslsoMqt7jwuI4gpmMVGJRO3AKFBiaw3GspI2s6ti4G2vVw
w80uB7hk1vpXibY3GQnvXyGMA4r04mVgQln+hc+4CwBxSfGBZcYnxJtDlFea0bzJtjW9Xuy5eyUF
Tla43b0jpMxBgj5rF6ORclhHJs06NecPW9yyQarWrdHNSMgWHZjle66esqW0GquxM7SsUwGaiYuX
7gXnYQzO4OrQ4DybUmYrSU/1LBy9nAb3LrbPJV85dlMupppNd+gbYOI8ruqFb2Pu8Px2WouzECGv
ykaO8pyTYsDYafaWY89q7oHaTMBnHJX3Xx3bPoz2qdV+ZpHA/xb2a1Gg7dtDB5jGLOaCzvjXHnfL
ofaVYn5nmUsAMQVrRXrhqaequ4pdBgypb5bRZ7R2BTQ6Sdgpantp0d4Wv6Nm8x4+4rNptjOzzAuX
rpLazqFubqdTek3Jus0mjNnzcYTvVU5AQM+m+/SrjllhAPRV2wv5FSsi6viXhtjbZpTCyqKpcBDM
iHT2Y1x8D3hB14lG+mFuehcC80mhiQdvXIKDhXvQSJE1F/X5afZuxpR3q2jfCxjCtI76SgOLE32k
ZVffjwuDHeiV/vpiZwH6/kINrljEaBO5EudZltYa2API78zzMEBQCi7+37RIh8qv5N47vWktpVar
hGBVxSxzBPxMfWLm29/2z1qfhbtrxHKj2ZNqte8bT0nu/sGaB8d53uDMK2BWju0Qbc3fDWqZ5mt7
awGbNSIBuMQMdXm/J0JCZehF0KwVzDIAjapLKyXVJjt6EmnwAUuAuHOLPlliStyIGScJdFP5Ag4L
EShHW0EUEPuBG9oHgRWngJ5zvZ994Fg1Fcspx+CoUjOlbD1Mbu39usrpiMNNrKgvvUUNRZiIPuOI
yMJjx6s4n0HKV2+cjlsFZJ9xiwXg8A7jWjoGfs9vrvXCUAnlk5Ka9mK3qvauwYeehBEZgBcmUCta
9N1MDRJNROjTcKUuzkCYMWnO6bQePmraVh90wPfmSPJULlMfH2Pl5EjwnsupSpTwSHejGXmF+d6C
tfQl1Q6Njo4QHUPfs2deMzs7HlClsZ3gndG5Gg+C3PfGBpi3zMx50OKy5/y0C1WNX9vCH5G3rVwd
Gb0XM+MHWkYdHD33D6mBCrRXdokbEkxxBvP8OT+pL6io2TxWcZndP04eFr01eNMB9pReitlb/uYp
k9GzMUMY1NuwmHmwEokiIPnbmc2cBTDDerhNXX1LNNWy/QZPHaM8yPaQYai2pqfuHs39zoKtdeZZ
PnZ8bSMsUGJYmGt0D1+gXMMt2Bo2HSD6c0CqdLPhL8kZAbUAYV+wnTh/pOrCtfp7sSHSxy84yuO7
jsDIrWeIUEPAAyXsJMkquo5pC+E8KnkpQD3c26IyK2pjzvMo4vTovvU6IzwiDKUcHGum1/nsNfk5
/d0XECt2gHbJ5b/wpfPh4fSg34pTAc3UQWlgsOeTGpnLD+cBi6334l7Z1SJQtkyy70pxmr4hsmJO
orwYoASgUgf8tqfIm4bpN2BSwYXlIwR6fJddEPJ4pRunWQ0/NLK2WZg4FkmjVAo28gGi/zo1J0b9
z1kGahQ9Wg2My5WMNFkNn9T3nMrGAPeQqelvobSeCNSMAOcM3EykNCzV0yIbUAjsQ7+/CNvQQjp1
idxUtz73FklusnLAXg945xp+MVFfc2PgARa8yf5OObpN38ISr9SWOgMdy42u16WFbBWWIe/w2cY7
FUoEQhlP+N/a2dSuitiZo1tWQQEFYaavPFSC+h1TNeceLf0K6JCVGnzRx73cIF5gbhC7lNQD29ej
m4uYzVLDbNlqVxHhBPIKYje/NGL2Z1uJpH5UXVzqhFTSTyCvB3CdKjYwHWY+aDLI9CXuH9gorxom
MeVVYmAZqN4OtG44vjTmg/GUQyaq91O4/UCrvoXJRE/V+Rf/pIwhcooilOoLfKQjGcTJVVPO7e9j
NFMez3/W8k66k2cGb6F8jw1P9sz3N3F5JtIW7bzLUh6vW2WZyxZrIv/UzUyYAsqvC/xAqh1+h6Ft
VAyi3iomv1moyAvGbD2O8Lvtbc0E8QxhK0TqS0NJxoe2ejwPIexPnjkZEglp59karJSebBBZbx6y
6BjmILCaURpr/AO/4gC+Pos76+xZU3bjkXinakOr8i5geKOrWH44FKZiDuQDwV0JESFAwYKvzpJt
a58H3HKYTuvWuYF1XKnRgElm+55L1FN5FniskzS7lzbkyZCWRTl/71jfotwGH1VHur7O7GZKd0+u
HMZYYpbaEx1knhvWMWy7vAkqOmKr/4bYOktEZaRCuvn0iqbF9/Ed0e5NIZveouKi72iNEJJsRCig
G27AwnsXlqw0stSRP3ytI3G/4lhpN50zTFpljCw/I/rHNDqPXrZsJnl3STlenETYQmw7/mApkO5l
Su6OUfB4deDw3XyRsxzZhQHtWRYcJbMDVOMyf9XKrOwLPL04b8QVLcfSOYpHOz7N3PzMvlSY0NZo
Ve/aTtCV8NDbgUbUbUsw6TQt97dhNZItcKaU+1W0SJy7dPkPooNAepzkXsZmrkVxUjTtwqB3Eysu
FblwT9/QolM6noV0Jfde+i67JQ2ziovMw4mjiHzCBaEvVYcssimu0xa5SOxauskIC6x89WxCT/H+
oT5skEufEqOeAsOlDArk5muRkxMegs+2ANvevxb5cjm0fIHqtRw23f8beB2NZ8i7faUzvgXVFdXo
grnE7a9PCLYL78GNdlkGWw+kV4uP1yqMlSwSNhj7Y1swDSA0+JRKYtrR3mr2DQ/RIYAouPf/oDnQ
KcYuGBVP/E4bIzONd1BLRQYulcnFGd749c3TUpVlUL8nGh5rYkes4agQJurd3xW1rWUMV19Ka1F4
S1AMm21pAlHU4v5KkLeMlmpqGx8/Vw9BfDyBFr9esuXL8Jy6sxOaL8TY1rgL0+Rwnq4gImrYGqG2
KztJQjxbKB0UgHqSjDWR9tm02jcdHgS3/Y7coLIpD5K9C61xiLJH/B93Yp7XrD8g1R25eO6KFDzU
2SgKLUXMqm50YRSwXqmyUGglMb9AIPvm6saEjr/YFsHbqRvP9vj7ecDyKbceLs48BBfRwZaYmdUD
yxizTu0byKm7aBXEI3fdyRq8OhDICtqZbswkvX9xZk7cNrZAC25niocX0qCJhgQo+oYG2xYb6HhX
cqM1rroXJGfWBG7qcGkPw7EgH0+kCcFipDHN9BczFUBdcNcuwILKDG1fcQWw7/QYfLm/t+WH540K
luqTmFvi5Lv4xmSPmm/VDZoRaCut4LgYf9q1oasNY2HQQNuquxz7VBCzSo7wo8yn9ST2xmm7Pvlt
6+6nq+h4zQZi2MWJOh9LblRBJVKhZSTReFYE3ZFfolIRsBMosgewJZTiJ3Vvq6DOMNxbLB0SXfBf
NyMp+qd9CiE/rWop8RxEVawZmsq6cm9wfTcU68MGePbCfX4ppQuUnf3MFGfrFdr59/mwn9SgFXsH
oPQgiXN1MmwhYTaNUeBZzJDYZvUkpUwo1DSPYwKuHn4/MzRIOI6PTj1riitT5wRhBllx0ZYcSjGZ
qP1XMd9ewAo+fnDDD8QlFcqe3TzRq1XuObbBsm5JkjXbISj8TXGxh/I/+iLceYNdljetje1Dc1ti
ryhoVGRFayGsYWutI5qAMHJBva26/bhjn4329j01WrPoY6wsKfO7wTEn4pWhaZeVvVjuIKZVhI5H
RJjeNb3RdEXbivrrveyDR7hc1OEPzLzantEjyThvk2FuyEldLRiZD3Qe6NnnKd8uwza5vD5jvksj
xhVIg5o4t84zh58tI06tYudCr9FMMHBEU770yXj6lgOfmWgFn4UWmncBMK7kS+ZanaWwYatn4v9P
t+XgTGSvFHI6uDpDqDo+hz96tt6xOx3FNCXFJfbPPhyro7PyrKHwmMP13vtlzVA1w5tHv0JF/YsX
RnkarWyNxUIBg8gcBkb5hFeDwPnokmrSqOIprllbUc2U1tZrl0fiQqja+JYlv1QBd2CzRL9eJctZ
q8is4MFJOpiC8iL3VDOErXtzJ8McML+DC3a3DymJak0ePfFGZ9A0GPfAf94P4t83c0kdPiIDdZ7C
yY7kAhJZSVHBHoG/c5N7iL35uMyuuaZEqloYHFWX5fzxZVKi4tfVLFWwGl/By12yPIvJm4lEmOpx
p23kmeuSwSKkrerfyu/oz6+67dl7w+zTi9WPWS42fAQvegDFEdb+ydz4yvRE5LfSEpS4tp0RH9h9
qAcVAuU97GUmrF65V+vwwzj/8QY0MhKI3pLCNxQLg1q60ZZBOUkSeiWu5kF9YQL1OA49ZDsQgpX/
T5Ah6PN1+yKx8xk3pd2vPwnwIBMw07bZBaFsx5Nt7OHc1aE23N23qk8EtzysT2Md2AzPW/4zUmCn
I/r9TsVMl9dTFBsuAFHT3ikDCOEDJxFxTlsSX0dBfLSsBkE4ldXhMqnxiL2cbXINqteOtoF5c33S
OSbSRY8rAX5WWkcgkZf7buc8dXQdge1nP9UtMsFR6ph7Dx0i7x3V4PzHJEhSz4qGXm1WgyKK73I4
fmnNAppAHefxmfybwoRoT8rvX4dHZQVBQTcv7ehD0XFH+4iW3LEnvFgIG4d8S3Yg8XEgvZoSXuMY
L5wz5SZtMeSjvTu4cbVsjVNnVjFxY9+UsGusyWK3Id+GabkQVc0zmItVQqVr39D74JfoBWiDqt/I
DbH3Enp3H2/VPxsAJr8Gii8ekNBOL4XPx5peg/b+yKV780cF9qghPKduiGQVM6lChQrGXvIPyjFb
lSeR/dpWyW4QXO7R/ifPQusaQPmNzVs4IWkFZeSZPgqEAZjMLZXfGWXFJdgEol/4NVe5B+mxs+n1
Dx4Fdoape8hpjaMKyYnOwiR1yfk9yoOEyki2FhhYpbL9cNBZ7v98ZU6kWNHfqGf4g9poK/ZIQhrZ
sgJMrthfZjFsVLJ52Yss5z3i88axB0gCvx49wjExlxZ7ciWjepgFFqgnzYaorFHlKsLA3jHKLEFk
b/2G34A7rmAvU1Ft93wta+g34VSIukXK/k0JEsjbhBodfk7fIh3MK00MisEc16nnycEVQJ4NWRI1
bpE5m41VwR5JGn87aavxZIhlq1GCTOecGHLznVDBbplDEodMh50o/2s065BuWaQ8eJ+/+gpdk9TQ
8VokvN+Kjd/YAy3Kr7UbMQYKCzvhxPCyNI0qaRL8yVEhNu8Gasn5EuNkOpnTqESVEks2uPndsTAS
+9GgPb6Z1JGTIeYPKd1YWfjEO1I4zhOftFkXEfKEJt9TjIq7Vgol9Nk24Qm1giePPzU/Zia0Ndo8
o/H5+/xWKRNtmcWbv76t7cj8uLNC58acyaSe10rECG68R/CcU8PEoebqHfBZvnCv2a3LFJXRgECN
kl2SbVbBQ16MhzfHPEdbu0A4bipEzAISuBYn9p2h6+iVF/BCUesIU+Ja/B93ABWTrKU3MIJL8pSF
snaqj0JFgsy5pkCS9lj4mlf6dzzaiu/svQ8m4LmoA4IDuZwypo/Xk/Rfu0otrEV4eIg4RNGH1fMr
YFWZh1VXAwP6WDYC7UVv/6QGXaf+ScAzDUaiMeKhO2gE6f5O5KPpI087m52r5QGuBHKmVE0rWk6L
qptNXp72uMfhhmRniugs751vUPE+UqDA85FfbC3SdcGu13EGarmY4fjXKRKyKZgiBDmGr+IyOnXZ
rAytVc9WNjjo8ObiOSzMYa6E6SKg77f5o+CBePWxQP14XNYy5Uxtc3Uub2Lom+YTpbFf7CgdMNkZ
c1m5hsjrDvgaSK3K7RhnJLCnJOn2EcwzT/rDJlhBvm4AzaCC/q5O6bUhJtTuhcFd0W0bjLyavQr3
4iRof5tGcGcZ2fKP8ZrUkOd1wvBXYDwAMKpIfaW9gyFmExoAf9bSAHNTgX0J+18hu5Mo3hUH0E+f
qk1p97dKZ4aKWf+KQfmOk1NV9tVpIwXxb4mCDO1+JRY/o9pTAT6mKUxNd9PNP4bMW9L1QWiAWl4P
x3tgX2CaavcHQoTu432ysgIg1PT1PZmzz74w1CObO/2Nk8jM/KXg0C5b0o1xMOhktQ6IN6IQVqmd
InL2DhHWopI2plWGTNCK3HJAdsYk6l7gx43mfBJTyMiqsWmKBRMWw4Php0XdpwApBmmJZE4ufxAC
soZlonRcQhrYEE16v35WW4xYOKjhhWordxOLYEOhl7mLqflvlbyZb7mysRaBR0DTAo2HBMI0fQ0R
MAjFFrFm45Ckh9CqXYstMHkYc35ctoPMtLpdwyckOg38DwLtxpEM4Dztz5wVSM9VwdZr4w/ElSrV
ilYYgsyaLO7Dp1mG2it32PLZOr0jcwqwIMVDAJPrbn+HfkjOIgpRkqhkLy6aHFqLL4VtmSx1ujdh
oTpeWrPXI06UQUvJ2bwfUg/0DsPNlhO7rBHpIi2bgQBuZhPh7ZP/v6p8bdabEyrqXqKqtSsgpqUH
I32bZhQw+EM0MyigSTE+2IQV5FkUC8YGl9dLLE/6bvREDOBaI7C26hGOZHS5FwbXccABMkt0YiZf
j3CQwuj5lBN3xxAXO8vmZ3d2/mx5QBebFcsu1VhBYexmK9mDtGKUpYtorOsjaW5EVIkBSbTi6LBV
FB5nDygQLlrOA86TRT3N03H3Qjmq0vNfG3p0sVdthwcqgvZWUGHOg5tqAESSvkHblp5l+iBn7VOk
iS4nsryZeBkd0r1FC7f3LgUV8miaeQ5jGE8nD3KBu44eybuvq5XKj7b5GQuOKrTm123QhD6nPU5Q
leepgx8ks+4oeaH10YfwPeTIv4ASRiwzQjw9lX5RZpjZKHFnjkrTSs+79n90C7AHpBMnYKKbAzYM
dXPrm/cQesXVhiDOh2Njrx1bdqMpQrfl88M2NFayfvGtiVZDJM1hKaYmwk+XULiai5npqrJDAMx8
474T3EeAMKXGLrRaFGE1L6egIKBWOeE0dKeNOH0HbCTX5v55RR6iUsx/a2CPBKi075Y0G2moENjK
HF2DSBydeiu/rP3OgWHHoPz/HAxxPz19iP0441rCblSY0/Ivco3xVY+lAmEpnxIolHQKibGi2meE
tf0yulIZi8heeSoJfwSZnM7ok5Wth0QV7AzlKlff4kdHK5qTsTLkyOit/c8heEdQ/nAq1L2SdFkW
SyxVEcrC1th5I2GI8wC46SHhoWNZRGVC4N6JMjrR1EcE7ltAf/cLnjejglZeXBkK3/vslON481CD
qeDwfDGCT4hz6tRsl0DFPl2jKVZBsAmwXJDiPpoYgSjoNAdfw6dN8+/jp20MhkkOtBxTUnYyzVoN
PFJScPoip0ndn772ceiFSaUf9729X6jmr1KQwYbZPWU9+GJ16S5sW2MuD2xnA2nVE07Qrb69X0mQ
wy+4ql5LdMPAuM1+tcIJQ4C7GEbxeX48ynFEGcvqgthtip19MxHq9l20TDi6trKwsM99s0j9cjIG
LJisPiNhW2UGyVliG7pod2L/pQl0ikiyQnQW+UkR3LqeKSzHEDCtBsa3y/cGF/tTnA/sR+sRP5Kz
yWl8yDCJ46QJPXpeXHCnEaA9FBNqXCHgFIkcOJyfKcHYK1kjc4qKVOVzrOfnfyrVRjfYjkigXIQZ
7cYrfpNVoblPBI9BT4xosVl31Q4Xg89b3zyqLk9Y02voLu6tp+88SlqgjJADg5QEfmnGmNUADEdV
60YieqDvsz4LHKTyH5pjyiGo444ugKRPj3dLvKCeIilVh2wHicP7Bjc2Y7bgTT1ZoaE5ArYLVaIm
nvCxdzL1LvWvIXLPJ0Bk75zsLMgxn28K6TELG52RgPUNfGGyjqjgDaCxTcSCfUt1th/4IXSyljQY
ySD6E8bfXd9SeO0KfmLWs+GIGpUSmaiPeMIrbvM4yg+CkflBEEBA50EtTojmhVNdYBnffDVeJwoD
cKxYvP0I1+SYi/Hl8BsBuRkIBcMv7XxXah77CBvPqp2dAkreEGKdC1gQp6X5XBDJFjDijbpJe5n1
BqvrlguyNpMuKUKu7dXnMP/yNKvjk7ia1/jrT6MVh4NGY/kFGBL+TT6q5BaCEm7IGZHaIQB5XAF4
+vw0f9DvUefWPoiVzHAN0E1F8oL29FxZ0PEDyEvdFbOzYIDo2cIsBS/NArMLuKapGCBJkatwF1CF
9OzbAw/2zzDFmJeYtTC7IrNAxrmremuwunl1X7B7UGwGYHx+twEV9p/OuWUko+WJROdt3pTw/QKU
QNOMQZ/491yZ3bC6YuB9L+INnBPoM8W1yX/SiVUiUON8m2+iv7eRmnx6Hj68vI80T8ol7VkK2dnG
e2DkBLbMXjEPfPlhPNwxHoocD7RPA5QF4f/AB2RfGz0IrpgFAbdCrR6smd370e0MJhyDBqCdsmBk
zQnVnTew/oUA3Iu6Lvj3J6axbsu1mZ1ge3tNnbJ/ks8y6dFPGvrcSbPinIckP8Ydg+BZTRMCvGIq
GawCjHPt5X606wwaLn2asauwRnrxzoQX4nIC1gPkXGZTjVCqeT1uupGiVI2pYJNxPD2P+Gpvzbui
rzPgTUi7XPm2wzKT4ksVCOTYISjtJG2e01cb2fIPoLe6T/5giX4L1GiywvhRTT9KJAB6YdIlNndH
VBQASEieRRqf1LaevxvXXjo9dc8wnlclkoemV6Jr+q4yeMT0qd/amMO0YLhUtTquGHbOvY6pOhWg
eQPFRTDZbAGa3+o2tTcNu+vAY4UYGK9lZjbQPuyvt4cYNys80CkkiQAQXzSPcAaIbmxtt1DqVBPo
flqYCoRyIGhEcJhGdcLJvmzvfP0gs7tXJNx7EHfG2Atiu+8T1epc1tVs9HjoNQQ7mPUKxcdJEF8T
SRnyvNIsQc26sMVXYr9dCPr9sVvzE+I7OchLLoITzZQWLAmSkl0ZJUp2J4SKQpbgpUiWAEOe2+db
WEt1saDN807GQesbQEWrueBnkmjMlT/Bd6t56DPA3Pd9yKo5pEtGBxLYTHf6vXyNHtyf16zwpSn/
XRibfCriTatO1NE8z9BSgMW5Yg5Sko5BUTOiwXmGYohcf6je8Y+vfsh1+wzZSuPGiNjBSv23lsON
khYoPy6VonSKRXEo+2GHMpDykSRwTHP90fKpv2HsDaW6TNHCC0eh12DihAy3EIrB1bCA3zzIrUIj
8S2rAQUUGacJshyuLVGpuNBwZlmCaQgAu7HlWG6kBqZdBAcqnABAx4ajD6Uer6traL5fbCxE+lxz
lQqEZY2+c5VVWBIRNptlkMo9kmoE1U83pYNOEeDvyyvgeTjAfGNKv+LCcjRJc8H4cg7sqEgq+YRu
Q/vOW0L5s5PqGwdhObU34E6bWcRvgVACICYlaaWFz42hB8zQYIPPUKnrNApMEnKBP5kiZ1gATYox
2nf+1jRtumeX/RoIMN0veF8WLH6ynuKdrxWS2vYs4wV7dXofHN5LPTYINEwyg7Ns84/drA4iLdKc
yugHftQziB4L4J+h90LveeJfjFlU3v53gP7lowFS9n0afbs17wq6kgkltqWHXXO7B1+LWw/pCTGp
zI5xnonu1adELWBW0NBGLINVp+qOn00qGtc8eYcqDSeOICEaSH/zZV4QMN+Bxngo4Gnf0Nvjj33J
nyrRGbnfelglR0nTxj1i9WfdzSVorkpw9/Z05xn5k4w0U556wO/usGkW6Vy9ZzL72c0RSTTuFumh
zKPhkI7AeKJ4Or+1v1OXYb/WMHJfNKBTueyb0IC3LaOU3WJ46JRWyxk8E5pRwDpbl/PEg96SC57i
s9eHJl9BIpcdwxdNfH5GuaznFgpbYi7Oe8oUxJO9Rfk3A3A2P/EzeY7dfufJ8d7EUJQYjjAKr/Ph
/cRNXYpa+U+RntQjydnTdWRSIxvTH4jROAZAdkE2D62RHn4r4fJvRlI+Bwd+r+0ZGOKbOG4r3sll
/rU+xFmTRLV0CeOGTlXLRDWjBSKouzoUf5nkExj8wOGbpFSkbohJu//eiJjbb+RdkmqTq5ajZSAn
iRExC3H/WpiaI/OMErGejHR1FwSdqDtc+ulLjlnt+Q4hjL0Sh4jrHfgdok/y3nlQhmvE0NEAg0so
U8Gfu4tJb59i7XGWbiLAcqbowyPzaDAZ5Ni3Hz4nOvHAUqIqtYGVCsh0wE+F3rVtbnRKdz7yVXP7
rvD1yPnzXomEboJpG4ecTns6lyiPP5Z4JcwIaV0JmAm40+WkboMVOcM1MFDoGAUkIuEFVFpBncYF
q7ibtG3+BsS0bkWwRzsd2lu9ZXrVslNXQWH6Tt6rIWpxKXmBnO5w6IK+iaAGD25GBCtYlnfLU3tO
Vo7wD9xB3eToGKQMVyfnr9jt0d4OyIcemSJj/ixdk1lgF6zPp2uzosJNb5uFoT6dJGNKLQgXWLSM
0Am6AgIR1SXTxVb98wN+YepBJooYmy4obh3hnIbTi6czQEwNVcnLmscirNCqjqsAYXckLPnfUZlv
I2uThW6+Q8k/Q+9m//TI2XWOo540VmyZK0VfRwrz5/FnPJrl6ubvjeELkFNPmlnv/7xaf1e4UdeL
X2AGbWkYHrsb+o5wfY2AJDf916p9G+7TwDpr3czJ4zjpaYoKGF/c15XE28cST6KkbLCW5f25DTzb
KEx+Yeo6qk6fdDXczk3sANjjZ4kFVvhIOQqgR1ydhqTNuMVzjxjmaSYtFdA5bXSwWW+U9CRU6vc7
21V4ImhbdfmNlH5JLhVwcZilJVfZK7n7IMj7ApntJZFfIRTBTG3bhNqkOb7u/fsdzpcNST0iipZM
C7negm599GM9Ww3w9GjtVK1KewyUzYsOhh9FtGVhjvgzXoiQ2HnMpgdeCLrUPRWfy5v4HMsLb8cD
nGVpmVBHHFUD2x3EAQrmiDzqcRAbcD8dewdMTunpOSiZdT/2voJvXVZKQq8VUu1hhzj7W7mJEwp1
5bDWzcW+lk8vFfMu/xXha8QxdSY5mQQWLm4ZqM8Gnf5Y0akjgNNDaNBKNAdbkmTyzKN5F/zWsLCE
pG82ZiZI+qSQbFdWeNHsem+uQ+iWDZoxr7S8FYg9au+gJ/OKSpXs9nAiu2PlKFtAshJQeaoy2++o
Fx1zmgYtttS1g1aD9LAyjBSvX7o3KixXEMyyPfbztxwYWYbiJ4prMK5KbJHzclOINBsk89MYJYtQ
G8xpNyUFFdVrr+HJ9wJ+ySGC9s/d9P1cke9WwdGrgIsiYUQbt8/LWk9od/BmuYBKfPrRmrGv8Uvf
VqgLEmO17lXW2uPnNaW1DRtlovREfqSEXvIai6QRQH5Q7/BQbc9SJfattpaTjLqbGfjajnnuRcMf
IIt5BXSziDkAx5voLkdNMt5144AujbHotPfR43VA5YoXdtl8BUEmt6RYNIqM2aChobVuA4bvSm9S
CJMXk0Rwu7+Ud/owSUlp7r/mjRmNR6nk2yP0GZrP+EZ4ALRZJH2rugQYr39q+frOMSA48b4r+mcT
wriPGP5j0IKcdgWSSA4kCH5D7vUt4asx6TxybabpNokGXZV3lsLbN9yocWMrSni6TlB7SrFa+ZTj
JqxXcDV7K3bnfJgFYQbGfhmTgfliPI9bQVkuHQVgV8CNGfcoawbJ/UDo+l4cXtYynFa0yP+2Y+Mz
Dj9q3gs+Zoo2Sfj4cYzV6FNwSp3GlS2CHtmRVo9XW21XxeXEW0c+JDDZvWyL/BoYUqRhxXtMp9wa
c2l4XvB9yjhQ6mXQNIENKNEOSeRf42DsXYO8ZT4a7avm+CYZTGWq7eXDEKHYV1JohIfA/Es+o0iM
wgshYiFGNLUJGhR+XYkrPIAwGoEyIxSLnRgpvVwEBXAgRTLh+HMD0hcTIdAnEkgBWDgQY15U6ycu
KtjQ+Z3Ya9YNx6I38DoviPWvzPB9zr6Ea3mX+/7iD2KGu5TtgVOnx1WBt7PXIO/fLzUxpGNwvOyj
fuK9ECGyWtrcRtEKZAlJpooU7A4XDFyGGt5Mv+NF+egGDEAGsdGpS0pIaHdhylMmOBZzcrij99vA
UV2kPx1ej/qTOMqVIcCyWvOc5NvY+D4FJrjrgO9FuKwYcKtUrUYhwpYBc5aHU93mBgwxZMYXmzcv
aCus8rTex2TtXk1FGJz+TQiZZOU6NuYXZIrrValtBmx68EiKYglIhg9srlFyZfPsN9WB8QaKLY1R
FJkk2VGbZYi8i9I3qaoJB2vUY5DFcXm9LwK3qagD3GC0mu0W8DVQe72S+MyyV3Ph36azfvN2+176
9KJ+/Cqp8spE+ME4/RdfLl/MeW06SUenBm+8/941sJkLL2PAe3rulUNZWjjfpDYZmqlp74+aA1ID
fBFN/W86scvtLuVVbpEIRme4J+Sts1fKwl9nJ+ACtn7L9dZGvc2NA18soDFHpHX2fl1SVOwK8n+7
cKSJIBTkRPCgJtWX2o1f/g1x6hHzpaeAwIjnAdyFT+jNVWDImA+a/pZYM8ZYWLSrKrD8t0sg+KN0
nwY9hCvsyKRRXgJfOjIlYDRRpQpxrZfPpGrsm0mGsFDzunBdgZEgoQhr36qxEbQpkxQ/e8rzl4Ic
zSTJnhp/H3Uqw046p8QRxlzosglHQb0jpz1221rQc/hKS8cor3yJNiiZn+J71/k1njj+EfPv0LHi
R0KgtNOQioml/BFvyV160jbDhTJXdLlGgs7oDr7yAC9Y9lSDPj2KWyqeqvaz8nrxNA+RTidFQJ6t
STsu37pRyRIpsis445rcvjquAvx9nRgEh9OE/BQAxY+z/P9XYqXLTkriFgFZRw3xDivhaKk1/Pe7
EUwpUIvxBAGBMkUOn34t5WIJWXhtX5mlXrrSJr4j3nDPvAjxnwuclBLOekHqicWhHJiSXX5X+2rf
vaBxoRaL5P+zqp2kgzANiga6hovIzdxcHiLdAFDfSSQsFxRl17x6eAAKO0pgoMVZU8SVSgZPon4a
TpMqMmMaFJEyMMO+pcODrkgaxHCvJAccR6iqOo0gXkXSSB7tBSJ6ZAVzt9Qqi3H76nsSUExN1nYP
IBXKc8tA0opeC51JAPMfmBfdasxxNhJAhQBI4KJkuKVgwclmKVjDGnJ0elp6ceCpui+nlVooVhxo
267WUHxOofcdZUEQ27K906LOfpTwxabmVo+gK0Kx29XtrGC3gn/MYtV5SNZDkp5cn8nG5tPnvF0p
HBae9aGigyuA7gYiCP9LHkKLsMwXhjVZZBdjjg47ryEotaKR1Es21rw739UpbguYfRYcEP0uRjqf
o6lYJiz2sdw2zw8t8g5XleOOR0Pz5kWvqbMq+ANtV3bcnNIn5Ggz3CBVZ8Kjnssr0UWI+Fss6Ccc
JJ+kEIHkrKc3wRjBZPskuhIP6Ho2u58kFWdDmuv+JGzrBFiBZV2g3Vz2DOZ9op/oQ9RrcH4Ya1oR
dcCKgXco2TyZ1qSvWW8mhKLj1L5ZKu8fekeX7KqPrpoq4NVO7yDt9FcxJn+msI2JftBjJajUt0Cl
+1jMt3xezf5/Qm1p0hKD8t+CtJBvLg8WCHBrEV1MnawHCgGZvoD0o4QaGg42Nv5WAMHEbKNbae06
0B1u+T2QvDhUZXJgq3hNmHINkZutZvOvmqqF4tchdxtLhHOWEHS2KlmLdrgztxsNNpEEnD/j+Atr
YICNOg+6vdwdBlwlu7waYkylK+eaKrWOVviZxCoYkskPM0rr8xw4SVT8+T5Gm1dDZhqKaJ5h65vL
PNCgsmxa9UHCy4eFLKkvXnipdWCh5ZQH40VJFnCJVnyoBmN+kTy9poZiBcXsQ+kDPce9v9EcTG09
bP14SfuPiNRI0+nGWktx2AfPx7Rs73qVtPwVl5tttobdW7rN2BSJ/JJ7HpOjvILCYafIatWcYVO/
qbio5KxRjsqhi55vNqNM+qmm350SefcYUd/XV0UEdJQYeJxlkGmLI15BjngjgQOAflYpkhWOuT74
TD88NWumWHdZnsLnHZvux4D6eQwBq0cISFXYDK9Ae3KSaz82LWJu2xwl1Ynl8lPcPDlayhSQt5x2
DvySoB+z3vOtnYIq5eOLiVIu2s2HTPQOKd010bEo8MLnt+tfVq6H9cTSSdKUoVP7iv77t/jM05NK
Qm+fvAeRTG7qMvia63XF+MUdi34en0np6Eex5o+TyfFX2uM5nQt4qLQGNkqVuYzXFcVq436H4las
b/wLkXQSwT81WtD1/Mo30uAK08JdHNvJ4I53ZGEglKVGVFkxQrJBZv1BsNlDw+C9ldI0pa4L/y3H
5+y/8ekRouon7I+TgzfjNb20nPfkBiNCFwNeMUUB6z2sKzVo9SQL1NllX7mi0BvAuz6kJ0uEDuy1
wfv+7Zecd3qjQ8rfSc3EG+1y5WyGobEoiPEFpP5FQ2guMTu7cGeOoH/hgBB0MRVbjJUAVL1AlmZ+
87WS29GxPoMgAnx5b34EviLU3ddaBilMaaIx15sUC2Uv+3UNZTmzX5RDju1ENyZ9lvOxsyPY4XL3
1jAPe3gLiSviCJJgAeVDpjVqLTf3mzwRDyBYpFHkDxXZOu2vtrLUeMpcJYXOntIaCWdQ5IaBtbcd
Ai3a9jpouzcCxDb/KCR75ajjMXqQndt73bHKCOgng1bdjnW7ZnveKtx4JCDtpzMJGNsBv/Yiq0uZ
484Yx6bi91otn0vEhapqZ76SSrR2PL3SdALXZ+WMI7vuoJ6JsDsOMbqq8MmGNxeFq1DFjI5yKwvm
VzD2xZNLnM5kKlG+W79Hnf5jV6PtBARjfWc89k6i3hnhuGc8SpSiG6KbhsxYQXEIZhM+KsL1dgTM
jgOMbahT71Zitk2VwnHFxoG3iQwkKDVCmebZJCw9didZaKlE1aALmQteDg4vSH8Kxk/K7Yi4seyr
CqgF+jiLidLeSj587LThSP/WUupiSr1NpCbHRrWfMvP/bzivm7+nJGyMnSWZDfTUYn7BCuoJwJ0p
+RcrAzbgiy01lZhx5JVhl6bW9Uq3PuVl0BCebX0muDltf3qQ9AwhzKtl344FlTo/EXgSpAzr0ZjC
8muVou/couHK+eNxgdaniyWvHLeYDmRfXiaj2ESSN2NZe5j15RZXfQDRLOZDps64FW9mXeBKp497
O19zbNG5pdV7FdRXVAudTa67dc5rbIV1DPzsPxU6p/q8AO83WSy7BfKg/0smrkLTVXsLoLeaqSpv
SoMzTozWmeQmW4Sw/sHjl72jgKnK7aVtdnvSlB7Q7ELPxHniHbOIYydgcUOW6HLYdenwqa3WEn1j
HlAq9HOm4h1BdPx3yqtxIxE8wcabzMP9Bb9nJf3OOYWmh+CTZADahblwcxX4qC4GmIobwR22Vhkl
GqwD0sYEOlvLAZOF06Kr8c33X7A9n8dugHHA4RGHhozKr+VnzbF2DH6UDl5Zva4FktQub4zQmA/R
eUSXTz3cOVdhpsF+ECze6yyt6Sllur9zAa1PgTIeP2+q8ISklxJz7caln+7rbv6sXjvNIAAltIHi
eWvdxgOcQPIqWxBsPXg/89qFbQmiwC1mPeYc4D+UqWOhDxHmko6Os4SsR7BjTL9R9qSurULm3sCn
E3X3CzuqQ04ZDqQYIGG8vl0wbrIwR6AGZrtrGuQ3bMncPQW+vTq4CW7V7S/Y3hXhtbjhOCb6NIgY
3h9Y1Z2EyGF8y5KfSKAelMhB9gRk4aADwv541xx3Tzj2AtpmMoUnKxZ5+kkJX87Xdxw9NteYWJTT
pJ8zAFota6kzwdF+/dfgG5Z8UGL8qo5j2SwsU8LREfdnh9bz54OB2jzFD8Z/Z4OVGoSHnHKCQXST
/fPN7hPY7kmHwkAoiqa3ViEVTeygzCWYeNNQlyXb2WUlcsHxAJEv0Ct980LKPl38VoN2HMK1F1Ak
qFLzk3QMbIZWFmXxQ55C1LCN7c6nFeKKrEKL2EecVW4+Ld3j03m/kZdZX93Oh7bMhY+w1buSZSlz
6TM1sjRI57uVCOkuHT4qSI1jUvxBBcVyD/9/eYcbi+YSkBV+fxpcAF7opd3+lfxVCXRi5c1Dsk5e
vgIoVB+/hhr+hjK9p6nDpQdrY3XOS6DxFZWESYj4DECJ0cHgPmTKZRXhyh1wPbfF1XsiXeokMgcr
FipU7Zodo3wmDYTRptuyV3q+ZZVUqA+z3+v0pgEOPQLU87X3ig7irR4reYo744Aor//kNnSMR4QI
zoy+beCvOna1cEMxvUU+NSIOGPmdCbg0Xnilv7tHD4VFBi5BzgeWaQknLeozLQSHRuXkwzLJk1SI
wrDcajJok9R6rMPeZjewsKye04BXKnl2gtbXvO3C6v2a2XChc9DNwwH5FXHzpGl3QuUEmkeWn/Yb
OKIrGvipne1kxUEhUdqEmfe1k9fPZ7mMxy0fG7g8vGOXSrbY/O7ekRxwZgxuIkmjFHw3tXdIZHnh
9fE/+RiSSOd2tPpUS5rF4voplOqmG6atPc/sgrpnyOJKwseyRHaY8TB9VkB1UHeDcT/MHf6KTS/t
0QD2IeI95aKieR+q6G2LU2hJL2tPiWme/X5WFuAuT0my2hOi7OFZrqqnhs7aU8IB1tgllwecjb9h
lUaPmB4IjRc+QaUHIqomgf+CXWhdB6jkHmf9nXXTObN7Fb+oNsZXwV2lEebJOQAH5B3ainhtp9wY
T+/fMgnM7pPqPXSvnkZf4diigJbmGE3Vgw+napD5PSrkumysMBtPGUos9Xd41lyp7PXqRZ7i1m5F
M8IIZLTm+0w0jm1joCtqZBtqCkphvOZtfDbFKFE6VA8kYyVVs4J4JIj2Sxbn+EKzkST1EQ7qFLV6
fmGRzO1zzvyrZHKdzZb67SAA4UBIZDpWavU4s9KWfEj6/+stVSsab4DHEooeQdc0dj5U3v7eUi55
FUdDQxqgeRSKpAEu5z1oVpWuf1+g2Ky6oPnX7uVQrHrldBjhcN1MlmsqiieZnKyy763Jo6YE4N9D
0j4d12k753XqYhgB00JnmylgJLqhz5VS1sM4zI+xs2uXJqPGPkPYSyQn6BUbPenCvMH2zKx6DMX/
bz93pJiSecT06Lm/DH6G4Sd8CJCBfrrs169qW3X0PrzeSVvr9aVOEQrE5gSnw1CmZNBvHp6Yt31f
RUUptI4jBkqzEV6rhJQPjN54xw//tsxk3AuBd64tIK0Moyefp44aaFWluJ78FAXYD5ELTLo6GyK+
8GF0dPfA9qBWKYKbis+5EzBwxR4DVIBYtH91h1H8wF0CraMAGgxtQ60+S/CQVdKBi/2JAOVbpV6T
WctiS9U/gJYv6442aIilsHW5A2M0A+xRPmlOIpnhWZb2yACaH9IhzdAL8XwR1DeC+bLC+EePuxIC
dx3v/sSuTRR/iLYkG3Mi6837PcueJpchpjER6y95MCFC74Bzcxg2uhRTN3Zu6jXGqahXbxVU5oBC
WFYmMHG25GF2HsTGhsr+uMxitP2nh5TCrhljscrApXZgnK+2lQO2VCa5xpv9Lkzm0SwSZ4ObhOxP
59v7Xnb27UOKgT4Nb5IUs8H1Lb+p4clgd5U0BYz6rZvNVp8Y3MzcpCkW0rjPkS7CQ41Qg6VZGJg9
s3Tk09VIhdWm/WlU6coTl0M7+lpuQQkINQ48hXa5+YIzsnGwbPzhXqJ428aL+wLx9HvW1KAUcwws
MCvUiBneoVnNdWCSRn62W93WI9CzInjrLjh0VMRxXfeQk865MdZ9SxhKAhDpPot+h4TqzkE7l8lE
DRsfnpKSEpPeBWzum/Tv/LvVtzqqhaQDe/Kg30RQ31miLhT7xW4S43nbMlDjcPdcqGnjuU0rtmUD
bBDB3dbcZoIPzcivfgYWFDbO9OphMt+lE1QsBBrs31pA0vLFqpk63ABhFOvSzD2ft/NA3K9Oy5Np
gBdjWGX7rK8hCuqfxKZtmTy3k6K2RhxuJk898lDY5FtkoWpu/EZUiZPUUm0ov/f4lonJPOBSwsCb
dqFHAksFPrQ434c3EMW/wIMZLLY06JxIHf7BSRSwLkmE7t7aM7Gr/p8D7/yvft5oHZ8t5vgYpiwK
8n28omde5IGvv0kk0KYbPtQa+3q4vG8WOZjY/CHFRTssQTYjXn1xNb48SQvFebRvpZOFwUNBjsi7
98DBexqh3wnXUWPQdRSDQp8FA4d93pcbpk8rYB/3M6cNtSosvKKc/gRm54ASRHBoNAYhgKjj3GaX
vpresDYWVUZC46I8UCtLLBhF8uAmrp0cIK9OeJUwE5gsGSlBCkmWjF0C8x7X8S/ermpBgiMLI3N6
xs1RUsPE+3gSHdU6ZktaK7v1lXrAUo07qoi6uvvgIQwkYgvgh2jm9DtabGO2fcbXYASz0CasTGdj
yPhklrkA9VvagIBe+ezD6D6I0VA0aWUDC8wK1aCjsm6V/AwGizmNhrHgutgolu8KsooSLWLAjKei
iQwYUkKZHiQ2onq1RHRs/FRG1lw+48p+IN+H9ywn30Odu4U4wsZ9R5NLxROdLwQC8Wka8gAxryKK
y2JJCryxHEPZXBimSFMLSd5jFlsEd49g0asRDi2AGcC9iRJYua0SvcsXW/SkF9uAUd7aFLNw7r0I
cFcd9A8Txvcy/i/mMLeYfekOl0Y7xbpYUeF5qxguF7LDj7EColYqnXcEvEMweQIgIqO7utfBGqm5
nRLIJZLoJqGg1b4GKCNbjnVVxHelTom98RLO58/ZTw0lhL4vR3yO2mC0QktVfab2K1o1oQ/uN4KP
u41c/Og668EgnBX/Rts1yWuUcmcm4XYyJnK9RWfxQOZqJljjtNtM+T6fZs63dqf5nL3wVKl+mPaW
OiqJtgkDAxsCXzjf55YrolnK6DJ8M73Zbnfevj1NO46pBPqRy2WupbDVTZqposGwuWDngP58nY3C
sJd5CgXzsxHtUTYMWwlgtZh95BnPmmJs+at9rFIwG33ny3b8hE+2P/BamarKzpmdpSrBrJc8d0gH
pKSpRppl3JHTrJ72cNFXgLcX9fBzkuII/A++vBLLdGeJfwSRyFUTawSRQ0RWdWoIL746vOVWJrn7
242LsufYoycTVGIZhV3wXpBAPyqX55F9LiXiEBZikEXmqkM3NYWiBfVtrZPB39dxhgYZyucp/Qgb
dHiXAdlK+NixBKLp0dxUuW3VnkzCvpRgP6dm2jl5NmKKoOMu6QDgmwk60swjka9Cm2hjeeP8aOqd
RfVznyN+jVuifvP8nFU6lrYDlpNDOTNpQV/S5eRt5Tph5+Qc5olVOwlKnm9XV9+uWPlz0pYJLg7G
f0GhRYYVDzCYxhCO5751AVZwod4COk9Q/KhfVbGgpuTLR66Lc0wrAVO1O9KgjaIDE0QOze3+0NDw
Pa6Gdh8rXpCHEzQe5cckajW14iNGRnL9meY3SOV15b1lce4tAxcIZvhTi2XBdyof9WkVyv2f0mcL
OuOS8Cx0J4zS3yvqLs+inirRZ8HbR5uzhVF5f2AyWF7MWeoid0vedehRshQlxrjmJA5jVZ08/Pie
HwUq4IL2e67SMs5DTQmztdi/iXtNV0mlaYKomGnAV6L85KWnFZA+QDvywnVAdw4oH2i0OXi+HgAv
9aMoHBwUIIH7vW/FQm0nK5R+JN6Xq6hHHdxXTohUdr+hoiBNtypJzBfhNELR6diGOoUKTVLbBsUY
S1zXHq8BAUOQpbVLIkxcG4ON1cfbx/NSg28YRQfc2f2aEtXtHtTIcKASqJjIxyPuKITtsqlT4tgx
hAtB21Za+v8SFrNn8aVf38NrdjtK/TJmT6zNiNP68YC8zo1X3L38B3rovpryzAXyA+jIoNcoqz9N
sE9XfxAJo42eRlFPic2bu0h1qPIHkM5Y6OJtAU30BDNl5uSIb2D8HseD/VPc/LjeGwU0dMp7YmXP
t2MjSVeQZn4VfCZLIKwgT+/rLBnvGNmcb1TYjuw25QGxxzsdxLEOoH6plgGM4cKu2r9RnuW2GOXH
NTbwfDASqFUiaXW3nSmovPdJdT+zxfM9RoyOhnjVxiBrkXDdjsSfInq2M2oEMKvxQb5QMBdVOTYl
DPXh/67cqsAhf3m9d/DcXLOSNptMuBb58Ep4jDOkR0qlvBvFutBIuIQq/GTczLKAnW4ycUPWml0x
+PRmNU60U+sroUjm3TBo+o0oZoexQjcBv5G595VIA5qqLCZp57oL+XGZfPYVwccKR9Hq8CjZzNiX
M3w1HU/5QKmK8/tXzTDcHbK4a8twLdCZh7+38FDTX7sKwVRJJvopO9ZUp9Ffk9VpCKtrRpLJcojD
66DOMXGQQ5VrC8DmnCfkA/4gcEJWtkuu+ek525m7Xm1WzwrUplqC96YqMoTR5tSgleyIACf1YlDf
ngXXazc3NpmMx01USkXGp9bTDxNIzV9RlR05vm/LSkxILmZvSA/G9FkyIWzk0rSTGjTsGRZ8yStc
3FS1VFVWwIHd2t8zxdl+aBz7OKkVbkBkk0V5Cy9HXnmqNo3Q0pO3dVumpuTM4kcDU/zh4xI/1RVH
6uvUPkRR5X1eY1kB2pN99b8gtaeGgbeveg+ObX7MLCUCtyZgXnb46MS25UdL9gFFrz83hR0McyeZ
ByAxP2onaHZo1aP0f+pv6hDVJW/3tvEFXaSzLwkQXKb0wg3jAuvwCaDGQT//dYtdRTw2h8lMiCYY
sUHKutMeTr2QK+cQk2oF3CS5FkHZR7uOSNyKti/U3hEGv8qqMHXvGYLsDghJBpYh6klH8TgT1n7B
4SVRADKms2KAs9EHfO0gtYpk3nvJhCm47Z7Hfh/CnCcxGoN+rL09NBNWdIaTbsO0Pea0Umo7GT+J
IZzm4YAUfy5Xt2kF7nDgmO5blZDdO+ZOJbvKsbEWM994/DrhjMGFLGAoTto5R9xlTn8ZopcEep8U
68iq1I62WTQJ/Lpa8msyW3Bz+83UpjrTjsDlTB94eU/OLrVWRcjCouIh3IpyO4JiZWnTdkhPe1PI
UO7+NapoTlQX+zUveyO6S2fj34cuPn3gIiGiqt96olxhmhuh4m7ZsSxUshXtTLzwK6NJdPQITEVS
JALZSXnHZFsLhjrdRGF851L0TieHOPgY3l6YIa9ithj7GRJLYffegT37FFJXVlcpZIudy7OvPmnH
kuklUm6ZmR6P9uRWf2iTmDp/SZE7k0OBDIBex+mOw/LV+InTwq/is0nAW7YovbQthEtNweP3X1Zh
WEhRX536qc4TMxjuwcGuSytFedh1QtSwaXdRNgVugRGG7usfNAzl+J2Y6e93NA4KKVx7rpLaj0zb
z/0ERAKXplcwag8O/+5ACZ9H6+1T9wVkRQpn+qGkmfaASwb1AYTpDQ9BZmHBvH1/ho083B2oHFlh
yOOoBrM1hsHePEZ1pk/XsX3oYsxORX+VFK8HHhn5VMM0zykyFFAILJ0mLtjbknq9AD6xeb9rb7qw
JBv/7EJ49gmJDm8rdLDvU0tu2J6VZk5hOr3YVGh4R2zL3uysYDDupdNHA6XHT4Bem0CJXVRleK15
Ya2A+14REWxQaTfpdnHP57Qw9SKvnBQyZhswX5ZIWP7IJjut1gbknZYrfUNtnBvGbgyMnyEgzkar
a9o8b85JjgZa2FSyWhhzY35OEGEWYXKftv7/8SmpiQ9b2IosLHQGqM5XfOHsB/eGrMOVvQ3qUCOn
ueGw+qf/pMKz4xTuFrGS+zvE1BkGQY8k2NtyPo9db4tyix/26pm0SAm+QWYL1QL1R115WbxMLyK0
8qaYSIaD2RQ2RVdBKewqzBr/hcUVLHLR+lwnz/s2YcG701CmmLCdVZy9U1O8/Y9LihYPFVKLhN2+
JoWxcrEUuX6iDc2fJoYCdWSQMYwerK1AOXsKgz8G4EucVlcRdB3FpeQ4hXcF+XHlswGVqw2c++uC
DWk3wOlFTpvEc2Smw6hMIyotETBwd1wCDsNXDrZY3SYeg6hRPz/KnrS/GrSIErdDnxpRq2br5O5n
JOlXZmPgDt2yMd6ousHuCSpRobGl0e1fSdX01nBD5DWsawFZY/dx/JM3C0DKMAhqEXHFDq1qvtZ8
ItaaKfvGKNKqE2Uup3HJb7nSZcmXjenH2XMxSMK6jx6NiP//c9sFeK5B3EN1riRSVWinyx+7FG2G
7gKiiajrJr80m+jSBnxnrDvrab5Sy9TqLHkb5E5r9h94QORrK2kgs69yLhNcYng8cR6y3Lv5hx5p
PcbXrFaTXL+am0FcFtdqVv1pVGkFk8eg7CkTJlwiQlS4Tgcd+DSXFrI1CTe3E3x3VCLaesy6zVlr
82eAYlVPFOdFESC0uwmDFOKhxy9YcFcLy8VSgVJRJJbHMUNSpWmsYYIaXNvmhSNAY38MN9JEveuS
r5gHhdwEAhqpOW5gNotFxRCGVG9XyskU2wRDRuqZC4Mgo2bfJN9TdzRYx4ilmcbAmsvgSMd7y5a4
jn3Knh9S8fnyj2sx4i0J+2dc2eAUHvLTfAAXXIYZBsynNbJOtXMrGzodOtcf3+Fffruk2sOxt1GK
sMZbySgYpofexAlYOqKYxPm0t72OtwETEJ1SN5r2zNkMBeK+4rJzE+hDmSmCNKGMGthDTiPwFL3Z
n6+gzQ0uoMu+3pQSsItCeaT4ujARd0iobLwV/SEbmR7ufvTTuw4sPtYbrGnp9aZKEa9aLOKcCccO
f6EARHESchPb85iNNtFE8dK98XzNyXZmhS1YipmxRDJjTff6YxGF66l/YhEFFU08YReKYk9tZMRa
OB0WdU5fP12y/anWRbRJkALwpv4+Bevk4+taS2bAuEBRHRx3hDnTEF8a0q8fn9p3IL3dZqtAnlHO
mgfVo+03D8RGizJDnifKWeR4HEpD9DeZLReQuohrepuP4/v0EmeRdhHgFfNOUU3zm03+0Qdn8knq
m9u4GJUocmigqU58v1JzDKXr5RM7jblzZZv+LWKv/mC23L2c9yKYDNJRUrBEWWjTXpJmPlo2UxLm
KWDAqAj2aeWLKOJQlm6kEgXEaNg+tS7C3jl32wGRB8Q+lyzRPNYP44ql9JgkMnUTBBPIlNatmuhJ
mAqixd9ux2SJQEEaJ6kdDmHHPgMHq/7sFwpK4hpsMuT/CR4MqGAlGzulpDF1iYJS16ntgmKj8Y1k
e7rUGX0/KlkQdGQdBq9TAQANlegVFj5psT746LLMZE3OqjAWlXQ+rShEaIUU016E6iPenXDZdph5
gFVtYAEYPX2FXJa2GS3tcMXXKox4CH7LwklJ5T04bOK7V/ObyAiPKsImb8k7mojFP/zZyjl4CNoV
ya6stoT/BQECrEzk/JpkQrjurb7znFvJBlpGqWh1TVqEvmUXiEgKYqVz1U/ka1LlDUqK9ThdJQkw
sy5iN73uRqQk7UyszWgaqzYDGmFcywkxh2oMDskoFKX0RPfA1ELVTT2+kcBBe4VIGSPjCm3doyW1
vrzrZaPBXSy7ifzY+rbJsrXVifCWfMvEvhv0fJbzK1JyGJ5IKUw4syvse1a1GBewp+f1Bhl0ChWn
UUICXnwPkLiXwn9cV2zlwLxKN8KjSY1A5CmhMVnMzf+hluWM4a26aAdtYkLwwx0dgn/bSrmKQZ1O
k/Dyc2bbT7RIzYlMbh6GQfz5WEv/c3cuPpmXvBh9rk1QIpFrZX+MOBwYEi41UFdemocREtk7a4d/
AjK4/AV4WsAmS0NntfNzTbJe18cyC397lzr5fiB+JFUiSp3K1yi7lt+RaXC01bwSZ3WehsKoBRAd
e8qeR9F9SL2Qzl4zj8j3S8MO1IkHddr8AHGFylpgcyx0Ps1Lv/gKex1+mtXWoSZhpzFNwyYOBIQC
FvhrdeKmk4o+8g4rGeyxqLtwQ2bvpAGjNCowYxYom6XI0I0gIf8h7CryYF3nb9MpvxzaDB2CWhC0
sjSLAZPfYbMTyOoJJfmRJBxQIOI7jjimWTramlDKssYqSCzSsb+4qYVDSvUCWy4poukeu69AcjnS
AJu41gxGC6iDhTgpnoZwbxY/osz9ZcrxO0W0ruo5zFTykrSxf8mkPK9UJ/WpVpg/PH+aaGliqQFO
xY4Gtb9QOMJQRIAadCIn1pz/sYA+8CyuDMuWIYI3eGUDISjsPPJ4R0CxYjnWywdnBDprwCo7iKGI
nK7HTZFn1ko0d5yqaJj5678j1SxKa0PmzM+gCkHSYm70S2Hx+Y/BR1w8w9Fh57krps/1F4XhfvXt
F5tUKoxIZcXiynIz+yjYr+nhR6PulfaxwwQvDweLTiuQQbmLEfNSvtTBm64/j3PzxP4ZTMzCFcCp
A1XH5oCMk3XkrgtszZekjuM70nV4MW4evKIYF4rnf6OCt1mkMh5ep9E4Uu5M57UmkFYcv07eI54s
VW0AMOpJyEnlNfiLeQTzJ/21rJWqxEOo7VWvvJKzbhURQcJvpYB41ZpJ/38dQigx2Ikcacza3za6
ivAtagPQ1WpbZByWr7/Rg7QmzsFUrgSrpTmam2lKrp5N/Oh5MJKYydr0lG3VJbCGWvmsZ7UxmWG1
179ZPhK1PUGItOaSsFo93MCnTO0rXOWoltcAPOBy1udoanpygLFnIbcYRfyv1RVLLdBt02IU21hg
atKNU+JtloenZaLNcnklP9MgSkU9oWW+v3CTI/XfIUM/rEPC326ccB4D+G0sOCxC2R1tahJYUK0K
u/hF8wjA8+eYwm5rtWiJFnuapj0Sls5rn0CQIl95ZGZMFtDqIRqU7dW5sBIRTE/bZnP2YCsK/5rb
jX2GK3+Ccn4tFH5M1VpAV6hT4JQUtWjHCuAg6GX4vP5RDBJN2as0OhAD+hJN/J5kcsFCnKCtnlbb
dnBAgAikZPuLOfXzykXdJHTxDfoy4offRYSi9VGvKYjLqUzE/mu/M0AqmllltJzzKX+rI0a+kmm4
Otox/lcuK9QoKpn955qL0Gqc40HVqdVqL6kf+ygJR0zO3Vp3fohg/tMkE1VTs7yd1rcd1hwYOIgI
jo/djorpebRHZnJ9TYJ1PiNejr41ynhqP5bZh3Aq3kJapINsrl/Pow/ZJH0PTfCzcO+x4X/tBBrn
tCWRgXBm0X4rI4ewtcHKV9pdTK61upsvn8pwYkix+WANzMbX02+3hl4dIIwlkgFkxirDEKrYsaTf
QdZ1ItM06A2EPA3V/ZHxTrQX32zstF6hQ8swNgCq2mVJyF3FNrY5RYWLdSteTwHcAX2gmNDtIiMV
jcZMW0BIi17LeSGwI8zr9GUCgaFYe1MaX3uPU+yUHoxjpYmcEH3VUvFLBkQMM8TuAetyuvfgXDZ7
SAZgAZIbcErisgrC/wHDGsrUnzlgqIydAdfdtu58VUkkEjs4+YvnK3d1LnDUzdCJA4zCDTTy8JdC
gkg3+yeFeG7BqZsw+uX/GLD6mcb4Y5E4cIhcxG3jX5qwe6MUlluUYVeW7MBxfXJXir0xeTwT/skJ
cL71WKFyLMEtFZnBvFFP6hqhz62DtmJzrRW1TiMSn37uNwBZ2+AfWQZ+M3j8ys56CwpxEfbizuDv
nzgsezdj2pQMlmRLHVSrqtoYZfSBn9qIbUYE9qV7arohv4u+qqa6AeK7NXiFFwWbFpxZyTrySpq2
5xeMvcrOrvkSjP1xqHPw+F6enCI1ldGq+9FPqO86N0OhtgyauD+m4CYPCziU13qDJeMy2jYK1fBj
hsjgKSeS4T2ZWj2uLZsITl/B5xouipC052314XQL6CUPW18dfmsZlHRA2iSwK1uYZ3EDCdTP5F5k
z6kYGjk3iNsiZdiaQxntgH4SUR6r63AZe6r4U1zzNUG+aqyJdf168gu/G6dscDWQTwI0kYtKH9e+
VMtY8d0rHmGtuF1/mZ11Nt/2oF2kZBWnHJb8ozMOBM9SI0FiL8vlTNhc/wVNnJHB+0EvvyL25yvu
SdUwn3K6q8Mk9klIqqhtngO3sGgXnNzvwZJ0TJaBwnr1M6uDLIVnQkjQAI59mt52D5lGdKosFLE8
7Mwb8PKf/onJX6TFY8MtSKUfZ9VUObtKxVG78d7URJT9AciOlMb/sHIRVfAqovNHreakME2T1oEY
KowcnaJkhRI39486BUCbSJ9WZcoSTppSicZvB1HV/QKFZq1TJr3OQIBrdenahhQg2vnm1pie++oT
Mc4X7FP+omB1vZPqzrNQUHg/HPYL2Cw+KjMI2tRc4Ef+UA6xeAf1A58kiqRMQGtvKmjKid6TLyrN
SB4mRxMm6lRJ6O/FDzyE8b8TGZO0865edaZD+TF4e4MRDqT3Ow8vvctGeiUeOEcLHtVCGDuJo+AO
XRG3y28gqVJ9f6gRT1RKYz9ak5dtLma5Y/gkaqyTbl4oiOBeYor3akjIjmUytqHvG4p2zhHBUyMd
QBBpECn0tSxjOJlpRESydq/n8cPjSUQyHdHJJmEJX5uHfou/HYzJOZyC9wJAGg602xhWVLwb6aAU
N7qZCmQYRqvd7+HLfBiezizIH5vb9C2/z7Na32+GG62Wf/EJ19QyLOzBpxMt4zBx8mXpL0UKvxFJ
PEgYU1ip45iESVigIVeMEc5DUpXayafZCdNCEHuKI94NLxPI/I3PEEsWhliN3fOeul1qm79nMBdQ
uQdDSydpzTLHY0sO0DGngsKB8iwTGT+7bEHri5JLAXGPcxyRvZyMbFTkTg5cXYLbykkPo5ah5atB
pEhWDxxGQYdXVRyCPjbUpX4fAQxAwtkHRauA+v690iUiX7n7frgal0GhPMjUGMKuJurV399n+E7N
ahjsxloVOq5u/J7g1T4LjDsV61ttRtR5VuHtJ6fo78nEZtVMeEecSSRlIwAy6JHojrlwWifCkF2m
cVmtsK8CQUARJCNk+k3dORsq1HgURBuDDEmGOZCC9y2rfmq/plEyHz1HQi8hcat35BcopZBbv5ar
vpkpaonscnMep2aBpGqBX2+h3GpAYpKEQth6K40AarMsJBQFzEJIHmt/aan7lEpNiG8IL32iIuMv
OgsKpDRP90VmkwNtNvQ6sM6IOYOfBtgrtyhRyWN8QmAOFBbcpAoJNEiXdHfd49hbuYla9EUxOJE7
biK3HJo/6i2vXvTECozJPk8oHRJaIIueAWEQ6V8WW+UfdDUcWAQAoF0jAaf7eZpgG04LaXRYAPZv
4uc5Swu5JqRyuMpkyTvgh6MEX7PMkU9suHnzFw2NboXyW027gMhMjqW0CLf9OBXrBDFilhN/njYL
lNY+qYzYggNMmGLEXV6KrJDNnRXthibM1g0T+17eX10V7ZZRiQgCOUl3PH+XGhdza3ef+Z7YyIbQ
vzk/jpUi7SSw5kCeLBzfmLiWv1S1RDUmISzheJG3/RRD8cnJetU7Cdnp20Zxq8pCC7ssQ0/81nQs
76g+Fon7LvlA/Oi1RkCxhXOqJ68u5Y/cQ7JuQa1eIhA+WhZ5irXvOuftlNBOVaZUSbFi2D/Ga6F9
+jEKnfbPbHo4i6wuJfedCxpe9vOTI1c2mzQLFUzyI2qHCweZ7jeaunsm2X8o/cpdsk0mxJ41mMQ4
Ooms6dVmuimFrHwQ1RdzxHFCwbxnImnjiZS/DocLaS0iNoJprWPMaBLf4LWkZ35+VWVwX67J0U0u
NDBIgdKpbj457X9KDxVrrr/TMQGWLFsgme7gYiJObwJNwgI+drsN0SfB7lrISdKBg+6wkrTyfdcO
dVCKjU03kmCnuRzTKOHDbXn4pVAZ65Gm2epb4xDqCcKUbG4Gx9rRoavch1T9PpiUAW9FbRFQ5FN+
DdkVCS2Aejp1K61c7mCTYGMCYdSkTdkJfFkHB6JJ97bVMnUDzxQKvESQ2bK6DGU+dKbDkKKj4fX3
3AJaqnWmJEReRv4eDPLOJMeA98hcgl18vVhLBk3RePsLVD314IPp0+5qdsE0uz0qErBRO8MVhKFN
YQqwNoDZHh+22MlCl+5bJ5B4T29beg3aSmXs9bgLFPt6gKFf4IvwCX02V7D9SJp/vBpSWo0/U81g
QxtdbLiGr4iVQrirMSN3s9gyYxV4FFQx0ks++6iOhSvHo2ogTSPf5TXlDslvkWJtEqmU0rgMAchu
EM3bqsxEUsjSyh8d51UZ2kcijwjPZU0vut/4sWVj3UZYSxtPomNXrkB3rtBfdTrFgVlZ57cWTGnj
23QOOi7AID7e/VA2GMuh7BSJsv7QGBtMqZgA/4xZWTaS7mZF0WI78BhxxV7wexxXa+zgfwWGM/+5
NZwTQIEvyJhwlYmLMTDUqylcoMlCchfdpBUI+j5ZTxe4kVNpd9Kz0pcIEG6YwnVzRh8Ww26i3SO8
1wEwPOnZtiEKWq78Rp+i7ky6ArCG2XdeV0rbRVnPiMpYfxTXivKiqR5I/EKDmKXckfCV6f0GuZYG
6wAL08yX+c7wQIHgMclAD4jZX/6AViHtvPEhRlMSjhNpnKclfFDv4vGJIZ8/LgMY61pdfRmmTgM9
cyiAHfIEmdgG/cBXYwiUM5nx73kL3B9Y9GJKIt7ibYbSROLk9cP4B3mApW4Hbrk/9MokdokFaoRT
poDyGUGaZEHzhBNaVW+JStQvpvvATJF5GYKTy9Oapl7I7AKk5yNuJ3uXNy7GKayAh3Y5IBIAmhRS
Gig7DJauhAbbhjwVy+1VmutjwL8jipWwFfjuHXDTB/jWgducCjaIZoDJaJHWpLtuyDZBu5GgYYCN
U3lk7VxaTbOzAk2K76qGUj+jeuai36E9Kto/5TkRL4DWeupBnRwKTdK+v7net2Y5FUcZsT3liobx
zLzHYX1vnCrSz5jeI6dJUhwAjl1nK/pD11HAmp8HDWZjeZGfaC+fEA2OAppvyblruXG2lmWy9/H/
hfG3Zj4TYvgd641tYBvR6DJ6cIU5UxH4UbjBizajfgZqrYiU7yegYJvuiYwU6KOhmEzAr2AQzPqz
ruGHiJTpMAoQ3ioSrW0QrQKYXmSfTDEGGAu1cZaIw6yZUb8ONed5Dedlwf6Nt1cHVrsVsfC84FDw
VmB3zKIMu4NHhl5FYuq9SJ8oGXuzUdpKXW5LyRFGjKO0jLl00pO6jSpZaSbdJflmtV3xg44EsrFq
x/uB669WS1Q4Bq1KAaqDFpzM5F3B1d+KZ9fgnSKku5InqrtQEnbXjn7axHsqzsJKKu0M6BrOOq9Y
ES//1GcPWfWUpk+J+DTpLQKJ/Sj1Rd5qpHz+u3NIo/nVXsj/yf+CE2CIhI/XlTDVUygxZYSP13bz
od2pZB22YYnDnmV+lAl1Yz/4y5XvgZyJF10YnWNHOfRALTBjz0rjcaJ49Zh8FCOserES+gNYSpcL
R/x7A86QUmePuBjJAmM7Po3J12eRX5BuRoLcKf9XZkM5ehCpi0sBLPnnb+eVnajSnHTE0PxDH1ut
9SdzGY6fqvFv/jJmJ8VZynlNmRkoiGkWyXlfzazdiEaeU/338q2c8m+7LTT1dfW3XD552KNWIlDK
+pQ98JdMGlEPJrLEMNYLqsE37EEV8hLU+joLERz1pEWBLMZGf205c4zaYVfJd5fIwbxPjH+iTv6H
lSzflvwBP1Ts2xnCOxdrgqaDwE9Rkih4H+NSoToP4hi1HhqhXfgfGr54C6aU6tLns1FfUmoCgYzH
1DqaFI6+yI73OnUPj5mONbmvlgOgO0+2lyfaDI9XSl0fI13LkXkfBlrmJ3jYtnG1I9etY2Y0lSTn
y1zheSSS4KJ/aRLaUQ/6qTBsOpGJvP00ZVIxxzHaeLMuyMzZQ27QJS/W1KdqzmriufjpmPqRe7uB
bFssFnU/QfNAu1f7mYilHwABx1H1iqkQCk14mV5h7qkuMko7hThI2OOuZRghvZqwhzq2otf4/uel
yccg5JWY8ozqcxv9kQRH7yqWNdMg3rrs2SIB/cssKUp5JJOKNXKKY1a/y9vQ1cw0JNEz70ySjn6j
jyY2JFhSDsT9DO5CkHvxTH0/Qpv3qDwOtug3Z/P98wj74FdRzTirhwQEXJDsHG9IjiNsj7wPoUca
nULxZcDiiH3NeOJqyVfFA3eKilTJ6EZ8UpbU8uWgFRFkw5qjHXHos5leTaXQW6IgnVypF2jVdSGH
E7X2BHgXKKA4rGFhMyos8shbMQRBl7+dNdJGhqYZ1CaLHO3VRa3fHiMJEfTjA6aYsDrfTPGDBiuD
uN4QbCUT3yCv8Py78VSRRkD8IQdQz+IsPpC9cO2TMZ3KzbFRf5Mwx1Fmai9t3J0dobt+lmXp5bLT
6QeaASy0LRpL5fsomQyLdDGExfWdUO3kpZn5W+mdDp38L5RIMRulo1ftpZn3VW1JaC3eYTkrN3QE
Gs14b7S1AqkL/oRo9FOTi/vagRXy1/II7ldaa1840wvOvVbYD+DhIS+ZJOXOmNT7uhgcqqS+CsqI
bIeI9oOHu1B5Pu12IXKCE5FNyH+Qtl9Pglzp8i3OJInI3wRRUnMf/+pNsCVNXLSA6Kj3x6wCjeNO
3LxyzwK2jYlZ992X3WGd18CgWRF6Oo8pmiE0jRR/pjsdU7lUOhwhn17T0Ouk2/dIllzsAxg2gLTf
zC+DVr8tV9L6FeE2NqVwmEnYOqMldOxEZL2y1uLcaNy7kdTKB2BLBjQf+duZFa5tk7somc5D4DFQ
rebaQrIPHHYnFM8+vQVwuEV55181uzKBO8PpLFSUFW1NhZV4140dOD9tX5hfCcVXojkA1pw66bTF
k6zMxl0vxBgD2zFwHkjpbNYi1q/2yTwYY2ML8+hxDpJB3b9HP61Rf8maMtaE4aJmZP6519cjUlnN
TZguHIku1OhqLwNMfB5QrWOwR738dom9H6Bm/S25vSJsGNPfx+Dxj8SCmnUyBFQt5cmkgxhatLeg
O1aBXhM6OOQmcHFQBJ4XgpMmgG1ecOZC730+fs0KRtd/WtHHtnr82bfy9v2nCKa+H/7yKe+RXX/O
03zYPDd4Pc5cpRKKWEawMQmEjZDcDoa7iPgv8ytXXPwlmJD5L7uEQVVTU6VVM0Yupein3b/GO1G8
6o7ZdFEXrTSG+wf1XQl8mXHOQrURldc8GzU9PxUo0Am2o/xJouqxmd2HbLIwrkmSHXKC5HABsKw2
zKu2pYJA69f0iGBcfOYTMKWMMC1O63Te+s73XRAY1UK4KtXL11FAGQH5xKcvp7QBAMbbaw0nzV2U
wwnNTeL/BR+9a8Jk0h8RXeH5jp2x7D9kmWUhVp83q9Gpgzz1/B/Dm6eb3/vdG7ks9p+fufe+YiBi
1dgnbzPepmJo+Cgv8v6TuLLdtijAxtOj15AD6wx88PANXvZzAu5bWOPnxNyLsSOy34eXvis0Zihp
dIsX1didKvUm030HMVDLGckcgmJago9IatZuBKe53BIzRL+4HcIUXGZ8MQDlP77tcsrhzCv+xjs7
zahPYY7HEI5OWsciDXRM6BiuoO8gK2ktglp+3ry3RgV+JUJwiXnY+MQ5b588sYHUe2H69uyGnipg
IV2E+jvhvxYmZltHxSf6WOSE6o66nQROuTRgm+fWuvqVsTQhSRExtM7lTXsygnSXt9Bk+/QhahWd
clvK0jEsxtir5JS+ZQDZFGRIGHDfRs9kiD2nDyuAlVQnu892TGbjX3xIOR743iJeSTqs9iW97rzE
PGzZTggRlZT1QLKAnaeQ2Y0OzMQozkB674+Bjs23yVY5gQOQfM9PeNmdNYqp4Y8HMBKtzIxPV5qF
AncUdV8CD2h/rLEGoch6w4LYwjY3amAydWVCSdnW4f2gbvpmypacEMRRLToXNzCUlYU78JadXVLr
e+M1gdK7p1cz9+ImRQiosIpub0SwJtQdu8uhm2ac6lEGtf7E9B+J5T0wAWIoegzQ5spy02x7zZo1
9gXx9Y8ming5f3mE0GpRxcG+HDAw1bod01/huWkbBOj8sQYccvh+VwAQlHfNGMVPXwhrc8xBuBt4
mbobEJN72/A9WviOV5bUdCiSfHKHnJY7CI17p937Rpi22DTPThbkD6GBG+2PGaAnDHvey3VdeSdk
mFndfgvxFPjrSo//FbI/W0lN8NNsNajgRUbz4AUeeBR00BzArLMzZ8b7ydsCaozs2aYyal8NiUSc
Rq2zp8HjOgrZ1uvwVfBsOsA71g4ByHC2csiXSbXlhx8I//+GGrYr0lc/+6T+TL8gvndokoFq2Cno
9Rl3mXi4EChgeODwd++7Xc1QW69Y5Qn93kLAxI+R0oP5GcismXl5nclIhUg+/5MF7+hKTKTJxLkO
4wYrnQ97lGQlIc2xS87ZSY83JfNuMWxJXgkJDKDbyTPVVXCgmNy+IEQRPV8IdO4eFGDR55I1MQGY
laUggWc5E1i6fq0SVf/HrwTsFsOAq/SvxJSU3SXe5E+VEtJ3ZG9KWXQQ8X7yoqhTLEoXpObUpFfX
xj4ikp4UnJN+qQxAAgT9ouTXkrPz/GTpkQaIY1VGJzxoqpDEEL1/7l6tKy5Yb74CpgS397BlaWeS
Mpgi5agAYkSI0YzYVNyilVSWZBvCv1hC+unUpi+tt91H689But8yuyMiHGjvyka+fUgb1zstarhd
VW+bpkPT7Q6DByVjwvi8psi4fNQMJdZGtS9dCau7c3L6InbbYGTDxrpV6uORKWom/R1okcDjsziF
RnwutmDgp37kdAqxLThFj0yP1A6jCZ37oF/1yvKH4rz4YcQDGKv6TUMO7V2OwtIdlMH1lznPWbFs
ya5+L0wpfbcaguoJax4I0M3gIlRje8tIjFPh3ezdKiK4S+H9LYdnanNaBwxqjkCjm0/BiE3hE1Pm
f/4WQFbtg/mbyWOhvNpgJykzoptDdGqQf3zY1DS3cU6T90GDrV62s5A97Y5P1Dj37t/6IsiGrJ0F
bhdQFbwaBzvfKJCGpoRY3ctkhMKWzIOF4T12XTrPak2ruuxqMksizDThhVfq80FbYmEvhmPKvimi
b7tNHYmW7hYfs16/B/2piI/BEVLOL3fZYSNR+eaZhFc/zI5s1MKWRGfnaJ+RzuSsvHPLJ6udEfrn
3ph7h0i9oans9Gub87mi/xwndvl4B2lTbL+dYuFxER6KvvmUWD+OICeRGA7frD2RQ1wlxcWLT3tC
eRwwXV5QSpqsWTf5H/rEcH+UbEy3M02yy6WWdcH9wu1UBLqVsqblQT1RFGyC8aWIH5oWTvNl5UBn
ZWrCH2qHdiGzy4gtIF2jDrEm0kZq9Qt7m43bzZzR5KNn4ll4uuP8VsBokGSBWj63URKi/MkTJNiF
kwMEXqZZT/39TiliIPY+kycZs/+79sP1/koI1eniQnAHKHmn1ICXZxsydL0NSTB8rXgCo2mp6jz4
FqPR04w4B+S2fTA7ZwAZDSTmRk68EHFvo7+i3ltfb1aLT4zPWWeIYOGRI2uN2rkFuA1t/Dg1nd4n
dgqflcOM7HfVUrlFJJtr/xH4R/1l297rOtGSICLIZbfal46GmN9/LroraWD+X7Ld3dtP3byg6fPz
uY03HV+ypujftpSCB27ADwkcR3RcudrZ9wKpW1jMGZDpFoCdKZSJdTL8C/U8BYoFvoxtVbZji4JB
JqxWvDqgKS4SrRZJdCp544zMZAQunVjw/zBv0E8OqTdQdbquNh3VBHexG4I0c84HE8SY02o3ahd4
CelbW1yrlSD/LekgroUzy86v2vJy67B1O/0HwqAek3Joeo6JQpcJxhkngmeQVX6k7ywCzSLOJx74
Gd+1iY+L059w5qCC5bmCTxIdrcHkmqRkVQSI/ONhuG0SFIT9gaWmKpoqmcyLa9AK6M5Ny7CSDYBS
7guVNsGx6vB1bmlDu3zCf9OTzgiIsZDxKml3cakW5SWAj2PyWDMrV0vUnz59rYI+f1nkyLQ95sxR
LlV3/M0UApkKbr+O5ZjjsQF/7CQ3xt7PB7JcBCUku36rJxstCyXmzudWfZfqKymN4BvZllmpMDTl
IbtNOuz7Ew2ZN2nP+gWwTu6KQwf7utB/6itNzGVf5Z6qO4sigoAMWIX/LwBxkQeKJw9JUned6pvu
P+u9OSlMJ/iytG8LIPdDla66R1PvHxys8Hjd6SSkFLtXnwTbfYFzNBB1DrwJP6olSdiEa6EbZPSa
gVmNISWmuQ0hjA0Esr1j4iOROOv11upNU9CcE+MtW+2Cg0DsR77tHesyXir1u+5z3U1WyjT6suk/
Ex/VWJyXA3gWchNPfNRUxbX+GG6646Acp0urYbr/hMjOin3ppv/bUAFM+xo1QpDr2L4l3s+qioDn
q22TPNGgmuQXFkhyxRZcnyzzBGffpbIG+S0uKqrt45hMbxo1m8MLjnO3N0s9LOR+mxaFOknl6elZ
mqTUdkFbldAaus2xXOH09dE6e3haSaVqSShTlbHT+t52US4E8t2LtHcNC+Kir/nT0eVt+DO8AuMM
/1Zed3757aSyO5qrQU46w9pf6+tJaVnfzu5vlqy4ouOAJ8qg0AY3xmzG8mvUH/q0hdlh60rrrSI0
Fnwyr6D1f7BYDm4CLMGmnhvG5FB6Z2/UwS6dMe16nb8nRAXJJCKp5SpaNCjcjnNEZPj0kHODrc5g
MFjjq6CAcuZ2wCrVyR3TKDyJF7T89d7IRyHPbRzDCIIAzTFxgKC2ke2hqD8oiji4EQAihYBKci85
rwf87q7HNh/XbyrVue7Z3VL1qv0/I7L7g+++KKPI+LpzuYm/1o7O00MMUScWeirI3ShMVwuWk0qk
xowaiLcKiq9ULrLhFNf7B90N+YHUfpEWefbz2oKu98AnJ+aPbJ8lGjtVeyB61nfWNsv7ES+O3yGR
eN28l3P8wy9m5xrePGK0HGZwXK9Fg2ZFCQfakCAq+f9+8rR/3gO+XHIeYc6y6Gyc8i19nerXRdxC
z/38RcvII7by4V9D35iLcMRWSP+udfvnPMl/RZ/nfmknWsuQAV0qell7tktljfa2DgtGucZizvlK
y+4IBtt+d8Fu8ESycOozVGgcTozbmxGDOGKoSGPxB2F/obJo10ZHvSiU1iSdoB1xBNPFKdE4/+2f
mTzkvXIE5JxLwoDCwb1KA2CqrC3LivA1hCDOI3m/pzUgl7fTg0RhGRpogTf0KZ3ZO5UmMi1MASA6
L/TTqSB/5J3/5HjNtwLcli+XF6NgQz5dVBYxJeLvHVmJBZ7ZX0z20sTcS44zimm9UGuFPYTHy6PS
w/myCEVUCnSeeRaReChh11DNoaXAbPTnD5p5IzSDBtzf2gtZgJnxvHAAnuvae66pIh64XAPBYr0u
uCThNITHaRtNyDkiRTZagoJ+qlkwsnAs/8dXTPhGY8YI5X2asKJhF8RwstoWnwKPxbyqp98Fl9W4
6NF3600OuL3P7tC06sr/3llR+Eh+/CFN9Nl+dyurIGhzuUBG9WrEvACnUc3G0eBTxDewqBTNhQY2
NZ47kA60qfBHnfyu6kzQ38hYCvs0NR1uDD9r7bGI8bLlYGy7JrYXQY1XlXhUUS8EgRn5nB7MBEmy
YSlJpQeSRG1jHp1SlRLPbrXV3iai92fsPtTNiv+0lpCBeg/kN7v3Wu4QJvQIxlDRoH7fNWTreBs+
8jtjfID5wRAzyDhPnjhKOcdV4r55+Wgw80LYpANus8SIVwqGJ1reO4ojXWJKs1ZlUFyhz/Xe9wLp
GzRqJTf/2GBR/peEM5G5z9hAQHE2F2zn0fV5lqRLPcCD5k9m5m9mrKeb9eOze38jCBMinMabFpGr
tWHN3nlbaHEeRuWs32Y6kSZraVICLl20VEO3q3oGJrvUK22Gexyd9KuWjDG4SJKbgIPysu6PI7aA
wlEsCHZ1jdeHeqsw1iA4IJGQ9JPMTrR1WoddgjpeOnGhuPTQd5sQCF6yEITLkuRUXw5GVydmCn5m
53RpV0G3ShU/XTyAUO9cn/IpD4/s3wMjaM3LP9UqNypY2KdD7bFPTr9tB5/kuO8u5WqBTL3GWPPl
DIob2en9UN57X1G0nZ8ARQ+vs/N0hZrHGkBYsLpHfzcfhzA7RyrCwbcyKv0NlgyrMsMzIeObkzBP
ve31YM9L3qSXl6m0iYsDjZTeXF6Cj9pVA7Yjp1iX1Yn/Pd2Brw216eMcmjek7/85wNySXTqo07cu
4niwvfbyMAM2cObfYGuZ0aD3WebUNeikqmnpcajdQG/sR2Mbsd5+QELu1Lb9ajCymfHVIaNsW+aT
YcJXAl2I2DYUTohwVBiAwD1+E2dpXKx3eXBJz2zhhkbvNrGpPjHxV3HsoTTi8ftURMVty/0ndwlC
m4cSPZs9WHgaqGhv7Qywue4kUh0uLrbU3tNukj/HQnuCystPhCuZCjkjT0vJGbh9gsbNqx9qweoQ
rkpWokRcEUBXn35Qi5tBZu47eijAhT+qbik1J4c9QFuj/HWIRbow+wx0KC98yZryEUg+4QmdWuXg
k2kDGTR37uUG1UZ57u5cqQhkRwqyTsXp/7Ik28IUp9SQFYEkMwvs5GkN39uN/Wb9bfLJCXDbd0BL
X6IShaxRCxFD9Cywh6zEAwqU6S9MRq3no6AeOfrEryph49VvTRkb/FWPUFlWB1m7FElJv0t7Ua5t
9E5iZaVaJTAaiIDmnvE+OR+v7tWFzhFfnbvF6QnBGyKPTuooUyF1Jic//mn66aakJaUECAK125c7
rsYjiOx0zKRupTQdNvHPZGWCDfZzyippsOAXgWzYuqpJayVbf3H+1u/ySSvKPYlxMoTuzjFXvQ5U
1IYtP3phA64U4ZaC1Qj6FULoq2bFLsGfJGz7+0vgaoWNL3SICqkqVAPq7zibiiMAmry+FMK55ail
RKb4CJSFWjvt9ZwUyLa9g+D49AHdx9ODKyzKpNdQ+oOIw/0gFyvaQnMrgZB5/fIjwPR1gT2POYGQ
dUuHEsHTTB12g1BvpJppq9MncL529R9LbYzTpUIfqy/tGSkVNWaCD532SmHkpq+Eol3l8r0nf67R
+ApUU83UoOFAqLllArR0YsJ57LIchfprYudCfHTNR+P/cAn5qhDth05Zgcd2hhK8yUMtlYVHg/uC
IfrHLF3ltFPTmLNKmHveCA3NY7r8l2rmH860+5nmZcMNhs+5aHJuw5uTpXQVT8meGNzEZRNdTDr1
/LPIV0zYva7ZbmQfvAmZEJZmW51YMhkt6QXJ4y7B3/81xYvErEME9HeSg9rBN28c1+PgJ5VYtBcC
UOYCExmfBfsDNqxXnPA0F2drVWk65RTtE9frSgLsQon8eM+rbZ7QRC77Xn25jmZsgk+Fl+i+7Qvu
DQxdXX+M/KWT8T8fAxM9JZ70zU9GS3Vs70pCzLs3NCoWUUjYggoTN5KydizjYoi+PDkqsc1TyNyf
FtCOF9pXoSFfzJxgGkp7T+vrtJKkKPkAY2lCNrvIPuXjTGyA2PRapIQVZiXbLhBicKOgPHEEJTet
hur5jSXpvCOF8+w0JvTo49VpKeynIuZupG9YC/CCYhcMZ9wNdVnd+3UWLJ/uDopAbxTan3m7t7eF
+Oc/4Keh7nn8ztfjO0vnCGabbnhBrAb2+YsTpn9zgPSzMTSr67XvY5jnGDjm7uY8TTNQIUTmGXiP
NVaGKMhiTxJSFhYRCfii/NWBDD+mDukeLFaQ062VaPHubN9IZ85O3l3OL+5BqN0S4L78+0Bw7ZGL
tksN3iKM57lLg43iZQ88P9/sKcQ4c4ltXaEBAglOSfeVb2h8FWhsbBKvYL8zJkt7C/YsfPRkToPW
ipCHCVu/tVshpC2Sxtf3w1RYguma62uA9BYp7o4tsBo6QQ8vMLVA3pCVSKDC1HnEE2oPTcDJPNTq
HkemIrT2lfoa/DO7f6y+6FKk9R9yXNdzo+YL8dtCvMm/r5CZuEcqPKToyEv6obJ5ByxW5ZSNH73r
6lofaYJqHslxzJr1aSiWB7bxVJkK+gfY/INxjesgEVQIZgPLpeMINP7qlaG+DJIopV76JWqgv0l/
iB2eJauclzl7MXNUHg+tojjmHmSuLwIo9F3lMxCU4c+KEh5iVuen0gcuTzLQmiCI4ITHKs5MHldz
CYe4t77EKEbiJMtA4Oc3CRW4r2CPVGgcfLUXBg4qClC/NJVDCqYh/2bvaGTErDuEvhOwfxoSc0Wb
KqQ8tQZv/5VVd7QMq6PJcZBzewBUSzzdtkSC6hlXzoY5DVdXHwPhtYd2cpJ9JgGVMhWtbpIMLK+y
cGrytEdC4fKaZ6VUaSluZuMf9KxN7X4JqS3v0mCCp9Cxj6pl8aiNuT8VCwmY+SAdqHQILQBkEY92
fUyPha+xC7MOHM7wcBEUi/GkSQ31WhDxTl1neWPFMZW0d2+nj2VDaPbSjFBikQyWdPa6gpn9xEmz
QzKndnRdNpUxHVCS5kG4tmkZodyy9ny3janBb0N5nXxrueRR24/C1ADwwh/08kPiQ9+Pl/QLQ9Qk
VNbGuEiqfVyUwCJ+Bl+76zs2g406s6TNgU4eX+XT5QkNg3VV3I8YNYYqTY9S1vn8jrh2z0oSk/Qu
K3ve5r4VKatVSQRblvFQF1T70HU/PJfAYhqV+UiE3FaL5b9y9KliWePUyV6F6GCEckWMGmZOvtF8
+B6RZGSqVfUaud0H58hw4RDhmqc5H3SAN+AIIJAwJvMVLe52o3m+5MFi4NpGSxplCUQCfrX1+Xm+
aOyUfCAWnlGUMcnOMJl2cERg4LjDMpxP86GLuELW+wjL/04JIjPGJjJiExg7ZPytknqK424Fi5YT
6Fgyk152sHCYBzf+2IG3Qg7pZncHxxzcOlcGxYp/EYxQBBZ++OGjWB6lnrun/6gKnenyq/sBE8sU
eTsiupQ2UmvqNTp4GWtxTDCsbhpOlIwYoBEJ5SN7MVB3tGAIhp6rzvhHWHr1aq2Z7Br/+dW1Li0u
DZOzXqbA+30NuTsLhGNdvK2Vv4BuvMgBkEbf+/GQF7CSTfr/UESc6tPi+LCYfI3aEZIDcNtBUlSI
Z8kQSRyZjyAAtoVe+ZO2uqUElZLq0VOmXC1L3fWPHE/4pobIV5di2wDHLQrBAKr4nOGtX9WhUQN+
TkdvqKXha4e37XymUCbeprjDg8v2ullHAM+hmLX3Tz4LoT2clplqCBaWdfnxwhWc8BmmuB9XtJ+d
2QeW1UdewmPAx8mgcFs0nMB0k4bd0DKJVtRklZHCi4YkPOGIVovPdZm1SV4+rUbMUIxY/1x9M1ar
5fpF0xtfsXXHMgX+Z97U7CoDdfglbUqHH3vxxcwE4Vb1UF//UytLgEMwZuYLxrZcKOiBhoSwvUjq
qpb9BT+oi6c6Dqfz7bu4tvn75N+0L+IXuHQ7sxoyHcaQ88kWKriFhwLNxn5KjxnHua+u80iEJC2D
+EzG5j4RwB7UJ1dPn/rcv+zKQCq3OfS9mO7ZSwSiG2YU7evepd7cOcrm7zMju2n2OvvAR6TmOq5K
HrSTMAYvZmecMjf3lB1/ANbKoPBFDsr0Iyz9KdjmY8JyrUhD0y7yfGGZC9tcuA023YPYb4NU5P4Y
Eo75HGojCDy5sKuhor7YNww7ytSGjoofgLfExBR5KWmFuU8ROzygQXnYek1cIvRAmbFJMUB1RVAN
6pN9vrilqmetYwKCMmSBbWrG0WmXYQ9apxbnEMMnxpBrHweLhrZjBdotg+C/IJbU6ufn6U+QLPqJ
rNo/wkfRHmjeGi4f3YbaFNOEHF2HI+kPdvH69jVWTn1rqljDZTjQFS8zAwnmxifNc++a4+143E2x
QkAU336chC0KS0g8KtOXxXP8rsZEQt7frV027HGuae6wN7+Pj5dh4mgrLWBgcFqQzPRX3hnMN1oZ
oHefufgSZjttEFMgE0Xdu86WBvkwlgoMGfBESj0bAw+wYKp3RfOw8Ige40f7F33mt3Mq+xsoeaO4
7MNs8pklK3IFa5qKQFE+ErJ56kGa4VunaySZwQVNyxF+w0uGJwP0q/gK2H3ZcbRyWUYigSaALgBW
Ni9fE77SJpPhXEZpaL513938EiFbvtnAIPVYfvRZ83iSGJ0SVu+8Ul6NMlexRM9EW8I7H5WfOwkZ
TcnjoXZPdoVgeOqfo4AjzO2AMM4jYOiLKM/3YpFo0MmrUoQvVeABWv+bl/9BHLrpiaIhGMizllw7
ifCTTlKJxhk3MqBvLwOIU9xtyn5w9z0OI05oTLp1nZ+0/bkc5fwa8mnjMqr4T1JDTpJ5pv7AC24S
qoCPBkQcEWHUdSPdndc5+lSNOuFGQaXKylWgjiz0kvQ/Nrn40FbkZ8o5BQSqUfAdI51HA6fG2EAN
c2H91rBjS7Qbah0fYh2SW6VPAWwuAO0YHbMCHBk+w2U6oWGzZ4XWV1Wpn9arj/ke0yHzKo80GUR4
IGvhBNWAsdmKqo81+FIdaaNvsKIrwIDVnTxbf11bdnr0+sbuBsQ7/CtLBwtPs8FPS2VFNzgCCjjO
ho/4vdP8VLMSMhdCpcFTnG4RzLZAsCo1dMB1fH61N6ewXEzWDETmv59tNAirFy6esOQMNVhSruHY
y8jPS+GMCMfY0mKOeSlz0pAgEhi3f9qPE3sjMX2q3WcPX1QTzWrGqGJt6jWJ+b5SSKjuVamg2kfN
1kGp2yfyaGzFl5F6hUfua5+A4mOI35gJ7p5cOEcsQUaojXIkgaTDAPZV3ZFf7Gg1tHTBCUy3Gedm
/KdCSK/ZNfIERrUorqWofeEpC9B/TKbtZYuDvAN1gyZx2Ph9UIFrfJBTtMEVN4P/8mazKd4Nxgz+
5I+X3V+RV1RA2oHDRkBI5iBNAxsUkimSLscXW2JXJbpRJugWmBo/GBrQdQVk03bU0qGoNbNvuX6q
K9SFMdgPia7NBFsh+oGqlIJ+XvqMYYvexvej+HD7qUq9jWD6N69QSsbjswFzIqmFcmVV7LUvn5b4
8RPJ8PL62Z96ld8QljimxktljNI9zwlFm5fxVGkkGufEGAUX1e0drXjy80gUjumnCWfu5GAQXZOW
6VdCNlnFDCwkBUfHhMdGl9WqPGyV5GJr275FsMrdUNVXxa9ZbOTLxlUTDgbg5M+nWXsWyv2YmOT3
4W32Tu7ykpIsXAbyKIVrO+jeMiUXNF2l3z0F5szVOQ49Bn4GE8PRdNnc8kh6iBLFi9GdYRTLWk+Q
x5vdTgdQUUEHwOVLS0QROqMImE+2aUaZzREiqTUBCbVCfheJ1wvA30BHfKWsO86GDeuWRAY6wkk0
jueBQ5u95PWnkUfc/r3dh1QnrfMHQi+09VlZzz9mtJ+q7S69PyxcOCi1NgDkIOVFE+hWKEIc7q0Q
2Au/BXY6c4/BZBXC9q+lafIK0FY3S3M+yxQJqg6VCSiiZBEo8W+u1cjX53NTqi95tKev13TZ5gPz
nSeJKzZXtqWfq5ojaK/izqe9TVy3byRVsxW8vw808s72Yzmkixub5Dar2ml4ZvEwv3Xq4t5o6922
Op8MSlpYZDHnz/ttCJTX4FxMAB227hZHZIeMdzQZDX/14qD/C9AgvB58JuryuwAXwzzA2kZEUraI
e+hAZ9GhnVnSb+IRT6dKCkxDwXkHT7Sn0yWlxYORw7BfEefM5KTR/F3p3t3yg5A26k86gd5ji4gZ
r4ilO0UyxvW6piYRuASy3MNFE9Bp4Bdsq7xvAmhOeVsBF7ZoJmgLnWLUw0Bmd1A1SdNo9i9FrAHm
0GFfDqt3v0gCfM2G9+ZKY6b75LR1l0UmVd9z9hEnGkUkSzQ86MtletE2jCejR7mzdCF1N1ylWvlo
krH9fV3f8K9+uT689hQG1yW89ukIsO19UjQprWQuSnMHJqowyMO9SwbJFfDUUpgIzVgmX/3rvr9j
0QwVVD1BM3HJouSB86kRrrMuWSepA89b40i3pHMHT6UgrOc7apoBhh0DWZNG3fe+pqIwqzfdank2
bS4TP4GCTZrpcFHT9IQYB0/SMRawLQBwrqxH7d5Z9H1uv55rhJa4ngan9yg/bWJKiyhS6PzmrM+M
vUNAhdiWITEw3uc+Xaubpidf8zvcaTIxKXLUdWvwOaVojkOZCK0nC4EDELiyBKjbidC3y/TFNgVJ
hArLtj5YfvM15mhYRpBWLE5gypz4qYtCHU1UKNY2mf3Lj9QM+2MErE50e6g0DnThIYE0vQMMXQUK
a09YrSrJQ9sgGMFvsGqjfks8+S3Y2hUbQNDMPTtblZ9ppMLtAZW11aBfWLARk2k2fK8QRnZhO4iR
eYJBgNp7VTrdGB+SMOxKHN7SpH8AGTfrx/Ek42hXgsMDuHC7DivT9bY8SknUUa/l9VJ0O0zu0rYj
xmQEhRR9Aqt/rsb70IQMRYj3CTR7NcKvHDvTlribSY6kKD2kA7q4aimLyRyT+9mEx0sJSOUuNG+5
te1UKKL+TlWwZ5Th30cU1BRBhCrDe7ASEXyY3BF8wx6UQDzNqtlgnih/pbDfY4cfOeR78rIsbf1s
QoFftSSqL9i5pBQywQjy0b2lL7BXA3loWJRcU/ToNfTQIY9ADADyt7pLvkAVJWOjiUZ0XkiHdAtT
Slver/x+t2x6zQ65qbKSqMaVYnbWSIR5RVCmMCitCPM4hb7ruT1oIC9zRxKP0NdDus4fL6rdzwi3
xrik7xh8oDCbRP/Ba9Mef++gw2We+EIjO5klrpN2G6TjVNXI31N0kXEWPsfGLhsqigb2ZF8Ih6u1
8ZXuJM1Q+c6g9PNqtFBcWbhZ9Rknmmrl46qBVOVHd3J9jNr5BKWp5DvB6FMc5kgZ5bTtOXoyUobS
qVRS1D7bJmYBdH33AajHQlmbkX5qH5csWxa1nEuEuCYsS/jn0XUFsnrkUcGq9sxcW1blH4w+wff6
JC8ujsSCff9twcqNeG/QJv5J6z6onaJQfJdBXQLHu+BRRuf5aGQLebvsNgx3wVcOckL0l9NbbEr5
DtPO5ugCfWwpgx2wMKQ45iYojnZVdwRV2fyvQ6IhRXMzr6ahT5bm4gyrqX+8LISepES6C91adL3E
CJH71yFTlu41WgqhdpkpvDVsUSSAEK804FvnrdM5zkZI3rDVJYqLRY3QGW6IugORU2liwWOttscQ
AA3/bDuURjejjL6D7ey435MdgaK8Q1kpJ4Ntdcbk9ffMTcEfO13QwoKDL54lqMJAbZKAYkbB35HQ
z+8VpCosQgScY7bD5udWtAy37WxEutN67/ewBPmMAWsiD8nKWJSvakazrQEgZTNZePF2nsx5L+O3
h14zQKHtjuMvF3K+U1rtc+bodefGY564GjYV+i8y4/weN0fza4x/kwX2uArExeDb2Y7flKvxv+aw
KvgHjkUG8oPC0At1TdJAynYi1Jf70pbU4PWXihdCOXCeW9ALGHt4bolCbk2BrA8a56/H3GMjpko3
X1qURptMNo+i/YiYSh63p/BIkgRfnSqUQjJ/5JudBkEdGq1thdTPiIc/8u1pg0//uCtX9B6mIz18
bKUJFAcu/bYyU7W1Qxt9nLvISsDtbRGfoe76FOZwU6VqHBCGx5xONOnzcNC78SYuff0BosYrIsIx
iPd9jOoAHjO6GXABQT9NVY1YNQCmfT9fpFiAnHVM0Aj4bS/mr0Mf2MO8+a6S8jeIDHEuf+3x2Eql
AElbhdx1bM3ji23wBTIHPGNnCM4QHsHzwz8RBX62j7lBlu0eTEjbuVPiZKZ48lE8UcrIJQZWXRjx
6WwD260fxf56PhG4Dpz9ma7qF2nquOlaRw1zrNLVMfRBL6NmUMl8iNrooKSfT+M6s5gJUzp+Zh6A
mSAeVf1nRMZwxuQqREyjiLsyXtUV10Japf9W4+SKeQf2UokGwz9OMtnbf76B8bWBv5FtnboC+gPn
bEmF7MT3uGRYTCAXf441FWgBVFd3kQNyRsZ2k0IpOvYQEdX/D+i34V9ZuKU/cWUdJOnKsBjPwgRi
eK5rq7CW95eX9IOfCbt0zWuh3ob0huek2r4EmPFl/VPGJmUCDjcvtMRD10waBFM5BBW9XBin9TyT
bO9dU7rX2pLPcln9Q1gkXCF6MxZBwZyCR11eUrZBbUh5OgBljSpHmhc9fBtbouQRPINl3YT0qsVB
uQ6MPIYah/Pny+qT7Re918GqohTEZ3w0oZ8uMDTgBzqRDGZR7jsQPiHhEuEMxM71KMqkBeMbP1+g
J6yOqzMvP8/lVWLbNXx9XpT7VEyvMVqb1D4XJUoQ7w/0lEGuzbMcSLXgekIE01lhf+yJ8OL6eFUU
fs6rn4DvMD12cYrdec7ZuCY14tE9wjV0Mxp6TjsMUX0KRpAPFVPfySfy8UwBkH0bHBchC0c1zRxr
/YO3qZVjMsrXsMR/iEqIh/kcic+nMeaIvkYIzm13gKiiuWzTK0t7aexy1V2TrbECLdO9KQbAzNO3
WLK+RgndxAq2Qr3JfFxbnXeSwmI/jhfpy6GUGxgWb2j125yaOZ0T511QX13nSg/Jbigf8IPeEoVy
h5cm9xBKoND5MoEyxGAnO1yfL3VALnl6TYc8N2lQ+usKTEIWmYeMwzAMj/WNkES7VLkkW3djbZ94
QhzwpkvKQu+KpPfmIxIcd3Q8/22hctY154qbTJ0ExYP3WAPxK7MqR3nZjdGDL1VsHR0SKSR4mn6O
l1hvieOqvkdT8vF2XHD2JgJdnKDt7YYOgH7ECnZWPCT9CWTqmH2bin2FARURYDOqV/H2AOvnmi14
Yrj8K8dmC/bqUGQ1lVnTLRBfWkp+bsK/tDh+4zNkOZgkp2+RCKq4gue/hUez8ZglQUSylJX0Owvo
lkScYZ5KhmJTG+tVAmPw3Xwc9XVyqaKz8h0t12Bmpbl2qBDSd2DYwdgc2mWfa/h/FQOuL/fzzMBM
eMOX9OvRmRSBkC/+0MaLtWxZObW0GJwv8j/W8OgKKuk8k934HYFqC77noX3Heb0EdzUIeu/KeuEc
FRNUDBfQyP6D7nUQDCnr9unFvgrc2sK/MKyS4lyZmSzCpuYHYA2UyULBHjw5yJTN+EnqOK/JfcsL
FUfnht6xwCop5EOBqGhpDr5o+8lFYW7K0K8PvppaqLo7071MLpPN4ld4G7phBZdTykAM2vq1W8Ng
rv7eobpWXCTQ7ttutRIimZ268exABpOhKX3UCadZHhWzjWySvK4MJ3PZRywDMerRbHxrsrRynaVQ
Bn9YxPkgbGFAiB1kGV8yfmQgexGeGztWzcOkcvXf/cVo1BQ9Drd+kM1FQ0hmGfZlixN7fWI0y/Yt
CAOTcrj0EPJ9w4t8TrAdCIAd9FdU3tjhmt7YP1kp5IJBJMgJc+qwn4RoU92/IfS2PupyltOYZSEn
7dEOvBbEFnDmsc9D52C9XJ0Av4FLc9UPiXwx5WLeKehb9uSohyjM/oQ2sYttugsfgijRP2wd9T9U
q572Y1TsdvtTxHgsIGGeYtl6IZh68vAua1qbCVP1Z0AL9dnJRDkFebQ/YR17AVsuRZyTGYN0fw1B
C7KUGRl1dw3n8RZsSOZHxrRAPuyBCIx1FESXN858LAs+VNOj22CaZ4NSB0SBvPQjtNiXfeeWzJho
RL2ZB3bXqohMKloMpClvci3M3SQTCCkQgFOLo/+KWyNbG3fSaFXMrtK4Y/uYDPtDlMWtBuK49Agj
o8bpl90f1g/ix9af+Oq0AwrTXcxjXBc4XfUcrHkNdQF6HfSRfTGtjyRXED9c1Z1QxyJSfYkwqKxg
Cg7dgdyHiFGqlS6Ullybsdr4siTIb5RMl8jZaZP9mDT/j88tPuPQrevsDf4npkJFdBAqtnhqqAk0
bVAhUZTP5gsom5uTHb0mltwlFG4CVbyZ3h6QOEyeNBiMZDGBSRGY+C5mb/vy95iQWS/9IFpmhn07
eeX+TrtKAOFFYSklZzAWtjbPM7cDTIpVaAyrqkdiPhV8UQIjQ/iTwgHQc0A6HZx9rDtLJfRSI4RO
mLWCQveypye2EAVJU4Tc3kQ64OTnEsbAk0XDs4YYN7AcHzCE+8f+YXthRA1utt1UHeyjFzTh88ad
FfMNwuKgZym4WTaooxrzasJHbrLSi1wqKwSTQGxoBqAJWr+JX4GFDTDv/J0QBmJ6rQzWbcP9qwEl
cgoEpAmWeN/YHM6FqW8dlWDoiEAT6oIYIrAVxTqk4Mh4fBj5lRkPysU6H57r2cReLjBLEBmMS9wF
9Xyg/G6cIaPdkZxquUoQdETrKa8R2vlmJsYue/topxVd+8FPJJRUPhbPqnG7bgLPqYZy42h8vioa
VTTMlAeO20R3nLQlmboO20+7jvmqbsnuZYBxUHQdygnl2KwT85PnWF2WgJRzOAoHzE8p5WShxcGy
1VYOs29Fx08T9M93AZctQ678elc1w203XQoOynIgQFRBTOwXU5y4ywbRDhLL5WVjUIpMmvbqkWn0
ikqjop2A4T9GkE2c/es+r9M3d1csRDvLV4EYaTBB03jUQXjTH4kzX5lUzd30wAZXpguNQMWybHJy
24s9iXftccdPmDXlPfo6KF+18ZkF+YR8xBNsuDOSPMYAt8yy0X7WMgcaOaVlmdK6QMdfh4WpKhoq
K0JVWVmc9KL/XFhXcc7OijOnBhvn1OT34QrGYN2sNHOMuir8FaL3GMyRt60DKTQPoiInqRglZjOt
S0JjSa/hGkLDp2mWMNgXNkS7+xjsHaAhwu/0KpasK6Mt7O6xBmkwff0Ecie9oSFpTRklByAvrIHQ
7BAw1whOretpZoKn6filmVP6Vr335SrMaCEi1Wrg3Z0vlmkZjA0Sth77zGY2zOepbzT6aLkFX2F9
dJFhIdJ1rpDd8LawwnzXoaR4IKEkXTZ8VagyEfl29bh7BqKrnXdbmObw17ux+WGLMke2lmol1H4T
GxdCk7VRdDOdTsOX4XPAHHwGxxQw+7C2HhxgHDjg2oU/0eQFQ7iv1qCQOFvqFHo6W4w7WDNuKZGo
cQ0c/prujcaC/7+xMa9ctaieGOEyi0+Q+AXr512DarcETcgSagP59Ht8iTWp20CyzStw8wn7HmQY
MVRXjSeZpUQEGUXPeVeI5k0RjLehjN2B4MuEfv7QDj8q9/tEQj2Arn+xGQ19mCJboe1inkJ/WVKJ
DDDMkDwi+q7lZ1kH0KXxm7UpkmisPMb32AnRaCL3jLu55KpZmHyMhg6xQQd7uh+40sHinv3hJs6z
sMkobjYKISr4YozfYL/VzhsqV+acDYba801ioFynxOnjtFXm7eLrPc8oWB1QNWYJOiPHWp1O3V+V
g84AJitdeIQ0sv8XndHbdNTkJpUlTupK2v6+WwcSWCldzg5PbUmXIaoJxfcrEMsFrVm8HNnX+x8a
cC6D5AL1J9PYSTryoJb2+zi2aS+p1mkizQZ50ybz9f888i1sUtI8iQK46QKokmpoz55N7RIFFkR8
s03lP9m5zpifkW3+ywh6eqPSrSuvf32KIoc5XCH+N8EW60EemydN/Ul63vugN0r3/0Ozh+3oZkzu
RncLnUShjxBsUs7ZpI0au4GQLK9smbOeilx5evAIa4yDwWtWivo4eLHKzjJWGYVtPPylfvnmFVnZ
CszWtnICeNC2kPe9Lot6Yopc9KtJYK0Af/TAcuKmRw9Mxx0elgNrLUSsH6jTegniGH7PjRas/BYP
TAmnyB7XI1UFuUKT7tl5V5Q2TYnYMgu1nsCHWRWzn6rs5HbsM0OK0dGbY6Z4Cc7bccvWP6Z9M/yR
gRAAMvFuqTndQ0r6VeVtnDiKbxg6W4xEgax2pWped8vopH6E0AW4c3Ap1lJtDGe76WNlxGHtx8xY
vWGgWzioWd7OiVxZFolbwNSPrwu6/vsNJA3JK4Y/NWL5XqoNQ122Ertn7/fw5P2Y57tKu1QwujBz
xjM+Ol3vHcep3LJM+OA7nhXEUfZkNNAvG19UalGSy7fsFfVDwkWI46XsCa6PtfJTa4jH2DlzUuHk
RDt4ONte3JEO2/vkNjWgxqLSMVe/9BEReFkNrsIYb1jXdkngCwfZ4P8x4lgQz63l4svNU6GB8+gb
BaoTjuxPmy8fGWPIbuTt/6VuP2ENpXAoEBkjEnv79BFZ0KlgQS7TP5/G2+dFYmmRJwhN3gpIkYwi
nsNJK5ydJl+QeGtMGmXKf0zKO+gTAcd2PeWf9XEVOIBFsyW+DEp2fpTFalHvtD2wq7Gv7f6e1Obf
ccEm0zzvvFCTbtmnVNXjgJnhtm5NIFyXId8q4LMHki0VOnS3JgOisXkJy9frP2p5J7ErsPnbiYXG
SyOAp3Gbyv/aqLcCryLHyljW50tQH3A/oLQH53zzyuQNqN+Oa9lsMm6gdm7RaIUIh0KQ0XpIog04
yjUL7UfhVaV+jpfAfAklBPearzTGzbhP9PT/UBudXKk4ItLUXmj2cZ67PYUDSbUr6ACmRzroppFX
Rsv20nXd3Bknv3eUBmFQnExWzRFVPfleMJHtfAhRaBFYAsFzNGt8QNGyJtKMWjY0626liISBnGK6
i/GWbTmHAxcCjiDRRy9h4D+GWkzxXkbxM/zKM/N7Fxzg2AJNrnHalMyIzIAmUlNsJRS+/jmn5axF
YlBI2rdV1abBq+CdWZbbfIePsnvzL6/ZPLaJBSKEVhDtrhywTDgVqs5mhmMkRFcTuttQ5cUU9up+
kM4e7Jknx9E59EmjQCfCPLymzn56GeheeZl5x48gAkl61mVMrS/1sEY8X6zFYPegkJqjBOKmYNRz
cOnPmxlckuQ9vQng3nMHxL6dN6ze/M/FOc8VIJ9z5pu2ArxnRlwm3JULuCmglqWFOv2NlL5LEUkZ
gbKGXbNzQsot1BYZc4ciH3iLsnA4SJCcwTgJrw3VbcaP3mjbgDEJMhrciWtH28A+tiq96+gofQdN
mmQjBwRe6vBLGrUPK7qupmpg3Na52Vcz3D1VmjRnyTuHh9SKn338xii3jec9bWWY+HdhOJ234MxW
5wJEi7PJz5qEs1QjB2He4wQ3YVLCIJLvKzcjmOOI51UfoAn1PytbuKUKcBVf8SrZycfEj82NF0t7
syIkw0JObcIRh9MZj2HBdIq4QKqjuc6rND0+GdggLf9uHG+SIGQge+Wq0rLi/DFxAWQukyLKMrcJ
O08mpvyoBG+sV6ok06zJFVMVuoZDRc8zvb8lpRWvD4f3Opj2NZ/C4KyisvaSxxlKHmr+N5Lmdjv5
VxxKmeOOX8i6J8zDme7bga8eE3G1jxFurGIH2z2MHo10pJX6pM3f+8R8B4fnj4+qvV3TWMMcdDsN
HVi+33tE2Ui5Y5UG/KrnyC5H6Wv6UXJCiFuzcjZE5v+cgoKDfiXOgFdpm1k22sjvXZ/k8h1J4gov
oys5WWnJaPsez3F41gXHoVNEYGjHHuy6lBFQsUthAHbwDbFZnzDIrVwwmkCE/GAvqvZgbht/TE1r
EtsqPdn5oUedNt27tlyO2ZlR48qheaDZRN0cHYHV7eQ32Wm0Qk7NHcC/xtXF+KFVdhdWLQNimDE9
Utr4rDi2ZUn2I9zMV2i3eNBnoEJHX3aWTImdNSORr4fUMnaJq4VFznvmTUOlA3w4S+WkWTS9cEoW
C1E5apzRLDz7IOZ5XKDzGbjWy2hHAPawVGSUEzj0MLyD8ijVUQApGzamqXasHrdkC70meWnF+pMe
Q8OMFbDqJ3w84aBHGSri6AnqqxVXbUTISg1fngI4k3L1KILT5WebrtxO2VVbiaiN3IjCaF2N821r
MVdapOMrpuryTtNZAnxyjIOoGOcMW+O20RbyrV8hGNxnyMnUZiu+3FE1l8z1BBk483wSMIrphiLq
3g9i9SIiB2fkj4P+ryn6nnPiY0SkuOHoXP7sD1JMGk6e6zV4kGqt1j8N1T+ZPZ8Fv2AgPpnH15G4
uj3UIQ97JFb6xvGOx8mnV3hvp4aHQwmLK14/U14Hku8dZ0w9dZ8vV+exQL2G6HMiDMQQmhNqdNch
orCzCWkkO72oZg4QqrDC5SuJ6y2rkf+CU9nh3QCiesH6+sbXX8hkK8pCH/84VWbdGUl17FjBBoit
XQTFbKYF8MMypFq2Zg+1evecWAkI+eiauzDCHnJIkxsYfe4gNjbee73SXTTSYOlq6EYMdH+Hxyd2
IRbM75GE6Pp15vLSXPnYwiPAXvLDTxN4xeIhRb7/0Lfs8rrEvJkFbkv72MJCZUtqijbW2o0hyu2W
pyVppScJVSvYZ5bzhDKDtsMOymj7lZTfLkoMuymsxs0iM/8yZ0G5wMxgaVBssPYLhxxYq97C7x2e
fhKVtRsD9Zqm08g5PDVQYfAChwNEUmsjhL06jdEFP4nMqUczogek1YhQLW9k9ek8QRrz7bUuXQRh
CM72DQm50gWAYV5j3UtjQakvjE2hVidJtjNkB3mCbxDlRaw9Jv6K2K4JF33494czzzije4uoCNb1
JNQLdVgXGKBb28kuN6giaJlB4AhkndF0SSkt4ggE72iRbxrx1al8N4ePKRCw/e/a728nK46Q70lt
AD/JiG/TIAq5Fv48nmjBNKH1a+/OPoMGFLE5DcHMP6dKAWXr7DMcRSGvDptBtYzcqXm8nBpuYk+q
9f2t73OfrvDGW9mtwIJAG5GaFVGZWaR23jG65Q+eVM5CIAio9K2YTezGH1YnUZYbTD2XXyrdyUEd
Kp3csfgznkKKWdbyZSw0w94vxbnSCXnxNVQSPDaOQ0XopH6XGyLT08wr0YnW1MvvLJWudtKS5tby
jY81RJLzOzNYv5xTXJAwckWiUCciESRkLjf3sJr/Ldid1IAAnzbfLTOa6FV1eXbUloz8D29Jn5gd
hL8tp1knZOegcpFkkJ6y4EURVIa5RQLpbGhNp7R+QiTrr0ZbXSBHsw+zgcNefkgnqbNeQ366leaS
g/tebazWF2vvpDqyegCuuO5hraMLrvOQ09D7WthvSLqC1pkjphHo8xAP9IdrqkrhadvnJ5QJb3c0
EmE3eTICJ+X1auiWKDUCztjYLDmdsOCrMkwZQKqcmPYiRkQO+MD+wL2AyDjKJ7vIwGe2s4LI6/AI
N0abCOb3uc7aCgb3GOlcJyKhJWQ7NYAbkpnSvkfPPgVIembb26BxJAg3oduznbGfBs68yWkZvfrg
ZwsjMmCpcOqwgfyIlYiNj5paflSkBeLj2xsoGEH7aCkAtLPZztM7jaCh8lGfPMZPq8Bozw/woquT
gd1Ope49wOivwDx9q+WGLAbU1nTKj3ALZl/lc8mLH9nwZMx+Vduh5TWOFyd4xcI/0VgsLkeYbT/B
Co9OOHYpWaMCVvcAfXuEVd8T6455HoEPo/yaNtbimIGjdVl1zNSrOo8UI23Janoh7d/bk6REdozy
Gd+uoWG98Lmfs57XiRTJbjx31WU3ASOfXHqdT7achbG/TC8Nlikvz2AXukMKsP+4DqnlE09LDMbi
Sv4WV38kPopl7BgEKLLsHQ7GqS5sQ2woIniqWyMqRcmNzK1BsUbjxF+TvMbFiVd3BO9DvtxMlOWs
7SSlN6LK5eboxPVRD9ozhTFVZwGr2JW6oKsHWe2+xN6TOfsImYCmiWWhRQtlO7p+YDHz9BbpYFvK
QgmPO0IvPVPejKgTZAQL9IG493Dy9BLADkb2AoDN0nbH/C82rhyZdKPZvq9YkDOQuQFvAF9w9FVi
MYba9GAIVFvWKInZS7pSb/jyAhIp+yM7giV1KIqWDIiK1bITmq6yzAI7E94v4vGiB50sPgLj6m1u
E8996hQqXJbcCFu6LgnRZA5/OPtUfJmgoE4YgkM5TeEhD6fm/C1O+/6jY+mgf5uGy7B+gWz4Pi//
mQishAYMIulZEu3Pt/7tvhubnI/lPBKpfyxqhMFA1tUUAjHtSP8siFSdCew+ttuvGGaaXgDONHO+
3Phmcp9w0B57u14qf2B91cGggPHDqO9Ja5nCR8J1G7DHWWjYyWEl5eUe7Lptav1pF8Denv4n009s
TPHehb0VqgX/cVa1M8vHD0NopXK4PYbzJIqJv0qjppk6HwLUYthNyvLFwmB5WJPAMyViNSjRdv70
581iNzvO/qYcit1LwbtXkjVzO2J1DDmYOSGnvHr2QPC3VLoQY93u3L3l1n+4YkFLd+6ehWUXA4BE
NbhAk8gwJwMTC27Jxib/vUQza2TjYAvW41i6KCAueP03JKEQ+QBjfrrZU2RzySdyOOwJi9RRRqQS
4+ui81U4tsXhMFRSIgP4JMT+UCswBoJnwZ14GjeClhoFavXZzcxooxi8/MKzn4/Hs0GAmmtvb2CD
nwpuQwA78F7UOXAHAF4Amnru+UnfVU31nZO0a35GdYxH8tUjY+FR75ooquwXaBbHRYL2ek6Uxryl
vXHC1nCJOiGMvyEng4yqhhxBYYblSMavwazOMfLAKdlhTVG3K3rU7GqjnmYFSckZrpH6XpqGd971
OB/R04iaH965mTxrof2Vfctk024D1DQFpoOQadk/P/QVnc7Rqm3Hpn64oWmr40pT4jyvyuRpJnxM
5IbZt+AuJxw5rsbf8CwXDFKtF3MptnLgqo1kZTZy6DmfmGyE9nd6cA/OWqQOUV7AVDf6W+t98wZ+
y2Ua8npI8pOnvf0WXSWgSrdtzBLuLv+KUws2QR4/x0oTXza0blY3jtSD2Wau6HSFgj8W7wMEpbKI
ZkG3Z5rXYV/NwkJYOcLZxbdXVHup1qxQCao24bynu1dB4/io/ZqYAbnaxPcyi00xeIn3gVyoqb3a
8SxiOOmqWD1LFiE168PSziwv92l0uAyEoOh4DGO2ztVifVyDxQ9/fNpeVSqpFCqcMXu6ki4bRhqt
8cfn7bZGjTecMIHgAz8Z0UJryIKHM0XylhmpfbxGTxzEdypGVDWaAFXNALGaj9LLmpJQXlFDv1Jk
t7cAzr3yAwA+5rPpN7bY4iQVStJQ33be+AeHr/x/zcHHYd5nJDbYPxilgoXQIx4lFnDhlJkGcHt3
e+yPW2Mevtd2hQl6yNnR7gyAsDqJyoaxwdrCLJk8jDcbxIu3Y471WhX0PvlVxGzHRruW0Gv4nBgT
WQLDbtOKNvm8PPQ6B3jqgghmVCrcc0PJo3KQtvEXrA+udsFbc9vcPuFbwOoWuPPH1gQWTMXfy5q8
s2sFgkPVOdQ6k2b28eOrY1v7BxjrP2mfZVvJA5VyOxH5lwjfBX44Mr6TelmLzDnCHRGNXWAIpLI1
YfrZEScC0mlYImjF02G1oo8/+WeSLSzbLu541evKbTpkariCwSLWzVN9v1m0/nib1w4hWN6i44Nu
+frVZYwy+vxZdm92xmTxUdVCEuvOya5sa3F5MJM5DF0h1tcnYjdh2L2QmxiZpc6wq2rOrlvYYglL
YMJAEcKyzw2MyYx5bl94RAJUAK4ZYzkRIx+MSOoErmgA6tzI14ur0mtNsZg3eNOC0D0o2+Wm85Cb
oK7QGWBguoVuRTxlHvHRZlca4bs7Nyz/x77Idc31US1TmzAcElQc75rzfbT88OVopKRo6HNdjJT/
cM2VE35xRA+RfQtp941NbLvUp1IGTuIA01MMKMDPwQdwpiiYipzYP5Vro4FeGbt5K2n15uE4fRnW
FiETNWEa39tf5EJu3Kwo3f2RSPA+2gM3qwrGFbYE9SrPtcNW9TtTTUOIZUoU0ohZt4mbXWLwi+t7
Ais3UZpBqykB0miyToZwXrK8O99tmfjiatkulRNDjibWl2yR8kFHqXscvg+AR07iSr/8bwM7KK8H
cdhUukN2+V1I3dvXtPhU69XurS8//AzM+RhTHpjmzYKyz6sPZmTNEKXpKlYpmxTBQAFWijMmhrBb
7zGeNTPhPMAiKUTlr1mS7lBH8SfmXim6NCTaWAsy+2fy03NM3IfRA4YH4i+D6iR8t8BQZ6DV/knu
9pr1T63i/wuUZAv/IXpBF1TuA8BkVbQIUOb0KYHrHn2AYdohs2PVrwudN+pm11lD5mbjbPuPiHkl
nLe+dw78zlixW+Z9hcag6B97NnEdzakdMbVtG9GoEihLcjJ+n6Mrdqp22T10GV/qRoU45zMv9FnD
/dmZw3TnRRage2sh9sW+h9UTLzSoIG9C4XhogBG5buECOpDnbD6n6ds0hSQff39AmLqXDXO6DF/t
Jxc4E/rg6RTOZ7XfZWrHNspjSWZzbphZuLt3ddhxdPnV5cUBnPOXtvHmLf2DhWsvX6nw4eREm56u
Ho5DQpVVwF9I6IqoiVMlYellgpziaHaQus2g/OOQw5PhJ0fO/oTSgeTso94BEMiGg5/L2+KV9CH8
a9sUuhVFDdApDj3F95pOW3bUG6ifGGjbuas3EfowKI8zoyhqFYgFbol6RTKMfcX7AFyd4Q9zp3b3
gLHds2d3rlwJH9B5xS8al9S6NMsvTJcH9ddASjMbodYRWuEHjFrWZ6jV3Ym+jJPyAZhzLQztUPj/
YwXO0Uw5LGx8sc8rLlpLf96pU4oIJsl3mKLBn+FzuwEtkn+3tv+KMWGZdpeYWIxQTfBRWGxPj1Ba
6MvByYDGLkrSHk3M7RgMgx/zQIfE0NJPSC16yq7pkYCpHIZ81AZ7/bLr7md9BwjdCAPRRwNQJs7Z
U4Yz7rmztvx9cEZGRhPSGgchDLtC4yrnReCBkjyEGMkZuiELzMkZKrsbR4ol6l3CcKFgjsBasmI0
z8g130ZqMC3lp8VDym+pzNRdu077fkmdOed0+8XcM++UBV/qoE/Eimw55jiVB5ySw0JKKRiqluXI
hnN957CRG5xMy76U9GJ9QxL13SvMkBQcTRav47WJJpGVpr+JVX8iPni6wQBEX1iH2UKrlOpkvtyO
NaxGz56z5KF563Lw/Na89sIeFpyiB0x5u8m8L8rngs0fi7SSaVyDwMvmiARbeERNXInxdSZ6xGcL
m+h679JdIzq99/dpHxSvwqWoCTf5hCqZe6fl44NMBuyjTYR4bzs7kS7RPeLpRkC9qDBdXeT/lwyv
SwtE17qGh/+nW6RoXrJMKQ41GgMr4QwD/VOtnCTEUboVibX30yfbky6AeEyG0ol97VI2qe682LwC
xUHf/dpY2KRrpHVa7DHINqkWvnmHU7Eacjhc/dnTTCqs8vCWSwbvhLEvfevhJbGVVcUuv3saNP3E
s0J6AR//LOQSVo3JqCPUIHcp2hW1fz20P+guSdWINjDOuOX17pWAvMp2mjuNTXdI2eQYOA590jUQ
SCzyPlhoNPmrNOskohgcM2kfEktZsNRzJejBAfxbALlTaAFDs8RlO/pWHdSbZVhhLyGwPXiuQglS
5uMApn+tYctRnXoZmYybFvz4yXU4PPVcuBgoxHou+jzra7DPfSssa1iB5EmFyiuIMykWPdJq43Ud
MVvx5ihLr0eZiVRdLJO3gfLbz0yCMvlSItg2v09n3IqCQufxWde7Lwd3aGND5Ogpk+q/HRfMYtwK
W2ytJeABFUfonfMbwnUpLmMaKArLmiTb97/PHPoYC7eyFsr8Wkmf8JC6qlwvW/1MuvQM/opq9l0r
CNNbh48UXgwWFFzp9bq1EKpRlqo5l1JG5EkE56VnHSpostPUOLYqhNGiGK2C6YzzU2ARtqdRlo/y
YlbvEGz5nacnMFp0sJ2GJ1/j5tCAqJO3FMMUfIFmVyouKghiGVfPmTeMzLNX4HN7sKd+oKSTstnw
uFPv2q2GEYDPnFsxZfJMIiJsk35U9G1qpOeuPhFZ6S/D9viz/KsdkyivnMAp1oxJoAHgjSQ8l/vm
BkhITnTr+vaFP/mZ9mY3bFlFhlpUNIdzEu6Img8vMRtsoMf2ewekxHsSchgwzmERgUKrLYH1U6ox
sJDYmFzAdjr3rCjS0qO0FPjzhd7T3YxXGT2nlpe+f3PIELbSsW75/ZHSFKosJkhzpqpVTK88hqjw
G8wIUKPC5vOoV6zKCXpuwZS0ycH1EjX+COw+9tq5K+FCDrxS4nVUHsQY1ZAqKXOZqMH2yfAgQVOU
KGFiXKtwq0UFjtK9IKbg2XKEgzq552a2orIuHF+YZ3D01VeLysILL+o2GAIOCy1VsbPHYrAyZf35
l+0Ld8StQY9F+I8+rYp97w97TH07BAcV2PonUH21GNlzn9+x1mtaPGU5/EHk7uVwEUqEtjihKxA0
bhp1gmmu4UUwQ83hsgIfk+cK9FjUrFcwT395Eg9ZwVGJCMKrzXywGChzGA2rxNCv1SMkzmJnrOTU
PUlutCJa4WHEdPsFiKZRlIkIq9hYND99s0YGH76XlubTAqdULSpIeFDVftEekPtxPd+xXdaq9aaD
fUETmSKkw0Is+rJkIOHNd44e3FM3JlD03Au9+YTutyKMFEDZLx/R1mWEt0fVpn/aVkLDdRVDRciJ
LB7bG/qYdQchtUbe435HNwTYM6547mwPNjguSnOYdO8BEQ86v/0rMec854YjQFH2zgHPsXDd/rLp
OREOtzxKkXQlcjR19cPCBVlAuZrnXV5QqsDB4wFM+M0DxvW3DuS06qWOtQVPpnZymjxb8nho4XBD
oI9gL64vc1pj02LxUp7f3SSqL8Wth8ypT5Fu1InfUwcDAJp6SuS4HijwwGE5VReLFpbacJmRaEcd
ZWaj6Gh2u7hNC412lIlmDmryBio1W6ZMrkAv5z01U5+C7IblxLywvQPEcogfmPbJ83nJZXInzVXK
9Lwu37NEnmoOO9xr4ZCotIzR5l8AnwkV9ntYUuLkTizrISB9UO81qiWXjSoVDtHlDRya91055laH
DFrGEj32m4ncZGS9DvR/LHh7auwJcx7swRugnn2N/6Zt7oI3aVIZ/M7QJytm0RgZpw6jHDT8sQ9f
krCUr8zKVi7XbOxDxMyaVlwn7k0HgL9Hu0egF4XSDxrMhLVkNrMR2A2key4ZNAG3Liu9swRFR+d1
O2nrexb5P26FDCefgctMkQUqZ0SnUvdDCP5Qgz3JR99m1DBQ8GmOf6n2S9EesA2Jvz9S/coPh7Qu
Kp+ANc+mqJjQWGwXf2b6/hAp1UR+3pgLMzmIaiW+T0u92cnq3cfq2XALNzC0bf8I4w4iJs8+5rfU
ddoZtRTKGL3cWewFZxNeROENuSSsYTG7QfO2qusV+Jtcf8+SeYJG6f07AMXV+AcfMwrUCFHhSLh6
QJkfGNkpH2MTNZbeClTn+DW/Rb3m3sflba/zy4/oANSbljnOo6ZZ5wtmQYgO4Pf1wbu++OBHxGUE
3yXm2ISK8ypV7mT/I9p4PmI5gUzswpoXvDD+DiDf3+z0lvcieQUmcfNyrfWwdztLNkSTKrxJaMml
kTLf7AD+q0WRGrxFOzefWkcDmcyjb5E02FnurIgcObg2AuzzfoZ7CHk5V1mNYl9dpw0EUi8sdFOd
Arjr9c/NNqLu1OdevBhpgp1OT6DdZAUlGTAb+dPF0h35mox46cA21CELXoFu+w5ctjGk23KldXOB
yB6hoAi/r3wW0UvR4uWKWqx7TiXBeFMgtSuDPNKD9JvxI5XNPJv+HN+GjhMrwM7tzvBGAd6hM1ko
WDMeXTy85s27ppufewL4ESaJR3LS4ZRVv/LLxtPKJTuJVcfavWH57PU3Ona+MDVrIMVqquv3q1/J
wxfxLECgYUJG+CaEO00nniCfBIweuR/pRPght/nP3YHdinum85PHaXyiZKqR2Ebwcqnt6Dyq4c9n
ONpsHYgIFROiMjUBNNKpurlVVdXbV4kioatamuNNhQf4mlUUge4TzSEGDuCELGEb+f2eeNCTX6xt
WHjd36h5HRagNf6Ws5mbdsfbxiET9gfHdz0epj8VQl7UyR24NcA2LjOfWmmzHYuoOhYZ2F8e6CQL
7h6q6+ztyWjkNWugcQ5TpsDZxn43OSK73zL+rjrZTxIY42MIlpnupvH5XTTYu/hVF6kpg5KhSpq3
k7kB+vb8tXiy2piKMc0HyxO5k/NOtfjLxN8d4s78bhPclC57FZaFouD5d3GnpdWxCgmB63Z6pH6Z
FYuCks4EDgt1jQugF93XFDpkarw8UNjjtFqb6ykNKmvY3D8GP418n6Fcbggmu3JUOW+Sfu7n9v6p
+xq5axDpblHyr822U1h612PuiFQgvK0tJ2Qde3VzDP/4qPDsS2zLbt9s8YoJ/Raz4tT7Z47QLzNx
LNYIM4RK5q5QA6YYxL225KCzCBb65vsuUKPuX7q5Zc1yqm/ADcZy5bYdvLwLXyDM/jnMfll6sQ0o
S+JDCK2E5FH0LuM2XVu+MFLiOS32IlaSAilLpbwgUt9HHK2+Q4gUB9Aw84axnULe/XBUReK1/kbL
wfY103ij7xXpuSsLdDhXldIS5l3lPBHLVV/JcKJRqvx3qxTGnxpyBq3/LnuoMGOKqLq3TKXJLc0b
gQe9QKChgC07Z/MmqHasI6ai5o3DZarzEPsp0+1wNai9fQLnb/ibI9dwe+zLlWwUMyCRXs0TydMo
ZXNSp0P13HZEeWpOyq5v4c58bfkJceItDpynOlafIo9956E2Z0xPZoTJ30/SxMHrOcrshyX9gEtI
AK72hsd7RE39fhe5Cp0KbcHNDCCJEtqKhn/c+8i3O7TExdcUHx6SlUKcWtNuHr5urhO8PQs82II0
4TH3s9vpik9bZvCCHLYQnrgzPuvr3VlK953bDn5szI1STplV/FKW/u3yxoBXrVcmsd0xtYeux0FA
C6Wy6oMZQSSJj+4TvtEoTa87fst634kwoMaIMibPHIGwsgpUXuqWLpVOB+/DWcfbR5U4oO3J8H4Q
bkVxAScsJBiVffeLYEqO/aKxc4BLnj3lno26rr2q7x/Kt2SgGa/iTWQEP2pd+czed/WFYwwSDdhz
8hMZwXauMoeV73vbjg8ytFxbNXNRcm3v9G/dGuNzOnl6AaEaZXTPXyoYGUGbvAzq4KWyx9uJO1++
tLEPUvJUYpKnTXf1UDJwqWXAPApjrPzKqLXzkXwWD/rv70XHSviuj6vL2A8fczrKhQCSSixngo8G
I5t62ZfHE9SGbTUNHw0KKHfL4B3Mbt7VNXmX7vOTwcHz7XQcXT6ZAmoNUScv2pg1wupo+cJLk3gF
ii2Ed5s0bAfe/2iccljqpJ7XYJH26eKSLvAwRPyKWT3iK3wuS2Gs0mGHY8xkeAlS66CBQj6za85i
j3+1fb+5ybMIvG/fJkH0I1OIkuvT5VMo0szzeqfujbkFtPjPH+xY3rZcQvMMU8siZpnSlIbdEBaH
5NWWqN/CA2NFQXOdx+kKqdnPiboRrH0rmRyEPYGMggsSaAEt9ynjmkVoyMdLYmjzermsIFC7EXWo
Wp4+KbgSQwj3bkSIOrrRqoMD1ZmgI//OeG6WmHXq4Qzil0+6LxcRB7Z4fysEkK1+kO+VIvULCtr+
Iv12DHkCvPs+Yd/4iNNSEbIlp/kyGwy9TjjmR5PLvJSnsnqTmmdjuAMNTueo8G20F6ZS+jOZMW+q
fPbLU8lOCvQpW4as776UR87R6+WhAoX0XMxQdrL9egrp8iqJ8vCFfD66GaKNMwdOkxl81lldXqQz
mXaO+5iCI9tXfWZRZI4GapZPCbUuiXzunkAdZwzI3BmOdRH0BKrAT1I1Qtf0D3edLyswK5X8AnyK
TCjHrDcNBAzrLdRr4POn16FoRSfzo8ZZvhDcjqoJoeJCoJDEcavX+CHCathVYwKlXu9UEwrXvxon
/PTiglfUUTVZ0NCvdKYFw2PZEXmNLIBVR/+kvwKkw1RkLlaEbPZM6kGsoxrY0mbNtjenUgiFtL8o
TQzfPC3BVAw6YkbRs7uzf2WflxcLt+Ugp9W6PXmH9OJiZoR+en1xAw21ywFQzrj9WudjYZj6fnaJ
hTpFzEKmAGa8Gk2wxZyJ7IdJKX9n8MLgkF7cI96VuiEfgiR/IT9l4MxaQhwQGXj7uMNpKcreSdRl
vFwVRoMtCgbzLvYuxnifNsPUke/eHiWuLFHyvhGzh8/+EPGOB5UFDZyuznPuYNF8JUDaTvdDqsJV
wo0CQap7vQ8Nv4w46JhteIBlz30WnXKm3SkofUMxIYXo6F8Y0oiZxHDS5n8UYJNa+Wxwampy/T7E
kceEqJnEaF5pW7I/3nj/ymIJNCJzoN+z/YMjw2cSjeyZeofnPmnYUD+Q0j59pgLivBefVsGjsa8I
EPgrsbo5deYvot48Y5q85h4Fos8tydBTQ07KKy1rpLv5l7O/5ut1/4/iTeNwusp2XSw7M9nxegg1
Q31o23CFO6yobme/IyZvLiix9idOQ8bMI3JotugJZQLHnDDIEiQ4BjKCWgb8C5ibK5z5ikwJvNR7
5PixtnnLwMe+XKK9bhi2T+AhkPwnIC8NbPa8mRYhBM0o+Vkq42U6+M8DZqRDfW/OT1Hw10Qrq+3t
YYTY8RfkD9Rsk2FNgcwGN60zi9fW2vC8O2j7pE7i8pEsXl1pJF7jGFFYMJoir1CEuSxvY1WG2aTL
ZKPjzPJfyQlcOyy3Rd2ENsbbkYJK0CtBwiu8Y4ONnVLLfbNV8OiOlHhSHjE/RyLwzBi5J+CkkzBS
ZJyiy+q4T2n+qygb5GcTWc3v5Eu5TUHM//FgMbjBV2eBfb4NDMY3o+MX6UNX67NeTAT4T2DQC9Kh
hMRUHtmzU0jS7atuBfcwBJ61RkWEqFXP6Ey4r4nb7iiuILMq9zw0H6TelmhKvZAK1jt+hVPyzD2I
eoMwl3nJYSc3bQ7ERgeEuu5ALEE+TRTRgyqrvCB7wd6Re/cYSXn1xwcPlZ4W5A78UuzwpSAazftC
KDAC/L9D3rboCO6xblSi/pxZq7c09v+Uh1b0pgjJlcfRgeS5LTCu1Jt9LbGiqeZdcOltEFbnpXL7
0X10JK3XUsSMYlSzsZi6NkBEt9e4kkwutEbBc/F1HMrl2OO7ry36SHgRHzUTKEC5Zg5qQ0vWsk2I
t1KEvfjxrUqY9KWr0fcRpuOHoIf2XuVjXs3X5r7qD7WPj1v/gm/ABRni6xAgprj9bwXfh6sV0BMo
6g4rUF+CmTEXGqsSAzjMvxAWKSqBepxcbhS30Bx9J4fVrADNk8rFBXNMZLzdlSj6XtCX463nWUQo
db3J39gaWwvpsXN1ffPaEfdgMY7KLHcpjxiffeYz7tQVf3peTQCbXSAmG8EN0mcsES5Dmz3SVoVy
tTmNeGp6uhhv9qBRjBC8nm+IWSWiW1vysPPkMsjHn0tfd0sHDN3ysOgn5JYFc5nS95JQfOH2ZO5M
agHgItJGpookl5kCu+X4Ux2M8hkDIkqz0Q/1wvoUVTpm5hOnp/0g1qHtuS0jR07/z/9dJRe5GJgE
imhbnN+H2w1mhsbCQNhfttsmdgKnYhwykmcSLguAxc9KbDMuaMU1QBhB6026LPIKAVpveYwEvja5
YHODvuaPAgS7ZPkTuCyAPxz9LS8E+tnmUPSKoU8mUkFPjDmVDzKSVq49zv5by/FlHHDuc2YUFmR0
iA/vTRDoIVjUjgQPCUgcJqKpkGPxoDjCUnsX5mMljabv772xGczURTzucnxc2xcs6FRRJ9BX6J++
CbJEcve0sMrAW8GR+lxJIgBQLfxxCPdvnMy4zyfghsUmoWz8WO5vwRYwH0o/HP/4r2Tp63QFbmkY
fGj/pgoNsGLf2CVea8Y/7JlqxU8tGAjF8OJWiPMI3xldKzEy5olg4MgcoxvV9kNK7i5ughxDqg7J
fhXB+uzFL+RIs+i1i7dfPqlfKzG2lpuQrPh1qc8rx7/0NcRnuY8R5vBJ/SAgCownpErdhkAzyUpP
3Ds/jOWMPSUD9EtVfjF0ZpYBYVI1OWYyokzcJ8MW/mPidKRL9C+reoQjcwnaBwvmn54eZpGV+n9i
iKhObKCT1apgbKESg7DmeyUyJjzaiUiQ1i1jobNu9KgTCFqbh1E3Wc2Q8J431QsH0SNt3N5hNMNL
+GrnnZeie28x6LQm6O743PcBQC7lQD7WWroOxh2JJ4Be6sEmL2qxjjuLvv/znTIfseBuJxdJsmwi
n19IsCsOYfgNY71fAxyGAqA6f05FHDV+JcOtXn0D/3074nfWWfGgOW7pPfUc5qKj1t4lRDDMIavV
zGbJqdQGf+tt93/k/lRZZjz76phgVVUvr1/MOUXwyRfjD+y589wnZ6BvGHGxwYJQ17M84JymfKMN
CDgqjje9TekmK1607kXFk4uP3DtlqV0s0WG/U3skBe2wOCs4QMWLvLewEWxXsYwAXlm2hO+J4Z/+
5JB7SUxNtJ7L8wpVqBF4b4a/XC84cQteURkIg/OiSZl9dxV/jPIhGdDD0TBmAk79Hf/B8O6ZZCLA
nI08g8TQtdwginr5qkM+UgLobD8lPihl7yjDGovzW3SC3Zqkme3ynCkQeOcfzlZrgUapF7N0qF7t
3Q3h1/6hXRoBnykDRcxXU/ybPYtJOk/vUlIeB3HHnEwi1/F3L0othCyC2dQEC4R22o0ks2lWfY2C
eR6PBWJo9a5G7/j330mFrTjLnLDAxnSMeSIdLIS4E06wQOkUnaTvLAe1mZt7lJ4vVAQTpjNfyE1F
jyBhb9M/ncYYJ4idKkBVqKeNQr+jr+ssL8TryNcBa77ir4+rWXEsF08En65+q3fHAQIN0aSWS1Xm
uWy8VsCzETpWXObEFThKsJ1X6KTYbJZX3ETCb5UWwL0x5rvHyrXks33Qe/QViZjhChs26/iLr0gy
NKq0P6nyonYzkr7ereB45ZTapL9CS82wefvNANybBEn8NweWr89G7wp1/tsJqsmQY3dUoxuYFy3f
X2DSFcPtwzap3/oSvVIS4NuSlyKKx4gf3M+W8dR72kb7aMTZk4igZRTpn74G6oIRXmzAk3idFXeY
YKO1TVNOvuYnSjAtaMiEPt1VjFpjEtd3ZNOHKnm6soxtlJ29pna+fXQ6jQga1QDm7nw/NKk2GbyK
sbJW1D2IsmKuIhBgQSBmid9dnnziswy5xLzE78LyKVnMmYISRxiP9NL5XxC61K0zH5QWQYD9rPYY
tfgycmmlj66FFphBOwlQ5lYq954TcBM+6zJsIipZiWCh9uOZR1rohDFQ6bM+upiQvjUelVXjt1ls
B59E1fplHi/DPignWA9oyi2wdQycvxo/WbvEzDfxgLZbeeuqwMaAYThrOwI44hEigMuJw1cV+PNO
mCXijCQVorK7zeSEqyZE9mdCA9FU0kIyM2i0ru/Ke5ntcCjgyG5yr0elUQT1AyBtyAhpvUYu+c4o
SUZbW4+QOHhYHuzP8fVEy77IrGXWrSDJmsulOPeMKXdnw+HKDcrvlWqln4HKr1XWLdzTOxJ5sYt7
fw6G8LgZQsHYvqTdWuB4QuWSVMYdy4ui6ld0VO/Ih7ehCvNxlRByFT0qDxWGvBRLQK6OpVV6xauI
WJeD6GDHCjoAq3npiK84wHbqlKQVA5FuxrR/7vGVYL7bL3A8j6S/wshZSXeUAM6HbQ+99p7QKr5Z
sR6+c01pyjZQU64lxUJYU13pPUA9kqbuht5sqKZyb1gQ80Pz0D65pIvY3/seiiHlxBPAExCVbSxp
GSbPEqL6yyRQsM4WkQqcilY0WtzV7sbpxX4wA395YnQ2BD+9IguhFUuC4YH27FYjs+K4TrzFK5Qd
XfqWDRUXQbvYWRnJNY2eTFFUli1D0OXI6B+4HswOH0wMeoIxddJ0ecso9BZ21jn2wKKCfFtYKuRR
vODZHH56Zm+dreKAjWSy+jAnmE+/kTO0MtSSeCjyTgsIfg74t0Vx4Slv1EmcRoX0h/ubcNRKXDCv
BrazSQL/Z6InZ/MUWO6NfiyP3n6YGAZIAUNpwE0dV25Dm/1K3DlJb3z67HHcoehAbFfMjJvx6Cy4
yY1ub4Mz7jp5ciAdaplrTFLAt465LjeiQCFoa9r8W1r8KUUNuC0DTE9k46brWGe9RRBM8w8Q+yMI
mmo/jLQzNHXN0yckgkhVB6qsXoO/6isMWEiq/TdQvWefaVsbwLwLWoo5PKeebubWbEpH+vGp/IsT
6Ol4zP8vSjci4DT5nvwvhxVvfxrGC1BZJqfaPNtFm5zpjh/WvlmHHg+KEpq8CEZPweyoiJzstIyt
/WDbWczDPV8VLEJU6jTkM3sIa0KUYHJSZ1D7ibC/nrYsC3rwuW4GQ8pTbJ7kL9JGOiUarBeJQ/VI
fkF8ByoRY126LliMwzk5ylYgCXA5YpeB5QycT2+XtUFGBlxs4a781nrg1OQiofO8NJo+iffjd7vu
025Xaisk7baTy8ofFwEZbbrOuiHxQykUnjb5rDERThmq1em0trMZQf9pFzJAnUTf/uMHshnbM9os
dkwa7YhUcRTqcTavWxr8CxXNNVAE5A3tql/70pmCQL3neucMvhhWBVxXOgqo2j6gT70KqE4QwLX+
/ha2LbWggf0FFSZW1MHDn9I9cwhlRFcQtyQSIB0eTNQ5bnD5h8n3Qpk5TZU77gcjjPAuItfRbXNh
kY+4Mx1txbsNTHAjBCUzr+Nu84nTPPD9IrcwzDfMG3bXZDMh+hFt8GcqVNqXBhh3y7xAqkZDRePq
2+gTl6pZt8FgvCMYPTa55AHtpyYRNWS6uhUQgSaBs1rKl9ROLMXvCZxW7X7X7qEcZcwygOMwzqIk
0puMRsFdFjFJsA2JvR1VriZsXKhxiWeZ2AWdOAhcirzRZUeRvWXREw0F80cIM6o3bPagpZ4QACch
DQls/XJNba6K8ab738L/GeOSwcFVi0GDpFAh8pLz2UP11zOL4WH4GoLiyruY6i95eIs/P8+DVRzO
FApHsMPqcWZGxLUCIHuxfzp8zYbvtxuMIrINOcBSVGRD0VGUyfjW9n+AV94jdsd4+uBnzFyDAX9V
parpT5XsydNo8ZehWqXc8R/Y5tbw4VSnyu9X0YscaU0z2X5TAe1Ocr017Zis/o+/hBivECgzrKSc
tbzlVeeoAKD8R9CPIedIF0OcVvT7FXe42iVT+zmMn617siXejrDYFIoIdg6FZu89aEnSghUL5yEv
D0Gb3GRC0XLpxu6FCA/+bJf7PYswL1XKI3v9kMX25qHl1mRuDjC8H3cvbu3mEDltifSeIZT1vPQZ
P4Gdr9Ym/g0IA1CP0H3wdBne2zdP8yAkJYWfWLnIOC9Rzf7QVhc7z2llvk0973Ge62+YKXJeo1MX
/eZbqWgIMbHEkAvyDIj3ya/528TRx/5RiTZC2eIZpZXWZ3Ltkv3HcHSQVTtqRrnoz6ZWUeQIQ73R
KFqP/D1ceJMcR1VfPgM2JlbBT7qRkhdA5IzvJTjEMKfBDFRQ7cvJkXL1BseCeMMvGwZMoLY13v+H
Py3LRmj2RyJ2uT80DvBXrh9k2TpY270b1aDHp/KSef2hBEQw/vxPH0ZbnjK/VjkfzJ4gJQL/mYXx
nT8PKcAs05gvN4kfyNsTcviHfnq5C5FZj/ZBPBRLZ3KyV7juiSPLxatpEvFfNpD5GfE7DPgMRGPM
nF7UaR/WQLBW8bPZ4So9+lwn9izqqJ4174LLIADVJSC9suEo2fDV1ShUlCUUEsi/6DpttHk7KKq6
jPpLSJ/xOw8SfP7Hhh/vG1ap38d8HfYiVIMCTg1QsnfG6eBM5hdTsogS4s12wdpz33BcaLpPe25f
zLx+sJN9DpNx99TA1EJcheCpOyf0j1vRIbDTzJLR9Z1ZSJk1SzgLnB4hpllRh4/xKNauMKxoEpTl
ZZ2ePgd0oxVDN4MQi9Xl0QbACFRP9RAAWHxo9BckleqknHE4ec7hN1SMgLyjqbQRByX3ep6mxqvE
Q3KqZpakZSuorOWyR1HGwH8TOXGIuq5P1VanxEl1jaVDPdKOT676z/kbrh5/AnFrDowN3wTCQfma
UhtE8YpNWZ9vhQQbzflgz9TYUop/Y+iCfSgbyTkdAx5BDqDAkGswsfS5E/NwXKb05qT7roNLNq//
ppYP5c/y/BDjZc1IK2XxpPxtz3dKDXXv+9FimZB4yJCFA18uApiQnAqz7APb6sRk2gfnT4w+aQMf
xZu1713Ajg2MqvF8TYlJCak7JLZBz5XLVaOddOl6Hzy72vWkjIcIjylCqMhccRNZQWa51FqX4tVC
VJmNt131ppCeLQWO0ttam89MkxZi79I8XsfhvMAZXlE1wceaR/oLEFJqheJiNDRypWMZDZowoLna
gc6nX9HI0f/trdhDBUKrOqvSuCXnK/+MHppWwO2dxzURWe/yU/pQaOWGnijAKM/sOH/UnESIVMe9
gQfbdegB8IBX9ErKLJ+bfMJou4BmkgZoF83Y1xbtkPOx7PB3kc9XBKfNtKgzWrFQG1HixcrAPEat
XTwhFvqNBGR4mmtkTgP9DAq/dkPqhLEF5b7rpyjFvV2tpBWiCiew7Kf37RaiK4VWIlHhNEpmHUyB
scjPTAsKzYNTpA+8TjPrQSbD3hu22cebVEZYec0mLTLm4JaarGT5CTB9McVb1xaxzJLNeq+TukFc
eYIlQ3OZMZV686o8ZiyItemvdw8W/WKmIoQzELgjcSWU3seWzfeGoFDorBwiJk9wSqeqzfzIv+8Y
MqKGQOP5iBTAC5q7wqrJCamfZUI2tst4eI6g7qpLLiIadJ2RHiSmGfpdCIVdIJ+Xp39qQTIe0hW/
GhGfN06ux3qc1oeZuB3iNjB+7UJoicPZZ5GgJgsuMmA9RlgFXecR2u9esZOY+yTM7Q/C7fn0c2bE
yZ4GiRsm9ojME3+NGDZ4IAoNwogESk2ZkFRThaNdhRV7AqIiBohezc43EdczZGFFgO0LlUruN1lg
llU+5dtzQ34u6s7GTcB5/8ZM4wLQWov7ilwHd0GHztKFOcABLUDzX7cXto4XoslNdxMw9U+boj8S
iTgjaeOReJQ7G8jPvi2lfyRxNY6vtGJ7hZ+RHJEe3t7xNCYDqc0VQNMxqJ817wosowALFhek3Bag
UYTDKmEQmeRoirTx5QfbFychlIdbhi+v7MKDkHJb0I1im/tJAVHh/cVxfS3raAFGz2++N4AdpI8B
ptLQAfQnGjyHqnINSV90EIbSIuoxefJUnxe59kJjdeadWwSbp0HwrRnby5GdCzv5i4Shc2WpKeR+
q7kAf2tz8DeS6bI5iBNdzV/+blDBugm2Ftkgx25oKEz3KAO8dUqjzYcLHVCbqBq41AxIDVBw/En/
wpVHrbDFt/A2n2twGBY9/9aI+IV7BuCVPKD+Nq3H5L7bPtoDUL7NCtNWsTs2KxgvNDUTljbZctKS
9BmoEUmZulqOVAtsDLiIyUqQuOys38uCFu+R8cyMcb/h4Z/pWNdnwUOQelbX0GgXamOWQps7VJmB
qGrhf9kwn4MWtZlh/tQh1945Nj14CEcaBylhgmmygC+Ft7QsXSDnp8tHoA7eMjdT1JuBsS8X86Yf
sm7qjN9PkYosePonnktEO0jPEn7NBn4UOcaweH0xrzGr1eoYdpjtjiHhG4RatfAZIEzjkp/LhGJz
jI/ZaxLGueuSCkcdRUAUAveAwxDhM26255i89Vt2GXnOvyP6wKmXTjWYGhpjSAzJWg1qLSPKNu1m
iE2SNqmptYTUgb+TAbMaV5RlB6WRgGNEoykOQBhsrZ1tefHYGm5jcoZc47DBrqQGxQrFido21JKW
HgnGQPa6OGQPvoydOVcb+tdImqyYC+reb6RU9VNbJw4Ot9aXgbAUmWtnDYC7E8KgTR8QZdriHrpB
dfy8U83hU/n8O3JsKzRlg7mnBDAhFfa3X0QbtJKhGOvlT8G1+zi9l5SUqOZiTqX2XRpqR/mcJLo6
Ys075OwiQleyzKDs+az6Fs6tyPG4MHQYsUxcq/GmkmioBDCUdLKoSLAAgei4axZ9j3HVG+orxZW2
hT/SmJGEP1QXCS3OIdoBPqrPbL+udjd4Tpmmza/dMgagsxlDldksgVqu8Mz4Ukkse80PCg5B/U0N
xCFJ7s7xb5f4wv0m14ZyHVHDHA/M9lm1ACkBUm6443WYDoA0SEnjPTkw6I4+Al91of4N86SjQtMX
jst7hMk2V7A1nWULfRJM+JcvZvlGchs+W5d4D8UfP16eYI+P+gOGYJby1hE1NoCUevakWqdDW2Cm
V/M2WAyPP04F1H23e6nN1e+rMMghXlsHsQgcT9KcZMCJsaborDMGRDfnKkdePjIjxnlHdXTZp+n6
J+lRC/sxuxx95Zz+KUz/gD4HJpo8U/jEq3czt3bM9XPALGmjpkn33VZet0tf/ZrDaFUcBheeetdP
88I1KdlDY1iIL6qstfC3b/ZR8QdbhFsCx9SXaKZIRIYTfk3l1K828Ixsu1ndsf+OCTeEShD9C1oj
wGx+2t8UOeMuwI3C32oGqXSAzfaCSTNiBGgJWDVHPswUVjDrVxb7TDgOjcwm/kOGEEJxxdHb/2Bo
T25DB+RC2vP9dimpaer8LtfZ0tHQBborFynpXn1ooBR5X66YdWzB6Hziljb++TvEt1PFe3qWxnhx
xCVUg7HHl05H+FA793J1jmrc9yQ/1XW+osdQ/G//C8H7WPCEg0mmMDIO3WOLYxq490A4QEzFl3wu
o5ftektph9btdbC0SU22sDdAslcKdc8Avl81S9Izs2mzjbSuSo6q+dJcqdpUnCtmLq1hxlXrlm+4
PczgdXsnPbC2DKPoxfJa7piVUGHcHR2fVA/EG3oKF24OD6icWbRKUh+cinJooiC/hGYK/+f+g3kA
qrUoS75WOsXYJV+PNsbyzi74dr7msoirZJ8oljHXn5rbI6v5s6OOLV7pKV1UtRI+D8z+W2L6Eh+0
n+sEg2uioG3n1WhLWxY4wgBhXx/JHRTUMKRcE/Rrt/N/hr9pk9aGlGSKg8907lPtlLNRxqYvgqRZ
KRYLU99VcF4AK1yUTR/OMCmcvEWqB+heFU9ObR6onbAcJVSwNtuamUOVbaKM62S7QQcVkUpvlwPB
GWFmoYTo2cloEA4QzQkqBfO/QeNY+3qaRHR2fEv4Yecom+hlwloYYWCQtOUNMYzOfIhzyV986P1M
QbK+JzKGdaQH2712ywD/TA8oq0jytKZCDD7TF69sOyyF/o2IaBsAAE7ThRoJuI1qc1D3VzuglV28
mCTbZ/LU1Vu3GDvfUgCxd6ZfeQAr9xTCIftJ5T6FnosTagKDLlyPixznuORKE+XnDcPWFuerGWtP
VK9jKPzlBs6JXoVPkaKEcuWVdPxPfFkDH+qR6apx4vfoTRtvZLH9e6dpkAs/TRsXZNuC2gLBmEZd
dKAKrMfhpd7d6iPTNWZuMVZChZCBxIVYkblFH7VPPXMSVP2WCbrgTWEXQuXyuUBs8wt+LcTQmU/H
6rii/UHJc5OwBx8aJEzoFB6ey9DnE+5LA3m/yahuetOkXR83jKOUiodSLof5Vcvk5By0eCsk8Iv4
vANLjDxnZGvfreAQa2NSBPzP4ZNub4A7WIoH6cXVSCApPtfPnurJ2pSOli/RJE88is6c+NRkpXEX
XHT2WcVcRlfX4hU0cuHC9XLz3NqeeHr9kUYyLErFLK9Cb+wY8heL71+Wy+gE6sSrtMXbKEpBxVEx
NHg8FktOEgK2K8vmL+gscpgDvUjxRf8MdxzTpHHcW8ViWL5NdPjT0EGCjYI2HWiSX8yCR1YFIn5B
pxD9HhMz2SaLqFCTYmKQumEP84zYRwraOPCIIDIWaSRwSf39bEATmCqhmvsQsj4UKz/0qcHd/gaA
EBIFkj9Awx2u4xcSfwqGj7A4vtI5x8WXZ2jdYu+j7qu2Z+nFlfmNq4RPDjUmjugrImNV01vPeNSW
ekXPAk1HD+Cm0lTdPMcY81lTD+Km7+TuUtgt9QXqe80ty+94radVDV14x8jwqm3WkqCUa5i9tkT8
g1jBG3wF2OSv7u8j6HRYJGO8ItUjoNmWJi6icQEwUligO6qpOEIgZA0a0o2wDpG1SPJ1ROXWoh1K
GGrlH0H86mriO1BmIMYI9OIRXwry1L/FV7GvaAo6jcETgehUpXiXyYKXD2wORxbvF52zIFlSDSI2
WyjTd/gdMYgkaK6jCvAcvtqjTiks+FaJYcdPhxk3GsozXji7N5GHutjxPjy9cd/ljxf5SEg87//g
35hNdk1/9bYHtlTi2pM9WBKI4ewhWokqWahXZdmgMZO++yESEtEIhaxbbCnVtWvI7rvzr1Wk/5m4
HkDCCigIJcRxK/4zdgIJI63xyrtCRNZfSb9o+yizyAnZhRz5eJpQ8iYX/4N5sJUWu/tEvF5wz6CE
4d/8HKwipoWksz/yYycUGpxDIGjfmkWGnjqhEgb4G5t/F6nr69hWeb+EdGn63C5uYj3MWueUCIKY
mk6mJg7GitQSFhg76hReCUjsrr5nF8SpKqyhP3dK8QguqHulMH1ZYGxWbnEq1STgrT9lhRT+x6Kq
kPO/h0V7YrBTvtLVCVafap1XlgBsRyBIaiGzZgZn5Gi4tmx/hXp7QWPyC+hB1ZHq1GkQ/kRgEOgc
UTcL3QLJcvSjr+dSHQJ4w2+6RiYkm+AFAoVT3nBHQgb1d74K795UCtkgD+f/vj2ZcjDEv/xF92Zl
JcDthdlqNRkmqw4AX95A92o9Umb9lBwRlbzG9dI4ci9CK+EHup7nXSqZMVedXZAgbnGNH61KHjjW
a3QwgnbBM3ICQi32gBxqW7MBGZxNkEVs32Z4nphn5U0qvcgnAVNUgFireMRBvWnr/Wrzpr+S6BrJ
L/7CS5OSAp5m5yI7roWvuHnINiogH+PuG0IhwL8/OQb/nLiTR2enyKVEUkmByzyU37IfmdVfcHvY
lg7lEvrXW9uf2q9gJ6GF7hTaAvig1sMD/Awo0+EpibOm9nhI7bmIOIYEKy1QSOUL3mxFLH4RkxqB
DywcwBytTpf+OYBNfjgz86+vMmm3RiKTDTPglzg3fyWC2hwnc8fWeJ+U9qb/drmqCBm9kkDIpNUM
KHSFqBPjjq9/osTxIwkxBb5wN8fOS0M3kvTWUju0C/+0+bK2GQ4tl2c/USdZbKU9yBGLxzAXKgrl
zoZSXxmu+ShOuLbG9NhW3mV+eqjZP9suIpSUDfo0qv0f3UJbowTf6RdoXt5hgHQyBD4BMHIjVIAj
m7j6/ssoV5/Ar8H9MEVeTQC3j6bA7FQN6yONk5EH5Yp6tcZfEXNJZI1EJtwgYkWTxSVT10t+NkYw
MBqMRF+szJ/pQ3vVXLIBZJzti04MIt5Pny71nDsrzEvdNxwc8YX8R6sIUEOYt/60fyUkCtoskxOv
th9VPBGunkYq0ScoY35tZ+mAo4J7cYfCDorcgx4Xywh1VhofYj9xLSNjU7uAICVUYd7dpWM0Zm2S
aNqW8YJpdS8eIRRqKamtVRnMiBqOJ8osvWnu0V+VPwRT+gh9F7QlfTUYeRL/XTWkfRokm3HI3uRj
DgD/BCo9h2wFBKC7jAZ1OFIScoTjQk2UAhtNNntgFQdZGujtR9vqSZe+gKfksANDm/949dYcOS14
7ImMJRFt53V0I3ikLixOkPJukI0qB32uDeCnlxhZLHVTeRPtPujYfLCMNILdlTC/99lrIef9VXzL
RE0s8026Tcd8vCxKMVrzQKZGCpWDqT67dEYtNvT+cDHOyl7uenmx62vbRdhRNBTyOeMH+pdjwQdM
sp5Vx5Cy70U/IrNnMSdqR/UGAPnedhe5HufqF5KpulMXkfsLtayHhvY4bfivY5A8wC+IzTyhKDIu
UfylDZAzUR+3h/T9wWRahR1G4FnCcBDz9RVXal9HdgULzgDPFxXPs8Keqap+KC9injiw7K9t7fR+
pNRIuxuXSE+QMp81nO4mApbwTe2k9UIOaZdS0wSS9o4G8AR7sJh9hfb2kl62+KlzdEy9284aUfmf
Q9Wf8hvfXGOvzci3T/WIlPxQj1YKiEMWVUUBx8yzuAXw7FNNVQs4wFLI6b96k/Q/2nNlLT49rhSh
ZeK+Fs+0mbU1sTqphTw6i13TvKToi6VFuyUW50nPNgZ9VeOnV/2S1aajapa4qe+uVKEwVEaEnTLe
+F5danJiXSvtI8pIvc/+jRa1jhIJ3Ym2C7TbgRv2LGU2+6CXquLmh/jOVWwdjXxgH/V+GqUEU+kD
RvyYg5+L/9bDIo9iUE3yiln4Box251wkRrFNAxRgYOXFSGTa2LQ26uQJ3tbxnTIOMm9d1ATK6Wbo
ZTeEQ4VF4Np35ZLl0emQ+2FY7xVhuprYrThVJLfhVjI+KZmTkzYLcHXhzxSMnZA64u02vHpQvGwf
zhqHFRKGcgMbDPeVTo2sirQIzDZCXis7n0mq8hD21PXPkg5nKmJriSexjyCov1nyi3Gsuhz9NKgL
PcA+jC2h+7qW8XCt9yCu9tlMTlEPWBvmNy+ttx1jJbueRbvQIRNVfeIrxxs4Of1Up9MFdidJNupf
eOu1ywY2+pC+bZYvkhDV/LQJhosJpCcypgmdkYtsrE1SHek45VtZ9abAE5raHBYPn4faWnGFBAai
4nGXlwqXLd56jMd7Z1CRLs7yq0nI7LMSTIDyGfo2m3K6k8u8pn1lDIRx5f4myGmQoLFp4rV/1QJ0
1C1JiqTAi5cVYlie04t/aXWFGn1PIZCaPfsG9a0s7UMQZqj5Q9RJVm101ghwON4ouYllOFa34sXE
XlQ5KA6VbHmPcGh23LKU0UMPTEQHhA2arUG6EZw3BvyVwdXmMiYDm1F9LK6fvFNnkTFSPZeTix1H
gIKn8kuagwCDGitTYarcdFRPCkl3HCCOto3BWiRhUG6HQtogtKetQyCnY+uBqumPcODNluv2K92h
BtPuJHtPnbdMr2H73NTcDDW7fk3LwOi/7X7Vt9s8i0arVWKL7DS7wHpDv9EKWhQotDOxlF0wHfuC
AeP45F88EQGUCyky/xVqWZBpFNeaxMLgoiYKJRgINiaGg5HndRpTy6rS1agJc7T8CBNpGWqs40v7
J3t1J0575KMeEYevaonPyW+eELcEKw2l+6KbMXgrHolQuBneYrEvKB807WX9mrS4VrHPJ7jgeObi
YcthcaLefB5ZSK6cbW+e7/867uBvb7zgab6XlUwjnMa4qGzg0CaLf60y9RGnat3NV5TeHtjwCwUN
SC0yyR4BMy5vUXCKm9Rt80IVDy/FFxADAp8sDBpTI8kfe2XdulETI/jwjzoLYL4jvTyw5SrBhNza
56BS38DEknuUic93IxLKhU+peGE20QBjkRrDfiAr50UKn6jb/6hK0nDYgD3s9I9pB9yVuZKom8hD
xOrH60h3acWWrZkgA8295nYnfE3/ERHVrUASXW9yaMqVnwSiQdwGtKrt3xNcwa8msVZ+myAe+oz2
otk01Dg4rlYNr9oDbw9HT1R1V8irGm6r90rIeQikEpHf/Ie5mzS236GebUKKKEZrd64JWx+dZSoi
qT/5jFKeFMrytAnI1XwQlP1U+RrsNYff1walZF674iZl/b6KG90UYKc/qjl08PPJQv1MXeg5jURJ
vdUDV8XNI9mUUNgrop2nSxVVUocvvSsTYj1VULmulj1hYoS2F1lNYTFzuRLek4RK5Zmbkdx7+ShH
/bjTOsUmf3Mik0Sh9QVADuXZwmvF2RgaPuJdGcnWkd/aWI3ZDlmErrCzUyJL10n0dQBhTixVCR4h
q/jdjEnp27afIunWLYF+gIDUm/jD52ZT+e5zN4LH+bmxz4NCCwFbcM5Ym+jXg78DnTqVLNqwdazU
PJSDXaWFrTvGq8WDxPgjMNcsDmbEc8lzCxH54FrW7sJSXE22JBMMD8EI/CSND7EfeC74a52yWlIJ
Htt/oBRRdfjurUhb6/sNVQg8qBlVNxDEc77F6kX6iPFJDdIvvCKS3cbPow+TDD+6UZX4n3hUBxTj
aKbfsaw57m5AdYf5gxxg8t1lBbBUUwfCG/pzotgVBFjZdQTqocDlr50bk/zHdmLB9jJ17SwJXi/N
A2Dx47Y3hEzJ5V8MfaPFfrvmFQn2f8htLgATFpYY5FGjxQpBOGuukzXe8waW94B8Oe1z4JyBVOqh
natIoaF5Uf8LIGf4GVrCA2yeAOUsoGowhEsZg3DOhLgHrkVx6vR//HOSgG9y2M/6f51WC5VkIVBE
pX5b0/xw+ABZuRY//9RCrUd6LY1lSDxUqAkTnx2VYL1KNmVE2JDBrCUQ16BgsXODxyJ1piCcE0o4
0TBeOAssCaVwd3qSMNwvm3npdUmp2VPnk8ZK31BJjBUQRoGREon/sXAE5nNBOMoV6RRgnYn3C4bC
g536o86WCxeAnzPqGoWbuRChxF4Y+OfOXw42yP4B3I1ZS3snSHo7+F7uWS5429IEOClqC6i78HNl
vhkL05moUfmHIneL4d3O9z7MjZxa4c9gY2586MG25iRyQ8y4BIW/jQkh7ViPQjEmfLtHWiUDTjWX
vebHHWRTRLU4tAPO97bBt5hla1qe3LAWD/qYTsKfTslSj8UzT0xJu/3A9+dkh5Erf69xdFrTqu8W
hwdU5XHmBqqW9NDIyVVFV5gA53LtHhw+PsD4PYhMpymFAWxUlYWm8fGBw5n6Ls9a7eKQ8/upIIzi
1a2JVMBufkubfPECcOXTi/xOxrC1L+ObmdXlJ3s8D0kh7foekckKQ0Jf+h6DQOTwesu1oPKmcPSx
GisNHN4cuO5/MIH7GRHB/Zghk9RZFwvSaGQAXnO+LIDL5u4lXr9qU61ZWh1uCBdjLh9AJcKrNNvJ
ZgIplRWxKW5lgMf1dVVh4g7TksRjGMQ9CGDq4ZrthMfVB5TMH/L0sGHvM8dNaiCAVdbfyOp1DeU0
Cb6WtC7lxqAuQTlz+yiaBaaVcjkcS0bDmv0N2pfmHuWzFVf1hBcfNCFhyOwGJ6Y2VjYq4D7j1a6s
luuEYF+XHHBjQCxDM/cXeQG3wPMtEXT6ulN39Y9yJEyyG4XWjdViYVmzId1ng2VldSOQcMowl0ZJ
G2wBi1A3PnNXICMrs/S0GphDy3ep/wnLz5/c9ECHXvf61uol6UtVRtoI4EmYWYHWI532o8AGDRnc
681AOZogllUr/k/fkbzeX5u1V5M77qmvCbmZ8lpDTsfXSI9ugzrUnjbhbNeyPPW/7rgGId5eOsLi
B2hsfI30RYyXlgCkKat3g3YvWdr1lO2v9dSFU8eJ9QsdWzLcW2oT99dC7PMmWX01cosg7Yh5h5CL
48ETG18+4GDXAHIrWsD7bEuYg/ZruCNkHdkaYeSUL8h53uUUUgRcsetL/OBUe5+ALoIDdUUHwfxy
hI084R8qJDiDyXKxDopYA/R5xGVTT0itp7J/R61gHAumGgycfwNN/S+VsFn6ums/6X47yh7gxN2M
T5r6LkBEQO4GfNmm9H22qQcbxoVBkXsfTipWF4P9WsTMKTZp/QGuzPm5VOAorz0iwuEoTsriBFJG
v3UeSKSHrUhA00q6BJosw2tcZeNXI77NQO16iVVDbia9cGyRMRxechuWApI+oEeyXPm2aRx76Qdr
8ZwFz5vzJb5FEWNlninXuHoWvCcxmkFjM7rt6cxM8lUSzuBAbyBB/p3GFKHbK8rsDAfljM0jtEHD
AFhVayw0fJyTdGj+48L0JvzmGZVDOe9aw3uS/Yie3ixgweXvMP8sYhTVJbJJv7jk4/zZCpJkAN4/
Wg4q3cqTbVPiP9xCaxs3f+LwnK4TlGN7qqlZzUiox3ex+xgckBXWpibQBN+wNxyfyxiDO5V5oxsY
jofEp7R/13yeEKY9KnZqtuZfQn0lGoc+a2wtuC8zNCRsYntOunRLm7mBMAEnhL+JRyjmlzc7jdoV
6OrBCRSN37/6JvAXbCTkSjXP0nYYwfxxZMWmu1T978i65uJCilqKFP2qTp+GiwcAcdgzXh0LrvG8
twY+2awogKFNqasc/vnPEuqGO2Tp0wrncu76oFMTIe7vawr6S2nloH2z4Nkds36xhOI8y7fwDFdy
+26Ok6R75JofsZNSPIYiqmbxV9mtUtprbk2vPxzLbHfDCQqndBmb2Y7CNYGBIeDJ3VrEYnaOI1PK
/XxTzLA6GWPqLMPPaqo3JHjlKUOsRU7VL7EJglafvnoQsxP4KbVapt2DvaC9xsT3tIqd8sTDlonM
rcR8zdBHs6iqMJbFxe0qt5uiGQP4UWSuXR2GGbUVnVCvi3MAG920NSMhNGIj0HayReBDupsvVh82
wyrHqU0oY7SktHILgwMxjYR8PYPFYNYmGhAVuZh95cDLNr5JpWq6Hae8BL8Oxz/WfhWp7CBOtPn9
ybZvxu4egoV8p0/U1VuBI8dffbHfeQHkvF40KgABWPtrcguzO2VVJ1n4fgdXkkz8+tSMhRjt9sqN
qcJwp+Tfmkz7aC1MTAc40jjE9T7pd4+CCKrVztNssp2sHNtwQ/OGqODqjpLsCIn8Ph0M31O1oUoq
fC5nDRmE4Wn5g64FE1pY76b6HUr7DkiyXht5Q8X22jVoauFvAqoB8uVwf4/ygxmXDiduRcYuzV7w
FXP35DreCnca6w/3bLzcHcqpTd+llNGevQ9XKidpaGm5PkFd4OUfi+nq3eL4tPZiWX4Y83AN6tAn
vOyEG3+FR+SenpA8ka9fbjpIDYjEwtyxrZ2R0PKtdmO9cWcoEsVSpi0g64Z4bk162ZE/HaWwFwgt
tR35/sh+gxp13tI/znaBy7+u2HOGooWfXv470D+yBxMi6jv7+5UrviWo0fARzxeZ/PxAZ6372lqd
yXcp7w50aAsd4lrsmcZYJznNChzEAi/thjPSzrW7M4YLriK+0HzS6bTc+Iwqcc0UPZnmKq3odCLX
zjrxAGfJGbdPXrCnlLM/UT1gunJg0wHlfnUGQbnal1tQ5Pa1gnsneIZPmCQkjRacg0UxbhmJRFy9
ttTA7w1quRSqkoh2KcQkHSTbC8UDMGZJzoQ+edRvaIxmCP/+MkaaLj6ajHYwMr8qXreKST25on8z
4lFqX/wjseGDWZbS9JwU6RB3v8NVrk6O0aQD8M0Z/jdNLAhedK6BZlVh6F9xD0VmM6MhY3+JqTx2
sRwK9r2SlLgdQ5QvBTmKfIzltXkm/oKsTzUM4R3wTjPUGIskqX/Ts6HA/4zz2ew5pHPh3bp1fMOC
dhZerTzrQBVs68JpxgBGCCkDOw+OszTv2Hp9dafny6qpoIiMzDWGeFJpUSNK/n7xXNfVGG6xp6vI
i7ND0VPyyXnot8IdUVzzYWXybNKb2zGD9ThFn9D9V1EqU9alg1H18eBN2l0c9aqNTy2y1oG5Ptj/
M5IhQFncMoWtcL1ekL6dGXhbnECE/v2OjuEiO7HJKoYC1l/h7SXeZUFwJsTKEkxP0gCWzO9TEroA
vasPp0ihs5zIZv69YFUujdKqMZPW9sqfU6Fo2omDjRAIp6MhuS+uP71pyuJiXVzHpuDCkY92AeY6
QoEqnqyhprlYXewmDxBcbHaixCWTMfGHpuLPGrnhcBiLRh97RuUlQcjb/EzJLvCIhJ1sWB8eOijs
jyD2W+KPq0or7JWk2i91pCVHvxtThaVj9CP56U3lm1RzCURmAeV+9+JjKsHPIuKMsf2TwvYqR9OU
HDCRD0UJK2UZ98ZD7R7dRp3sC4zXmk+eB+hfjv7hnRlN1Jf3Rh3lx4vBTEAiCKWj2cHPB4boMu1i
lCkYpNrfSUU/BIQjATdPlHxZthuNRfXaOqLVT1drpLqAVcSHP69mKRbLcdkefdzOGbaKJsvL0cG/
K9/TXwvuEqdN9YvHLwaph1Pmz5bdxsBQwFu3d9W0nOe1wFztUY4pzBKFMOht6PcyDO5QKr3tgJSZ
tqrZbe3B+M4atwHGXYCM+mJHLl9rJtbETvROY0l2D5wi7xH5nNVanVzArOg9KgBwMYVyWh0BsmyZ
mJEDRFmA+6LMLLxhYWGf9cPHBOPkYLij5GsRXJe90jQiovQG6gdOBhucuB38nx8DMqnk8EkyGZVJ
XvuO1wYBGP1fn7Tap8zg+yMNgFqpML5pK+Iu3epnWvBaiM8XZG3cEW7NYj2cVyx7GC6dk7DBsQTo
2biFoBBBtALJ9Z5nwqJbX3mt4KcCNS+QLxu9VEljLzJqTmogIqQTkBn6cw/SH0PmfmFTY1E7ryEr
5Zx4ob76fzMJKIaVuIJ8q6U7Ji23DLsYIkDneeC4yhrxUamdGgcjZRvkOH/6s6l/dQdTVkBkpBVt
Iz8yj/jZ47kLUOb9PNBP02/rIMVYebRDtiHdAtjbagNYb26w4icgXAC5yvp0OGosWiyVdwYZpP2/
p0EatPJ/obYP7fTfQs1LwF4dW08LwetMuTfSKw40WruONtUdWpGHEFigJyb3EUlDxvffpBF8++3g
RR5N6wo7StcxBoSsK9PaxI8O4k4P6couiyTui8OBNn2QIuuJ6JbhZHAE7BOBSDnCLYGj8Yl3fbGw
oA4fyFpDGeI/Mbsc9o+tUFUVHL3NlRdkjUjQClgCkVcwBuln0apf4Kul1Ta94Vyrw3V0dJl+QSrP
u9gSbVXq+MWvbzCNlbYwaofqX9Tzetaqno7UsHV4tBB68uwj32JLuLk+V4u109VVa6Cc+8fBFQdZ
9DOYzf8LJr4owLUHmRdzeBkjIPdhyM5sAsvDrX+YQ39T8hA2orJGfmBAetMHq+EOpLDmdnszES0l
6MZfxedWWFsOLh2+iMOmuxeeolBASlpdx0QY/lVMQtKERXTOxsoB/rPTC8/XwrSISOIjtitPJD97
ATD+kMKadhGU+IvT4ojRVOdryJD6MCKZk8VUwQvH1IlXrbPZstk9g1mcrOxEsGGjZ9qzWAprsPGh
4NYHoXx/dmwUS3gUpAhQyuWzzubOqtBeNFt0vvxIykRvH/d7jndC4KSWVJREwwdfBk54F6kenjP8
wYMh0XlYUhaBj8JyiXxfcZcnX464CWFWPbA4CT8tm6TsH3rzSIlEMgaXgeMBHCOqYL+vBVCDPWP1
AEQcMa8KNitazrmiw2p8ZUiZiYjFdW3g1Knqd1zWYtJ0JQHA/rSIm5Z6SfPsaj+a1DdZSt5tz4kn
Zcw2q2olmQngseiq8xN6BqOSqDCuXiTPcq2ANNggSgvnKfP8d6kRmorwdk0MhmZRUW7btMEe+2xL
EYOqLZUYzwL7FJdwIedEL9GG40Rx9u710hFgvHRWyg2DNKi/54e8oYxZkhmLguCS/yZ+bGCOnZbs
/waPc/QXv37eJQylPE9huUBNVzIKbYNPBAuSzkCNIDkj/r/2WqNgfsI1Nt10gPLJMIFALEyMYXXV
i0pxB9QEbApqM4hcqwRy47u5GRahpnuZCsfCttvfKHKAyImXj6QielV1rET4FH7WKXcaIyb4fboi
6nsP/AUDZPphQilCXcQ+WRM2WL/NY3LUOP8xFC3dZEFed9uDMkXoj1WOTuh1BoY9MMRDeQzgd/Ul
htI17bBPNu/0PBuWa7ewXsKHDjVJ/8Cq8xMTmZEiBGxAZN2QTVohJdMEdLSmevBdPhRrB7c2R5C1
unr6or3dKbuH+laO5Lm7A2NiJMiho8NDy0t1ayjtq7OeyszzPq+aLxVXslnZxV1FngQ3MDkKBnPO
zanjDB+C5mO+c6cXaiMR4W8JHTCeOxDzpMtijHth0RWl4+CJklw6sMshGdjORFPCDv4WdqgN2oK9
/Q1EmpQfkf92nuHMZbE0qRt6WcN7JsRQoaJX9Xmjc3lUszijziuUsIPJ5GGykO/wdcFkFJqoKNJB
nFABkrWyVDk1DMHgpIBd0tLm3YiljEPKgClLSVAxGu9av/esXNtZvSNzdSjSqdGCp77/AhIqmdZg
HJWrH7E5i9xsmxKRfr/4P+F4YCVARd9UJLnaTncPQD5UiD3/yxzkAhinAhg0hgrnFhzDvqBtUac5
8DvSv3dfUbhBy2O0ozWH0ZoCRALx7A/yfID4VfcQgPkYzdAk8dKOYFIvChf/fTMa8cYMNZvMb6Ju
g8HlPlAkZveVkQX1OQgHKeGqUS13Oq0fhrpAqPhcnjL/JYvC0HXdiq6UwEmEemf/ARQmqH7V4peB
hkoHeFXyezZNWniVK3QYDQHu4TpNSJYqt7LB0aYchMtBtWoI0tH3lTE2oYHVtwlo2dJNIKMx5n2s
kZK0ja5VFw5cGjuNvyKJXHG7rXLn+HV9D6AcRU4DtBrs2J9kyCnfGiQ0KoHknTTh8svZ0QjGBTRp
rvruGMTMESNRmQt9a1UOxCdGnB/fHpNhKcCeThTgnkqCyscDqauvSS5XXCdHU3H6vPLAgmXiEdks
CeHEGnB2//HGqN/YqiKUcY8ZnOL+hhdIgE+END4MB9eiX6kTn9o8AuDacPDByp6XdMIrB3EbV3hz
jZvNeycirXv13sorUNe2y6fqz3O65Ur0eYxWkfBMgZD7qZ+NDqYqM7H1aClptl8SArwAeJYJ54go
d2N+b0tooavcPYGoAhYTcjAYpSbzPJXPzC1yxCVujCtwfODg3ooyhSMrbVljw54D/z0USTxv1R8H
id1K16Npq+5E7rcNV9LaAwtUJmnzidu6/eaimGD8/GOIZCI97CzDG8mO5vUji6FgYtYqR33MxqKe
PiYK8VY6EGJl6avhFjNh3Zsys/mV+ABZ1w+atvJ+625vQWs1ADD+RddsoTjmszlZvGL3GQR0VL8p
7ejMnsm6CJxkVVfMuTsVePhmEEtI+wXCYJI9t2JmJXuL8OZaVmoDIEwJFrShllkJS/vpbFsULApT
cYAFMCT0cwfGpLxgLjygFU8gHPE7kr7tnloIqRI/qEQUhMtWm+2xoKV2RxXDsMwwkvEKYrufjfJd
kzeFhif6IGtBgmK5vZ8ZXBciVj9LljfIjK0HHUEmey1uWVpwUGKBzIhYbnRZC32DxT5Wz6/rwxOl
a6B8yguenF8NhhElSgw0yaxyAIVf0wp2c4c6wwnRpjEKW1NEV1Ba1WV0yQ3PIg0WERHuxjePvaLh
ol/mLpJhaw9W4UIMCC27q4bX/CzDy+pDd+4MleiGovF8R7nP2jVbFNqeljTV5KJtZPnjoowS38/I
S5DrG34ugH454llo5Q/bOjH8MHCWFHgeE00IeuLHVkxYHi6+WeWD7TPmFXUw76CgD8L0t6niwtIA
liZxzWpVmrxTzNFjF9kkWOiEhQaW83Jvyyh5PrK1Bxj6xzlAEJujPiJCaKKz8wA4IkxLaftk6uZM
XqjiPf5tj6ySiwDPw9aUpVBQcWZo5v3r/9I0D/1HKLws+19uFC+smSOWfawhmYlVW8qpt7SN5HE7
L+vTHGdT7J/V0+cWoIs3KobBhIECT+DoTmJyLxfpcU0076ikskVNZnt7VhXuZh2c7M8F3jNm7nJX
MJHvu9IzDgrLH4iWSj/C4CKInFwqCIiT9/gk8BrdSimH05pfl7ufmuVz9Fxl2syw9AlVL7cEuKrC
iosh4jMOr6bZKQgXb7RMDt3GfYkrw9De3D4840HXc26YEh/nLqHpRT6HDygSUBvYb8J+eEZtONW5
auLaVX0NnceZh5Did3pzj/yd4tHbax16Hb0iSSsZrtIvzfvqB/cXpKa9N3z5RZLS3IGFZXKGCali
gMtcWgS0MIeSEbS++FXzc85tPs9dvXjaK/581tg/3TireSbUmen3oW9PLBkDGBvkg0SnlgDtfDiJ
V+i4SojKlX+QCPA3RKSlTT6D4UmaddCleEtKhADcXlGWugflzmNJ9+UUgNoiolguw5jhfWE4Z1Hp
3bzKO+5PVSo//dQLlidleJfLfVzCPfXHFVUj++9Uu7NyKU1aykYTEt4bvRiwEIeVpap0pvQZ/8/M
jCGm9HnnIb/A+C8593bJQ4SPINpL9mXhUJ0QQBFktE4P+pfp2HCdr0WB6YwaRBT61T76IQAjN9/H
hlR76RgmPppsvLrmLbaJsJq3ZVxapYzE3EebkKOMfQlEY4P6ri95oMjeF36OxD/kkWfeSvR7+r3n
/YS6iK7GNLu2y8DGAz3R4i1r0xfXRV2GOvIRq6Y7k0I7gg+HCHyjcRl/CQIwCZhezZyTOXQMoV7W
VZ75tn4nzhy2dVoFlsgroau4iji/D/mTJrqjAJbRY0/Q+vGJJa5TbTprBz11OfT8OjCcnIhons6u
6oTN1QUpqgIKayLdfMPwmblbj1Hv0JP8Stk2HQVorATMSi97FgtMKTAhxV/cLDwASJ82Ugr29CGW
0c+N9WI0v5FHvYWrvrBszNLvfuJs1PThxIloUl96jXWDYinanGR0R2+kjG+xIYdYkgUg5PRVgyWr
/sG9wCcoJTSiWe0RjkEVFgnlh9uLFD7qAJrpFS9MQuK+4FpaQhNjzc/gdDiV8vVKVjAUt1uM8IQU
NTYxslBIl8/2brrfKw8JRASjnWCCjhhXwaKCpYDxiGJlg+ugjlNo/k9t3oYvXsTDMxNs9veExVjF
lkiaqkxPTKFAjECIt4uifBYTZ/uJDnq/hwIVmNLUQCpFzyPjs6ojH++PygzXsZWQ3L7dVjjvji/e
dXW/ZZSQLiMXgzL7LA+OvNv+0JueXuCzzDoyU+G0DhhP9DQzTjQgisC0hC9adOfr8qJBveG3Olrc
FwR0+kLM3JfRCJtAgtCv4JOlJmhRp5a0iTBE6W6LwcgYWXZQvayDueuA08Rp/rQaURfNt95j5TvB
0YHqOBOcBrjCKLXcloU9pV1tqCWElbYP1Ut/fBTz7bIt/Sl5X+lMOeBLl5WB6Da6BnrqxQM3KsXC
wmqGr82Qcwn+W7WJWSJyWDWWojltiGwKIxrglDbK6xUwbO7/8HOxLwFAkLDKV5vU9R9hdLeTokn0
m0m6wbgr8b09XfHexpPeou4AJhXSZBSqL5giVJhwRyX4UM2LBWyEB54QdumBjzOl4glsMum6zebl
H7CQYTMer1bieunYHKmYsPD8bGVAIW+D6iGP6P5yQPePQSWA0tw2KdyBcxFv76jo25LpmzqRT/6v
8FsRFf9xj/TpZwwcFFH1mBd9gG4k09B24CaAghUFIeWYackFevk1JJFDCSGtAlL+oyfANdPpYCzc
06xBT7Qv/T2Mv+d0tqrSeSA6vWJka9BK26CWfD7TrhuLiBTQRT/GXfqDw3jvNI6V7G6fEFBJ5RL3
hA+NP135WDb2+W3h3yeNWyFBH0nZe0G8XL4zetNtG1m/VdAzy4FB9cjJpgvSo1S/xWlcIXEG2NP7
8uyjC69o4nIMWPvh7aQYQ5MMo1DB6dZyR6b6OCe1U3p/AE+TRFJxDiDViARD9vxswtTco5n7tQrL
zdAbD/tcbdzyACPXVhU4Mi6UUqZvIHrd9cLtzAZ9/ZUVXoYORMMK1byJyAgmXOxR0mQTThfhJ0r3
8SY0Dp8wbrgDJS91gozLN61dzOJblYjCmbFmS5ODunP/fcu42KuDcXv9gWO3UXMT3WCqh6hDH7zF
lpTA7njksg+n7n+a6Al0FpFgkQpOwwlLJd7uVxaJsuyrV02b1iPWt28nSVGYwMCd769XSWOk65Ei
i2hMoxhiIJ0rwjV84hsJSm725duAG5WSH45cWlPRdDFe17R50xoVI3Cf3ccBFNmkeGkMuZUUQYs8
2W6o5abMWyo4xVlb67sZlPGofoFZ++fn3xfvJso6I3IEX09oyKIVQTvCHSgKzInzkqLzKePW8sX+
BzeDIF0s+QUL/f4ouGReKvUrhu5prUdvdNezYrdckmTG9jGkwNe16SfNw5lWtnLTICFWbA8Y/cUf
xXH8QWQC47w91bJjbeFH5Y2z7TArJCU2fhmm6Fb4WXw6GWTUd0wdkjVnXp72UVmsEd31jYzm098h
hXi70ETSIX2249H+b1tma6KlEEOAJhF+g8fubEnW8NFFEw4zbIVklZAAuDb1xJziCpHmKakGT3j1
6Z85RS2PhmdJhDNqacBJJ5QtNMBb8S2WyzxmJPZOv7dB7iQYmatUS0q8ej7fYvPXlNgX/FedhfRG
bMTnWgcG0DM6t4KafdOx3ln8U6TLzv3sphVIKYXtdLMs6pUeMrreFLbjb7oJCFPHqzfyO3xCE/el
wl+NRozGXxeyZuE5xr0R2L735WUhAORGHHtMiGB8mjzSRaHUvRnkWjv/exEzq5CyhYMmAc+Clt4u
YDh/cOMRM1ayX7arNIYHWF84Oq9r52OI0ByqtYJKzxnj9SUXlMKw9c/dS/oyImtyfwqGLoFqWKYo
XVwxdfkzYEeRiRtP+8BU3ioGcnOg+ybZOTaFNMECp/aHaoYII/BpcpcIN6i6CkM16FlZgtKebwZz
nwDWiVQAPbATgl6+NINf7mlLu1Irp4762XBZVpe+8YvwZJL9KVvTDMjeIWkjbKZSOdvfL2mGbhTY
8BsgMHyFiqe51WjmUWZkbWgoZY1qbGOMRbDAZ9tyMPNuLwFlqvAZySE/ARjvOI7dTjs3fieqWKCz
xGYzxZROuBBi/cIkWRj7Qgzua+hA2VQsKVBmGYYG2LjDVdAzfHRpNtgKBw5PFPBK/EZObaRdhj2Q
sOuFiTIGnfHaKf/0VzXnmNTFZDQl3NA+yaZV8QS9gK55kVIwisG3oR+f99K8971iv3nukP7cWdB1
4Ym/2r5RB51Cy4YFWS0nrw52ehWBussnX22qSXsGPctI8a+S6PDhT2TFUGnDm4uiOxtspDo001fw
qzW8xQ3nvElJ8zPWjLUtGsBcltjRHoRyMVGrPnS0AcZQhmVho7uJKjnkC85IYlqDbQuAxzprqdN1
/nH7mymZGWaD1eTkZhgFnmvTn26SR4arbVsEJMs8CO8BOMfHIXnl9ELeYPw8VZ2dg7xsoacHV0ku
DK6O067NyR1H8FfGrGO9uX0RZs+N5KS8a5jUV2GqyD9vDaO5WEeiD+omHnOiy9WxZ2JUyxODTFHq
rR1PXG2I9/kJ8ycvMZ1L8XQI5qdjGdsSKBH7XocXpZ3dJJY04oCYoviePrCYY6PGNxs/Ut9t+tbT
gT+9Q/XpKSkE3XNiiILiYSR1wLQgHrYi7oc5i0yPOmSYUmb1StiKw6BQ73BN1xxKrllOT5kbqoCW
mW3NpAGwsbVzQhpVG8x0iD+NhxBhUDZACk7KwIW7TTHlaqQmgtmBhNEo9K/JLGFUMGeya4m66Cms
qQMcO4aaUIGF6mKaa+McHS4iXlhYb4BPPVlzB4/fW+HV/DHXCJBgK+5/ScU/4AWJUk3+sw3ownEf
4ycvO5h/88nR9IKvch3B8eSmwye6fRFBwKTLbt5bpSr1MFrpe4gFlI2lp9U/3iWOsubky80hNUc3
9T2mDMfr33+wUPRShSj50lqjOYg38jPHBea+znFPU06giqb4b/2vJZXaNkjhNBR/P5xW5QnyG5r8
qClSaWhj6XZTuHsH+F1F+2vCQwcWfS1hywuAnD2pmaxnuk20WdTuShFUfON03iGUHar2Ldz93m8a
3ZV279rkS1n3igzuy82zJyBvYna2l9lsW2snbjwWGOWxyc04i0ocpLaoFs4kRxb4T42kaeo3vrxF
bnEUiN/q1w8gqPSx5CxFLoRDDfI9ysgzX0kdhkFLDu4WoxTHgMW/r8BKHG6uBiuMJXHckzL5a7qZ
xO9EznH7U96FSFcYB6s+F+sHAzf4oE8f5bJMUm/9i/nZoF1rwnc/byHF4HTV8C2J5rP59j/2Rf9o
O7IWxAABmRYeGut2XNomL+qHODgryuOfYCIfKHKSjMZP+X0wqU1QfiJ9+kFRnN2nyS/pfxF1vGLp
kM1aeM2ovNbQYkIc9nxbQR3sd2os21Kb8wF6c0n4lVw+ktfJ9w4snK0slqOQchMwXBegEdVVilBU
hk1OaR5/3DiqMA4CFTb2cZkGmYRlFxOfvj6dPkDcpzA1mJzTbIvMYOhV6CS8+yc5+HwCONFQgLJj
mjMeYhlgcbu6wONr0Mb5tQiHNw/TQcCuKLFLi8DgP699OsahRtT7dlmQpKQCc5LaINENj9QaCMta
+ANcp1qkT7i5rBwAMdxy73pTMxhJIgAiCuGEgr8pALzp8vWa3r3PHg86S9Fk53tbST4CcFexi1vP
6/h81vLHsFSNbtxe+f2i1f4H5ALq2s0BO7JfqtBne25/jYLrZQTJEjb5IM7jJRiYyY8z1zewLwVj
2wv5gCqpbo93xRzHrj79mYTyY1qAkWNDIzmRv9AwFBQUrUD/lP/Wm1IZGRLSx3PBzIUrOlz4nX/x
VissrQQrtw4KNXstI6bVGQ5jvcTRK3DCSW4YBM1YCDH/ATmg4YQtEPRGWZxWRonrLGPE8nnQ1I18
U5o0Amn+IKtxTHZNMM0wg93z6FFHW03ZIYLiIk5YyUP+0GTDj+BdP3Ldwm2ZUZHeilC6twd4fc/2
GPH5xj6ZX17SpIIxgzLkz8drdxVFW2BUy4kSzGF7vt8pgLkK43r9Bz6sFJVegBiNkIPaAV+xEPp/
3FHzSW9CEZ9POO1ABrV765gXM3E9X7FfAAkUwGlRZexxGqZGkybth1yOPK6Tb4BXATVJHRgmuZy4
ME38TE6+4LferXP9/6hQRPLy5x1Pk8FCULjAfig/cYbwbxkFbOmGI7NW9XLMWqswe4MMWC4+OknN
7xzEX6yzjURbdP9FS+QWncd/5GkyT5tDrA82Zl3uupApaNN9GSQtlBM2QEEMdtyrGpjisr35vKIy
4Ih/Y0ou71KEeCKuw5HVHSs35nfA3Dbq3HraRK5FgSJIMaWemSf2bKiCXnzUw3RUDGkHaGFUBy8/
cJdARq+WC5smXuvnK/c5oPXOtHbWncZboxpc5YrGx/FYAkU3LazDMl7XMi43hMxL5GqhDwzluLDq
H7CVcx9KKuijIwF4t7/rwMy1GrBg6cU0qob1sfwZIeYWM+mzfD/lceUKeQOmzK7+YWzLvu7SGdQf
+RVHgDTNW49/NA+1ARVyJWFMzq5FPag2mmNyoalXw6BIdnqQ6cdwnvpDn+6fQWJHmCEos0r9iQDU
b21wXH2qjy1P97b8MdfbxKw5J8XJVuEKuntqTo11UlTUvuD6Hn/RYQuAh1KHxrK3S8lYgopduPoa
xLHRAxNzwLAkKUeSCRn/6TUMcVLchYARvN9YCzKM+8/Nzoq1fBd9u+h2jvyOgaSIz5s8yurfVKls
l1FwXMkLRUjASlknixW5g9sNIHfFh9XJZnlOM46To6mrmB074uyZhZheGz1U5x284l9u6QA67Hjj
2yGvF9ZOw737ruzDrxQi6QFmp+m3FPA/uWIg7xSXXJwm0gNcO7jIahJT0koCs5iFm67wLneoP/h4
Old0BsODHlq3t9YF8uxfGxdseVpu/lt/KKQj9YzunCFykOCwGnxo5S3V+8sLBDPCr+mLnqL6yoII
Wj+rIZhBNlM0Jhy/X4v17vWFk8Hsa6icDOCxHUzQvixHXIAndDyek1ajJWnLzXtkrx9o/DMAnXcq
0JSmU6oLow/N1w2oK07wdjgIx5HOhQlWJmlDu7gxHrmTr/X6OlTNS7I7qfx2v5NamvEBq6V7/RvU
wnztdO33yeL37U187rYtN5E7WnP4fjX3Ir9qLg8YYK8/ik4xrfMdRERXkPw7LGLF6jPwYK4W5+L2
t/+L3rHi0A7e57unEyu5yYsfUo3DPkBS9LWa1lbZeB1rf/yJz9LAVXBHGsWG0RPuoAxZ8PAaEl4n
hP5oeGK5y6aId4HY6kGhV80S8fXbRx5RRJ8i1iR+i9fdkN9D2riINYdSMv6Tin9aPipkw/pV51jO
5/DNTDiJFXPCC2R/MK2mFgxxjRoVvOV3xxgj5PzyoLmoURHzcvwpr3laKMf+eofisWvpr/X+3l0G
Lh/rN/eSZmBxeozmQnz2WXqQ+Ht6HUSc1Npt0I2cef8LHTsIoWJdqgCK8VXerreVfAdmjSXUGhC5
5v8LtGyuw/LlSz7D+MoLydvmnwh3OGqV29OPAG8SiRt5L1WVG2lMVcL4A7yqf79noPH68eQGIHqD
dFD8byBhyHRG+E1Aw5cJYphBBkPQqLeONuHIVbPPYcRii/NJw0KgfkFMlV/SjofhYhQhbvjYhyyn
UzZQwf1C3PKbQUtTVPCJKmvBEtkwSbdd5IGmWvmklP72y3Q0+MKPlXLN+yd9+jWXipGBrul+AnpE
Ndnkqug8eqDF6dPNWKrX12GNFtH6j2urYv1H7ft5+Mxj8ipdZgEU+BmfW+syZgzAQ50V7siJg67K
N6mlmktqtq/ibK0VQNTSqsyLqr7gzqWOC13JA4AmBp7OI4nu1Shg52s7/SJIFuPpNe2LCp7KU3/3
NJsGdiehLkfDBQVc1jwmqoakorug4hbxGvHLlg7Q450jF/VhKqh/bkepdKNWHIwa8Ga4Ua+rs7LT
R9grUplHcXILIhX28OtcGbq2E1o8CnK/gKAGHQeYjpOkGdbMOD6exbhaI4M8WuUAXIPsBkcR5VUz
OlZngQqvWeYkamqQyRryZFYwUM1mIROPoUZDqYSSESQNJ2gbf7IDtKBiTvKOHJo+1nJbiIvJkje7
NZOep8zOW8tXuqqFWsAuaMWBArBYP/YSbAXNq+tD7bE+qyJGk9xKMkJlKBDFjY2pi8o/OQc7sufP
jcp1nqB1SQW+nLhovSuE0IXTWy/CDl+jftnKJEcpZinnL2OwWPE3rHUT2VGCNNH3y8gJ+9j+upDy
i0TTZud72ehxllaJLWJDfSi+NnAuHyQHgCEZuaduHtxj4GaDIKxvhjpaOsi2laVgg/NdAU1KcDrE
G2gDL9U0saLtpxeanyg0p4/dAA5gvhxx0e8h3rBAU2QAU8ym4lGBZmDxr3jtnBPMjvolmdPJAt9g
SmDMGY3ZAjsk8ISHPrhD5sSCc9fLdvbVZZ5WD7m+gJrHz2OuyiuY9Bs5yMyRM+qypECtLInSeS0O
pQVwaVLmTMvGL3q1inLLlhgwIn8INNvLhz5+DRbqxc6N5X3GE3PC3s8NSfOq474dJ2/1QVGUKSBC
lHuPYr4cN35XaQ/uX7gVwaHonsSmd+MW/4ABb3CyE1RBCtsap7ajrSX1CMSSRs2ptpJkAIE1B1Tx
KXAYbRUDRtj0TlAG1vEpyjeKyc9nS5ajrGXwsVkHLT3V2DpOEaU7BkimkbBGDkxzdlP4ysugv6dd
MtTPpDMs0Vcyqri+Qly7+K1w9f9XK6+WQKnz7rU0xdAlN+j4szNMBofGyHb0UAV0S4xq1NVFXwxp
6QtVwVQoxu9nSOuxYH4wNv74fLp8GaSXVu52HYOImJD0kCnhjLH8zNCFh0iCwIWhxXATQy9FM8Zf
abPxdz/A2DAsrYbBy8/6A9tc9G09RU8W1onNuSIiHfu8VDDmzeQV1mwg4kTlRCKHE2PqjjbMQfSy
bDQCtREa44VAHBp5EAWohr9SBceHwxhny0jzkKEjgMX6SasPelqUhc8VZed/06mMHgMfzjTxic5k
y0vN2Wnoev594CwY62G+OE5tivigWogJtKmvmohtjKc2aKkaLnf+heUpKm1bVrGrYZ69j7nkcEYk
s4fEMQYuWIZYFpfD2uaoZjMLDkSOqkqxaFfrHwzTImkNACdDBc1/MlBa08lHexQdv9t8Z50WNaZz
awxfNW2dMYegT8tl+pNKieQ2jIALUsVqc6WK9QImL9KgRZs7djIdu/e0CtCXEg0oDGHT5tZXmDMl
IOdxZdw/wsSU1v6+6eFWPSL5g0pfA+lkDr1wZrHXJzLU/0eic5KLfDo8nGJUAJkCPVCkxA3jRfYi
XU5YUldu8a9fLsF9BwSrJmUs4dXIDP+agAz480T5M0gNZQRxFSFiTqkS2xsGIQa3ygmAAs46hOTa
dl4s2zvkp1ObVPPENtZzmcxxDU2cexBwRJQI3hopICQ6reJ7Ob3lOj1sOhwpL3g6RidVNNLwEM+f
MW3Ux/kJQiynkFrCNeEcAcqjmlE2a6hW0GPieTUkAguHJgB5Ceib3vmAw+EL7a9i9hvOzNvl6qg3
kDJc8yEnCQxE+OzomYV6/iqImhVuKHl3FUlYevQNJvDPBxRl0V4w8b8KMj+Q7ylCGjZ+d74dFsQ1
janxn22y3LlUIFt5rI9WbiN5qmcYPb8WmFcNVpDy4rqKi/lfITPl3/svzSf2z11yYlfnZwGn/L5x
yRCi6pu2Ah9zIy0lwsx6JABwoOZtuZ3Tv7/+He1BkJvw1tOy9HyVITjW0R+nM8/XLOb5HRC3te8X
aPBtbQ3RGS/TbVz9WlVoOXq/f1jWyw1GrLCmwjMK4LvJpdl3z41MLbTTKg+Bw9llanvyUg17igu0
s2clLV40BTh83VKRDGTQ4Wkev5iWw2QsfszEUoiD2F1Gtnm1KaU5bbPfyJxC/TfISZfwuSibjNcM
aKHQRsj2ma6r3BBp355amRZJpNZPgFwwu3AGVFEdHMpXw/uA0eFFTaluNQd9w3uE4JyZVKVV//R2
vO3ihrz0ddg714awHk2uEjtau3+u8DNruS/H8/t5ZVIFO4zsOKfQNXCGQ2KUkNDaZ4cymagfgr4s
KMUQ+T5VPsJda2Wbe4FWki7zVJY1/60if1bMIURwQem8xo5u8ORrEY13n9787WiIvq+NKiY9WLk9
IOZbzzjnmJgqJpAgyEBK7/TcAIeO26x063exOHrUf+xYXkzIFpkxhrdqaFyzc8OspI/TRmFEX4k9
4chfUHSFttCfH0JSKNw5NuvIdYy2hzyHWH7TgMwzqpZtJrm7bS9muuSxppB6HufUGV5WwlACAlXO
iCEgrtDimDi/ChzZ2yiQY/whH7QIGsHIu0hcsyuWFOQYd8dzRJ+ERET6wIt+rcnKq64YHOJYDK2J
Tv7guQu42DViRVSFrfMs10Kz37+39NLGpMLOOceDWT9OTls1T1GZ6gNufdhRzMXmez10/8r5h4gP
NhaJvpSgM/db7H0/GRHZRF2EE8nUtHoTn6lVS7AxJnStsEfiQVlcn+b9jLfF0j9Ux8oolDjzatTJ
CgSHhb9xxoCvxlbr+bUl/z2txxbZjyV/vsOxN/SibPZgRnBhYf7Vqy/QVm7HfulnaUDyt27rQKsf
MjYxp+XP/nck8d1w4Ae8PfnU2lybSPTJU4Cdn/O9xuBGGqWFKYrksSQmjicJtc7/QJC04viX28NW
El3qbgO+irj3Odw5KiveOOOjBmENSlCu4ReymJitvfZFAywfp0QOiM6CqGtuWHxGqCsg4tu/d1su
26JcXX0vmIKBDmxrDrLpHxbgcxlGkG06uSTng0bKXY7Z1MdfoNBKI/rkQPckNtjdn2Ti6uExL2m6
jiuKo9Ofggpq63T+Y0RBYrtmWza0O0Y+zAQr3IOG19IeSNBojwzeu7RLarK2QKbgAMisO4DeeYo8
47J/R4kLpvk+rCej2I6n2PLsnb5IirwTBzfFtEqwk1P/f3WwLfiv4epq6uxNygdyfaxRZ5u8EpZk
jZtIIBfVrGgxNoSQX2DnDf/luhZX0XHapV+zQ8Fp+3NiJ8SivNGdb3Xf3RdXanz4ZXdCARNCYf1+
ptQ7ZSv4WB4RWbvaS+l4u0Bcn5HCid/rDs5JItfw7ucfc4RpX3ZRINYzfqPfIqRwghZZmFynyZ00
zihEjtmCNNn93uqcfW3VXfGs5x4XofBVuS43G7En7nExWJPTcUlY5huB697GeJX+JUWq6K752raQ
3Fa4cmure2xxI2jc10nISkrOTWctQvsgwhH/vmSO0Tp92G24uL3M9sZ2Q5W0dpBicRFIvUWumn+x
XN+0u5AXCf08qUWIeVyVfBuj9R4rhUc2Q+pHqpC7/arrMj+i5s9xdJByk+Z97nav5ENrzsAJhxdY
40/X8dYbO/SDYDu0pgZCqDt6aAZHdfEbyTV7GbQ5lRkfJifXmCJARh/mUKTX1hEUlG7zS96aJ6pw
HTxvwBfPT8s2YMj4b27BSKtkZE6n1oHN9fQpOrXip35aturN3G6TeLB2F9V+Dblu0+446uNYKOxM
McOX7WimrcCLRhCfQnq2+c1eDsRBdDxJfyJf4m/koQhqwOkTGNf8M253gVqNJanxm3kLsIGicpmC
zssv/S5HXfictTwF1C1BHkslQEnJmVrKPMmoslDRhPA2yq+Ie9od2S8mZJE9DYYtE7BM3ZotiNGF
061tKCL2fxrgexasbPblfPxzHQgik0OmsbmKKMaRynVTFjQT61D+/bFbrJ41swVQOEMdCds7SUKF
4XXS6vjXt47zIBy2X73t+FN+bznCMx934oTCkco7lG6au1zMZT9bQZhlOh8YMZfTGWVQkaBB/9wS
D6bbMJeXbYqJXL28XxNCo2BkaNAXa+6TEQw6WZeYzIRlz1KcHqK30I1iiCe75GMe0xetA+eTB6gj
qIXaaQFl87m+40OPkz79WwXs9Um0Jqu0MPG1D2zd47nVQvfU84cmSIYh3ywnXyHFKlgql2J628oc
3FxXwDQpLmHgN6Bgbx0vMqu8HEoUj4FglyTZpwr0QQR08KL8UjunDuuUdTihOPQOjWVOSVwsvjrC
cVCZ/u94gGJWOMskzco9Y6Dfdee9JuVTtF7D8Oh6EGTktttonD19ENFhcnfUQecC/p8A+PO4Whme
vnHCZBn18qBBkjmGLWr5afiStJn/snHH8AtZ5ncdelGb3M1jEiejmfO/K9bIc6VEg7l/Gi8Myr+T
juEdJz8gTBCOQO72uSTbeQ4orYZEBLKUzWtrdxuLohkiTcBphIl0duMgCZVlFTNmJwrmxlinIKtN
VQ5uOzbmDAdnVLxKRrcWbniePUkeBTbeWDmdngPFEcoLhaGx4i0s/uG0brnsc1VvTJitCbMmzvU2
W3NnfymaB3ViJ9e5d+mP0Jf4a3aZGsB817OuyrNK/dUyPsvoHdYpegaTLw7x/IpNOxwcf2gL7meQ
h0jPuM/89Uo8G6vf0mWcoCl+/rkqFKjj0K7jRAHShOeHZWi73U7FNGnl8Kx5R2IuS3fC64Z7zzOJ
SvIWO9kcB+MLuFHvKRHqppBAgM1hyLQIc8MnZ5G9Bk61BIyLcutz4fdg0nsJUBvIazAkPPbCvSm+
KAJVfkU+iW0AI6bQ1aYHA162HE6E5gi8KJj/OETLpFFbSRKSb9nnP+KugJdrmTZ8ZjEwZjCnNwT3
d4acV9KlmoaL8Gk2zc+nfI3qUCwZ4MHXneC/5glfR/nk5M+Ik1C1FjBGBU0re4PGKrVPA/RTi12e
e1r//TrcZHcKMyQnMoLYgkqunJuuR1Co714R98D8EQcrc+eTWf2bdz4ewlLxrAdT8y3ewcoxzbrC
hbAj5J7UMJ1W8/UIi5uqI3/TR5YZQEDN1lwmWqX9+s2VegldG6AK5w/cNvw+55L5Qq/hfd09355A
GbOuKE0iBHs2Utf7WQofonCLqkCHRjYZe48RlvZnRw0i8Pqat8LsSnCjjUwuG6xXiPD38GcUfAdk
rlyXyN04e+SKNwOfyzwZS6oSnRqcHbuIbm5urqfJZp1lYPR+X1Z5yF19g98y3evEadIPxK471nEE
tqaXum+CdtqsQTD4g6zo6hspvpKwsaiYtE9tHnuqfkpKvNpHVU+My4ZDFo9pDuH3ZGXr7emQq+Ec
RmBwcLhbLZgNknIaduFmANKzMwBEvRsRUkbJCwNIS1I0QH5wu088iEphzhYgkTTdqeBreJ6HUV8X
S4DGrv1tXT9oZ8naae+jAn5dQ8bwytO7AD5W6YqclbC7VRgA+Cimi77fYyRfKmK11oVJmkNBfL3B
FWodNWhgD3dl6S85G49mtYEqMDG0FQQRdhBF8NBpBLlDE+hOMAArKM0ac0dBgd1vgI8c18pCN5Rg
nybsLrc4ZXtMi0pj06CcRHd9DBAOAyEZZhKVIj/s7WT+9aEn26fjh0xjzNbWrXS/Euqlx8Lz249D
2PMr4NbHfJ/LY36QduSIHeIs8ro4mgOA20lc3vq4Y6OVxflmuzUXBLJf1o2UQWPJ9GWvJ9V3pedE
UtfeVWeLjJvw6TRxJJ9sbQ5RIhHokeCT0+qh89dG2DMnlJgJPjnratDnQ7wZKa0lzfib9R0fCBfr
E8ZOxjWEtoIXdHMNOWTcuOtjvhYSENIdK4ZF/owx3vCKQmlbM0MT9htc5VLO5tSeroNcNtMNZaZA
DRN/ha/KK9di93bOVcSC1TUT3xwFs0mu/QDdWynVrUmDOjKTWmtKZu3KAaZorrQ2xzXWGw7ChUmJ
QUF8M51FJP6SDp2Acqs4GdHZ4pUczHCBpNanzFPYicmPnfsYdQLPoUZhtcMNc2/5BoSY55coqnna
1ryrkhNYCUTiAtrEZ7dljd0+Ft74UUEpFn1/pLjsyIdthZ2OYTycg/zn0ntZagRrfq41ZRhpv9zE
DwqlIgtgy1ZWrE2t2WhKt8q7CEo+w7JRLNBhSEuYEHfBJUJLA9PlRfGIdE90JUWSDRGYMCS6MhuG
+Cz9vvg+5un/K3JaRSBWRcxzwkRZn+dUf1FXeHhHz4gVy0iywavbI64LuNPu/dPA40wAb6q7sAU2
jd6mY2rkPr7B2heZIBC5uO5bJdz7cd2slDkC5JCBDv9EB+QqmZ05RKreEcmLqzrusBxzZPjq84+7
uVoZ2GD6oDjQsl+R1wpwkWAWdoAKj+FueFVIyilRMR7QO5jSSLvq3J7ZiIANOf1zEByN6/9+4xxV
7cgJiImjgFSsC+Pi1groDgcUrnZdIng1QWQLK/35AHT8hG75k2n9XIyyETSqi3JBMJJ5d+v5hJco
RXt9kus2mX44Nis5iQMd0tH0WFxgI5Ly64evO3HDJydWxROGTPH3zJ5HKfcNJsfzLCz0GotQLhyy
NRfeRu/o9hDxtW+SSTTais6JlLOAQeQp67VcadtqjCtH/NJ6SILZ/gd43uzDGmpmsF/BVnEuYkci
7sOpjV7vfLZyyN539ACHUrEyQ/xh/8VsJNbDyMP+VxDlg8Nq9yfMaLnKCXF4WpQ3K62Px7BQDEHQ
EA0aJ7NSwO2zYgLHz327bG3Baqk9RGuwTT6wdPYU3goJCT/G64vH+cMFnsIFYaW2KENUxcOop6gV
OKwi3zBWlxV4AjV5X1/02ZLu5w9aPmm9fPLV6F1PbZffbf3y9La/1yNeH2BI5NKEiLej/Ghsa4KJ
CpZ+ycwSMRUPNSJjWYuR4mFnY+0F/cp0pkjay8j/l3+bQr2X6F+p+AezmyIbHY+9urdxwyWeJQxQ
pisxuaOaFQJzakXi4O/r+tnRy4H3s6Hb+cRVYtsa7HU7TKQdOHmZDpgKtq3h/2a/RModrcvAkIlg
TiPXXriCP6P5259FkIcvMLs7ts7oMJl9WCJ/fmKKBV+d9PEDevCutRuc477guEXZMmF8jfQtqNJX
saUxsvZUVwUFJP3DqfDEHgYTss347UjKrBwlolE+KGmRyyRLLOIrfl9nUsitHQw5tiLNYbjIRqOD
0h0czq3J71Pf14wcHVm8EBCRcsfrrlzJQDOTn7sicrIUuicrhfH0D10He4w9xCGUMJq5Z4gNbWcn
Zo4/TwL4VLYekjkRDLkXs4mEVe9+C7MvxNOXa6nADEHYN5XcwG/3XOY4M9INyBGyGsn76oCy7vOM
UQncBO8ZeY0ntFeTgUQgGwnve8EmnVPqntKF94oPCo2v0+ys5si6QqERYtWyEDkw2GpG48xQU7QL
4N692/JLpiV/j+oc7kq4w6OWI6EaZlDZJjTXmw64UB4fpMiq+6K6/B6NMFRH89fgNLaP/nuWf8kX
fXU9oW+D4k1psFzPsoHnKY180IZKTGDBn6v3mhe/e0RplJfpFo+QNz8yiAyW4ZcSk7KCTfwcY/MZ
KQwp+qTypWicinjZElKbBIhoSUj46RaAIE0likQtENauHoazwWFsLFZmoovLYb5waa2QmmIRjkHN
XuxvuK30Dnbb9hhK6ZpCWbyGNcdB4XTMiiBDG/eHo3piXkeRtV2/ZGe28BPGDrH2EwDFMSVECSZ8
M5+kGdzMsMgsnjcKC4EIVF4Kyb4cn9AmO0xE6lfVBGGgkl13eJHOBs5zz2aHdc/4ErRmaBm0ymnV
2uhHAPf8GWet9OH+znfhmvJb4Gh6uz6yKSRDi99zqUCkyHT2MOY+HeXKQngsF0tf/wvLm/WKp+1f
nYlL0Rolhhy/X+igoY6/c3aZJROIVxV/FV4DeVirqGejr4Q/y/Qa6cFMECx4EVoimOtoKQx78QHT
zwzhYVun7WLdGiqUu+g8dWuf4kpvBi8o6y05hmR9ruLmWJSJda3aZB8IPlp2Yed4bQGNJw2aXgqQ
U7QN9mR/BKRJn4+zR7Lf9XQiw15peS7OYtlUvU0/Xb9RokxB1UZe18/e+948yVAUqxJCf2JVHrT4
w06ohgvth6ulMUIi0DwKQ+BB76YwkHlNaYdg3pND/XIeIZ5SkqtmsrtVj9ZvxgU5o1Qn6g4jMH/G
sDjMbixaq0/NjDCmbgwqTamKI/Nl4BVWV8PxmaywZ5Zyk/Hd4sonvWgWG+xjP83xR+HdrcMPo5QQ
KuSimiM37/wuEbYCkdhH5JovsxNkKBvWBuSjw6bbsUx6aWkazRmmEP+p5dOPrZXqr0BiisaGoTSW
DDdKlm8cLQSAxfuBA0XE96gaYIZJOPhOFeVfUKkfVfk27rEk89NRRAhw6DncAMn1DBwulOAF59EC
pmT83kitzZYRbooylK6uUtCi2rO6WwO7FWhTZ5fb5XBQ+wqorGyRIwr4a7Kbm8f5mU7E4bfQNgjV
t9dySFePAHXmAskTTKgD8Px1wovaKXnVWwxMJEsm/tfpooVc09AwvSX/cgUnJNze3jBTwhqCLLMt
k7BfciO6JgkcUqaaSL1ey0onxYVoSlKhjs9dQ335XSuwRN+GEcUyyq5n10O8n/k9C8PCUFFCY/E4
xGYs8e2zSMUhB3XLFQKbWExj6nWyunzeKn+quMgoq/uXGBPNkDVunZxrjKWcHadOGOt/J6XE/85b
+DG30YfEhKRJ3hj26wNC+dU6jt/85H5u2xcwYMpvHjPqvWwrHTvz96/rQ9H3Fy+UCNvqyzjXVn2E
dNrMIF2qMiMJ+43xnP2XSvfiPxJuYFvuhqGPG6AtIYev9yO8dz1341P6jU3gOFMRHphYF6gDQETP
82/52c1H2CxmhredEw1/IMK6anB+RpIEfAhPthOWBT5sxhNXytZ3n69gqqT/HoJV7CQ4ko0Gpjsl
m5dowXnIdYqZcDw/U2xtgp+OdTR192LN0BSbp7OZOcY2qE4Y/CvOFYvktcGP89F+dCwfag4/roL6
iavtnYSO78PxtncBZ228DxxRci5kpX7VaAIc10M8yiJGlz8kreoFY7xnVrRECdRvwjcKyMGeySng
cY46P9+QCKhmRGprE0IyrrjRYRCN8JZuAbHMWsPgPanIjwZ4T8pPPWugeKrHJpYhejVkzWKowG61
bhes8KtHgeI2a0tIjYsDf6vqOEstasP2MxAp+Pkl0GV8CrpxcybIF35cmx4TNKaVPKqOzNvhU/iy
kPlIRQ+JCO1mOXlV2ZVYOkhlavsd+QepkXJAuTbsIdy3EGBjTmBXwP2fDYP8+MhovNOb4YGhW8N4
f9t8Bjsp9+8mp6x++fOvWBdN6yhZpl/r/jFYrGrw5yWrWLyvUHHZqpMhzZWibQ/KdnV3DGimGeph
0uDrxoxa+fCzQg2oszV5o2Pf8fSIkS2piLIck2m1p+SwzG3G6P4+NmREqc+GD6jLScAbCATQ2RoN
bjtlSeznYIzfT+UnYppuN+OvGOYICeRdvYAK1cKQCNCKohukAd4o8S7aRGZ3k10CV/rnWG2AUDMU
Ss6rCizTYfVQ18cxrIv5AmCMvbZz8uTD/JQB0YfVBxiy4IN+ddqOxBWqeNLPqyWgvT1y9FrJnOpZ
80Juch8awVEu6aF7Ntca0WtDJt6ZTYH6P0WPTTfLYogCVi+BG2gQmTeiJUX8laTSg5Ceo8SNgytQ
0ikgjOziqBEcf55zdZ/ILst+8c3PMJgDs2CADLQvpbeULPcDNRGFmmF8yqw1qCVgEPd79tYULDie
Rklf/WACteyVABbIeid2YW6Ru0rZ3jORRD2eYLGMwT7NsT9tcsZCiIUmC9G+PnVs9gkLlOdXXLkx
4wxXk9S1T0u4MFNiJul8wldJUmQJbEiwAnvYE/zX5nT/UcXF6plnYCQttPpGedKSkUzPAx5EoCFu
L0r9SrVhpngMuCoR2odEIqvW2b5tXcpFO1qZ3T0MALAyEg9dfGkEqWVeqZkxi+F9XNYySTWRZebb
GVfQNTrSkyd/3KA+ZquP5X0tOVdZVkElZ3YnDbYvkv1rxrC1XZrQc/Cm25xOmY4yaTMFoasRvhGc
yliTHVGDyYRiYdY5s/fA97YK3GBF5aSIljCJ8S9IPW4t2zzsY7agi+0ZHkaeFhVDuRBgZbzGw3OG
IOiCCj3u47B8RCcpn4qYk3ZwOr2pLhRTQ7ClQy5ZSu14HxfIKZaSjHaj+fLlVJ6+vy86tsDERmv0
jcKXGhh5389N0Oium+fOGq86FIdB57ZwQoZLSZ8FEvZ5OKso7OdtLFD7b+UmQbGCiaibdujnOZJJ
Nd22B+w/uxcvYztEnsRWGjGCgxhOGjsCPtZKtjIboVnpgNz+apt4yRLCVT9ucUMPPdnRhi0FYhS6
gBwoC84QXhGmITr6p5dQtmRqDcOEiXITRk6WTIEo05TL2e7aWYyVWSd9HPt5z1PhLLB3q+9pIsr+
MHkmrfBgDqs2iUdZJDwmmqqNekjxXjw3gdqbhfJWqZFL7HCDvsT1uzwSvcDg62KYLhvFPjmLCrHo
E5Ty2PqFQU8POs4PjxmWIVN01pslaNgw5Q7HMnE2zwnD9gJFbsJTjvrEysLuM4BFAceY39/k59Tw
HgREKEqsbFCaXmQvMQBScPhH0hY66GtB2GsnGU19sUt1VX2Vxy7mWvyswDBlT6IS6465jVcc5Fbj
Avs5e1PTXn4zMgm3WQKPgsshhuALHAHm/NK/VR3HSbqaT+ST+rGGQI3VOpUQFUjYohXNfPtWF/Td
WvoHYaFOpPaYGY15WfoTU1L7neRvEaYTktx2wYa0QJ0OM56ym6BoiuH0Aoq6hrUHCbVjdmZurKsJ
89PLOHarBgudeKG2IjsJQUef2tpJjISy+qtTBeGt+lSMqDPIztTDwBg1K5TcOpUZjSaPnRxs9rj7
83lB48fLfj90RxZhZiTjcS9Tk8NUil1Us1iU1iFyjBykGywcg17hXB/V2cMHiFhfFaZ3hDyDoKrd
MubSZSRSPNM6rZqcrxFrsE9NsMFsDuYW/sg6Hl9leTE7uGnmsq0uYBTH01majjc9NM2O3snWADT4
iJSHDTVSsA+/pImAKzGoK4TuF+nvxUaal9sgg8s53EVqBuVo/jee+ZIiF40Lpf3PJgeA2vUe1L42
K/8TtAjf8T745cWZ8+gr0q6qt8rPipl7SAKuRc4kvg6tks3yRJXoxAqhi00FtiiwHMYWfwHJctoc
lL/pUZ+D2FcwkIAs22QNxeYlzx/WnFQtUJAn0uSFDx0on9WOY6AAljtaR8wxZ/haEyDGKuYJ7fWs
dz1H8gNQg9QyrSoN1mh/PpDw9IsU3eJp/o2s2R7kL7QieuJGMEn6MPt7ge3S+yu1VOxysynrx9qW
rEbVVrl6/pghhVJqm8iT74coVYU1Mg3Arn/8cJam1qxOmcrmPkiY00SqMmeIHYb02bMW5YYqvlhG
xCI7Ds2iIi7M4LENFU3KRDtdlPXTdVSjNqBbUPvGRQopS6x3JpQZkhxd/3oHhkq5xVsivOUKpGEK
w+bsVL07PKQr560K1/GXHnrXY+SRH901L70HZsLn7fZw+KlvcC7R5AXA1TcV5416PwfcbgmftRAy
3KnvrsILsOX9to7VolQupQ9qv5e/gYRRklVkxxwansGMPIt35Fj9xBZ2a5KtVk7ZWnLCMmi0CpwU
tiB0VRl6PUSuAmJkYp8l//qp+cIcHONjJ5jcttnugbooSi4H17AXJ9C5BPhH+1ihvEzuN4x4UC5Y
D4dCcclyAO6y0SCcbREOGx+Wj6l4xwuksqb4Kuk1ZP3QUQVDu2s+YqquXTjuS9ugeLTTnIbZbJox
jAx6+7IcP8WaWjW6CLVoNI2bWg8iO8T2VCoU0nUUkclfkefwNotl5V6jyBiNeWqJIncO+rZxfGYt
zuJM5eGM3cX7cI7ZykRF9Skig527jztJn7PzHZ9F2RPPltDdTYdN3Qd8juvO5lTVoA2S68u2KXI5
GCPhZ1g1cx1j+HMW7pPjWX+rjwDnWm/kIiG7uu4bNECtB8hm7G9oNsVpJPdqrNO8Bkm6CJsWc6O+
evaBqouChaOjA9ti05zpZy7vVpnlzt30oDt+lhaNfp/Z3qbi3Oyelre2fv0fPQr6Unn23Pofansg
5XsD+sKe8CiMNGU0t5tD9jg/Fn8jwoTsc6Zqe00B2QUacj4AIi/fsD/aLvc8TiCfKHJ1M2uzCrzS
Zny60mdAe6y995elQWESbgag1e0an3b4IMF0N118KzUzmto5hbLQHPLLN3ipwy/mnUOHgW4yd/X7
4vktviS6ifO/jVLBWI9KJp1ONkM+jAEobx3R5ODdg1fvR5ZvYDFjS86MQ9p/AuZpRM6dwAdF9TIR
bl1Yt/TEup75oxdmZs9uWoJtHjoc8S4JiMuANYTKQAP1z/PvdTrEfHv2CGcEEKL3Pqveq5I3QFVv
wRbx3pX1DaWOYxw/6xenEOfD8PFEB06vXClQ7lUh8YwXJFGqtMdaS+NaJ7gEQEXIOc0N4Up4bsgn
VjnUVxpqjVPTeFwVtaIUHGlib/1Caa1vujoE2eRU/Q7wB5GwFPUzH5jQtVYK+u6makpA3H59GU2A
XwK/Ft33Fg1cpTazYXqt1cuVtu2paL45UwbzI3gppJ2T6GHzoIIdiDstOBs92QKskS1gatQhkOU1
FiCZWbHFYyxMQo0Q2RIbwXHxMexIVvz3WPd6AQLBa1aMGs5hL4iLWCwBVEcwEUII4S1vNLybVdk1
ERlXFI632KtTwGVitb0DBol3ay1I6GVs6FpRwFGXn9YlQ1apzJZkB+CiS6oSTAsCC8UDoFNH2GrP
6rA2IYLBWvdkAxEkweDcb3rDEXfK8uejGwu+8QRX//5ypboOReDTnv0aKNBkgI5ahwMATb5HzK+i
A32BWiS9TCrvUulUoyH1Etfm+4YdbCH9m2T3zbFXFi/bbNT31dElx08jSra/OBjHvwQBNsDlde4z
ny0Zdr0YygokRqFSiYU5B3zWp06WaVH/qRTVQWMzRG2M9FXwgi/1SOUBvn4hH5LUQzTFUSmI1y08
fU+DjRqT2GtM4zA3YpUUTK8u5MNLlIZfumSyted67dmNZH5xx6rulBIKXY+bAeF2ke8tdVE2MC4Y
JvwX9/OumSek7zpcbIUAV2n0Ewpx0vky3E/6+EyyG9A8f+iRu7y+8vimhNMgSISrt1tZCpwpkt9u
03VwG7BZhIbCwJmN66ni7e+wFRH3CnzZuxutQHR4GQNAXyeLemwOyE0q/c0Ikxk+LRVoxZbwyKxq
vxNzM963X/WPuD14YdWavtCKNWyK3vb3DgvXlMX5rzzfvkLLby94FcgyQMB9pT/kgCFv4CY3+cFv
Szdtk0fKr6g1FSAfZdx6SaATTaWiRulBFZWJrUo+z0Tbm/C0haM2PF0xxibza2IWlgUPhr0wBYYO
s41dQUKXweMb4W8/fu78QoYjdURz1ATfT3LxTgHu34A3aChlx/tTwZ3wBzBtKLeDzM3+Q/c59WJD
nXAAmRlJoIeX6BpbOwq9S8J+bXsXQsU5VHObZpb9ZtH1UIzVp8JKut6nq/260I3Ge6QCfKbKuPMs
yy5z3vSAxHuxaneAqBojHUHmT2w254RiVE7vB/nIUW2t4dbRiTCmq+P/gXMi/w6GeRODsyT+hnk2
VYadBTQGEVjIC00ZO4UjnSFj4Akm0nH5fx3oBU2rTMy3E1TdMgxOtaWxFCvJrkHz/OzCEvBVo0i5
GZ2hIUYaCyjPiK6ksx7oSDqdCjXUqUrPZngVfSF38Gvv1Zt8dHKk1szL65EHQY18iia8tIxyWwr/
p+KpVv/ZqMQKOQwSx3W/JcSt9oPsN1RSssQBoSYkX6H54flgDHg8CvZgHdodUHxpGGpr1woTA7vV
0qmOAMLIR9neYHn5fYuq9+zX3/QkUWc/j1KgnvrsT83PT8Aciwp1EkBZa3zRlX2ojCgTkAFy2GUg
xu0zJJWw69TVoifrpS8o1qzAXtP0Y9uE7rbMi26zALeigBtpk9murVT0giUa4N8AC7NRuAztivKO
kSyezNqg9OCBOnjjXubkQGHX2GEonL9aecg43QUo7P+cZ/kBFdjbPfUC8iHKEXC0rnRbBMIH462U
H31EEx0z5y7yNgflOsPJ0SpYyAplWXDAHPN7h17muoIhbD7Z/9Ww6/qkXjcF9UX6d2xSzpq5kZOh
1GSYWasdtPTjgsU3B4Z4ARRwfr6bvzt73W9aa4A4bV8Q4jkMEdcS+3KocEZZdt4ZBqcG4GPvJVNs
8tm7Ju41Dx0CdSNvKMQKGW692hsjSNoQTJia+Cdi0f6NYrz5xzun2XuzTUBBqUUybiT2hVolCt/N
gL/mbYoxN8w73EAXKYM6JmATSpYBYcMTtT8lPmnkZLNMsv9iam/SWtHedMbEP9Koz8bX1GPgSFuX
XOs/4OdOj08uuqxw3SpUXj+gmo2wSf0owz3E9lRbmSibtsajjXNpvFDqTZR/NRD4fBEl37a2nsAi
4G8NUF7nPuDG/7dm/TWJoMChLFBgTj4ZBO77/WsxXoJTGld/pNxVhcWwJeQAod8TMh+QyqZ1LCw2
dTEiRTFlbtCPIkNB1I16rPeyQXSZ/gCp9XrJBSatqY4WaWwyyLA1ruTMGM4TDOt65uv8JNR1gOvq
QB9UYXjQgKix/TOaa4q/c/G27y94qwvfjLZPAzPMOm4l0NpqKfHPpJHIWgJZ10ZIYsbCjGKyl6nT
C6FxS98jAQPiJsTZ+xQVPz7foPdoMHZyOKvcHe385dpUqJOAxulSKS5Ha7EIXiIeXFjlhiqZS1GG
ZlPhIYFQA9cBoyXWyyiQcH9xm61mklUMPxqiQMh0vzWj/qvm5MCFtzGcuOLGmIvxNpyF+hAGUneh
7j8H1r6badOHCIdA0LoUeHQa5p1nmkdcCEap7Yo0GMSKowFGCXx0H2JLi+QOhXyhpxX2UifVpjMF
32v8DwPcOznypHay2vMXrlNF/zMZtKzrkb9u1KWS5OesOd5p26YXsopatcwXwZOKs8XmUD336hbN
tvVa5PkjG7oTNAxBGbyWOXNRvAYw5D9W40ewIDfi7EjcU29diceLsmSQw4goEQPSvwL8rL2cUdEi
GbhtrS4pXDSg6pjRgbduhtDivcCOC+aYuh52nKBbzwoNXnHifste5pbGdQ6CCzuI/P0gxPyYz+tC
BvkOKZ1OSSdBB6r7kR91cv3wyDvZzHKqrmjCubMLLra3cSZxdFg4O4d7vSOfEeNeLbhcw5eSGnTN
DvHaSU683fZLywpOGa0t/a3t3EgBbf+9ogHDJwxBShOvKCSzE2nbWsNQtOMx7aYF5TnW3fbG38Lf
Sr2Rnlu4B+Y1muXmT3zBtMIZkxUpuBqYfMo0bwjKc91+lUlD7v+FWM4WWExYr4l03xFI0O2KgKxK
gv7yoFOYdk4rMsawNWXh1pPvQPFAXwUygQPYxDRl9pgegvblEAFmAa2G/CE2Oi781WK4As+aqprB
a3kgio5FNqUZMjzPJPJHnzISxP3hq4E/VA2SGAAiDjRJJoDY8LRS7BOXyGKPzxiBEv7sWScnVkZ5
9TPYBf7rW7Odem+6RDD/tY510Me9gUdH20X3HKytGb8LYMOz81ThzJemNeRp1frHX9w8IkkkTmVv
2Z544iVxmjz+sLBMTLc66pqe27KZIcYaeAH7csPD19ETOn/s0w1CMX0hbvfCHjuQemYEe53MSH59
swmhYC4TlCzW+dyIY8w9hY4jichqRBk+sGVL0aL+AFtUUvax6WHxV3yx7oaVXhZ5A+VtkxBJdhtz
r3/eGg6CfRGyhLA9CiLTE/6ovrufZ1vdK0oasFS+GHEJ2HthfoIFLGKaQVtBcqVrLvC3+qZc0KSg
RU5LJAcGdvjdhDBZgft+ATEUYAH5kuEkfpp1NWO1/pPUXS/NTf5jV/gmc1qit5GY6/gKe3jv/5Am
FrR1VRJUhtMcO9s+xNgu13si3LeuVeJfLY8vn6N4e6Me4V22YyumDyKeMq9ML03lb6DTRi3E64Ig
JysSG5dRAZxIBUorEbzkXdZIwXgdcKLiCLwiXzqVUi5EqNe1HbaYVZznPtVx2E+QLKb1XN2WffbK
caTprbiQV4znYQYHei82yZ6W0Kd0fN1DsduAILNL5znA4cyNnyG8joKD6DIJCu8jdP/9zmA6mOIJ
NuAead1t+sRCweh2J+HNx9AHhGc3Wb5NHXWoTi2rYtTOTk4x6oqTYMXaFv4uREGmUuBvoPRbemxU
NNa6l67M0aDai0BbXeFEFDio+mpBsF0c5Xo9n6RuD4lXMgpYvjnVhGTXfDbsGrTppsFXl7rGdFCv
Bl7SM+pflLYW1XlVpF0uqKqtN4clZRs3funLvDUzORPduHkYlXTLEhpZc+C00+9iQs7NQv6Pdate
7G7Nu4fU2aVwNdaMFevTQMu2UJk/Cjugvr06Vn+7U0y6MFOz4lRRAneqU7BFlJqZvLw2DQWZLosh
MaAlEBWeu9t5J/GXmOzMExxTlpN9o0mEvAnLVArgRKWln074O1vGLtSEN1qIsUQAI5CwgE+JaFnA
26xBOBIrwPn/r9IKH/xAfS67bHZDQ0R4DeUlBBwn8y4+uT6eW7Lu4ypx1HoO8fgFeBb15hVKKta+
igGWkABLJ4piNX9xl69njE7BiuqBMoaZnnkXdtq0T8LcOotS2ZDZMvtBipNR3pEmbOehEtS7QtXm
W7GvGljsijVoyxTtHE/83FhAp42xXeLo3iRZvTRJjpJne0Eqvt4H1o3ZVOPL0IMj6ReGFWICI2X7
QCm5Gx/N7XPO/eQF/PndJcEHCfsasYFhVUXVFue3Uq6fbU3/MT9ZiiEs+A1XoNP0SNXmPzTndmGb
FASrktK15946PHOV672AyQjuWb3hVlLZKDLEyaepUQMGz0VJyAYVQXUzp3nPoZsXSqp/f63o4xDP
z2wPFCdoMstHCDRWBXMNSf1dcbMt+GiG7y5InjZ1WLlZPvr8YiRjPSJYxIs/cZoSQv3ZQ/VBFvm8
LVqqAlDiPDRQ+1A5t6RqYfXteuWr4D8XXRoihRKTVq8DZE4jEKMuLsJIRSuHR9fdqcfCrgQtx+5I
BjJm4rDlPNF8lCemnCXKYoHh89QTq0ub+jNNXwzri8t7xveN2FOnL5of9qMTVy8uRBVpTNfsS509
DSa4B0/NV1De7HezYchlgKPzP7GhWIxi3+QV9QEAvJW0TzdkOfqQoA5X/bjmCtpmQs5pJeABxKSZ
C79Wp1WlRYTJMCKWI83+rRNXyGbaOlH8FHgZmguUZioQgsiXrDnK5dNN+XiZ36dTfppqMPZZGnkd
kRC+y75bELEZNgdw/LoOglaCxM2FYRXY1zsFA9ilT0RUc8qOsK94PMHZeEVHEsWgJnRjTO8AoR0f
bPrZetbM5soAC90nlmrj//vGcJ1QySzJLx9O8kjqpBMN6G5syzvqpTYCm5T9fhg+9nMICReTTu17
f2miYbT+ZL1DsuT7bdjhwdOrnAHbhZG0WE0iRWeYJYpHNk5JhHYCI+Ph+065Hz3em8p+XZkZwNeJ
351LvN2oH90zzs5RQkzJjpEcQM6VqwOLOaHNo0ZztBFKd39T4u2sb2SgYL7rL5sjDZg+H1mYONSL
7AD5m0ZFOkWzL+GgGRyFmCWDmYwwva5esk6XxJIDU2wXlYtGtxEJ5qg5bMydPnnC3tpjnlJiizgF
xLIkYew4Aja+fqsDhvXFMM5YcHnyq6zE2IsJo8Tlf4mTimcRTq5F0EzT7WmuvyD6HV4DaNliFeW0
PdBDXTeNKOFimY9Tq69wVointuODyx8jauk8/+18kV0Sb9TBlhWzp0YnmyJDbzCHx0h/A8ppYDvN
e2AB5dfBKetwGj+mNXWAlyXcdCEdcQnXju83G/vRAMKCG14P9HA9I/lUadYBB1uSqmWKu2E4Zsnx
AT58BiZYXQw0DSkxNVHyh6B/2Ri0fMbJ9qMcav+qwtyQKLnkUhuWj0h4Q2wkFIVzDE1yR2oN0bDZ
J6MVmP7m0pyBUx0VAwz3RhDxHGg2IwvDiw+ln1PS9/DbPgcDZfINyTHLEMbSLNLy/ZjoDSKdy5UJ
itotf85A1F0BPaiKV9Ni+yOAQJF5/XqeWM3XvawKQp3OW84ayxiAk/W7NdZsWbSb4Ea+sdEEyXah
CsQ8m2Vxd3BBbjBp9JxAR0v9pddwYGD7lNPHb4+c/LG0aCApZRYzYoyqNzhSmvCjSnDsxukQSRAg
jIBu+WTcO4t4OcCezel2kD3rFVOYfGOiw5onejXrYvEpa/7FgWn5mmNX4YcOUVM9eXSuANxrMBR3
Rnzpkg0ctx3hJ0BBznaR3jvm3EkbZTHgn5UAw36H3K70jelHAaPiEyT0vCeR31wvzSIciunNTi/i
O4bK4kvndlSQsdKNd6PfdgQmCfHNKa6yZ/vNDOUwAA4YwPXPQcvcnTkEgZc3HxPzuPi8lOdeMsWz
bS6MM9mSCfkKQxVVJ2uWPoU7RQzvPydhxdfTLzCv308jlwN4KrRedKExbqC4Q652beZsZ9hFAziY
rz0eMBqyQggjo5sxvq0mx2p5gn9q0GOcD2bHnWb3/huAILRChMV0caUoScFaCbW0c3RvHnqfLz7M
PFaolCcD8aOV/dvmUniX5d92hPEDCjyhBBmBDCuWrdZH+r03TXUySUy5VBkPh7DQOoO7yXNPedGj
ORs6H6rD6dVCk98tMPdUEJPM1oW71SjnrJIql4rivlPogqK+0xb85HdoY/zoA3GMU/VJVtifUwDT
+LTBEoFqBUs17Gt6Rx3qJi6pqx/e9scxj2EGr9KBCxE8HIK/OT1BTkAkaG64ttsdNP603UFvu/bT
8C8drmI61hyGLIIsK+S/2QJ0XpZBu2nCsP3fnc6zv6+Y0Dzz90qsiDQlZiIEtiNSqu4C6gMXS/4O
WSQz7Wzmt9tJaFatBpQjQTOyqCvj/h6fDiDBk/Jz+tw3q+09dx/Typ+Jo2JwgkUyHZajWClZky3m
MfHNyUnllOVStnI8wtUFOA63uaDnTk5F96+UbyKOm89hMiTqbilzapETK0tJf3iHhtOYRSlqWQb4
Bs8hDdixAAZ7/3jr5m+GfGooF84/rhgYzw7FZFruWePsteJ1GPfS+ON1vkxi5HsJH2KQ2tRhMh1x
T+vGlst/PP0my2b0gPvPKKqs/bORMgVv0/E6JTpF6zuaVGokWEWV/PaWSZSwWeZM2FCsywwyF5sl
uJYyOYpObIB6wKcQARLteh5mheHm42M8yG+Gn/DNrU3v1VjELh6USi284La4HYAfje36c1sHOfcV
glD7FzocAixHPvh34udChoWdG7aiqFFFUnjVllLIyjEDWyxTcSE2YjgmYh1TbxHxU9buVvqEtJuz
N9F2OfYvdvKR3mpSpGq9w0g5Ql9lvT4NQSIu97a6HBpqwym3RFD1QfKNop5SDqLCTkv3AKQbY7RV
hfEXHtGFOhaNF7jR2Yv4cSbAIO2QfpouH6ri4PTDooF8MLZM71YK5GQd5uwjY7B4Ui1z3poqFi2Y
RJAKtyTSNHxnBhqtueWVKfHyjClUTOW8FQdb1bmGhPcvyGmNKy8OMnakR9yWZIQ97NHEHOCaWb4w
av0K9M8y2N7OjSQ/CAinXNg6C6bPqlzO/I9SH3IAlu2YKnYifMkDIaLHHcVBBusn9tYBKvKtx+4M
wIIEtASYAIUBpFWYkHJY08Y+RFe+zYWF/UbDd5MakjiqFnPP03/lTQ3JY5AdpkZr3zqH64t0/1Or
BoAdKthuAIqh3oshSzGLcbZ0bHEbX2sqtpwWN5A4XsN9NR1DRoBx2c1rXcJGM2oYfsF4mGICphOK
CdUubz1FcI41z88USmnEHMw+ZAA0S9LmHZF/hVB82Kpgz9LDTB0qQKowbkSSdDmLCr+vjmaS/ngR
ML4vsQIO/XjlVtwUzOSvxpclQtg4/2oOFEkftSFp19VbS8c9Isz667lqu3YkgvJN9TmjDCkxRDb3
+05zB0vQD7zHxooRrioPtgYIr/2STV1+t4Vt62fDJXxZTzSwSn0ULGuHoiJMsC2riyyLXXYucFqb
lA3UtIWYg0eMhdRRyDA7RWL48W4sgOwnku8hi0OQnaZKZNqam9f3OnzVkfiYEYMGJvr8mOw/azCe
2/vrvg97yoXY5QUekRkCsgZrZjvzi84uqS8gARscG11d7q7Ndhmwyd3CdGsKjjcUFFyeL0J6lJ9j
Rvae3xZr6rgQKD1E3GeHCnqRVR3cBgl3hYty2W/49dZoLd/xcmAyJcmkQNB/BetgsScTiUY4ROWk
l3q77VfLXJpwTVgF3u91FxFuPvh9JmZUldSl2oBK4+X9wy1wTI+JuaXVnPpuuEGmt8ozl9UDuajx
fMzfGvkaDDrGts/d4Vs6s7D1zEYM5NhwqLfzEZK0YBIJizff0efVTp/GKNaRlLnhwqeDCUZj0oz7
QiPhTwrW3h5ZlyNjqYMaJE0fhK8BQF//CFNULW4DmUU/7PRBfl/o0P+cmnCrRh3/Ps8d4MCI54GR
GcMSR/MI0Dy8oRCHKWVy+9B1Zx6RiyW13/To8Fi2A8S29safiT/Oyo95INw3/FqCTx8Gu7hKd75k
vjK7DfST/ITIwieaqWIX0rB0kpPulR2JvVLUax+wPCFduLZ1TYLd0itPbheSmBJFORBnX7rdgFGL
tnRiabC0lQQUZfq5q/vzqDaYzH+QVS/3j7tHeG/6qCa9IYNXcFA8mrcnXK0VMlh9j7ryQjvsDhlK
+Tk/AD/MhS/9IqolhlTPhTsC6u/z6AyMHoRF0UgUNMO9OhHyYl3muC/x1TurEd7GxSOw27Z9oqX4
kX9EnKwkQDXGfso4QYf4v3B2VN0BK141BW7XvUl1hKPeggyyaz0nNcowA6aRUeO4laXiy+iIxFGK
bddq8QJTlGzMX6aRQUhoBOdhMaVAsge0q8O22XQP9fHFZFw7WDXipzQ+nh39U3KI7Dd+1V5pfe0o
u6CKOGAQrjjjhCSlrbdvGUmtLwrjBgop1bydqQ9PthhFGCMmgWNtoP1AWB9uskCsEzo+0yELmF0Q
b54xGKgvT6tAaJzByHb8fEX+0rLI4PECmW5CjjI2yYIMkkKbuky9O1glACGeyq9jlfmPlBsl5QMJ
PrReLbjtODw+ZHtpDQ9+p190Kf77I9hH5SCRoI1bn01g9/L/jH0dRu1k9K1HU4PKTR6fcpRRV1gr
WaU6Lh6f0pW2roQBJC45K8uAWjXh2UaK66pWZnm62/Vf49B1m6yXp2oUrxmxQJP+BiRkspRkz1I9
AXkZ06WpQXtjcAQDtU/ZaQKQijgT1jMkewP+Sm7Y+uzgxOPLaIYx+io8l45zNv4bIgkYII/14r1G
22NTd/ze5WNWNwaad9MgfmUlLa5n7eMKjingQUm8//joF4Pa7fhgKAuSZ9YDyTQjupW1OTtDvdFQ
eP855n3HLAXz86kuiLFkIOXb5EQpCCevuLreURSON+LANvcaew7MHub+ws+M16bpOkBZ2EJADhLq
q8aX4xUPz/wxJS0OdcaIWE9qny/aXnDVY9C/FPb9cJPxi8BxPjWlodVXgdpBr4sTuMYak2HSucfW
PUt9G0i+Ehbk/fjegIow4hQT4EJkg/YtA1XcpqpRXyuHMG4wpf+odwx2CUZcVjsVbCBLbexT5732
1TiLZgXbpJD3vDDuJuDHVxgyslsV2FIwic4gDE/TgHAXFlIgRX3kh4u/2jLbWFaxc0LYYnrX6RUo
ebKY0VMRhXHYEgkJsdbE1qA0SzIoDPn+hvPC77PKxfRRKd2pRupk0K3prHGlmxPFGGbrLxFQV9vv
oRZ1Vxd8hejnp8EA/3Q2Tu0WobT2Tqj0DvRSMAdRFP0jAngzRINS2TA3ylpc9Blan/S0jDn9KOtI
QcjF9wlpkBpdruL8/94OpG/14F0j6T3yMxMHDodsznho0xHUyKkdwB7rtQuPQBDWPscGSEFEzPPK
EOpfo/GhgHcuk0tXaCVpbDKeN8s9+N1ZdGU56KjFpaROiCAf6aqF6ES1G3aA8hfVOXZLkRMrkSYy
4gq71WNFRR7w1sQUJts8ZXwkUT1nETIy6sCWJk9HckQAZEbXDgNhjVxW/bCyL7g5Vwptt0t9uhum
UEyrTcCOeanfDYw52bVe1iK9VsXxwDOoinK0tnXRycQQgiztx9naBUBFcPjVFtqYTn61vAd3mgHu
RDnMQCU1hy4Hrpp+qqx3/n0zLE4ohv/iuAI6Ab1bSIQzXvNfHACeKW7y/vfDBeGBNOPgTvREKTkd
rTdUR6ZQOmf5pvBFYpJyoCNRa6NJko4sWurnpsQxPdPu3PaeaMNqa9TChiRjNhFWQKytNVFqqDaq
wDoeKk61/lJcbJH/N9kS5xL0CzIUq2Bk+F77UETDFuEsfAQfHf4TlY3iZU0xVwk2qFPbbyUV4Bw0
97xHc95JBHYhnJIb/2tHrDhxSwmBjg3i94MACYaJbRibBJeSR6YbBld026DiOWtPqtHwt9DNC6yl
9BaU5AiYEl7fTnwyb2g2BzDsUmh5mXDP1AUgUYp34p/nQpHiRk5HVN8e58ky6N6DYF1VXICOrof0
1GbGXz5+/nPTZNlrJwKC7Wy90si6wbBfpRtU70NJN/XiXnvyQMu5/Fs3tGMNshfYTfYmyF12JX7m
nVxN9vn3BwWKaS48Qs8A+UeUur4js7WnX+bzu7NeqiwSPAsoJsrmUeZn1O2z1JHG9CULPh67kCDk
Lis6bW2sJ4EbyIA0mrq3aqikMVbgbinvP6y0DHaUx7QLcXBf2midoQkXDYg68BZG5sLSCjth/jPM
do3DqWQdRLPyRZp/k0W+Q+DUxbywBd0t8gjxO628dSG3rX4bKC+MW3KSSwywLqKBT9qcrbAKyoXs
DrJLXC10GkqJqTukY8HHpyOC3gNzAi/u0QsoukmE6prWICJ/9YCmQhkgnGuPtSIaudGMG5zLBC6P
7ES92yfxRp+0akGDpEuXiWKu1wECRT/3UhS96QWoCLRJ3ysKL6Ct69tGtBS0wiNIxDJCwJD3VIzB
k5561olaagthYL7RRJ/HyJwDye5K87b9fQ8QhYTFi/cAw1uq1vFX9QK8SaUHyrM16lDVeHkZ7t8h
qpvFPGrH405laptu+Zy3HWpHSgeVrv+trSADgOzYpE3GPAyHv5VqJB+dJSWeQGIDgpzWGaMNE3u8
VPHrsr0a3lLGPqZ6HWsc6bw3caTBYUbvdEw0Rqvy3B2bPF5JF9iMrQhP3YTnigGvBcGZ5Pr9xQN5
/As5XyYHlkQ7JC/BGr2py9aUw5afWb9SnLJvn8cUFIxDpTzXygsYvOOE8cfYLo96C4euO5EMa2T6
YSYSMuK/avTycgbNiWaspdxhO4KI1jr44BDnKihCUym9ekMlhR+tsdMlsumDAkv7IFpSNE+Te5cM
znvejYQcmtB6ez0ESlAAS8NzOvnR3wgDQhl5ZRVYqVwihq34vZYLI2tIy7mt+Dx4C5qufxDwFpqq
hsUJXCzBvLRt6x3IbfIN0wsC75rO7DVV5J2I+XQ6jwIgn2FH3UG8V3VSo/RYJMGnUz8yG/C2qjOx
vdGpWy2DVmLuPLjTNxPZoGoWdnj/8qZv3QyrN7FZ7tg9JsP4/nBJzcTK3FaK5a+O1jot/9s0Vbhs
X5Gs17eaGG9H+zpkp/+zKcjvWLdMWYZEn0H4dZldfvtzVhOE6gYuFv/5T1Gj8h6UFRQytFNE6a6s
5+KeJSHP6Npk8rQkqY069WfNgYondiE1uJbT8UFMI7Ynw9lvIjWpzAK3Kt/2Co8rzFGAuMmOOvN8
GHp4EBMBmWkUrL1MsSTCoiOsvZPP1BhbBRBgNrpJPxYn9hSiyjks+fK5UmtGuAuCmXjbm8/e+r9x
jsWjBm/WhoHCmZQns7RrzcQ3iGpfn0ctftRegPiAyeJMwBGV03Nv0LL5z9/8+0vq12KDOjPqqIeQ
cJ9NcUMecR5ds0sozhLcvSmTi+6ARc7iji7j2Jroo05XIVXfkGQmXaz+mFKkXsx6Pl/R0AEUY/pt
0Ow/HPVtPkPMqD5EzrYCA4uMDifc/fDUSlygKKAfNzO59zc3u9iwmjYnrSzQRSITz/NCBw5wJxb4
dBJnRNtr0i+JjGlfbqXTotih3+s1Do9FtonzLHBz3t8F/4xVaAOJ44h111SozxZxHN5xA4hijQrD
SU/yMM+DwB0gaAwRJ8zGjdgGE77q0KBEEm+UysqVZ4cjIULDZiV1Zs+jdA/adYHMum7WZeSNkpnJ
6NknisXc6NSsMHE4TiXxCAGJ+d9whRRK1pFzrWouGySTD0QtDUPIJeSSXQo/OppinO1Ex3J3CAha
RWIKtIZB6aMIpHvJYQLNkUaA6+MkKW09GBzeKZJejeanOMOEt5rKfQuHo6hR5jxAGt7gB+oh1fiR
XsVALtvQ+kgq5o6/OmCSof+qVb2UtH20r0ORhNMvaBEOzq6sEi/dEkFgjE1AxcVnExeCSLerFfB7
KXBJXfcOQo+uwGPUH4u9mVYKD0FQKblrJWLU4ot6BvD558KegBify1iwOgeDjzkC7wimHma0QdV5
4KLu/G1BeqfAyM9ASCytcdD6Y4mIXYBKFWzjcFAQ9QNuTH0iYIG3r1rXEdIvo0KX4HnQcrMZyprp
yEBAOk99uO84GvDoe6A2RjIGUjRokw4xhmpE8mEoggxt9o8SiADecwvWQ8p2CTg2C6W4EvFWCt7z
NSpX6jH94kKs8ZqBtshm/3XSfsf1kiyF6ErgwGDR8IKX6MJDyXu/DHj+4rKVPPX4W3n1VEIxDT08
kAJHzRM5OYefz4KGVkDZoItjT2MKk5y1hcm0HgWFzN+iCkgs5rcSgk10S/jhW1JBuOwHKMvEpnta
QXNS84/qGNZYk/o/c67a/SQsdT2QXh6kikeEGS6z8nkCzR4xtgvaWF4Sjk2IVWqYtiRwCUlwZZ1y
QTy77ZvFi1yWNRa3qmYL2TuH23df4y75bO32rSG+sBXBZClnsvEYn0ux9Zowz3+nOyZahKIEphi0
Ag//JF7rZDuqZq0LcrAicBn4VKAo5q5CgfgGDLEnUIBSAI9sMzrfF0+LmUGLh9MSxs9IXNqqZ3av
vvK7D5HVNkBbltwHSKKbINnd5tTqVB3rDrIpqurBotZQqJ8CeZ8GdBxZgqlkil1L0Oa66hicYm7t
/Wuefz5gPMeOEC+wtgfX3aYLwjGFOJ9DLu+NKuF4EftJkUJ+V9uJmeMWT+tgMLHeBq305zDYa2HG
tsuWiPOlDE5HnZjKlDTk7oGceCsn5RPsndrsw1uIauT7f26di3lRlzFB6c3chUXtt1P0fKMnMEFE
NXr+vBbCIIdEcgLcFZwX3aX22KAM2M+QJY/BB/jchizIuC4oW9Fk2Lzc67C+3LL6YzIXHfE7IAP5
ZgbLU19oA0/cTxSfIiVLCUDyHGpXT8BP13rTgajDECXBxUSGsqTE+vwXOKCaFVE9hq+TLQSXdFc2
ozFj0JaRheY4Fv2VlzZdAYqgSM/WygrzaQFWVbyQHEak+wmwkPsoQsskOSqAwWI/2h+SMlo5SBeH
YcvzyvEPxT90LVTiXS+zsD2ebt6scuvmFZpYLwicxcBI/D9RKrUWkcOG127tHUNZSYkAGxx783eu
OvlSfG1RxJThohEL4BF3L7JZA+c8AGVJYvlHKfnPw2tFCDTUwrPCTMiskgmxGL1FA8mX+GsXrsdd
mXuEbFMJRjmDC5/ONCRgys29/cRZn5gqZCi2jofDpZp6m5xhcB+Nvr2GgjFPHXr4KQmMiSI5pVvs
fSPciMOAVQSrn18ZJp3PqsldFro/7SSYpldpqs5HjhqxY3tpF8EpMm35l4Rz60CEmyejTYuD3pyM
a/Bl8pLBMv2UQaJ+OTvJTLvi8+jbgSg1V10l0HbYwnJBTSnFg0qKmIXcz3ZaKUy/QtQgvGyqPqXo
5xLt2H+Z1yTyuvKNjk5TBuJFghddhNtJbjccfVBaU7WmQpOk46YrIY0Z/8jTI7u4CdBE08Ye9Js/
CYHY7VAT8Hqcg+1KtEy4rsEfT2g9qnbrF6yZooGxPhSRQqrNi0HqfkuX7VEcT/2THrkfqXNtIE0I
heSG2Gjr7iE8l8a+jwef2yspwUeEGCU4JSVGUsbnKqw388vDsuvOnDhkEH+QT4EXWluYnde68WOm
z/FGZogv+zq3fRQz8B5XsxPvVjo6oMYumHegi25tRFytMFrCXPMBnOtC0JQWkv+yChWbtEZUl0yj
ZnHT7eLcDkaq/9qyBOn6n2AZlrTF+gcouMQtoCwLnZcvnXxtA937Kjs2Rz08Gea05w5qiiP5/cgD
tjL6EXm3KztP7Q4R6vSRckGx9JC7V6tlle8N8zs9AGJfP28j7+1qBo9QVvUIxGfa71sXElJD29OZ
w9KiyFz2xfXE8Jtlv4FWTCY7h63y6/C5yRO3iIy8bwU0CZ7WeDGAnNeo1/9ezJTJ8WhWjg59mTC9
Mg6/SYXT52cYpoSASFH5jwXv0LoX3DGR9zzruDQuG077x61PBFQHj67Y4RrWB1YvFV+t8xLPWx6T
0ZeTWrpl5J8rG4toZBtmdBL5+OaBMPArIdmhNXswxiWqnMQfXJ5z2hmGmDYUQG6uFGvEuPG2lmcK
PXejxXaOEnp2DRb5wgs1sottFfd9uesh/KM3x0GachOnhEPlowwsCgL8oNwKM/7P7cxhEQTikNMp
h9Y4630Y+i1HgUCqqSchbz6AbGvIANUO3pmM0gKfijPpNBdbNXlwv7j8+Ejlyj404+SGfxvuul51
bTZzzsHiAjSwd/Uh39A3uDML+k8TzwBfE1UN/LgHGuHctPX5tmHOpyvS0dnjrU9c8d0LIWVc+wJ/
8dN4pU6+QFRXgep79rMw8UfL4CwQ5Ruixp5+uBLMqrav9Hp4iMvs1IYe+Qur4h0P1eUQRFKN2XkP
7icWaGs5zsk/cCQM+PvpnFVYKfHXq49yznMgpz9DNLdn1hg69NQd56JbA88hQ1wNUN7BMXshOKb5
rRrCNhIm6XR/EtDlhK5itQS/7bz9vNAcdcH0uizS6pwnUuP7lM813/HB5NLk7BEL+qF/yrLVnrxL
QXbZhrk9gvcoyGTkM1PxBFy6IbKuZLjV8LD3A3I6F2alGgAD0s69mYOFG+/zpfCG6ve2dMmooI2V
hwADajx4VNP60H+kwTKwbwuDvWKDPnb+EeqLlY14YByRtE2bLnKdVOeDkDGVM/SeiIrF5H04GE0d
TJYz0uwwukjoEuZ++LfENX7y/wr+R6RdgY8O3rvOPslaEsi+J6lMz89+uwF8hglTW0OwRk5dRAH6
mpI0T0xMzOMmc8RSryYxxXKa+b5otBTgpQM8t8R0/70rprklLXaC2H58NGJRiTIpFh8pKVgDX7Zl
p61+5s8SUS0YbcFCmwvzIUm5Qb03/hQAU2j8nmZxUmET54kEKLsLHuTmcBYRit2Ry+FE0hDknnaE
e7aTAn11kuMCYOMrWLZy6s7hM0ynDKC98a2toz4Mf9FxmOspDEsnSLZh855U/xAvZbjW5stlgKC7
Q28qnf+U/zXGAnWqJumr7NkEa6rUeIHdpkRCtA7O2jDGdkr3og2NWMgLQZ7TG+omzDUuipB96pUx
YXl3u2OdwDShda8+ArwO1j1aPqfCtleUleSeophN3FGAea8SK6NqU79KKI/LgcHqsnI3Ve0cZdRB
MINxrZ9KrhRWQuqtAa6+fNcMyCaB1slfu4gjwOZZYf3VeYIn2Sy4wEELZbWQGC+4zgqMZ0noeA8D
c08PjGh0Rz+wpFEbQewJn4m85WR9Hp56MystLKPdXlYJZYwxllgKeXSXgNLQ5EKqS5DRhailjxB3
W4kdPR3T3wCSGsa2XQpU+ONpE2ocb1zbpJhhTdcT05udrYMpO86Cyg+a1X5UH9zctJeerP5Fm41p
hSVrWxQo9BSK6voguJMDb9RwFNm/DOI9keJfx6a3UaZ4sKYYDbwDk83wLDfwVHUjDlA7LhURuwST
xRlsTVP2YCr84lfrHiIIw+H3UsepBTJrZcWbtP61Zysk3UeThzmGb2qY7r7kC8nFmTOqn/hwGxYe
AhHv87OPti2Mra6v8MVTqSUxLI+VfZPUUpp4GoddUH/acMRJycsjLqJUuba6EjU0pnbQPrrEjtcn
nRPWsZG8oOdNTPcup/xpW1DTGS2hPDQ7s0V4wemTn4aYgSwFdpc8iNuGPQjWvgl92HFfbE6XB2V0
ByJOL/7mqJW4wmX3nm3vs2ZaAqRLX07MLcdMPAQdmJbNIgy6JCxvjk3oFaL3YZHHi3fGS8oDoK7Z
M+2wMcbD2zZ+3TinFS4TDrTOOBHLcCQXbjp0j/IxueYpK0h/QAkQY0EnwVZOhw4U9+LFgg67sfCY
xy1E32Jv6C+zjnpEVzbDaxk1KcCefg/WsjyD1iIlbWQlY19HJf/fWpMjj8tejcnLbsHqaA9vJRcR
wRyZ/puEMG1w9Kqq4GUwVatwKu6FqClRnEsQc1hez7t0GZ1ymbWfRdEHebIjfFyqHY7izUgqC0sC
lMN/rD8xXJgJ3XKa+i5fcl9xij4MVt55P77KDFwnEKs3ZrHvIsa9/h4WhpQrAlo1HdIXRvvajh/g
pyNG3SI2aJB/Y3ggnuF3Js0Y8iB82kXhWgj0b1tfJi8dJk8OlQlyTlKKif2jijRB2ZihfDiKxhdi
DJLsRjfT2J66sKnRnT1S8EPt0Iy+784kNQzyQsKUTo6kJr0CwWsGlLPMUcp1LjKw+2QdSiP/5Mse
JTSfdkpdTExcmuZmZfPtgbNNw1oTK5kJ7WV9QOWMLw7XdsTHBVjpztg53ski4/1HB4KriC9NXuMz
mD6VlxFbdmwwxhL2iaEG+NCvGTbYKmWOKNJTNFrZZSa1pAeFrNSdt3gihBIaNQIJZ6nGdHBmbSbF
0SirQpfcFc6Vx6FJwzCKuHIdK1Px9a4ML7EtVFD3h8YDmm6VwwrG4F0wRyqh7HUT07/BfnVrAxWW
QDr3oEGj2rvyUO4xc8p9iiZJ/HLMFF5f+rK4LjIItu2I+eKX2mF/OxZS6mA+PxFjECmAZFbwd6ny
2bP51GET+g3HutNsbN8SmhfohlToeVc8hhX/kv7+pzK4m4sj7ULX1w8lUr9J+mhIGb8tmWjq8A07
SFmV285gkINPlAKaBXGtgGUUf4l5abngsBND20k0f7WVc5ZImQ4rd77LJTsRD4vzQnI5fyB4DlrA
hncAUvrtlBam4hUVx5yuBkMgg/qs4uXpwxXRJBGYRt1spxtLUXiccXivWCWAk1nS3j5Oi2iKXFBa
vOMCXX4z5BDCRNuzd2ZZzTdNleRFO9iDbS/7L29ZUOSYnme1272IFNMXQPD7kdRxP819BC3Wt64Z
YEEFiiK3q0ozKhZEeKT0fwcUeVSMhO/wYrnhJVSi/GoB6ptPyhxYGuc9Bxn9Ec1szICUgzHsVsZO
pkdw2WOhWitlyMscyeEjM9lyiMbaX+W7R0Zyrd1KbaCEGuhpXC5UwX2mvxH6Mri9sfmTIZOU1MP8
fT0sdQWnV+A4+Q4NqDKOCbhr+CCa6QyfOHu/8k/Ow8RkB4NaorH/2nMbmoI2HNKeqY1t0TZd2d1g
W7xnerwQYvoX9Bq5xlvHfFu3gENLMj8z0fi0C0gYrUaJL7QsuQffcFrR4RMrN+OyY7kSZXwozKgT
RZYA5FwnilE78jZkj6lN1BYBpIKeELW8eLikaPCPp6v/mcEaH5KoXHywzOeSho8k0hz+y6Z1HDX9
4ztu8GSmXbRK47PucUh7jHM+DfQDySmH4CiQw7zTxDlGmXdkPxpJaOTkNt9Pj7FDj0xN/zB/r1bY
ynGk6VJxJ1MO0UPw9rIAFLurNaWsz0IyKsQCJjPwPFCFuq/Hj7ZqEKC45flhMx3z7wu82vGcXKrU
yd/4Ksb6WO/B+IZE6ynRzG7A7weYVsVxWAE0enYvN9c2+9W/PIFVur2695QUL84sPMQ4jZCmQ7Bp
7AfEXOvwDI/9Z58zrPKEDjOg73p9vP/e/CWb48B74yn/mJWgw7cCyC3wpY9V3V8QzTLNG4e9X1xW
Ij0h5MLTP60NY67zQS2U0k95YkhLjGFT9LOwCSxKNEMY4d1hoWskgVKwxuyvgEJsquETrK3549PK
otLsp7NYqp4rajNoa+wF2/xNIrHhNqX2JblSFuN4oY5eRpRCr/X4DRukOp/gIHM4UXYNBS8loqv0
PrPZ9O7qkKQtLj/7mAybgySuWE/BfgKV/b5+OY4QWGkm2QOPZ9NUfzyjgab5MI07CT88U/dalz/v
OHIHOZzZtsqHYDxRbMdocvm5tA8B24OdxYY5lJmsipbj2wKRUrt6TbLRA3bngyft1G8LE7gi0Idw
bihlLgbn6iSmrYmfe5zUQkUrZLVzDy932Ok2F5G5bhdEN6i371N5bN06jNaNDGKgx1NY4Wn7hBSN
QXNfTsJWH/luiNondwXgBbPVh9aRUVullsv/B2Cut5k5/8UaCmkITmJ9XWX0ONtTF/zMWWirmUrE
+3z3kEZQ5MGPAtCXCuCN2SxDZXG27lHVa4+n5QdARmmsBVjsMy+wLriVZriA3AYKtro0Zm72XNTl
CQOsfkL/a2cup4oZVR5pLJnWFomMmNZX7ns1ExM/ldiOdkU++VetSLCyePCAoRWpK/5yzplQknUM
/WUDAXlIl9AYhneF+BI6CiEnVzzSgYLW3C/8pNGbsb+4jCnvN6JHZab1a2FWRU1T0+8SV8k9uwfr
YezGHKOOZZSBlLd6GGThWpsLy/Qckw24MQOhDON+2xQLD9e5wDntkBW6xy4N89Yfe2OdK4/B+k+r
cAml0m53mIQTD8e5SbPgDyyY4AGbNAlaNhesOLhJZMkTXudM94qcBZT4+S0k9MHq6LlTuGpC9xaV
wtGd3zRlxnQfRQDs5KaV8E/lhslaSI9rLBrj9c3wOq7zfXo8+8eIfhYZXoh2LnvR9ged2WKkLgvw
TcgZnrNnrCpgtWwOCj6BtQk8uHUqRxmOMxKbX8T3r47lt1Wc/CJ0NHMf6T+P2xZNYbPc1XHo8z+F
tDryjDctAzP9auAzobaA8J6TLnP8LlCZuXUpHNNp07qlnXrBcW14frx3623hMwkmi92wBcD/CHcY
4G0dYSrnVVDthygTBL+VRQZF8pmj/WI+IdtzeCOiMYqqKPW5yTR/8OxshvpEX1R7VoO2etRf1feQ
MzWc9/PNvwnk3IAQK+Zr5sg44WWWvK0JkQP3w5ch4edCmYCCeXdy7J1dUfZeTJ7SiYpt2R5XoRja
FqhhXWD07j8bJlW4dC7gnh8EG323AQIcyRlLL5ZXrfn8yGQzr+jsAEFG5fecsqLaUJuORLCfQBTn
c9/d65YavTIebIS1vuvMgOt3/CarATsVQbh2yDAEAizknPZ5FVeV8oa+aTLIF7ZlpAK4HX8/em3O
0UIuvgTkoaChEqeEEvkCIaN0M7NCrjnkUKWo/v4KNdBHWuy5q3D9Sz/jvZr1e5aB0zmBxPLzf9sb
fQNXuNd3A5IsDuAect0oiOVHyT8ipJiwu7DyICNPyG1fXZ0rXS9e9BKI9rHr0aki6gSfkpbt1dg8
lYJ083ZWSLGJRQZpDjxZrYTGdFjpl8FgFBRxy7m9D4bRaKQmiRvasoEAO5IXMjKkG1CtRuQXqfyw
nQ+4xNChoqSqg/eexn4px9Bu9/8sbnvMDXA2LxCqnbVmFiPTQBuLBJxOdrfPXwgMc3reI3hCCX5S
i4M+myzX5vNWp/y4zeQdPs/hZUCkX57w0KBGZZaSNClnBLebt6JAOaT1sAcoBylDWi5YwjPYcmAX
11VAMzE0fOXS6+lt0Xs3jt7ByKYhI408Dp0nSLC5fL9yt4Acyn7V8M7uHbsZXBGmp+mJxY126S6B
WoXbEQn5FYcyqX7Bn7ONrqYFWxe+NdJKy07OKYQa7+MJ9B36nExW8g1LHJcp8K4DOPO8nbmjqVjP
dm9DG/LE7lDHl4AcPfjmXL7qdtatQRQd2T2Na94Ex4D/Z31MCpu4UlOvyAqkFTjv4dAReFafEVEe
dT8tCd/zLX9wGF02Qqsk7JmcpbyzRvNYoh0ntIr29j561xdyStWDnmEJEngqV5h+JkSy25Q/tc9r
mk4LGw0pK2/9oUUuzatl4imIYVN+yAvr1K92SUFpJF4SsbKAqXqOav0d4Hy64019xTUf4eglJ5ek
xZMg4S6L6TEbZ7puRvdXNLcEh2496sOz8p8Erqmn6lPXs4vbscnoWCE3FR3Vm1iuVMNvziWJIrSx
aBQCTPDamrU9pkcAfuwyYWEHN04FQKzzdcvpyjTj8lx3OzTtDL2X2opMc2HHSlwiVyigPAnEswlu
/UqNRQby3K5XDp9l8wY9OGQYmjGdfVW39WWWJw62GlvRuntQD6iYeLRhtjZfzodT1M2pH0rSBBP2
IUHJxWiSgE+zB8Bpy0PBpnJrzcBy+9LSuWcerNec8DAAQRD+56/cEYd9QbV85aGDuuhTPWLrwR/R
Gw11RSXmwaBdl9Yvbh+AgPjv1PN9lbNM3N9KdEXxs36zxTj+DD7eXsJ2DAFXxeiFogpcC3eXPSNd
WG5Z8q0jdBmVTSMeNoHaK2Qp04pz+CmCfIkh3xzZS5nA0oDWcg4nXLpgtMnWTS7pcsRq9ZZXr0ho
oeP0F8ia+19zrRcTv6Ti1OGQrC2u8Byv+SKTrDh/EqtkzKxzUSWHAZVu7ejt6jUCwZIMlgnlDK4q
n+CAAbL0rpYRmN8+UlVaYVFz7P5GMh7PnHAEX7nYgp+BSHO9juH3RsFJtiUiHPjNJC85vrElT7RR
0oZgGzMbL38UjaWrMYIZuIW+5rNXDX/FQcqe+n1k3rxzOHLcEH2EmfOBqopVivvnWvYl43E65PxO
1jPO5qyTpN00sgqlJDTxZTociCb4ZZ8It1lw+94CehGA1vaAmpOHDtThSRgODWmLvcX1Rt4MM/JS
vmMwO9dQmzk50RcxyVsrz7YbdoqQjrC/Fu6ES2VTklowi6QRecDKneZiAnYrgpxZz8v38BjG4M/k
uQvrKVwg5YMG3KK0w22AAQpNpqYRLgDANgv7tJXdwo3HeP2g3IXAZLatJZ2iWWVafWPg02fZ8Juz
m+xqYPnQw0mMg/iDxgBf/tvMWgP9T9jdfTyXKQDj5ab3yho8+WUVt43yxai65awydJQQFvz5E/qC
e4IzGM/69KYMpkUoA7zmVF3/ALqSukS8mYXjqfE1W52CGgC5M1kFrnnqodbCNH6PH1c0dxlXMX13
XhkSvvXGpM0AD6IuqnABhWCVlWlLxsEe5K+OIC4BhW6EOJs8S3XvV6/M7A8Si4VCQWQYNmYGmHlE
CE6iHWUbyJZ0VhxPWpbQyGYhuLSnFPmYebyip6bUCt+ITffa9YFWNEeyCzOARUptjBAQJnSNm4Iy
E7FFAagEknL6mSglbskH7UrM9hUDqdqVqitaVcC/SE00xtlvBgWsesiROBSPK9FcrugL0+cxgk7L
p69q4+zB+dQ5uG6CnvzlFpE9UYk2zeBmtebJbPENv20sqZPKWAezGiLzqJjdt1YTJLSEeXY1Y1b9
CLdJqJhDwptuc6jJxc9fZm4UHXiktwnu5Y0e2QofbiDgmINrnkCW2c8WuVqxK/nKlCBmdLoGCb57
r1fx9Zayx+NrmHVqrMcUEwqFGCrv8YO1bC33NF16OiFscNO8Lqj/PpQzf2a49JfhPa8AoiuxZphQ
dLxvvtKUXa19abw5UmgD8Bd1N/3glGNqiSfQ/gaMqlCVI8QA8ky+dBo3U+gHJYsEq8hgk7GtLWTr
V9F/DlefsPkn2iH6qtysmhPpW3zuI1sBH9pV4jJn4W+zIYlRQ4+1SKpA+bXRfsTTzPBsBtvg0r0B
8JDa/hAt8MehQrEDc35igUqqQfgMpf1K5M3jLaygD/juwPZdjGiXTfmJYA8UGmq8P/78Ddk0jUkk
YZr6HYw4gTO2E7DrBowIIgdCofq4bIMiQfE14if+pl1PkFKbxpeZNXncunwZG1YHOqYKluwn3YJa
Pgn4mFJo3V7T4FZ0NK9zEdBM/LOc7X+XofNlweCiAhcSxy+TSHU+bvVG6ux5tTwlBL/EjJuCNkQP
1sKh+t+f7hnxKaO0+OyUqfaBh2/t9Hq28EteD2eFmk6Xw9QiR9D8+48bNOGHIxSd5qZW08RR22kC
3GdgNdi633koNU65xC8CZVJqJuV9PBbaFIjVd4U7WSx65c2Dc1CJakZM80RUUUYfITWbb6jhoGZo
ye241lX6xqJa2z1hHwGvwsPHtufzixM9s89Kt3raXxy7HOw85H4bjstitF4cJ+mH3xso8AFTmTjm
sZ8UVGAlUUBFBJGvF5Gn+NzCUay/LTFBXcT4oFP8Sc1yBcOz09q0wYRQrcaacmADmGsSj3VEaR1j
NMPJtJnvErBifgO3ZWHuhnc3Rcqu91cthcEcGcje45Vs6dD3G1BEvZPrBFQa4wLm5qOktUBVdfJz
e70oBK7GMXHYmjvS7br0AzDQHHsmSkDRqNsebB8TntZooh7lSCQiry93RX8gsqaLc+ya+P0EUEn5
FkB1+hEvqpIBdrw4r/AMnw5uQqTyhmpXQmiLF8/7WJZHfwPXVHEeU3txbilzCnsUU5HwrU6WP8cU
OOUJ1fz5ZXcm/uXYiiYAMVjCzz4kIMdtkqOt7iGlfBOazlpBQqEptKmXvyK+tVqdi/8S+3MNPFti
oOswWi1Nnj1N9Kbp0CXEtM8hP2M03cel0z2r44Zo2C44Jc9QiytdpA+OeqNOjThIOvT7zqhktWTA
PeyEBPiAgMYZzI8vRoVxGax0CeAuB4NIxaqxvWJn4q5YDn7he+9kKy3wfyQlNuLQzG1zI6ay5yZ1
4EyL4+6mzVLi3CT5GAb/BLOCX1YqWd57i0LM080jocq7OPe/y5u1Ig/JSsvKuZlP4taflx+d3hQQ
veEBn0SeDSPXVCtvKdgO7Nf8yuKgAlyPq9MB4jULJM9inb7YEYU3lhNOV4aC9G2RUb0TZGnFVLcs
HV4Ky5pSiIM1GgOQ2h3RvJkrJAUpzAHpSDqy1lflOqs5TgjwUGL8qqZqvXquFdeGbX0FeH4x2oSM
1G1OSB4qUDDFQBqPmWTayqBATe7Ah96PR6BCsn35Se2TPU8nKp5zkMKpQ8enhTUZqArVKl4k0+XQ
ma8U+/APiJoyaiAXFxSsrP9YHES1m0ToVPjaxPSfD4bxmeIyRQZc8b/CSLnutGSjMU5do1nY/L5z
8g+6LH2CA1CbEVj8/oCmzqKwwSm08g8sXO+zDwFIJxCWppYJoWQbU2OiiK3XKVnKoy3H5Q34pZuz
u7c2LI5Dt6cwpMZHq64ghTjf+jOhW+W/OU5Q6k4VPM0zp2DKyT0+qMkjlUzgIelqjfNZK1x657qK
40UvxFojoD6/Vofav13yeV7ubsSpEHKbo4XRzqC57TgG1UZZJQIF8T+R049HMMBV2JAO47EKKXlb
M+bochj6RKvsWdciYydFkRbrCyFr6SRTXTKYq6lbQo7v9CvV+PPswM3GxphYhmfl1Z1N84Rk06K0
LqK5J8rMWbcXIe8TpRgeYseYHIqg5q94nS+Zc3wI2c8qtvkblupv1HOL0b8YUA20FFxgI5lWNcya
zYBZelIp7pyQdoMyvMpHPD9+tWAXHJsOmqnFyEC/pIALDxODUiJ5yrysP6u626LinzuXhyiETw8p
GMu97yE8Y3nYHShIUxHCr0OG98R8cvPHScNYBVHM/yKvmkQkqxC7CelwEqaias/t+u4ktRWTASYE
SgFrEiv7BmKKS+UxCSKIGZsOr7bbMMM8PMRsLB//+dM75xMd8PLl6j3mIjxI89eBGOSnzbdIKORi
kBxczlefezICTzjbe2WcYE1XoUZd8DX8Ion/QdCbzzik++IKVnPYP8WuceWeoQfILUuJw5wdZ76c
uEbSTnI1MBTv/tFZmfEPGodjnuYu1otR0TI5U9mqIHND9Q8QsyOfrkoCuO+mbNURnpBkv2OY2MBS
7oEADum9zhg1+CmXI90mwH/y2NLSLJhpd5/ez8tIh+YPlFtnjcrEM51Qkx5ltWAa5nWxz3xcsBBP
trbopaTfkxDDVyCE+STmYFR1q3JgffiQzZDGKSHDfV6kW866+VAL8Qc2WMU6bIuf7WKadzUDBIkV
88IoxMUwyK5gQbBRkv2yJgP5s16DwqVB4G5YwNDOkbJjeqqSNo9R1BwhvnSyg6NomLrlg79unRwI
2HcvUUjhCXtVRkLGoTJ0+LStO0CwBEHLniCUtno5FoLPjeGGZOJeQUaxwaiyvUMUJeLrXUs0t3FS
h7+zMIRYEjq5PqVGoh79MeRmPszBAKiykwOUR5t8MjbkDFkmOiyDQhSRvyjIadLFNUmbDoELW5TG
eUxi6Lem3Am41WvepAObggxGTkxf74NRPvhWMDV9UBcj/1qMMcackhveXMqb9wd7E4C+OefYYgFQ
yrUp6z99Zu1mKllbyTZixxE7mw5RvUKuLNwRCgMjuFBhU/dUkPkT6sNTpjVoSyu7US9o/Y235c90
byTIZSUoGsOuFWgymcjmJzVBaHg465tmATSOW2E2zTrTpxPOPf0kE7oFRm2dilw0ZSjclIcGyiB7
TKpqVwP+bI84E72YEtOU2mv55PwBtsh5KVObWWbNfPHPxxjwCtjwwKh3+jQEw5piJirLZY3RS6Yu
5KVOrrUGZVSiMycLBiEDEdH1cjHAWe7ztS2b1OkFiRghVrL/6vdY3AbQqpraX00v3la+T9KHJm31
h7Uwe50aZGIY7rcee07cZ9IKYwPEonzlqgZ4yK6KxG/3cheuc8Z/MLv4C+0kU8onrGW01UUUuX+d
o/w7hmWpl1y+8CWbm9ZLH32ZRLUkFFtGf6vF3/H0FD7gAAr97e0KuHzQLjl/pPZmnOOcAHqf7w+j
tSALoWznZc9mJ6jbKJfRi3MvuHPz/mvsfGWV2tQyNkdrev5mOLdRDkKwK1eAUtRFKyEsgYE5DDhT
aGb6z2+wqEv0gMVmkTeY0KCvqvnlaWld5gTpZdaLZCwCMkGgF+eOrKyTff64UEJ/4WJIQvEpbBh+
G+lUZ9KU1HDE2aGc95/ntYLXqntdEh/VVPL2kF748oQ52PYdyp6TdtDlotIW6F4GVa0Z+gZBQZkF
ZDajmBDcacBl1SqdJfJwwZjRzhhJC011DlWmlL5LKPw3efF02DoKAT7hmYF0o+fQkVqyglgsbWYg
TyXzMMi7eBgKdpBsPzmasO4j7eicqSXUDo6900+Ug4HQEur5nbT5l3ESI/jcjHREBEXTvWJAZ6wI
3Tf/OlaMY+kClHZoXHeI7e6C29GyikGZplU6o6zNCkCLLzhHGU9kwXZQCNtXjD/FSiSTexoBGvOn
gzSi5tRMtcfeNphVHtA3QafFfRMkZW2Y5JWRITck1lX9f3EOGgsbXY9p/i5w6v7lMPqV+UEmehp5
9ltptejAauFqTBiLbpSfJm2bv3kbS5xlpzplQWhTErnfhie715DAjMAZUEyArI3bVlC/qjEdTmeO
fmydYBFE+2Gi3pCOhE3lCDSqDR0HWkF0sBEJGSb6VKgkk2pKV9W8HLf2hUFzp0jSJO96GH6Erg0d
2k7xv+zMPPdiyhiEPA7PsZnUYJaq9VcR1bHW21xwh6j+pnjBK0fFUKGbrJD/hFWjCrQV9KUdKgcp
LulidaVnoiBoliso3tNvGbZ52+d2YpbbIUD6d1p44ZfY6paq+VVWgoxxdipB+L0LOpByRUMTkDkz
zcMPc21W9MPu8gCz8WcbN81BFij2IiFsClcEfuyKZ76MdVIPhxyHltYkE1u+nPd0nDvEQ4ypQ8AV
+04CTuYfvtM9DfQarANX4d7V/Yzi2LPjt/BOiuLpbUGQjAbcfyXjoZYuRY7a4cOTPC8T4A+2ZEGO
YEP31Z7J+72oCD5lG76XLJDAdePqHONA4rHj69VeeUErnDQqaAYV9ghnO+GElhX1dumFnQq6Fe/o
l2vSLYbboDirkIWRzvIMUHvlFcVHhZvlx8PFl7aUNwqwG6RK1tCCr8X8P8CP5hpj/blyklKS7eC5
m9567Y2RG/A1JJvbKrLROAX/4WKHy3t4iH9diGHh9Y1qvc9NYdd58nieVW5sDdIVtCCjj1oRMb47
jqhlOqCI9FCRNdWQG+Z/XhwOMHDN2VKsAupCxXy5mpTYMwTHWxcmARc6ixuL99j9cyfm3E+jUQ5L
1c+FBSvaQzzC/VVrwjnE1XozN1zbeg91aNJqrNWFf4OY2qoj44/U1+J6QdRAZHVBSZhw2N3RIjJM
TmWOETCvF7uXvxp4cErAxT0CJ8nLYo/rUSX0LtjZUwtIQmGlI6y7em6W5vy/Qk/aax1yKH1OaQeF
Ttyywpczb4XwQVf1RDZ+vGoVUQD0r9icGpFkoJOT9ophzPd3Wif2JWVVdsBGwPQggKukAvuYCapA
vWfHhnWvFeknSfP8+Pb/fkXDQLKNfqZSKR5j+O99QR/i5hGfyMeehRDaALxam5DTKTurNcDZuQYI
1xGNEGwLo+hg6OMl1fBi5FbrhcqH2gpqcudSy48S4soda1qLOqt8ByT4pIhkCj+DrFJWzPScEcxk
Ss2gHobRV2AJ6oNu8Mi3aXzVcJeVesynbnQ2giy8mBMdJZTa/ghxsi4f9QS8TeAgxWx+DaoWIHHl
5MRzt1Rl2echQqxQ2n2qnTc0N3jVvI8CIRry1uEbtWDYeH0MhFd4Q20Ot57ew/BzW6ajBvqWmN4b
GgDFra2BR9X5saMvfVK4L2of4HdOme8rj04gMe8+Z+X0vx+rC5FE1AVQpVfgoWyFQ5gbmRC1S3b+
dvrrAnFF0KMDv+a8MRTK1J9DxaAWt1XBTms5rTzgX9aSW7m+Omxi2Vn/qQcHfmhYXKizBQzjy1BG
0I4hX1wxDY1Eg8XONRTI2JzT9TOGllXPiVf306+py6VpHPmJAEM6R97OpaZeZK8gCP7Wlyd5GA15
02R2MoHunICtJ5CXwUu2ufFjBp1pc1udz6CjZTX9V7+QjMwpm4d+xvUikqC9LFK72y7YlD//YooJ
j73hmpniXwbWPICHg81kWIQgKFtS0inKahtJOA+qpEq5Cpk4LaviN8v1uVEPKdQsSBmhgt85J62u
IzZyi7zKwHoiKwBSuN2598B6CabpK/rC75y2J5Jmwz20+JFg9vpp43wVquPUdkE8rQCkSu/H3JL6
2JeUvpLGcg/YwKMUmF2/RyoOHghZawONb45AcFEH0Dg0XFPGrvJX2XRDyZSPZkPrMchk8aTIfzia
0j6BUfGb8uCeX8uE/z6/SFAG7n2/FZM8wGSMY1MSOmp8teza91uuc7ocZLDlRaBr4kxfumFb9SSp
juP5U8ekYxIKUmoRynNfYYOlrw6Z5QBOMKE+8V+l9b/fSghfScy5Ok+Ib15DAdJ1NLf466Db4xKq
br3aDCiOpLXo3H/GqE+DvfCoZzFwqlxOTsTI511cP/pYk3Z2PsBMVXhfu5xuz9FKyZFhxGd+bOvO
6ZCwDmpftNUatIIOdB8oTy8ca9NyLveQriz7pM9iORP7cy+UVn5zuZVhaiEm2a2Qs06u5mSdZ9HY
IHjvu9lamfqDfSRNEogBaqHI/Xn/qZrOtM4hCjtxmwgohnWzhlgP4x7M07MIFDH37WfPfWcrmlMR
WOOJupQ4KnIhxCZMspMrNDkt/aRFumtfYmzx5dVF0SYmfO4Dkf5cx7Ns6/viFqqbFvOePT8f4ko5
aiedWwrZ0ReRQi/d1fm8JPSVa35C41a/OI7O+BqEskX9+MfvQTiIXuhN5sFsW9QxUjzbvs9AjJwb
Z6XkiTI1p+3LyIU4ONsk0YShqMdW3e5+mPcWSz+aQsR+WtBlSlPZzFDunJ+etZU3rlyinfDMVqyQ
ROd+yBCZuXISnr3eO3f75jVtJzGs/XdQbPOn65/jN4Lg+51BuXaT0qTlJzAV8tANxQOV58NDk0MJ
nVzd3kYxSIWaRg7Jk+n99PmOc+Bq7zHc66Tg4ImaozyF0Thkryq3ELv6uG58cgUiOtYVhKW4gLkg
VG+miGLkWkj+95cxR1qykYuYBgwEC81gs9oC8cT7g9um4KuGA3hYS/mMBFGFV7RAQYxU/59qjY0e
7TochKk8VckSDFMBXUgCZcPumOWBy6aNCvFgD7m3Z4unPVk7ETUaITMFAJ7nk0f5gH9yXZVxTQWl
IGPfODSCaXYItDW2GSWeOaU2XneIIvzb0iVoQ3Whr8y4WXuIFtYk6a2wCu9Y7bJe05rVDmM+Fysp
BmZPWSGIv8L6oj3pKjXc4Bjg2BeFQnpqc3wDPoXghFR6EB6q3E6Qj+CMwnRRBprGfTKNgpjRZmsf
Dcsa2u+mjsMhsQ4Gh9onEY5VI/GTmHqy9KfnZgCr7wJAigN1m78/YvLh+qE8H7z/NHREiXYNjrxV
rAxKwC4c8n2lEoZ9D8D5qtLF9nzM4I8PfQgZzJteLMnWafqEvnZXJh2u4h/0hEi6Gl+onjuC9MIx
b6AFprUMdlyJzgzmTstI8CHZwRehZ+TWTgPdc3yDrfI71UGhoVuPudaB6IDFvP9aG9TeH8HCskQe
BnM8Hny0tHtbC9l5pxIUIWPS/1x6ErfymGz2FI6+Zu846K29eGqr3NFqVM2NXcCY7b/LU2xZ2T3I
xSzVLCjOLUJau9XTYhWsqZd/WUWwYRJ6JnNrcyCwz5HvO8/pMnwmrIlWsVPEcQ3yIZkSzMevRwU5
18pM09oG5spCGseOZb5xyshAngVLv9WV63goMYuXKQzrNmblCS/bSa2W3c4q0DUQMfxdEvKuCXcr
08jGukYgjESySzJ9e1BamUgKPWdvAo1/QwyRu2tNfVwkIsgl6u+7VyKLbJouVlWTlvfKajUw+kPj
vfWf8I5LNUpw5t3Dn8ZCk4eMFj1fnvS4WpBhH3dm9T7eVLrVPTUBGJ6OSgPW8F/VhS02p20TW97v
v5tFIkJdDy1ttAaDz3T7Mogt8BcMuERtuhbtjMWQCLmpOcKOv06t/13qX24adlEFWox7IAMKnN6T
o5CkKuPFaUtSB4saueBRI6MOUa3GC3rovrtkJblH8pzysoiKyOCgBzfHbxsSBqHrx+zSyJvEDxvx
F+OuDk50cq54ccNG9LSMPxYB1SoZwfgKibOzWKq47S639HZJmqG79Bx7gsycnWp1KOkc2tjCugXf
L7tfbZ2SXiioPW1Huu1CJCxukDbY08KCyrqXxgxJVNrIgaqWOPuWN5QmuvxIxpKxibO5sE7V5a0m
ZsOtiTqjKoZokWkCedzq9kthlZq8xNwluk1n/ZrjAOfWhNwr9uvuqZVYkRFPa2hPs1IWxps7MYdg
RHVy82grB5ZjwPacrraX+qB0utUaX77aVaOAVCAuvpFcaAG+m5chh0oaWdQHc8TdLRjUAOtya5F+
UEhVcELWzTIJ3FZb3OZdsLIkTkUSId7fycEVPAd4X62vrnriUk58rHKQ7adny5527YqUev1zeOIA
LL0oTjGe6tuB2Wzqwmhl7stqLc5svFWET1nDZIi8HTr26m2YX7Ojg9d/iO5NMGwfS6KNp2W6RHkk
pu2FFeg2v8hrRrV8GielH/2ufbcuk0THcLikSUqigogVFaPnwSodGi4Pegmxsn12BadL+p64RYuw
MOe9HsFfMFO20GybaBZ1VfRcavLMC4b03yVh6nOCxrB3gkM7fWfezKTGit0oeJ8mZiq6Hc1Dxnf0
1XSNVd7o8YeTqptWLb3joHkS3LOMvXSUGxr8pBs2B9ENa+d/kebnIaofSCLA8AyblhdyN4ajCRxT
bCej7w3K09jeX4e0cgFEwMCHDHoLwL048JwoK7T+fwg4WagLOsKqSHRBDozn7GhvIPfzAq4rSBK4
a4aXD+NEP7QQhad0/oj2wAqJSLVHAKBaS5A07wDoja0SwcgR8lS5lKpIO5NJiLV5HP6PhRILlxvD
TSEi+ykf7rAaYWOPD5OgUMKrFNk7p5CVhkbxDyn4TRGtVHiEyFDUPJtperkI/wVy8CJXv+RDzY8g
Q9ZN1eEvCS/1T2K4+5GdahN8KwurKSMaYGc7qQ3QR5sheGg8xBndvJHELHlYwVvRyPJFDqqOVJsi
RjlVlRXCHOKn03H4alKKLYsmrC50UQowUNzaX2zJh9E0e2Ye7qqLhLanaHokNnki0JI8W8oyl/oz
gZZPv5n4Dz9jAnyf0L5ckOf+nUYBHhj2A56qzOvjBbK7FPPNdeWiggJ/bD2/Z1xoSoebJRmIcbo5
IgkrssBM9qCe9O1+cqFE8km6vLggpDYn53d9SIm0gE0eu5gO2NUV/Z4k6Ng8GbNtIIBzMte35xVu
N/ZTfmsdHLk863X8JHMJdhw97jfFoGWhvfQqKzeo+pRoXjginjfDJizZGZ/1lx4EvYR6G/rwiFEv
uNwgybTVfD0wEYs8O9bhaLKfNCQUeBVKc/1fGDaqdXlpzzqz7us6yomDUjMlfBzG9Ns6XMwolTi0
ZgTCJjyiqs9RBvJKQhgTkmc5uv2bOomUYRC+tiSXEyxEPXrR6lykdG6srkOGaM/nuFbFoWSQfjNQ
8dDyJM/glTDdHFxsLS0JJBSriYJdjmR/TKn3YyE43kszWz+NvuGs7nJKND/Q/7aiNOcxmo6xcKGE
QJoJJhuCjdGd83n0CPtCeBVA/kY2tualPORNejWAKSywUa+yLW/jfDSUtoyDwJrAVDPAElePlwbV
5J6LW6FMxGM9KN6pYaPRL0cjx4t/Wmf716B2I42qyyiRnXhd4eB2DLaf+2qpsrm0hRGTcfhWYvY/
DoJmdOca6MdMU5RUV+H2RZqkJHkW90HLx9t80/AIrpdzO3KwwV4YOSyNK6lrsTbonfLncEGFuQgv
tI4L0qcFUyDe4XyAfHCOsIsDQ0QDb296WocHuK4hioL4h14eBby1yPT6JE1791dyxUoc+SwrEbMB
sFgpptyZv7PQtQO2ENT5zjpQigHEu+gk3ExbiQcPOGwcZIHJAvzNbNkhbm/oieUoiKorMY9TEIOi
p3r/YeYAY+5w7A/oBaJUIITpTAsXIU9q1aHoak2RwT7PtvqP+2xyHW+CLMhoNmek7x0DvOz6wens
5y9bCeoGaQZOJSSlSSzbDPp9Yes1KYdvwI9yDds3Us1waBNjTTP0tJnWNKjIS9hnS+FfI9j2wgw2
gf9eNYoDkRgLq4yGa1LWberz2wmEHYxGygQCzXDgcLR/kvbowp/XljWAr705nsSeYbDrOth6pTlT
WdGD1jUnyCPdbCRYxFQjvzvyTNcprOnGSVU44AsJShYL086VKo4fvxp0BTRM1NTmxEXrSq8Tw7FG
PtoYdrHUQAgqIzh337H8e9aLz7BsQVrYyxiXj3HZSdg8u+u7eT6ci14OBvrYFe8obJUwb65JQwZ0
NPn+DvFQnsRl4oR6ws4Ad1yEXOn3+YhCNFWbO9beRbTArMqwCrk/RPMmiuKAGvSGSP6YD1HilOWF
CBIWv1Hclf7OvsV//Kf+QweTrbLY6c9Gh0175qEWZpKqfRSHcKPUvRpp3hfi3lAStRAjbwGYMpTL
T/RozFVVS32qy0AygNh5m0ULmE+vb2/vVOUjTSD+9cLd3r5YSZmAms2A9daFhWmLvnsYuh46mzLq
zndwEch2YZT867oyLpl+pUcGtFIBVzWkNKO3I40pqFVl2Pe6zz1oeCYsgCLuH9EWNR1hxvdLwr7S
IyntyYrLqp+vKY5xhO5n0FqHvedwRreoyImJfRJHv+99qHCVXba55JQ/VErwLxXw6jooADq0NUNK
YIwgGGTa9RgK3aMjme823/LRAiTvivkVvo1xUYuMjlfIS2tz4tEWbWdoibERiBsYmyhFpYD6dAPd
OHuIzBPyDWbUnOvpNcW5sUwQf8ZYc/ZYZhm/EeEAVWphxI24m80qOIf6o5d01jpfFVV8E49zg1Dy
zD/a5DFgLCVmTT5jg1yBIiYhu0nQw852zMyJprlldHvFrMcI2V0/nHRbi/BoxrepBB8R+dYmbOc8
tekXQivBPh7VmvdFTeJhPfIs/NWhGWQBXdCy5l7OQGO3kUPZX6Ysgpl/sMwI7QFzunYw1Q5WlSDU
mWnH8Zjjsn23j8pAsn0kdCZmvRE1eD9W9H0Bbzw1ka9jJ/9AsVWURRUspMompTmA0cHpv90QHzXw
FcxARKWZLQIhH3kANdKBr6pmHj0+wwS8pxvUE9gj/uadp0SovRmVNlmtLC37GRH/lv708n4cwJs5
uaOgm/z2tH6faXe3v0vSw3Hm6brANDcLoMb/YwhhyMbiycW89pSsQ3wOmhllGiDwhjhMI+KATOHr
Zx9UImoYh0QakYYOd802C1Pm6a3alsCplrYrn/ULGs/+9mOU2wx18UwNYMPMXLn3vdC/NrPCguoq
SoDntz9wQs9PY7ZU0jDjaDvYzCVoC1pA+MefAGlozmEzsJSxAhzWunIR85TC8ZCgSlJJOgWVwLhQ
FahsE4QEi5/FGOuD4v5s/klCRXCc9NrpVLtx2y+0IQ73uXngUxIg6Lt8/lRq9fNO9TkUrk04a7qx
G4IPLmcLqEj+gHhgXzp6ESSJr8mwMr6NS3UpeoUT+gRv4Ve7SVOWu9DhXcFMG96cBwhQAWHA+n3C
8Nx+ZKguXLx4T+Z5PpJYlH9wGSjOYsc2eKrjevNyBi3xMtW4Gq3dkn1Pda5uAH0/77eU3L+to61J
I7Xk6RMd1/OswuMD8t1qSW7HT0LTrOO+KSRtCiKv3Vfoimv6ToraM+cu+jyBiUv1iJmSb2Bmdc36
euvegbFMgmLLbCy1YGYTWMEb8EToPlgOdg1GSlt3FigOrkifczNh+FnMhXP3hURTtpD9iURgN0AM
BlVUFZ3xzr56mCrOC/5oLokQwE6GpPDyNWdEX/v8NyHRKVUP8bB82N+3/EGRibu9I26GvPPGannr
f7TlE5tyPJyjGJtgEEJvD99F8IKzD3nIML2RxY4ncbx2dR75fnjeaUvVGa0RXdOjSGgG48ljl5VK
XEC9Xg2816oVRNMqlyXb/ZAufjglPfRXFG1H0P2+zhoVUBM/BkSDyFylcAB2cvUME7V2H+EaMswi
PZf0BRrhw4T882f0A/F7iasctf20kQWTZhEkMzR1tX7JE+rcj7w1iDxkunBZlk7NgTBNJ8Y9+vd5
TDJnA7vCGtwjhpCIIEJy4YuOrxVidExiUuf9xCj8v4faLdPJSqV+6CnmuAesb74RdWA38xgQMfku
WKjfkF6ozCgaCKIzf7QV+7mLDxVjuLcvM3q4rYr72EySjRLE8Dr4iyaJFDNk0/cm8EsjS33WUAqU
5FDLuVoiPfLpjQv6dhUZGp1sLg7T2u/xau3ngIJi7k1kBpVOYt1DaLba0AdtMcJD8JugmbqLc2zo
kkqyYfNoYbjZGt1C+l5Xhi5VCncAxohLTcFqJyeSdyWFI4u6LYqqNhXSb/hYAsoMAzeAANf/RGZr
nO3OlpO1yfL56Grs+b0Ewet9i4XrWMQeYiKiN/c6+RDgFsDayXJjrYxaq5VFquKh6vRtSpyfr+Vx
FYXcXTrmxtmSlUj2r+rVhfiCbiOO3Q0BaKblWowkPLLG4MefGTAPhB36g60E6nbBLoPMme0ni4y4
LT66EnAetKut07Qz42jjC7CSRoXmuBpvQFA0iRVQspxSCCkpaHCpXPhKrdjzX1qBEHZ/fknRGAgL
WQmcyZfzKtmkt2AvGdo/7JdUa0+t5SYoc8yO2ecB98JHKWlnKFXzp7HrjiOdz9fZ6zABMaIzt9fR
3op75xlOles1Y7YZyRvKbx6oKoU4vkUrskiWMi91ySBAEPLLpbmsldinnA7orrxSIeI+NCqMXTID
KEBlSrhWztfzomEx1wfpuGY5MoKLFV9LVg9Bk9nqrfc/2Q++dNu4nOPlJvIZ6aVbrEtOvOBVGEaO
C6VQLE00izfDHUCF1vYFPwcvVEK6mc7Iywu2I/6m7+g5SNdSUwJW31qHXkbR+vVHHe13/E+AH9LK
qeaRwInKTCVxCWg1rTxFkd2PuCSpV14iRg/Rg9pT7TnB47Lkl/IfptnS5vI0ynHpF27NyPMhu/uT
jflXf6VL3Leh+SgKUwxyMlBbLbG1KyzOEDa491Nwc+/n3DRudyOxc1CZQ2AksJ5xozHbRbcFmZnc
L58D6pr58GfHKcDTA9ZX0Hy5qBpOb/29K+ONtf9wXhWKT059ObQkKPTBe2Pb3PKqw7IO7zQJsda6
Nzf5iiaWKeMIdSbOyUM4TWDsU/EiOaC0C6VjfzNo1cx6Vm7JdB1lrzhN+Oyo+W4qRZ4dXuxu5TEQ
7i0tXd3t0m4oBmDvALeztY11sNdcgqGktoZyAMHdFlGwQmPQf9do0Sw27yfXCCHPfRhaQRqiRs4q
b90s1SgnwT86LUGxErWcdfP0oedWsVqG8I5xH14jgfKI/UWOFXIcjw8MTQuGazsajJwyfY6plnPB
gDWEETbKhfUBGNDRlZlJiN71hx2HAaVvvNwwkLuB5jWa0H7qS8MWe8J6vMeFT6cM8rqC5NeqFHLP
IbdxcVx5yTJZejnArMpEAZA8B0uNQKH7RLA7J2FRTc9CM+b9lTe2y1zRqV5fGxz2n2V8ri0eFcxt
VrCeXO1I/bf1O/zv43ZliGWOjtHc2lSlAafayHggficnHG179TJpg0REJ7+X44u2yRPm0bAMvBKP
g/voxdDyeDx40tpxzd3LRx04KDro3b2x/Qubs4m/Dh5NzuSCpX/HckYAEG1siMeWZCOnJQ18RSlT
47B4yQN/1U8g5aEOetRwbM3QudU2VU1E7IZ8uCt83Y23Hl0h1OlHiqWo6AbMhHvQBHoBPf/9W8sK
jej7rS0A2Z7nA3/bI8fIPggAvXd363eHS3688PArKFBcHu2MAiFMv3sre0ng/FykKJIU25kLbUgg
pkKi9lEwAYe9TEKztVr9BU+kUsZr7yWwpz6v574rkD85kps/zWeMNNg0DNWmKQegndzkitH/oUXn
DCDpCVmlE8pjT2jRORaJxMBQ9RSHis/sQiabWCmcJE+/2LNUHJ0eUtqz5RlF0hbQdgvPOwBMkH3V
Cl98s3/1fOzMGV181Hw4RGt8A2tgXKfSue8Z69pKVPxpArwsd34ZC1RkSNN5Qu23GnnWX498JXHt
lT56KfvJxOK8Z8kp6Rld1PlX+zCOKNTIg03mQWlcKRTlk/y39HI1Do6ze3zdBUYWtpuXYT+Kx1NK
MYVQQLysgOiPzOk0oQsw5w24TSouQYEfX8JJeXWbRbC/D38l1N2C5tf4tmufywEYfKxsihgWnD+d
FYQmtXku97u1PBAYqXWh9EGhoB1AaG7H/LlFaFsBS7DVjaw73Kvcri+2+Svw+FznwcQ0Ic4qJJqo
EGEVsgPO41cNaPLaaB/DV6oael8n0oF7FFpcoIPdEBmywjmPCcWVhnlM7pE1VOt+VETYcxkwjYXa
S/vxkWongt8oth7uXxUQONwMfkSG/voj9y4Sc1xQ7fbEPxg1/KghPCHU0OfIo9Yc0mIqw3hyYoth
AbYtyEm0hF3nMDX8mc2KSo5G31j9NaWQcRcKE+VihNroalEM23T2WlO2LWYv9T/rRrU2/QoIESPh
GF9V2FfR9LxLvxK5vd21dZPC00YGCvWbef2FfAJv8K7vsR3REft6cMFbqj140v4x31uqAbsOxdIS
WPg7pAHQwK3acrAkWfmbHTK5UV7xyfTrhj76QThAofYI8Ph/7n9DcbpFDjKyenmMu3O/KP5SXocv
Ry4Uhj7GWzRYLcvUb3DNb3Sby7iDTktCFQ8lNSc7wrh4e56l8QRvLDqyEDd8xh6QBNMH6c0zgB+5
NChkSgEvlhPbywByeb7vsq2CelbwpcRlfX3PwTgwaZ/D10so9Ddj0Al8gBIn56Lvb/Ni6rwyp4eo
B/F4smR3Jq3HHZ+jtO4s8KNbB/vpqJ8y5lwKJfIclu4eKm5IkJ8hhr/1RBeGJ5Yb10yH1C2p2LQq
yZ60aVOqg+F+lg2XsojFCY4EzATv5ixjoRVkk/FoFg83ACriqk+lNWB0K1w04alOn7gg/+VTOW7l
liMORzYamEfvQ+pi7VoM8wRL4WrSv9sQpZXzd0MerT1agH3cSSCjM7lwnPD3zrEbytI+IUHDxhPu
+LuJsvrN2feCMJDPKgy4AWgl2ytEbZJ/3JZzKZJHR6sDfKxwcDSSyKbTOJ1dRIHlzf9HmHSlb9TD
oxqIgzaF7xUF4V9pvyVG9sqeEIrHlwKe6kaGXIEGpD7Qe5/mMThYuMbWNM+mpDpIXgWvFxBOFFSR
B3O3w9k2q5jFE1Iai8eewyYcl1YqwhWz/WwUEDh/4CDc+XCBkjcArhB+M5GGmNQ7TXHv4W03YEyU
+Cr3e9fgBvWPj3YPv+iDRMKr4v2iKNNTDTz+93LHtOxQB7ffAhmSuFB5Qybspw5GdOwqcmrfn1UH
qPt0wyyOIAlX1XHsj+cSIGwEajLHOcGX1RHF16yl1RYQGXTaGzh5cjQ059iM39IYQSc9sJz0T5KC
WiLlBqVuerIiPfevm5C0bECdNHTmsPdDONRlnaUaXelh4ovF9btSp9ti8MY0FXYyaeQeC8B9CM/a
9DRDMpH4lLTHMSVr05NB/Lj7K1C/v6QHK8OwR/0OyhZ+7lvR+z0y/Ji/uSVOpr5uS2tt04ZnpxAo
hGQgHYT7QvUcXwxXq8NN6/2MkFJRAwsiMH9XaNTB7s5jO2jGkeJ1s3qg0/XyM6UBno/MuSc0SteR
8+Zfr0ls2jh7NHKh+VU+9kNWSxpYW/5mZs66Ha5uq03JSxRkaoSZiDuDnmh+r8WuUyEHC4xsKWMZ
xl16xBy3zrIUvW6FBd1Fmh9XDNn9dCpAZAsBrumI0kZmjw7r7BSSPvVjmDWQhtqf/SuNLVHSn1S4
dwPev44BLm12udEcFJE54pRZUfCrIYmUdGSynWIbS6lxiz+xY6fUGRsOd1fDVFQNXmG9eTIbAr3x
QVFjQ/Zzm+j7ugi7F+lD0EE5Hbh8mle2DCAdecqE+9rZ//9O8pZT+y1cwoxGP1VubzpCGTAmaO33
S2nFP4F7jaxZLjG17jaKQwfxi2i37RjYot9fOFRu0WGX9G2VZK11s0pbzHcUC/whELxnmAvinIxd
8VSLkuRWvmlcmAIWSSOweK2PnYAJ/pSeiC/acUDVIRpHduQNqgfso8d1UzFbRHfztbBYiqBiiuvt
aAL/p5kDyxz2BV9A18EehTa4r7njjzFvJaFUTacdWUzia/UZDFeF37bx/0aV1ES7YLvpRCENxlvL
Ggs1UQKsm3jFJVbyurAJ9pptvPPIkPPBn6WXvzpIkF6JLlqygph3Keb8R12X3q0+3//3RHdd91k6
u5juBpyvwrtDGNqT9ZFR8xNed26/kmeAq9c1gASCiOUviGSiJVl5kg1AQ2f56vJApUkpovSK8jb8
/nNLuEdjdPDONG3FEZ6NxFAYjo/RGQgeqS/PPx/XIaVXZOMgiN49upHIAMXdXKBh8mdbQyKIkVob
mZ+fi/5jTfDSmaVWKmiPie+ln4iDtRVfiqz2WAu6YQZNmSu9WFA6c8Yf4QpXN/obIvX0fkSAJtOn
VP+WAql/aoIy8XvT33Q+bhX0oZXT+W0wD1j5R6wkapWbxhNFNYnjEeI5UtJexKLO8+qMYK/rAWme
zW+M71LEB7N5P8LzUY1MZH+ZbQXnhAyBnnMAMT02urQq19k6RRzOPXg++U0UbsdBAkUtK1YXWEKb
BLvH4F9d/Ep/peGHISB9uZwvpGeQFXf55lF6DTzD+JpBQSOTgvoyKWA7NzwVSkZeSEruHNDAWhTM
Y/c07knTyrB+hJsHTYQtnHvdtfrVoP34aEYdAxXHh6kCu6YbHxhHk1nsZG5KS8H4SdfcHlg2m86x
WiglyowfFjl2jKSK8WosYsINPUsjR+adhaihLktl1ixWYe2Cw6gFpmqvS9UzhWFm8ePN7o+z7r2J
qis4Owrq1Pryu24fQEMWN41B0MBS4umy/0vzOy5yYuRKEaclTfhXINiwnak/brH16OqWtjTpbu0r
kuvsDF6Iav1kv7AAiA1lihr3v2ByK3aMr0VG9Ah/7QFr4/Lg0if6gCu7QBGfrbA5FeP5t4ZodQE8
OZMSYNoXv8M/pCyILuTzJu2s+v9DFtpoErj/KAxZGPvBGNtmrp/ETxzOvDY6t9Zsfn+zPxpZR3wY
2KhTTk+q8XsGGmLYInz9m060udPyJlVNef1Vlq9K+TieHb1dKjW+a9E5566o6IkCjC252tq+ZpwM
FqFNkMrk4P25oIQAZ7ExM6DJkPJROKnfwMskcj5MNV0/QwSfOctlPWg400NSx2mqAWELxxLZHadO
p+kB8tCpeCXwUcbHeFyGYFA95VlPXR5rcIbEQl4ockJD4GH/aUlYth5jFhPQHUJrIeumFLzJNhir
fCBdLATsJcJ9EyAHSv14hqcIKT6SBYy54Nx82pxS1KNxxMxI15mEVPtcFukw32Kg5xX+7tMvvqOd
vN1PgOh9lapl7W0DSm5YsHX5WQmGWHkEs459vmFkE6czkfxef2o17SR8uiNm80Dpp2LhU89CWnYj
gRp1IOW/nwUDS1GOWw/ufuHY+MGPGcBFxiCdv4RadVkG5SzILJ0Ouj8orqlL5c8fii7TR2E/m93D
RtLtIU/9u80e8fiDSz1XBcleMDbxLydZT0e/2u/45aCpFKaONlPifuqGJ8VxBZnD20P1pmGCpr3z
HcwmHhMVyQ+HnKpuamgKH5dn8a6l7x7IFV7zOX50WxyWg7DA/MGwngycQBSzYwj2GVuTploqz9tb
OMjuq83TIMRQvGg+BkjcK5bXaUlIuGwE9D1IzmLaLnE9voBtGWSj0xK01R6fPpqWMmevhI5dnwbg
3+XZ6bKdptt85axnRYM1IXKPh4Lmh76Fo7/GqrTRLjd0Y5/zEhOoAlV4pD1lHSKMH4LFZyF5vuDF
6qlFKSAocG0jFYibPtX39IGWjdPlQ3wd0PtHAlX3i4tlE4PV9EmITCvvJaQ8Zbd4qQsuAOEJZFr8
SEhlZnc8lIesYHaYUkKk8UeZ8msJmaHYMiy8lm2eH1c+XP8DYG+rXQVU2/obyUwKI3Ajl8tRLc++
SIApOk9fKmSQ1y8vcg26HxtuDOUnlhU00fY8TThF9dT2owYCRnw5KME9oQrEKr6AATUcDONWKXHh
WFVMZMk/6XrsL2tpjPFMR+q6ZDa8PQaNo/zQyc0G5/ZHJETtgoS2UTsXek23hh7V8Z7E7GwPprUS
fXYUklTOFeSPloLyz6XiaUNcUscvhcgIOmB/0TSNJR7FlrZADXaE4RrWQhNWHOQxKyWPHoLs9x24
LlvkufUk0qCVQfZYRg4diZh9eUvvNWR6sH2uVHB3aP2FJOZ7v5rJlS2xXjcqy56Shr/mND+/zpSb
lOVSIWdet44J2wRGbChIdW/m//zNoMgZErEmJEDuQiFsd5DjXVFOpIVMKgCNyZHb1leLg4aUv1jB
FX31KhavHNTv7q3O9FwVAd32S00Wbjw9baqKkkVnK/2QwT7cYyPNCZ3qxekfHyuNt65d0Rrmklcg
Vmv2/Xtp43WKYD7zPzMWPwcXrXpprDklAHxIdXtGc/wVigqoUVihnLd1zS7dWPRYIq3stiHRTIsF
vaQU2mFoJEsKzmK7PQ/UKJwwFgs4BHlNyIcrZqWTELGqUl4ZKWAuX45ICgI+E94opdKfLFP3iDol
HKh95hH+X52e0bhvij/yAF/t6ldVFvt0O1W+4Z5xMDT+JY8gmPEKD7emPNu2FVGWFUOnutjmOtv1
K8bvXSrcbB1jmXbMe4+faeDaj4z1bdTK5eB3ThxaC1TImjSjWpoGjTZdIcL8ptvBLqSy03o/XOCe
qPRVRjLWPx79mL3S7oZWQEN6qhMIIGudEZ55qqmp6ClQhLdx4ZzVA1LelJ+mgstfCzP2dYftWEDG
vGYoAbAqyuyAHiooKUwKf4DZmN15McIsRzeZ12mHYOTqCGgMYNMCjVBGwyvvmWgDTF0MmsCX4YhX
VW9gw9f43ueInm9yE9fDvlH8m/xMsyZ1OH8ZIAcgkLCLxHi3TW+F3/Ahh7WW+1NRBJMO3goO/J6w
avnm/EnabptZDO4aTp1+jK6umP7l4h7rG1WaVBNhXK596BQUa0VXjACWN2AJZSunYOvnY1R0BXF2
GR70eCYkZACnYDguSzDCWzQlhowmd0GT5GeGdZji2+cy4D6d+XjLGvp/wJbE/rbhD1eKmXO/rtqC
VlReo/eD0zqD9p/gFxkvLaPnweXdYP1WZ0ARyrSZZuY+A2sjT9X5gj0+SfrWxO5yMsG97zT3Sk1r
IXvlq2Y5R2qrQi0HM7lRj/KpHj0sPkMCWFfKmUg2ZZao0wZ3sI0U7ryvU/pOf8ssxm9IzkCQC6Im
nFDatbZXI0OrTlaRugbxBwrOB7vICxmKSgtgAlp8XqOGVxtzAmxkVN6wRrN2H0g6tV08CS/JiU3s
7r2SWRiE83dNU2YdPpGUNrHzOg3t5kTrryaqKL3seyFHzy4P8K0yOqzW3W3o1ictipnR6ZqdaTtl
nsWkCMy8nr8ILYXjQOOBNw1DtuhqlPqMak/8LX028Dz7SHsDjvlj1U9uVp9P1fhvbyImrRjqnu4J
nyd3OoNKr+jeGR0mKGGd3o21ZvjCq3jv11pcbzPZCsBbxDlHm7Auf8B7Gr94mjyzfJ7FjbzsyH3D
WdyD6r8X3bH654xOYK83MYOnmJogUKJNN5NsbdfNQvoUUpp3wP96qE82Oghq77NYu23mgfuZhPks
UgDn+ZpZ57cr0kiwNoQFMcWy5wQNIPHKQlpHcF19l9mf36dZC2BDoGF7WhbSTdpCQwufKFy+ghzv
uw3NmaDfR5p722rptk2JT6vFGVHEzOUhanNEqzCnxGQxcfcQuOW7grU3jKzKDkG4ns4QLDgrhE9/
Ro2zS2qoPJBqudMoYtaQ/nFP4FUNYxwkab9fxGCQTs2HhjALw0QiNUBvVAKIZohWsPMMmLehGJIO
WcI0yDiJglIRk6xS6FdRdoU9YhO86inF3clsUYF8k/n9vf6MP/KcufuUj+7NEeiYuG2xRotNpOap
cQFQ+bkiQVRtWOzLMUbHWdmrNPlhDrEh+Je5+1NJlsWbD9isUO44RAfxe7DhA0T3Ii1kQ6OCQeoC
+DEXpWu+zYnsgc0HObCrCDr33JsOnvrk3H74x7OyV5nD7bHfSotQ7JaBTnBhnmm75AYCRRINzyKD
ejlV6DtbaVGtxff1DVL1lptbE8mEv7lT7kbBghyj8s8Qd+6hki/dxALxJyPSK08N8N/IqfzYcRvW
waAIBt31gqPrExR0GaI/kJEzlfV/vYEu+fAKriOE3q+mJ45zzLqeIirllwwImxMgIs8tk2gIrkg0
RagSKDUDdlZBuCGJGGUPPnfjhoZo4f7vP7bL9zLDY9/it3lpWVxOVeLXW+/SpF0pMBeqAJskEb5o
GmcTM4SDsFny1znaLEFpC3gssFu5Vj29QGdhHU8cAe6LZgy7orUBFB+FdT3jEbjV4NGhqrmRV3XV
NZQ622tlwT3/FC8WXqTJRNk4Cqk7uwZyx32HcBKT++5MqMwEz9YCslIFx9CqvOzktZ9hzi94QdWG
J5/60H7fmCz1BoCFO5jV/HGCPqfa02hAMwxSEblGKOuGWlW1QOqmbbPONb/v+Dw8i1fJ7mp09yXk
DZ+/EFOnAO5vkNRolk3efGn+V0aIeh3zpaS2q9MhJ7hHUjG79TEjBURqBQyio4SxD+w+HWMyCV/G
Mv7JlyTkydpxLZ7hXvGafZixQArlNLDwnheJH6yMPNas4Ddzn0MRMIPoUBBSa5tnU6D3IAAEeskR
YXr//UkhWrebscLRZXVq4HCjSK542CPmokfsB3Jh/xdZqy+IJv4loWp6Lhi0buVleTPOJSA3ESMd
cVSkTMQCdsyCuMeJHwbq0fEqVbnL3xNYFOL7IbikOEGRAykF8tg11MqX8rxQRCGjoXI4LXzKzk4d
lR5k/mXV/xJzhzgWYxAovtaZ+xpuLnOuY5qLNSWEYgH2iHr3zlOi4jx+wMeGuOZOU0P+PfRulR5D
mg3MPxDKARFo3qwogPhk3djIdVkhTQSGkl4Bq8PyEVugABo2Xch+yHkVMOpX7AVMHId9n3oBTljK
Ct5YJjpXNB+hLcoBD8dCG1Yy+l7tXydfAE3ncdU4YD2YrVB3IDs/xxJo4cGJoZvrCA+3aHujm/zj
kQLCt4b7ZLuoeUvvDK9t55BfCzTNg7O/9YpGO23t3xM6YxoxMK1JXtS8LBimegm7zye9TohskHSX
mMA+dB2Ho7//VSFBwKtqd9pakw3MXwMqU+e+0VJKKOAE+VQ7CAnAVrOXZCVJFTeBGZyFZvxsckGz
euaTossXZRPK0rWmvRpxaTAVcjEINP8cew0G9OFVNhS9/vKxSEhqfsvtL5eSStum0Synudi54XPq
+OWcU9Tfrm9K0ligRDoxEGV3y5HyZ3bN/BetZelsW55ardC7hbI/xTf6Aoy61alkbb4FZRiZdfbL
7kfqD99yOOfSE7chPxHZgZPn93i+3dv2qcX2N64m2OZ/369bgbOWGHFW12Ie8EjnrAWxi0NFk1UU
rQBhRL1grYQKRsfKStuwOKHTwX0pmMAdnQF+2XyMFohjJ1dKHX0WX4HQGBJumQeHp44E9y+UwLtc
PyafyJBEMwfNdpaQwM+/UdJmHN/zsm3UDvB5HJWKjwedK0nRWXNN+vwdW4U2gFJsjhi9Y9W8yiZe
WrVb9s28G9ZD1hP0x9kVna4Pv9G3AVYUN0jOADUX/Qz9V7fdrfh6+dAYM1FdtcEjvJQhqJ/j2Y87
uibWerZ6YIUeSL+hhZSj5mam/PI1F2mexBPlp3oomymL/PKAyDfCaqKITyirfQ7JNjtjL2BhKpDA
kix+itqwUdfJOKsRhRQQauLgzPHrEZHi+nuoK1qr4zR8UTYi+zLjEo8FAezvyjOvY7uCP43pbefP
ufo66nLGp0HwY0alLIZ+9Unbw9ofrjjHQhGUGL8BqxWWGZCW442TVgj1czoPTUw3gtln6P0iA70M
JIzrvebIfbggweSZTknItp4v3wWpe8akYIoDPe2rHSVOck5l+jpmr/tJ3N+DXuoCLTEcw/syvzSU
gLfvZC7YN1M2E4Fv/lLEovJhNrBsJ87WkLJ7LnWdOREkmLTnq5Jl/aFyEbx2IhUUkFpLjEHJWWi8
T2iMTRY9fv6XX1W1cF97YxQY1RQcHnEqW+8E9PdKSU0BV1Bk6byN2BlXBKgyBohdxHoLg2Fe49RM
BVDpKTSHKjT1dx4DaIfsRBOQdqbHXcHfMLCHrg5XBuHLVk3COq0b+7ApHaw90ZzioWxC5rCzfM9F
ShI5t5aVC1kC5Q6Y+prjduALtGdcBqYLTldnKSHtfOmsVKilxO6lhgz5N9J+JAHInT7RpOd8bUoh
HizYdQOV/pXTuF8d5LBFmni4YI6hobDqarkzF775zFbjL1suANsYR3hwWNemrLxGook8/F7TijvR
X3yyER0+gc0CQUK1oEzdPNdo4U1aI8iUbjj+qET7JkBCISz6yxhpwEpB/PTYp+4YsDh8p8WA6WzQ
HUZEf9vly/dxJ6KF2UVAPlYwgy2KrIReRDSDzsqUWzYo+ZDpbqLct4z2mAlMrzMDZeFtcYMZ4n+2
zWDuYXmvJLNMAk98uWFi2JMu02B5SC4XpgTd3lKHPg9sxgH06zks3yyYO6GM8CS+k8dRGnjN/KOV
d0DPEwQ7kmCgbUP/pKu/+D2nY4sD0qPGk7oArpdlZzjX7iYblMfOhYzebZy1EG32XhkTJR2pqA0V
vX9fVOBDP8DiTOnPZDO2yOEXadE4lhB7OdqfHiTcld2sPIjlZyCCVr/a2Dk+cY3AbjVwPQ13NTVQ
hogPtFVOFlZDZH33CQBqKWN3a4XM9eeiuytlvFGXD/tNY7dxTmuxohLADRLSMZdWA/cmiHXXwd1C
on2TZZ7my7TrLjIJmHaq8i6zr44DE5VR0fT8DXEGhRYcGnVcBgNs9IvQ/X3O0THnA2xMJXP3EZAu
ey1A3S7DH/eiBf1RNwIOLOApduKkKsnFeNkIHMsnRyYYbhWmAjUbGEIFChaZ0WCocNaLwMqrTGKx
bRytDdy4zVWksCF4pXSLvFoVvQXIetmNr7JC7RQNbfXIZztnizOQF6cFsrLUPdKuTHgTwXmurux6
MgLgSL2l4GH210e4ChxDrXNTu8VhDQYYMmKIJKwv6uHvSarFTq5jV23fgkYGqn8/0/0EIzKxrilE
bM+lA1F132AtXKtMRx7GadpvfgrH/3dCalo05jwQnbMgcPgoUblWGyPEeLGl6SJaRyBw86X6WOVz
KYDDtQL1eQY09zaj/XpbF25iQDU/RRn0B8/IaLhbnnE3ZnBUTNqQfHoONLs7NvkznJ42uHZJFRqJ
jf2NVdDKzfMeOM3fbz4J2duyaSYi34bLN2E+8sPpmTOG02PX+E7BJfyJE9f6zeBWlNb0Zy3zTb77
PPMtRBEYibKFO+o1r2PkYhmLIa7/ezT2L9uLx/dSQ73XsrkdOge1G8EyQq+AIiBQJkjjCZYdTgnx
mK1xTLNbSNFhr3Z4WhwEoyLjRIZW92dg41V8HTfBpNHZ68JgTFBEVuJVJltaSqu8B+9HUZEPPIhg
CQLN4ePQTdelLkftJ9G3c09547T+ByEQET3Gllc2l6g0BJkaXLWTsqIc/gAdNfolerOZ8xxZU6sg
ixOBeMdu9ltYJ3DnFuWs6xK3s9tNiZdba481XvQFcIe8sG6wEw4bU1IGF+/G1G0OAwJWbBsH/qpD
BLvskbAVDV3rF/GcqWmKo78kbhwWHvNuHelXWIjrDwhMi39FXw5tbTGhegfRqxrU/is84rOcnP6c
Z7SCNctBz4E6VVr704wU9ZF1lYwZEg4/q/qs2tj/sZlp+iu9ePPg8xEWcFwrXWhy1QmtO7Wv9d8t
WP1WaThOfhurlo8K4boC8XzH9Nhtqk/YdTuAjB35gKQJeDtQKrVyf0IttQwSayBQNWNoEuCweVKW
Ug8FewR9NVMoJ7Q12MhczCtvvYVV4v+WoNhe2ubZ+/YF2SOb185oL/y2hV/VpXnkCUmbNn1PCFFU
x5XI/QouZGOMBuM/ojF7j+JM/daNT6gXUdKI0aQ2DnRQC2gvt/JozNyt2+8HubIkxVS3uyFFHz/+
7DhT2lqm7n24E8YHtSgczeQE8J2oNh7il8ZKVLr2EF8mYk3FsV9QvWMNAqVFHxW0fhqTVHtodvRQ
cAC1cbanvFW48+DIUu+2Y8L1O94OG7GJwtV6h5xoBq+8W0CImtTFZRa/ejJpjXNGzBlaF5HJTcqR
s1K1vtEAlqYb7tmweSzjo71BCcdI6TbjfiqQEgmZZFZA+STHHrDdqDp+ovNkOj/VOrjeV32COtth
9OEKeXuLJH20F+2rarzxC0dqs23AU8X06gAq9f8K5poN2y/9NISlkhJG4/ZKiglwVuQJ2CwIadi/
ijf4+GV6uaQVmItgd4Ggxy2qKZdevYsL+cQY9u7uUGidCPizVM1YYmmh/spRv6XBlmBCDBsBGife
F1ahnudYo6WKuud6J5uMwwidLhIEwIy/hcPQZKvsYB76+7Ma8ZVSYR3uvr1bcBgdmI3gKIs5q9jJ
dDvYWy3uUiWT8cpZmJKSvJilovxdLTnG4afdQpvVyuZNSigy0TNRAmNcR6Eo8vwqtwwg9U7ORfLy
9ly+JSUkLvp8mMVRqgTafjGdUc110YtnpSkPThqoZDxQSMZ2E3UFFDfXaS4sgKndcGJlzaukancA
9cyeWk/4HseZ5c8fuB4XRaodCC23tAwHvvO4GEnoFfHqu5Wc/mVK2QTsRpwciVOsZtYejkcYh4Wl
otf9xO7a0+rWaW0alJg51SKLrA5PJmIlqznNmzSCWMtao5tPk9HqdJQdmW1HJ0MGzWmjlM9YMrVP
o0WbWDx6QTq9m1DNmsGtKs6qoUdzrBpL/XwsUjJ9xjGeY5j7+AAK9FInK9M7DC5rQGqQwbGuW9xD
RwZQ2FstWzHI6+Y6MTHbFncaoT1rnpv6HSbWOf1fpFXcFT+E5y2f0XWxyd7tEjBYosJIC24N8M0a
CmnqnMZbnCBf0QqACBQp0FgS1Q5HyEBrUVE9F5TFXae6SHR1ootNp5rkQAp0fc1Ixen5JC/KmACs
s9u1yaXNbH9b53Ru4MWEvCJkzedywrg3AxOrUPP9WHlqSt0vYnld/W9fos0PEFg+mH3PRNYQDDvi
JInAK5ijZvmA5CvRw98V1eI7UU0OcZ8P8qbKZ3zv8+AfdOVcjNUzVwyqJa7ef1BPMrtMoLk7/jom
RvToUz6nA51mMStFqgvWLQLv0nWfS/YWMJVyYZ8+vXPB+WhMQRB60G1bq/NFTntHgQXOAPv3EM+x
XBwdI+p2mHZXOiDFdWrnmhWZYaaTiGFqYUY8+RL41egHGvr1aA/wvi9gtKu6d1EL43UygW+O0uCa
gXeg6z+LqFNlij1ZQ9M60zjL0449eJLaf3dWE653v2SqkiGmAmJBHHSfmeEFXdDxNuUkbnoWZArq
Y1+snK/JVmm52SnoC//KZgUWDZyOcvzWwluQA4gcFlZOEksY9J91fttsJ5n+Rdi9NeNIUp8BIBpM
xqEx7PQXuawRyxMtmj1F382YXJx1gER7ZwXluQuxwBWDVAdBFx3s7Wm8hhOU1XtmTaD7TbfUhjNB
lEq9Uje13UlNqVE98tfya3aIEfwMnVAdkBENVlNkU7mC4tfUVv6gP2OvEbWpLcGXesriBhr1fwFc
oNw2vvP/Izf2tu3+JKPK1J43rzYRMyiW0I9kyyJj/DDchOCaaGbMxLx9lMB8bwtd8bBp7PU6nQkq
tSenygis2SHH+5kPGRuw4ixKPX3gUkd1btUis5/mAS0wb8NfJC2NJYA2WD3dyjqDSU3RaRTcoXIg
snCircPnkeC2VHgvYlFRQRFayb1lKaVnQnjeLjdBReuaeCqz/igeddjtB+f0D7pbBu7Hdm/o0ncN
VclLsdZM2Qt0ONLYRYZxNWiGMJK1qnaJkgSJ/JsbllS1fq0wdXh7glJc0uNs5EGGamSYxpuoMc/R
9nyuzP9kXnsMHzKOeNF8FCNwdp/wxpQGgoibgxV9pP0VAMLHuWBtH9uyj5+cSnBtl1dYe7uGGYCc
u8w+xvL7QDeXt2BMUV4hpzZoRg5/Jo0GGXfsul8LyZrrYnFROy78LWLS+mZOu2x3EHPmEuIOV7Mp
FS+pPKtKwuYEziRkTzfHmaZ/wxR+tBVu2M4l00owZxHbX5tqvSjmKvlrgwD8jVgLXjNBCoy38XXa
GinM46xqiIPCE2cKkk3tKX9D//SipRHNwt3DbGMtgriCaX6/YzFq/2QSWQeaok1puzQ4/OnC2SlC
tEjABGYOZ7EHZ3XzDDnQ/+DeYgtfy6ncdELg79kfwSnSC7joHplEpyRGl7/NfkvyiMmpVb/ZlIWM
56HoBxxjYcSa6eEBKRmRB4WxHEmCwTQbBrteZnbc91stEjpzwei6fAsAsEzsUntmtNdnUW51YgAF
QvjdPru+FYJrg/pFgoTWAALGH+rPsE8pNphjR9hFXqS0h4LgviMrycIuDDa42MapQ9jEXZn9ZxqE
Wa0F4U9+N/oAFQV5yAQ1sWQJDGKNwdtNN0viYdHgOdKK3fwLfiLJXu4v16cFsX82KGUwn+M+Xfav
icW4f12hpLgnt91ofUslFnstsPP81zr2LkHQwitbz41hvvVTUVzaRMPwGWmSuiLgWTv1VjImKjl4
k47SJQw/o9Gf2EZis1m8KI7ZdiWihL+Z6gh6rTfyXwAYDhRPAxiOcR7Fq0LeHmEOEw5AqXJPIHK9
T5wmM1JsR+jZXMEoXLIYeo1yHIRywOxkzuRGexVpRSSzVS/jVwO6lpxt81Q6wvKCtOnsKgi6IY1x
Fbqu3cF4fzg6RZZOfVDlSNb5Yi8m1n+VS7GUWJ0Yi2cNeWqkALyMqgTHnE/fJPxHEjY2abBW0WSo
wSXMdaOxoptJzUOFY1hiZNlpdnir3KUc8NpfIHGQWruLcke9Dfg+PNeO/M2CN/PtLU1ICTu0gZxg
K+XKsuwL9txRvKTdOKbErb9OVu8Cr4wJuZMTZToxQ56XL5nGKjf6FXjPvrRKMqS+41NGfbr2hfBI
oay9u2/djUVrGuXCIBtHgFSfXx8qkPgNl9kVyFKZE5//ExImIBc395ZKd369IoSVYOkl6u1CCJhd
YfPxFqtWZrkAo9xTRen7nGthJfsO+yKqaULw+R+rd7q4RDxHJQibcvdExkkiXykn+WylCkkRR8Jq
4fJknIoTLOtg3g+pAd2hvR1UBQpRsQnoG7qdZqd2g6wCfSOFfiqsKU7sCanfjQEK8hIVLq6+wwkU
AtNyCzeHw3XLL+pD+3uXitj9W8Epwpt3dmVS4TZA4KObWlJAg82370bcDfvZ2oD45UFacoTjv6nP
UHTqX+02iAddTN9oUeii6dJ8GDD3TxSm+UZ4cYclaSczyLNy/DAOkmC/eYJ3ZNEbj55uvQNEqpJq
fnbilynxYcfjw8n4501w9+PbLht7Qeft0UJ/2YERSQPnjhHCF28AXrGjRKLjcZN7EywUA+fOtFOI
LWFrdZSfYK8NseWC0jq3nIabUdv4XfOx/hA+e6H084i7J2qhrd0RCzeu5hSLTEf3tP/qTVrSdY58
yqIqcmFh6tGDFpCxWtODg9LzTe8HoAPvZ/ewx7s9KA9vB+Gwcv9b/U4OUPCioFoizPscx5oxj4Z8
7O1p7cgCWjX97fiZzKxJsswYWmOlRUiyVGYtVyW/rxfhKBZj2rwEJ7QsazEQv+NY8SkEIXbPgu7z
K17a4SS141TQgDHtfNXivW+/s3mXQfESHG0sP87ake5q2wp631t6BySymwYf81f0A+XLw60qRoy4
V/kyeQGvK/1YkYY5RaeiflqUdISjjJ2uNGx2DB+O8IUiS+fIeuXZ2/ZDjYfMND8LoekllWMoMBrt
tSazCSl7VXa6RkEthxTfuHJ07+kqgMDls6gzno199CRS0yk/KJ7XCI4tUiwaqQj/7hAROjc2GnHJ
iiBVL0E5GeQk7820F9yhfqFaC7M2fW31unQe1U7CJ8lxlwUFSys4M5uAoyl4d/SSEgjAFtWemffF
CRVf/l72ADPJiHqijPcwMXD/BRNGHECu73SXPp9dgm5/zyah/+fA+DxNQ94Dl6n82mUmCwX1qyol
cG5gZ48TLj9pUKgbKWjlFnN3IQc/oYazsHCgIHfx1a2ScUUXMXVsd9nVH0fafKZ2EyozdM4xQf4x
eOEMRc9mu9OMUMSrsj5+rDO+0aGttJha73SE1/obBq1Hp1cVq55Aj71FmlaCIPoz/BtexQ2SCKjh
1cxDa9F6pdpl5DZn+LYybYS2SSIN5ZxZfVZ4ZPNA9UdcYSipb3TC5CHN9wiIa/aqfIEEOo0kGb8F
pIUisLnUAcO15Z06cInaza05mTZwVbCGd6YUpzuGXBrzlkKnIRXosRcUkofLAozKzankLfYudEqj
uPbYINkP1WtxIy89z4eHFAUWX47i29hIpxuTZ2i4XBq4FUlYkJ0tEpg/syghyqjVVIIS6HTbWkdd
hWmdQCFaYU58RDCCCw3NLODCaJgzeMvEPeKA/DPD0A4zVLnwpvdD81yJMOfqN3gihcGCopmR9G/1
GzJ7IvP9UZeWKnly5+maHRkWM4Fm0Zu3+kMkTqiZQnVi2LzyEFpZasnjREdNhUlGHjzPKzN9KNiF
BvY2SHx44wlntlAYvuGgQNPte6b5et55QFBeDXESKso/B8pWdDeW6l6ZnpL0T2iI5MZ3IRqJLChD
8Zvv3e/BC6fBb9NF/YhP954qBKWdnUVTQwKfqH8sCgIuO2RgTat3hrhMOTkOXoIkdKp7Ri3YwBB9
epUVoA2a4+JywIfx3fsCWb7E4oOI4OhuyYKhNLNSfUr5YKEuxq5FWsIcYMRTZL3EsOrTRYqUkpKx
ZwE08jECv7qh5QFeMeEJfHxfS1/PhLZbGtjOOgl67vsEVQvZubR+ZfBfcbKfYk778La29T0TGh7r
OMJ+BQTIdWnapqcBBP7Z/NlxJIQb4NuT444QVjv4WNKael4ugI/Z7Mlwoa1rSZLin5igOMIE2X9q
TGhfGU6UU9rx+gbkVJ5Gt13wJ5QCfYw8Ckxbe/G4pEflRxNetLHVBKZaB4lSeC/AERLHIollzVs2
hy1kahA/gZdW+fpstXGLzqxcz6twWXhBz7BcNjYcCQnyND08pd2er023XLjLaTgEBGpA++PNcfQ9
DC5priSwdwVUy0fbjvslq6akztLIBgAQDpUaH4/6auLVrqtOe6VRi22XksNCNQf4B30qH7WnioXO
c00YkrewAl7xXYYgv5cL3WPYtFmyt0WBzDHp68UV79HSPlG7qba6fpwR9HaP7j2kDIbj7nymQjQh
02arHZ8msyrBSlFBGvJSJbBx0GnyzjFSx3dEXegmYfClSj8ndSSG2Z3soHMGg0pREHkQuXCb+Fl/
D0OIW4G/47wyDh+awzkaabveoA+lx2xFng9LunNwpq/t+Uujii6hCXXnxsbsb2HRfE2igMtm6t8N
iQdyBv40msA6I5RL6HXiQVfYYVqwLqQMdYyxiB2WzHZbS1gyCfPbwisbPCW/2aQNIcMb9uaetX09
I81wLoZ0EbPri5BRl3i02tQ4KjhiJ4PVP0b/kQX7ngkZdkX/f+NA75FaxUOvYvHyx0Dm/G/i8SON
m+dhSRATWjoJS2XarOJCqEKsSbHVQFDm3/gTPVDGYcfoPWLfAHbuOb15svMwHqLciGUtrCtCplFt
kaCVdFCli+NKW1oCKn7YKX7xUPmnIALKI3t57KORT2bp1GsTYVtPwierdACq1mfMCchWqXZsGUV+
MqoXQYL9I6iZeKDBfesYQRbZDxnJqyJF1VPwdWtedV7NHHddG4YAKwsjHoGw/RI+3AV9tCHrwl1D
G9c/aWqaPcPPUiGJT9F8RZx/pDl17c5l7QtKGMlUn7kdBqoMkW9ijm+iVDA7QMvoyJwf0Y9X3PxF
YfPeV9PmQD4XZwEJLw/1zb3flpx10NLLOLK+dNXOhYHvuYChxBFPJxnGedxuhg/utGxNxgYMrXlo
9Tvma2KnsqNXD2T42KhqI4d1c03ysUBoIMAT2MgmlzGi7uFHJC1UIHqD2ja8uwpmw7hsfTmXxLeK
R/0139Op65oAC2dbmjbsgvpWq2U2g55I+s80AKFutS3ys8f7rxMIz6dTgrPcKiDB82z2MfNsPR1m
0eASkS96Tj+WWqp2fyNjM3msrhlSIVpodnqcIumbk6FkUytgKqCMv1K6HrScyXaFemPj85rTM8fZ
iiH4TelUf0vd5M7BXinPtN92T8sUH1wSJ2qpC5VKxzCOwPPRaVcsen/9qRLz1lRmDC3Fx+45wGb1
Lc2auOdg5GHd6NmFVkSn8WMQSoY5dRSrL4mBjkjAionP0WiZJvZ8qprK2BXSylunFe4qv9/KVow7
br2/uppTV21zkucuPMPYc4OPZziJPmvtfgkZBjLWvYJeb9RzzC/wHnV+OcKX7rD3pI7qC6arOSLd
wW3EKb32QkWOpgQoYM2wUhNsE59zlYrvc7vUdKzWwZKXPsGzO1QxZR1gZBm0RYPsCm5ZJXyjqPPG
vB0t5vK4AbjFnjWvIcOLqZAEPiFVJ4l13eN0B+qqn8xK2yrY9cqZtGqG3kcyzW806t69bAy08tTM
2IQBzmx9ySX541Pmb0wuiLFoSLkGmVqc5++jUIgHhp1lw+QIFkOB36ySCRWQs6Di4gqkdIO8Bidh
jfa8aAqzFpjCtVUIWngwCG8n9lk5PQdN2J6FZdeqEuJI4vLGa13yVqjSp96+tpzGf3JXP8S1Yh9c
ETg5LSYYjzSWIdhdu45UDZNl2KEWnX2Y9XJpJ7MN0vw0xRJTGntvjP80Kza68HlDT8FHRtG2opJT
8KVl/0MJO/AoRkV2y+AsRvCXXNYrTWxwgVC+Fe/ef7/DW+8rqArph5gjxyP+8UOnRFdPaWCvxwxk
foIsogoNlBnybzWPOZcP5tX+ipkRRhxxH0eJuEQUixOkaTwm+EUuuuObvmddw1Nr8gWva0XFZMkN
QjAvphkPzmGPK3JIY4F73vC8fX33onf5ncPgVU5ju149o1I735pYaqXyQYHuJBZv1bINw0eDGeVy
ztSAqUXCEH73gZnMdHhYJPivRwrb3y1QlhYYohkG+ZisreOEqs1eAje4m6oV5K15rTmg2DcJle/V
gJch/Rsv887yKPJf9DlhUxb7A7DAZ+HPyzUMmurPXVUOVbuYwih5toKvhAKWrUdoZzWgA++KsrTz
H/wwJ1gs8+BkJTX+OoAGOA3A8HvYMG71LCJH7wrQ1/3PJmco3rYyuR/+RXhbrLXVab4KB+fkv8FC
yjp7R49uuhmsllSozEo8bFH4eqDUAS9LVHfrqvdWb8CYNY85DqO4jSmec8wMKxHdRCFkZ+38SG3D
P56nAc/hCE1gMLPrphhfkeT5LqVpzbs9aPzhPtgMdplKSThj+YFgKcZN7yuDbwl9jW2wsWuqq55z
kAa65IG0BDZGJ1JFBH7RxUK4nQQal5zpYDvNu4XSMgDQTtm9tf9wdY05Bj+8HT3nx/53d/jN6EN2
SiADvfeQxFv/psuYzTj3EuMQ3ms1tQ4a7aHPKk3mZA3N2pMFjvoK7PTSKlYTNnJJKMxOWED8TC36
9A2GSt908t6wswVltr60JRb3iaGvP53D5FIuW9uSlwRTlaQx8UQt15vzBx4RcE5wcY+zDFB/NzkH
jiUpb6vWBuWAW+6PUoIkdoeidqicJ90HIGLOVrj3MAgMib884nYCzKytIYQuEIsh0NNF6uuJhoEH
b7WLz58FpN4B0teb0eFU6dCjASZmncwzrIYnGmipHQKzDy2Yw4OYfcKUSr+mvdFsCIDxB6ApB0Pq
lzzzPo9gH0ooJVVSnmjYGi8vuyeO51BMdeBhwf8xfG2p8R68sys+xVzwoIU80fVwXCzc/wIi9xVP
wrlG+zuOGkVMcE5+z4454bVcpn8WKveQnMiqYQnYAh/ViU6mRyPniWy14wVnq17F35AmEprcFZa3
M3xmCTwZ2g+PB7LLx6rM6sdVfZR3j17sYQ/uUBV+DfVbn+JfwgYgX5Fs59t9kV6i7cnncT43fCrm
QvFSyUk5ugaTkwyzm44xDzTzXnxx214yLSrN5TVE4oxTnRUXZ33g88HGaELpL+0dv/hbwzOW8ybW
eSg2vKvmzcnO4lGlhcuIEYN9ZfLcY5N/pSe5a1YVVWI+fHAXBssKfrUsPFYnGr7uVdvr3tIll9FD
A5cnh8TuxEIPjSGxa7VP4Pwcujhl2hb3jW4vD1t7FRq45AGZDqCfX/nDoxkjdSgt8aF96B+G4+M0
Bm9cEes/Ze6BphtlN7XsP3Wcdm6YmlJmPrwP73cjefzU24BlXmqFRLIRhGiI0FAKxpn1Hv654rzC
bqFHdldDkQmQxs16jFGROATple1gua4HWELAFbatGJ6u7mnZOVIUm3NKgF3f0vklwjDmC3Jftmjp
KK1NUXaYYMGwrAYV9hN+wEIOQA342yZCylDjZeQ0qljKCcRkPiDyYqF3VP8i96h2SE91tlTaQUxR
HKH7/6kIUvPJ6G95WFPolZZ4G6wRno0wPCMi2aSk2LKfrIW4bTPucEFdbjXD9I0MwzKnmx7CCjbw
IoQdQtMIRbxzlX4Qxhc0wiAHKrVRauLSiA8x9tWIa4VcJlKlGOHxDVLk/D9+U+6tRO9+SdC3AAXk
lTJqlAKEiNQm+T4V/xUIJd7bdiCmBvTHg5WhQjc3vY5Nr96DTWkLS04qJF//G87DrE9zzFzR7n2g
4XmqBuPg/RLc5geHaAQNgAF5hUqhXyvo2nwBjf9Z+9I/D6bT0Kk64LditSoWsFKra7/poWrlSV0z
jBotsZYV1wWfjlI7TZNOxPvxvmaeKcSqhWHnaxKBHMBIVushJ6+ee/6HDzoNHjrZb6GgUuRD51Ay
x09hqConuP1G+ta51Tqtf2MM6b/wNzmug7XfmOAJrOHkaQdk7LWgK98B59/TyGQJ6BzgltA6y8Ao
uFJqKVu6RivQKp/s0+JzJDJLRbgyHqFDYM30xhHJIOEvmoUNkv4ZfGtO9n+MXmnlncIiygI+U4xj
Sle21g2fBJWRm4Y77irKaI9NAkskO80X/CIknUHy3B05VrtxB3V13frD6UAMplXST1avDrWzL3g0
/Dz6EEMXY0YeCWzsUQxRnHl3s6ExLiLYZ5xOet2QcT/U7996QEdp8j3HrmNSOHsQbvZ+hPtUntMm
odsMRAvWxyG0n4uNpTePfkSrifcLwxeo7iVbxfjzqJS+IRweT0FyJYd1JPSkdauBbto3EnAgSfG/
lnUV+BD7lnvU4IiLlscdt7MX+NGgdNh/fMewhQ76W+EKs7uedQT+pOVTyv3+1S2mkvWjsUWMK3xf
0UaRnVdrjAi+AN2qn2r0tcNef3iC8RsA8T4qIAcWwosQ1ocAyMRthxz+QsT/sbpRCC8i6XR1zpHI
bFo2YuGlnMxKjIbnniR4N1VWGY3mmsB/1MbakFgWeiYhDFSq3g5qQ50e5E1mvk4VGVe46yQfj/n6
1kVv9pWzG2KYpeV+/om0WyWDHxkJQz4y4UiqZuX9Or+qmCMpwpjS7ectYLjDEgzzLA0v92UvCKUQ
YEFT4iY2aAKL/kPPuhxIah6NhBkttCj5G0IbkpiL3CM9sHijGgwgkuCjClYFDrzV0ZA+94IIE/c0
3dtjoy2CFszVp+IGox9KQmDQVoZaUjlCxIVSK+na7a9HXbn0M9H6Q79+5vI19M5PxwuDVJqyql6h
YULrvQOym31wjsuvFpSOLu4foBOLV2wEGKB/0oiem15UYAhuUzaoOlmieJWNvbxvcGUYrCaQvieh
P0jbfBc+W0oQKpkdyYPpEXfppIluU1RapM7Kc4aCCP+tt0ttxoyZRtGApSfcWKt7nAfDvWV0n5Ws
vPapkG940Ak+vcoDNBUl4oQuMqfVELXXC6wJBpI2tqtT6rf6AEYVde1JjBAnFS056vLG1nUIGMGH
TjuhYsdwX25jN4j0ri1TfqvphNHh2Nj+xnajUFriiHOnFZr/WbXhZc7Xv0gBNZ7or3Cb9micrhb0
n0oYT6E0ar5YBILK17NfiYHOv3Unuphed8P2KlbyTV/ppIdyIPwqXAVYX1mky8UE5PzjqLVoFCou
ReNJ4GgKlbMa73ySP2KoGgA/GjcoIfCRcsbG7X5WG9IosWpCWBMWLW/gG5nRwSSu5IWF1hVI2b3B
aZ2klnEVVuC56jsTf4w38FsQ53Zp7ECaoc+MNSST5mYSziV+B0MkNUXXSpRzvosd5b7q3Ob/XUEA
PlUQZmUnBoAL/SghQLt4YZTV/EsaqLvcXI5PKPJV8H0RV72AUqSBKEjzR6RJM1zKNc9US4fiyE8t
SBeZpBQdB1BEXaBIGetXlJGGH853PYPhXqU2xDU+cbL9SOcIuLNdXba4VJfhp69tvBOz8bQAkgR0
y6xloF6Xkaz/tS3lVuiSLluue8uv4K2jbDSpazupfg7cgQz4rGDjpQ5rSj+pOGqW9mnj+qCvEy35
TZ3n697QEqQ4aXI90E1C28XxtNBigSBXkbAXzKIxBUaLFAHW4xZvyfVbDYQ+HibbB1FQkSN0li9L
pien9KzDvfDP+yDI+lDLauSad1Xqf1/f8lhwj5tGW5tppe99mi2sIeSTVvgYYgKEzsAJZOTJRh/L
4xJdL01QmdP7E4RSRRawRASGWp42lUC/WNbFUJZDTdDWTNjOrNR+8OHb/QxhUEgqk9kY8ZyZ9lSK
6NNwam2J/xHhRAWuzUXZaYlXw0njv9nPsbbkS9InCif4CX935lcIeSNgqrcVyv1VtiPIhlII3HKN
o0tP9/wXBM9jsLRBkhL9zd9F2eKcTjCkArYAq99Qo5e9T4m92m3MM5ugbCQltBJgE8NtVwVmcxH1
42tYilgQOcLRDEW5q58u4Uaw/JoeXyHQOPi7S/RROnNJHzKf8sXYb86kPojkfHGoannhIXO468oM
39mZcZ663SINpbrLauiQWYBtMf0sQPCGuu5mwKI07dVjMxpJ5uhLv6QiaLztygMFgAVvZLicqDXg
RH5tQY9444WAyCo582ClzivGDASGGJUBavzpHNOWszJHr70DHNEhkz08KD6K2AJXuQhg9Vrudf9s
a3VcVaIU0jdaVx3plS/LzCZ0a6o5zHJ84cvjDY8JrlQB4rvCkmA2U2onQq2WOLV0EPZlo1kyS7Y5
LxS8fsrKbXWYZyO0P7W1C5SS6kI2EpYAboTP5K8mqjlEvJ4EANwCSLplZaDBFOV48HbFoGvRlLLj
sOI5ax/69p3c/IuV05u9pfBxRv4PlCvUrUZtic9a5ZEVE/ObZToT5XFIE3jxfBmLMwxKiJgkdxIq
NUmn3018/uDTvzYbueI2Uw9Z/FtwcWUrPg+9p0odTM2LSg8/fpCNwuKcrNy4qdRhe/lwLPSvyDjZ
sCqITFG+5h2hCYaKszCkQGgLashj/v0eMb7FU0LTp0D9Xw/LfaVqlkWiLZGC0xi8gfhlKI/2HmoO
n2GZfXTaJIDZdKlQ6o6inEJbhQqcAOBjtZzNvKsN4JLeJpCa5Tds+mgp77I+egsnsB2A1k6LF0pF
z/FlGdjuN3fFGEz2XMk0KwFCmy4jfhA5Q522MDzo8GEb3gK4URwtHRkmNNlXwObMuqy1N4Izz1ya
tSvwng8Az7JSP9u6ZEQuNbXh1KU8hg+b7U/TYVGvFGy8XYgkqyYhjQSPVwiSzH6hVCLshMfoahld
hy+RO7PEUN6WztoFBkh02zAaqepGIsQvHQxzg7ZSwTTjWvBGLenVs4xDO8sAic5GpslH5ULdyyZS
F04+iWvBFOH46uWa3D8exucgPz3e4IWZU/JeM3CTGfDQbko8pMi2OxPvgDs/H8kcW7Dop2VUNHdp
3WDMwDr9PN9/vOojOE9q2AIkgaUxbRlKvnO1QRtfOHTzmepWF9G55MRTDvKBR3tdx7VrdmLQ9eez
HtYisxCC6jTZyhM0JH1voaf/nkI9cThcrV7/iQ+0QUke3sGQ5oP0yblp7ybzWeVHBAB63N6c/wcF
ZQHZ37yFfv3ekYQhE0of8PNxvlZhnXxUmJWaDGQ2fa5kHYN1Pynn2GSYYj6n1+t7oLDdCk6SRXBJ
+pRCBE+hkkP4dGOnCacQxN7aXR+1+XRtnYEiU6ZNpqCHMXu+A7d5O7EJypjjXWiGaPygQK/EThul
0K9/6f9l3VvQTgkyjyQxiYq0makZ0ZRgFnhILE1Wv4T2ymF5JzqfIz5rNX6Y+xiRzPZhjnsuMAX8
Fl2HDBz//nKjAWM+byFcOHpBvauW3/RpWiN4WMbre8dw1uyzz01WAbYoLqTCGa2N0EuX7cqi07RT
U8a5JgzT8EFdhfhE5YyS78NhLwZEPdfOHVFostSpYNbTuDchON1HcK3nsHH0sRyt7kez9uEpiLcw
xBc6t4wcfwS5goar29aaFAihBk8+qCqcS/gD3njKm3HKIq7PAI3fLLRbJmHCsnyeOspQUelFpLvy
YYYixYC0vl1z4k/Dba3ENDpbZ4jEiv1EJKb42SnhKusYGDo8ajVq/XJ0g6VCqgKt0e06vB1idZ89
IYOFxTj+J/X/GelNVk5U/3UNaVsd5cLJdQ+kgxTqQL6s2yXzJjLxsU4c64aNr3cmbK6LZA2mUXz5
U2H/dIsX6gDwR89p71cybxaUqP7VOBspLQPP6w2Jf08qkxEKbTphR75JMeIv7MIhFcrmf/ZquXfC
1DbEW8A++RznKKryES7kEepybfyS9vtLPfjbzGIed961THi7s7rNBK0p0nMyM0hpcb1dfw0F/bHt
MfSShW1b0FUJvZrB7JuCTDw0BUrVEC4WY2wIuST2OaOlunEm8cerz7qOIpybPhWZZRfiKFUtAHFB
Ur4sjFV9IgokNrKP6RtKuN8gopF/4PR3R83PexlydNeo47AgyAsePKepw0/hNhwhbQJl4uBcd4RO
mmOwFXE7jvXzrjldmT9ZxAjiaERbKAa4uTA8Gyhcn2WEXxVRcH6ruuUXgf13sxA24Vb7VPzeYb/N
CvUP11dRnv0o/Cy+AWsJ/Qc/om/FH9hXGzfmzSNlLer0R/LOD65tkZCJncSFkCIJawcyooZQOCvt
iL9aGK6oDbsruwI1QPHg1xHkl6A7PVJeUniIQUrOyV4DV8vEVkE6bMgYq6SnBNd2+utFum8KfUvt
HMHKlxOr/PmAYk9v0h+yDkwj4i99kd0E10KQ9rGp5f3CjhDkQCkLOt+vcPHXytaP+X8I+C5YvtGc
U2O/c0FVO2omYWp5IbDxMFoST1tQekeHBdtLLklA+lEM7XvmokCWyOseq5S4Cybdw3Q8cIxgSGjt
cl0uxyujMvz78WSkne1Xn9vfVllenpvVqGtSLHDW9ZiMmRp7SSL9bDos7ntVEM0Vuub+946P1KJp
bcoLcdcI6yxT5GgQlHL1Peu7vUwPC96Dczn3wbGc6RCaoa9nWwGbYVNdr4ogQ1hXTKJiRr1wj2OR
Fcqbm1G7wsKV/zkXdFVPlKBu6vmDCHu3l8CgnZpKyyl8sI5fi83m3Ahm3/nPZGkymlWFDz2Y0btW
B7MQPSizKIWeh8f6e5UIrZ3J8R28ms90+ySoACvxmm78JtGv/Bp7sWH3Jww8ggYbRckXLRcQjSlu
+pSxDzs505FL4z837VG+TOWrfgjmmM+Se/XnPSUlicJfiluOSlXcScFjYtgLI0wYNdR+tnPZ7VLo
4K2nnQ+b5yIfLSgjNDmkpq/T0BkX1OvjEH9+Y2G8JKDjYUhRKZxlXCBTztGkQO6lh8QRYs7ZDlgu
gD3IflHv5weqhKI2aHfwslvbyrI+d+9Ab5r6mbkLqaqUQJrELcpy9mmcngYWafsAOFPwwUkktzZH
a6iq4yx8Lt0op9YDGhUTSQp0Xzx6VnQJvc+TYzZ358uq7WnrAdErSG+P8YTawO0F4a9JYt/3Sfyw
t0b8LglwEX0AljU0spxn6SJ8UdCnJEko1ZSicWrLvn06rAQSOnVzMmqKRA8L2nzdMqUYC2eQ90da
npDQ6k35VSSSMwjooiTpnH4hV1W3E2VDAgLtX53UhBR3l/9P57LYnUtUpdTJ+aChikbCfjtqrHD9
oNPjZMtCVhJyWsI3JxcclsQpuOSoM6hxhYUEGaEEa92UlGaxr1Go6C7yUU/x2DhtUlhzrdaWgzx+
lceYzeBpRvdPvymSYCl1d8GaHUivTtwqmrISRJYnDgfDbbx7u7AGhPl8dm4msFwq/Xy8wOUODKbL
SJ0BjHkVj3rz3WVMXQZknivJ0pHr5Iw3fZWg4iaqFx5u42oYbEOHAyp7HvRRWKWBtzTTFYUuJVC9
2zGo9cseJG9emmAjIdhDmZKK0wUkvo7zyhZGH6MIzgMSt0jAeBa/02s038poUO0vVXIdKXFn5y8N
ylVBXl4wB+Lu+oDtn6CCWFGbOY6HCt9sP/fucjD4gkrRptp3jpdxMQ9FX2htBJVd9A+SXrMGUeq3
h4lZA+ii75yeB8lW4zeqcve1+kWbTLTBomyf/EbPiupcaEovSUg57s/jsDoazPIUeoqUhXLJnwL0
smXaIJamZvw7SP9pGIM7e5IsdQC9jP2p+6bWdZgvmYli6csmY9/LHW1//KZzRbW8dh5uxX8lDOZA
Ob+NcVUk8fMZe/z2ZUc58ZdsR9syM02TK5mxnZGagb/PkTA/wVMEh1JwOfAywObEHIwDNKdUk2H8
qCqvow6a3iAuMkLWF+5Ju3LYzQCQz0Fuxp7Q7Y/3b/GsK3XPHhFqfapb44x7xyh80ivMEbuQLjQA
cSwW5NV2ZgVSB/vE8DLE5Yq5atNJgy3oGhd3Epu1P1OYN5FMD2w5/SiUp2zirMKt1+TVpefh+PdT
O344KpkBn53w3RMxqqJcBo0zA2PW+iDRTeDT8K8Sgm12b4yyNsSPB1phpbBb/w48DMatu95zSwnM
ySOx0uws9KLB0qDRoT5TImokDJn2bufQHMS5l3oxrDI95RiEVE+THa7k267bHOA9wtyKTZj/80of
phSWx4vPUJ3F3VW1ZTo6Hj3MSu27ReHilerAthrr05aGcuZsHgk1IXCZ4aHv9mj0VTOKEw5dva9j
escQoTrbZHQkspGHAgQxEi4UnVk3L4J4YlukaHJHvOAtZSxr3bF/dzSMPHC1HBD/HdKP2qucwmUL
nhuoj/B0ge+hsH7k6c4iHQZMpQsA5aAve11O1EARasS3GDAv7J9C2lhgvu3b5gbGT+i1PR5t0quE
LoYeelzQj7PiGg9wX8cHcd93f35PPYL7hUo2VhyapGCFikiqI4RRbCgOt5dU9JhO62LnDG6OJVRW
5BuNbZlE/5e6zD6JFUvdQhjk7UANuVXo3ej63IZ7M+CKtlTO1wJcEwkyN2acFf7jjaCWeuut7/UW
gbgdZjiQDde2gM7fyGKXu1tQcaB3ANmvuPxV+jxY8CTuPDr56p3ObLX5DY/4joQT1hJ/925YGtYZ
eax7MVUgr6jtXtN0j3yXl+wQnn6AMycLHmExHSha7Agw5YVDLDra21ZFpre4Yf0aUnTSMORUOsIu
HDGWvbSWB03STg5sonX20jVN+zyfAzFMSrPBih5cCckxQV6NJ1eIrpiS/4nCPh+UgbRxPkTa2ub7
aXVpS0L4EJsDPhLvvuUig6N//Y5OApj+QEA9Vw5hGlorMWWz+q2Ey63K9SHYOwIR+B4z1/WnB4Kn
d8w0/35iNiDiouZAymwj3a2nJ3Fg5OPSzxVLnuE0V6GXDCrBvx+yeX9/KH3nD67EDZepb9fPon0O
gUh8qRAjRuxleNqb7RV0qQ1yBn24xxdg6dwfecw6wbZTvZvc34WmO3Yy9eoCUH2WwSRsz7g9w/z5
1LSxGKp2zmgIyk0iqhXcAZDeGJ/vTw0zBf1Qp8YJ9ty2xJUr0nz9ackIof3HlxebEatO2TEPK2VG
EdllUw0uHibFXexSWf29I6juIY1Dx23ZZlqygix/FqqZRoBN7FWUdJCQxcXVPJZqOa11VEPQKbP2
ZCmLuH+ti1NNOWIkh5Bm/lLyVsu1NHFo9jI5lOwCsfuLMhd9ij4fUmmsLgFSolVbyXTYUIQAYrN3
vLujpemK4GTxTeiqi0PtIYn3DGzcZxIL+w68HL21/eXxcl7lyTGYZHbJVWLaEZ17QcUE+XjKRZDL
dJHQfY17C93uGMVbQg7cwSkW4zrTH3PA/vmioGkCDUDSBXSoVNCD+ThhI3Nqy792JpqG+EkLyRVj
q+wOOUrE7uqw773BJeZfLFRElAzzjZWdCv3Czlpuaqr8BZu2LkuotCf87PSeVBZ0YUeI2qPfey0f
1ImtMLlBMFX7+SRCZahdzsf79s3BKTtfz37WMdwoGE91Jsh1rHNwXmmAytJ66kQjZ9iWO5phsLrP
BbQlbSviy1WsB+cFciuCYmO6jSU0nzKYDQhR3+BeZrqZFkmRHlHhyRsyZs0mZaFRoSOqYn9BHUSK
i6dAmueFNXW9r4yY3rekO4N8HsTTsT+jv+TOYEJMIL1/v2CelJ9i6iCAzd9mIwZuNQdIwC4QMc+/
LhcAmSlwNDSVz+tIa8GMiAcLTa89/SsWBtLyzthGh5fFenUIBVVrmGwe2dkTfBFIpLhibzKoWa0L
nqe+SRDxOO652I+lJ5nUUjdkFvRB/STLevJBqajg1SyLxhM39Xc62/l0CS+Oc5HJv/vjUPE+WaZZ
Ycn921FwZ2yZQ4I+ywwlF4+iOHOMSemXI+4YgbuI6Dqe05bZubHd0yBYABu/Tk83Syb41cYQBDam
j2FAPS4NH7mXlTZZW6b80Amsapb9T7jdp3FBECcKIDTTGYCPEb1KMqKyA3mI+lLTqH8ycTLZBV0q
4CPfhF/QaCYcqhA/Fmsf8cF/q/IEeUSZbFoiphX8Czq6Qmrivq5hBUItstS6N5RIxM5Us57Kb76M
9LV3V+gVpjBaUqmEsMe1cxwMmbm8h4z2TBwSK5LkPHuRTvShXkRNZfp5HC8DJqc4nKnv339LZw/n
+PRmy+0NzOJfw7/QpTkInfJGFqnafbeuSq8iOI10KLAHJTpGFzPs3sNsu/4qCyUjp8IcAxjmV2SW
SV3ac0OXYbeMSUDfeFFV4acK3N9NPnzZajX8Yn1pX1SACXLXnWk023C/4tqhP3HXDlun6UrrSIca
UMN36WtIkn4pngIQC+M2l8gcDt7R7K60qZLOPlolSFN+Oz6wJMRUhE5H9UGih6U29PWHibIlWgl2
+3om3AETqSCVpt7VwiDgM00iIVeWDyso6zVNPdVMUskgJgGQu8xaqzEYG9T3etELMFzSxjRfUCYq
7qb873iE4oR4L3yp/VgIst1j227dfOXWm6u6kKt+rUOa+A471yJwcZOs4/cnw7hroEC3Xj3yxSIt
DW6NCJY+yYHRh5PZl98MZ+2TpoSn7UsUDvBBsEzqADB8yeVWRE6MJC9nqqYd3eFk4G5fl3mq/cgD
+Ktr6UJB0FaoXdmk8YLKmcfsNwxtgkDT6ZeSqGrBdjn+EsihLXS/oB1Aktqe6Uri8s1RMKPpDK1X
MN07+wbEQ4jCI5R5NeRl747totI9TA5WjwAlTgF1Mh22rPgNeC7vDtoVaKF3Ug+3bEUGB7wVHu5m
OYJ487i79tsoaF2aQdKc2o6Qo6dVlYGGaqdszXpCTRAU4cB9O6kpDeXNtyeqACwVyMp/2Xl3E/bc
LcZk9SmcF5C0634mKjljEL8yAK/Sem9/TvW3aOlk2k3DBNffBkcqn8rYIvBnbuuX/IZzJ5R9hc7R
zkWBhnB0t3L7eSV/x+0GdKL1M5NtK+ZdZDkafGnASZIvwW2uCKAJ3pmCRjkAvr+Wd7cZAG8+COxO
He9FpSZiBc5gxF5JRIp1IB5PIGDkfNJuZAeyrTipb4l1kQcPPoxWoI2aJjWU4hHqxzf+K/7goTgP
+LZ78VP63mk8m3m5ZsZES/bVZwk5pAqZXwfFH+xKrT5bL543T37e/DHnWMbOQHjDOgSccQVVmcbC
+7cGV0y3ONUaO8MTxRL15O5UAF8j1pxNYM/B12ssRZpIKNikk8DB9mFOafnLQ/1MsSMll2mlXGIO
L0P+iUuRgAn5Hk7Wy2NvrJgw5fLoRKplBbmLeIhaoppsGC6WtDOj4yy/Y1HXhHsI9ki0WlZY3CSp
32MHYooUnN7xdbk65Ct1pWaDatT/Clm6vV2Za8JeAToP6bbS7nX8A0LwqY6tm7T3oekDn81JueEs
QZ3QNheZ3xj8JL3eIMKWJeacYJKGrcgHlt1Dz+YunqE7tJcSzc0ktqgvtCP4s6ml5C7cMacfccFr
QMJsrPKoMOrUlZenDxB3N7RjGY7GsjjmL6KPc8Yb8B7L0mcNq75SbXME/b6jiGqFlIuEl3P1X3vV
+ovGlSKusRcux8iTM5hAVigzBf2iGzvj1J5Y4NSu85iqbEMkvOz5Mx9o9pj1Wuryw/4vjURs+jTh
zWzXFNjpI0Or4naRXtS0SC7Al8A2QDaVmZsAewiopwHxzt7o5YuQeOsROqP0HAZrtsJkcw4+UjhY
+EjA8sWV+xPHqR+O0GUWvkI2vQzpRqMzee9zwcxROibqlZgOHMSVLlifYOGRlOac+VrbQL1JJKUr
3s6C266HWSKnBhYzg2pMKPQwFkVfHmIbDQiOJmn1B4Y2+MEDM2889N+CqXBFqAwdoC7FMeirbGp9
5MdjzdWMCoQupE5pOeOnE09/8wTsqcmA9yQdiYsY+uq2fYKOLBJukOdIqB0c3uK0itxFxQYliDZX
/ONY/9ecYz1Z14LkONfJ4g/DdZtuv3MbvKO12g2gA7N07/NT2CC1KxFweNf4pfyOs/YQHwQnDKVC
CfmLmBB/5e5vux7aHXD+MiBHV3gRqTJSbW2KVcfExxHOUmIJK8uzJ0CY4UpkEQfKm88CFCf9HsFc
7jn191rP2qsxlVCW1fbaRsVmFcJ9ERDUwpIajscWnLOrmYkdKEaq5cHeBVx987Ure128H/Mg6xJO
6kT/tRNHUN7/IXiGVsgzJeql22J80VspOC5OOIGfwb39DA0nL5t/884/LA//SvCwxR9Vm15+gpmH
UGOoRT3dOHOahSm+8Km8dxu6Tdsa4a/an5K2iLTFVZ5feUK7h41S+esTZRmatymmF07NT7LpMM6v
+lxDTTUiRcTvBrM1QZ/DfxOujnjFPOyQzZpZu2nWQ/RWuVLhc4OVKKBqZoOPkM2prEgBNC8ja/3W
/KioluHK2FNp1SGVjpeIfk7oCnKxsPycGzqjXUwy7t7RhC8gJF+RqAmCMxObOqSeogKhAAST4Q1k
cBWVnR4O7l3c/G7IO5j/tuEjHV6uVlR48LqoyfCFSamO60CjQXFWXxfU/ZRP4jiC9HHFBsGcvaAx
EFHTIsvhdIqyWugUn/BssECMVmMtZwyiLUN72ges3GU58o30rSA8lrrUNfgm6UVpWaFV/fupdatW
IB1yy9ajyIKBgrOwm4cnS6n3Kmk8DbRmn/8j2YDVw44F+x8Wn+rkiiOH2I4v+DiIhm9OK3z30LNr
UEMBUUtI/VyLTDR1hBQFLWe+53STR6O+GK9fdXQgclDP+AjMphHTxYOO7QLofX/HpzSg0dTfS4gk
YzZCl3+SVqHNg+5FdyR3eXS8hyMxFmHMKDILVhF14cNztu+hGLNMBVu6lO8iZS5KdX15jweKGnT5
WAMKLQplsuJ/h0fsolVZcTSM5jD7oyGxz1CfnNxflbayH1PJd59+m8eziPO/U+AMFqWX/jGhTg8M
DFeFfkBNm6XXsQ1+MhwjUMTbed3hEAyXc+F7AvtG4KQuemjNWaxObqVgN8q9w001KJdOw+a4TrVT
j9orhz5AXFoO9hWKpVzWPl9fUjZoDPSCAo7xVQFZ6h2sxej9WK/is34rkLeSmmc4ZypL1NU8QgSp
U/Bn2eg5lrI5xMWhgQ8DqfEVy2B8VryQOC5xAvpb1w0hYl1BI3wr74VQOyXh1ycl3YQwHy4egvAg
fWT3Ub7q8n4/2DgZG/tMW0k9CdVMGE0svLlx4k1Ve3pdO6xDVCouoqcQzVT84A0DRheDi3k3QPkh
GEjuJ8DnvtQ+k9oBy3hsgTXI2PkV2eE4i2BuJnfrv3hzyvNKGeOrRXBVAQKsx8pwyydK9vbuP4Uk
ypaeFmmAYVmygNpC+wx6u3D9uzKUOE3+6AqsZF02UXnEg8Wy2sBjpadeQkhNTA7nwE3f0KDXTJ1b
ka7NX13S++hFZYZAFwEm4umkMrZZO1/gK7DxWeHK4AxxaLbKG5fFRoIUDaACdA5U9srj+Oj/rUY9
jRgaXKCZ744Gomm+6Lws3jGeeSsYjorB12ZH5gr5+4Hf/CO1HZKWwpDRAAN0g5WoZwJT+8YjWS4Y
KVqajRZJBWpy3u5Zwtc/y3+vuV/b8NmMsuYwCJB3jQe6pBKC7FswJT4l8AKCG8liMTX3dU73INXu
8US9W+Wg6a/rBwEmBb7m9Txy7LV3WzmIPreW2cIHvafbfR7+jHCA7yx97q3K8HFips5/9EfNn6Iv
zO6umgMDeRBGJjo6y4EuQ2H4w8QggxIPuHM/hLOBjAgR6qMJIDrru6GFT1qTHSqGb/+oNwl+2DwU
3jKz9ZT6EikAA/BBR1QQ4K3fNnvyovCKU4E5mEYNot3z9t6Z/9ux1/rCGB9ImviO6aBRydyukNdV
nDqIC72CfhV4vExtB4JZerf2fjJoPWCGGaXnmU8V1HNiwVSPl9fLVl77GCbGfi7ug8ZmGDu/gweK
x2cN1ffxYKQyHS7wRfoncBICm5dWc1aZn/WIvt3bFnF5aftV/wXgKssM4wnXKFWh5AivO3dyTdkw
LLzEyFSwXenPWD1WX9DZyXcqHh8K2jOOmODD6F0ENZHMnrAuV2T8nQ3Hq6MPkP4E2jqrpGzydwBx
NPfn9uioTFkUnIu9jkLwhyx6CDtQwBSobIGQ/cgTu2teDFt5Qf0l5ZE7ReaDbIrQ/Dz50b8RvQRY
66wdBtM5pMzoye5G5HwKhXbhaHUSqYWSJPAmycfBGfxj2TzKeIcnS0Kelnljme8A2LcjhhuMiPM/
yQR9uep/ifeezrA4FqH5r45acbl6CKd7+u82lcFv+LXgAQJ5R+Vc/PdB/R4g0zcu/b/eh1+ARLPB
dYhMBLD/WejRCoJXXztPx76ygGlWCFRNi0gJ4S25Id/IL3efzR+z+yd/u6r0xFLcQdKmZzx1U65/
SQPD5pkWnN8XUi82/EplY1JteQeBnEpPIuuaAGrqE/eDuuQAoScpjG/KrCvzS3boMFH0lHVP6AN6
vNqFwg7Nd/9RO1/hEGJI930+hieTgjlCkAHhyOdNjd73ahL7wqRhTxisAdh5obvUJ/HQ8GCt61MI
r++y3BscdCI5A+SpIzI6hQZB1gERZlJ8YrRTaw8zi52t0OUUKdyznHetXDPAC2G9Xkv6hlbdpJEl
BBQYrxG44nRYUXPZB53XKMx4SEaHRs2JCRXEryYalORiLF5i5OC8KCLiJgPurRzeveLkvd4bWODZ
R95ZljWNdDtvxfa4lxk96WAGN/TPKxlZczzFPXXf5V6Xy/ly1d4ZIrzokGQcXt993Hm+U8yLBrYL
92EFCHIAHwNCRkl7Uii6D+0aGvQtV94c6p0jPL0jUj4lRJ/taiSb1GDUW90mdyRBwQU8mzmWG0Qx
yd0nBhYGyKrvaSH7Cp2Q6WV6zxRm2iqQ6xrU5isrc1tKlOf6od0xXgSGutMFCY+IkXodd42C6Iu8
zARH1eaUK64OLTblqWveqC1rhT/83v0ku1jL0JlDI08hZqryGYsF6InVHH135xx71ehRYucxLFcq
htnNqVaKl4Y5y/zKcLweGhNpl0SIW+xos+W5eKWwXo6jcIEZ5UbTCC5DRzNipvZ6QsLwDiXQaxs9
52w3BnssDowbxKHJJja04BczRwyOGyE3RqNvC7gnF8VAIUMxbQQ26bEzGdtdj8icFhBRg5O0wzNt
iLeNDDrNLfwz6HSroXnTR/kC2iL0xtynSGVaCxf/9A2iU9Mq6lcRBgvSK/KOfFtOC6BWtsWOYouC
CPiz1hejeVMWYJHTqvx0Sj879sWnX36uNtcdb6nxVdCgZkNsHIbyS4zSXnl3T/wS0kXrMiKeIn4r
NmyhhyNhqpJHjUZOrvoIYQHkAYrCuc7suDP27getK7lg9eSxjqmDfToQCEVQS9iTeltFR0obgoTl
+zjEpkbk5zx6R79dvaDpkY/uzVgIl/yYHR0vNbRsC1hR55bEzRdWPzUnaz92/kSCtnZh5fWaV+Gj
MLeXoNz8CN332i4I94ErbK0hTS/KWtSYYGGFAMtZ5eGPBfahgwaGN3pifp2/bUOJdU8Il37DW4Hk
aW8Q3dBLOvPLdAcekpiFGdK/1ynTJLRJSkC9aVqFUJUKpTyCzlMq1e88Lo/16luw9SameSjPF65A
4cROtWt/F6ptdkDmZKa3d3sABTv+Bw+EFjal5ioof248GMCOYCpP1n0BKFHV32F/8AotZkK8HCBn
nOz2u5dAdPEwyJODZxthcicBWYbFpLOT8CoDvGPQZ00xaLa4Z1yOk4AjuIZ6AS559aMG6obLI4MC
Rorq4/CUph84bAUq2OoCksUbis60+R30PwB97KKSKwPsUyyzphAFVKvrY8PePfxlhADuFpdhG3nO
YD8jh/EUFX82znaZWcKviykmHjDCOtpsv8zR0HMnN/lIZ/vqFdhclvtXuCVDsdRNS0nCTVZ2iqM9
SGbMhfN4BtNjkAgw66HerPVr7rkaZOl+aHvkR8oAhStj6IwS+w+C50SY/8pWl0TgO1nU3ZWkzH7o
2jsqwTVvk4AyDXj9U6yVZXV5YiN3d4x8lVvs8AFrtS2/4s79uM15MluStjhvcvmkEqN3/P1yPsdi
BeT06V881oVtb76UCz18zl6K6NAJMhXSGBl85YW85hx9CCQBkxm/A7kKlKIZtPV+VFOXT/4W0GHk
AK703yEQ26Cb02X5S/gbcoy7ghSiW3SCHOXFyqGux8czvXEVKAAV+03t7OptYXym3haDa2hsF1DT
6vVrKBvXbLeUlEC4b6B0XhXe1CEpRuwGV3zGVI8pR25AK1cghI5to9+JuSLuCIPel9T2FHOpA6TB
bajOGNbs4qK+MfkEyN9Kf3cJAkb6LHwY2ceagIkH8C/RjcbFx1B6nDGN4AmV92NvIYfyy9mr26Mz
zb0pgqMp14JijjiPBCu4mCBW1nwhEu0AClA9NurBu223XCkiKFhwZOfnT9MWa1KpfDgvSa/ch89H
v242tNHmjt0RfSko9FoaVXsInZwlPcR3HJlN2v9X1r7mgjDCUaHkvxbFzDyzE7gIo1VpkAn1aAys
6Pb4RBeJ8CHS2Mf+wGrXVIR2bmOZYFq5k1mUyqC2ZRdoDDYruJyHZU8EmRawzqWsZK9a8dgGMrXS
+FkAWmZSXKzE88FsSxSEZTNB3O5MN6e7e7HnY+ZP2NRN3OLNYQBq5sewMg9cW4g5pvXdYDa0MZU7
DtKI2+9wjBYtiZX3kBAH+nmGt8ItEwj/5UhgQgdramfmnS08Q2mDRYfqn2F/j4N2RMpFaUWPn8uO
oOLJSPA891e8mK4qYXiHyy5hIfRNG7EsClOHmVv/tBJug+ZByy93WeZbXvKGxseih4xbjuA4/m1+
D74BS2f5Ileh3aZXh8ST7pPvHWSrEwn7hVjunUCs4VvgCb61hy5eC1vb11Nkmi+KuF+YnQB/oTQH
++mdOl2BvvJS6s+5DhSAHGqCfgp4Bw1qcuw+FJO5kPZ9qFFzDY1sI1ttu9uewe5vv0C8tL6Qlez3
tpK3Eh21bzjRUY+lqktgr6UgNxZ5ci0my05OsuiZbo4RgjgLgbpXmz0CZw1WChJL88+rBDZEiRZg
mAQXFUOYGXEV7MsQFaMEcWlhOkl2zKNPwiMoJXolH2xGP7ohplKepPwufNO2VtOubgTWjZ2yxXEb
KKa+JX2upA/GT0W3lPsnRkWSqqTgEe9Ty5j1uB2bvow22VCv2qhvTvjWoKpzloEsolEoFW4iRlGx
dlDuwrL7vERU9hIVHwkkZy5THOBDnUJQuIINXTH/wEQCwTIOUfq3e7RXHCw05qEgSyUEH8w1Ex1+
mO+IgswfxIZvG5Qmo5IM5OYGqIoxbThLU52RzCPUay0zJZcvD+N8+IjkXyXUaAgW8O0qy637hkOr
BodtfmB++D3KGgR82iAz0iUG23r2YI1pwF3/eTREQ+LNdWJ18hlE1XijD1d5XFgnZKQ5O6JFbBQN
OI4SDWSs5LuUkuC8X9qQJO7EIImza6Chjm8I1t8jqBq5NtuZ1ySSGvMWXqCmEQqYPYoiSeGNjzzj
ABOP6Gm8QJwJg8bu5+woGZ+kDc1LSovfQUpG70Y6qhyXPmw9yhUdX5pwuHCXzlUF3evuBiWwomNI
i3ARk299eEFHS5b/4mQr7cT6DdxzLeDbMWq5EPXlMMt/WzJD6VrPwVj0PvcHMFX+QjJKDRFDmWxk
YkuNCuEJlnZ57JRjOc/+Njz3eYKRlZO2MzcWeksc9/DJDLmPCBYq4FSRf5SOj1n849R+7aOmogWR
tQliy+kXdRRtsKjJhOgBu5jRcOGv3Rd4R9ig9pwRN7NVF35WWmc5oKDger7qvDRi7rQSBiH/hAxm
IV7d9BGQMdkI7G//7WvrN3erFSlvPi6HHn0cM2PecONtRffPdKFPqCCXEcqf7gN7rIy0wUJCzUd8
dcW4dwvQgZIFdBcbuFbHQosQYI2JwF4cRXtOXvl4k+H5IisXD32H8N3Ufyr3ECyr9QSfMsE1LN/e
0/EExUnvcAXFq1Ej4BSb+WQfaGn0nbDOb4EvJcBiFLysHQ80eUxS5WV5Uo/No8488l/O1XsEtIPx
fFrI5flj2LDopLhaFXaLNF2oPWfA7QpsYuDjdoaPC5YbCv5i1IYfF0HHYoAN9LD7neA6ExseriU8
nyecBNl7PZM2f5fQajviv0xdkz2L08K/EIOMPsrH79cYHemeD60HQ3BV7xwhP6v+cC1BaOzgK8/6
oNfxVE7+b6GXJ5CO1e6SpwmrwzH0OIinJxrnlOo4ldjYhfv3rgOqN/RZwQ/5dk1BMiT2o3uarNZ3
uLy1tUrLXtZbbmRTir8oTGe2tdJgxtGxjbZmnMkfnAQgtbivgJGencx4xb3UXjxm33lKUoKS3cHs
NgiBCZ990XybXoR589KpsK53rhPe8fwcRFBsn2xq1l3QawOA3aKPE/3gYKqAaII9jdaakmDRniij
oSJgwGW+HffQkU3DGNdI2JoBDp6woeNHrEeW831dJxUA9c2HOUDbOL97oPgB2DUucWGlFbI8eon7
W9B6zDptNb6lfBI/hwCTeB41mAhUgHR1ww8R3ySUhQ70hb1eaBAKmpKRmaJbBFHpQLDIMB1yufK6
zCnuSsqhb7AXrj7aIRlyyi3Zv1zNfpZS61fumqPZ2fBughuYH9yeq/Vowj6ETJZGDRnzLUMkLWMS
12EKpo4Duqd2DARq84ddT7wOuYVLExAB+MfW57buuqu4mSFPThkH7zSUQ/9076L9XVyB6RiN1OhS
z1ne4De4gRVfWHefFMC69RuDH7KiXhsTNagwe6G6Bnp6jcXR5XxcK9B0jQ7Mp7/jEYFsMEFaeLJ9
4x616dTFeEus3/+huHd+4LuJ1Qn8lYZOf/ucCDtTKJuN+c/RrqDJwDK+PX2987PF1+nrAOgWwIiR
M/sYaVV5248YqBF6zuoUlhIyJ79PolJDsuV+2I14Dx0XCzbYu1dhoDHKKAuIZ419qRhrRUa225QU
vdMG51MiJmVMjwnQ1hWJEeCici3K9C7MMRJNnATzWgn8nrHa4YR0OiBvtb8UINSjRwXp1w4GFaP9
JRRrJUUudlHyNaY8ME0FYjy/8a68crMom1WkR4+jCJo5I0FczgiN23aLirnrmwua14V9dPE5wI5/
eCZb7W1fJcF7ebiavQBA7pDvqiqNxgGEqutvQVakgmrTTHdX3q72YJoXPB1sdfGkaFHswPn2eXbE
hhs79Np8jtXKvS1M/TTKo9SlL2aS3U9baTqa3MBrlHcTdNy2gxb8NATOaHBZR+hviRbrAoC/kP/O
MTcY8AImr8HAf1x/3/VJyIhu1i/2AdAksb1793xErQ4sNKYEdc/SUSviEgspn3oz1BcMROSkEAzj
C3l1YBiBWfMZhOYupR4OG6F/Lx8eTT/RtCswg97Xb3+McxvHDU8nkDdB7EWJmQjHL8sJbhMK1oI6
rq5vWCsvlbOwxD97fWc6arlapqx91c2wpEyi1rMLT8ld1V4K1bTNSqDfK8+92bqLisjTir6Iodqx
cXgekV8N6ayeNXMX1lwDhMDKDBAuaCkj324G0Z81V2tqD5/bZ0MGZ4/+dEErFVSHYusBlZlZ6ABC
S/6txTS/sRT9xLtS2o0XNpmRc3JG0dcnJoCPjrEABO299TQh3girgF9Dt4Xn+gGu2tEEVFguKun/
U+59C2F64okfclvwtiKM/V42CDWOKpEi8Lu62O2SYuZDEf/bnp2n/Fx3MeszNC/SCf7RMP+sAI7e
a/2wXt4m5rtSXe77KnrxZnttMIMTTrhJGjNVJi6Ns4Esk+CkDGMt1l5pL/6cTyBA9Ga88adCMFov
ZITwvqpOf+5p8EpbKeGYlstWceAUpfpNDTVuWD0hwZXnkUidBZQUjraERCF/dxSCqXO5fqw5Asxc
/Fj9mQICPpy/NAXP7FpBqm7S6CYalq5sjZWla2dwXkfg42TZrWQIk5p9EvTyngipKu0OdzO0Afrh
CCsyZttUJwia50wy0wUe6T6lcpCAIU/VhryqNFX+9sOeKk8+Xc5Ru06bSXJOR8VbeE/50D4l0+ke
p6wzUPnX56srtJQu0qBCasikFr9mh9EwjAiwB+GE5dbiNMusQ97meZqPatrEpLzE0fpDEMJSfWUK
MROGEw9tjlfI54byQ+YKZ82HqURgVE2B58CjB00ZvMvDB23HBArRZn1/SV70Xxn1Yfe6qtZmMfKc
5lmi/fT709BewvCB+7sIUxkHhcnsU4PNFhHAF+QKJWVis8d9/RlYLKs07Blt+zARUiSxxvF6ZeSo
nyzFzbXi6ItuwTE3DIPVS/WgrSkzYWlBSLG5daw9hg3kGhJDipDqdEpBHplGBuh8JnlCDT/jPbW+
AgLIwMJW1WxuJDP2HM+9T5KL6NXNlmujDUyOfXdgEz1JYXUrIyWXdykMfb3D5DU4X4kVobrSXSfz
Bupc6/DW/Ieofp9oAkLpy5O0FOUGjgFHmaGU0xierp7yBEGQv+XiJJDj3ETOzwD0MI0FYIoRxMSi
mGsuGDM/ws2z10O7c927sCcuqqzc0c+NSqjYdjpQ8q8FBNyDzJtDaeIWp69+WaZeWsmq+/nHymge
TvQr826lH27u1CtWBxLpf1b9wt8RNBQX/b2YUmkL3nR1SlpjuV3r/7XIL0elyg3ywEeZps0CtKBb
Cl+ICEAztxHxKah/khniTG/LeUrzEPKoXnhnisEk4RaffcOOaoVz/paMaoPEdvctWA5vz5vAPy95
a2qgX73JtWZO5howPMbkoxOwwRRiEzVeAz5JZ5Qc16h7ZjFRW21xTc/ZUsD1lwsidGB72TGB/ela
F1HVWTsktjsbMBwXuJR5SM+SvguzjW4AmzgogPkj1QpRrdXLj+3yahxJJ+arLo/wCWd6fKi/Eb2j
o9Bdq2bJztkzvZQ4mVkAl6FXBwwxhcLTwWf96l8eXcZhpGlbKVEkiAPebYyKgiOWEG9yvOqCcrPl
Pu/+iVOk2/7dnF6X50Bz64BgHWti8M5a0CRQoMFSF9Ag/pYC7vRKs4cDTJUBkjKF4Ix3cQJxgmld
ulDHDB9GLCAAEjdEKhRtN3+ITUBgS0bMw3nKIOsgb+VgMrFp5haTPxEfvqEVyB3JzzSxk5tICrah
vkWjjvlUPthUog419+geeV4ir0T0xdxdlQZpMhZGn3X+7DU8gOr4VJfyKBmCa3AKijZgktm/+odO
02YP+Yp3y1rsqFUMMTB4n8P6+BJ2CsygHWIMs9LnNh8jhHpT6dRcogeyfCAZQU2Flwif6wT/SbMM
nvBQV353tvv4IJH3RabjnmJ7Yz9AvjEJKdr3vo9xCaKiVDQejU36ZD75ZnKLdEGgiDk+Cx7+ooVP
GJn1ghZNWO9KVn9ReZc3tylz7K7zqoYIMMNbzIKcfKZruvCXglz97JKrEj5oTOof7DWwP2IlA7rM
g5ny+mNgcyhD+N2FHCbhOQaUip6Xabpyv8D/B2TJMMs+R6zA5Cxq59Se6T46ZockA6Q7GhTm3itT
bRvcM4FT0rzGzwJ5ggOTZ2xa1VSj9gEd2SVKCpjtUh39vKVIyYS8CzThHJv99aOTRS8bTmcAvVXk
1RhIpXWKr3n8FQW/m9aSxHhkIxlkwzgXecOe8nnZl+/O0qFQMgLKLuqXGrtU5TaBTBIB9SSwtKPL
ux8SVCP5gCoaY8e/DsGPUAU1r6f3bTsWnT3PxGgY24THWKoG8avIvQkRHSuL+DJQvFt8KwmOTRjm
MT/NOC43QGPZ+yHQVWF/b3QKnFqE2LtCaIJRfhmgtbC0e/ncsbVKzILekvahFQSCMzLGaN2tqtAz
zBs0Ebbe0Xl1YuyTMsdwnc15Ig9/HjRnAiOcNu288BZPMuOqiklexqWeqcaVjgjRK4umQcHNxFg7
Lxocc00W4uNdwwZBGkGMeIXfsAZPQiyI2uXcj+pu/fS/1hySi/GKmvx7D8VBWFi7qUIo2LrZo3C6
EC9ualxiG7/F5oi1wR7sRWIRSUQUtwh/qMBMqeh7kN/S9WhnbB/uqVFaRWo61Y8BCBSwVJu9f3YM
yVUMZHEv/7YLpNlMn74NWpXt/iWqlyKRi0WhPJDeHF9CgzgsKGpkNw8G9R2WY03Ml2Bouo9BWlE7
mvYbJjiRxFtVtQ4C2uvg65yWMqMYThh5JBzqr3Gu0R/+G+NIUTMtiljdS+cd50nY6KA+AosffZnh
UFzmOHytYlO1pens1iJ+/Ojy+Z6w4i4t95eZT+MJmAjWZt3F/UJITDCQA/97d/vkCVcq4rdcl5lI
WpcOZ65dulgTfyf/FTpUwMRiDrYx1l6Q3MYxEZ24yAl/p40WQ1y1I4tdaMpohl0NGODgxLBBjAKm
VrisviytnmILgD/cfpK0/ggGe5X8Pa8K03koKDguNh9r/ra0aLoNCmPsOTTurKq4TQdStUGEsreZ
Yij4XkZ3Hc0Wfv01xVmdUUTvSA3wjuBRAB27AoguEke5yV/Tt3maLgEPc4FpdiYi/mcJEb/AqobQ
IupQMxVM6oOyzGIkvH9X6swh4ai7875bzYDTjYrtVAkk1RwaGuGy4PmIUlFJAemGHqW1FG5RQAp6
QeOhnsuAlnotUvvzhoLh1aaudri3WVdshlKJj34YBRExhECsFOUYKBcnVxks+CxWgazpH10TuPHD
F9QCbF5rPHV2vU7gq/u0PtBeA/QUEWaLg27Fnk0ESI4g4NEXG4bPw/hyCp4w2k0j9vZe6wUnkqWu
ubqjUQDJRfu+zaDwZ1bi3ilut/tuwt9fL/Xjq5/JyvAzOtEGuZEIt436dhveYld1SmqP16ed2FIh
Jn6Wu3+pOZJXSLrKcWP46HtieELSD/my8xPlrQ0xckQD2/pydT4zA98E/eOxduG7oHtFs2o5ipku
eyFiVNfpqhQLItPExifuuQFSdNp1r3uDHSTMZT9nNInrkQQLbawiQ7dx1FuzPHN8JtOOfqcG4/RB
HRY3Y2ieMEYHlq3HrpwmMXB6l3jXg6+BFUfm2B+RVpVse8CtzO+yKWaQ53CwSoD0s9w3a4tJKZJk
u6p9KEU9HoDJ13Lh5Zv+4eRw86+Y35/77+LVHjewjVQDpA/GHLCS9GZz68f1wrWdRQPWq4IVR445
+2b+6rO7Pf3rPhGSsicjEKAr4dqbqkN/2rvHY/Xsph+ZuofdUmIv9LzHya+1IlhukoYaG52QAMyW
esrvIlWNioMbMmwfAn9nZ1Ih3ETyswG67sCitGIQDE1DZXAEH/orOOjdDp/zJMez1dP5F13eJBlX
Kz8pPJirUck5ByMXciEYJlAxadNaWtuWJAs4fEjEPwnCW83wn9+e1cr1hxJetaRP79zWXoKTn+Tr
mUiSUl/tgal8X1joyeveLcOH+4USyeSjIHX30TpTbrzBwTNFC17odujGAXQK6qLDJ2Tw045ZPrTk
3aZs0LqlWAPW5cBaZ/SBAtPyCk/wqeQgpBlAOMZFmBQS4LwpWgW2KF/Z48a3pXT9tsbCFl6eSdUS
AOxWsJG+PFFGajyW6FzZIAyoRW1nJYoIQk3dBDcJY1GW8oyd6MbPJzJhCJWymKHutVVIJe1suzR8
UCcfn6BBFO+gqDp2TzJ4rx90aiMWmdk0wcZyEkyc/dHCBh7FmAsWU4hf/8jVTKEGcVEXaV3gb+7S
7Mg+jWcUeNUZzmDn5rttfpj+uUxeoaBPWGtDAqM671LC+KiLNO6iK8VQx9D2YAOcSV2ymBZ17XDP
ZTq6uFniycdmZYFCupg7R5D9Rn4sSDraDc7dHirf3EQEPhgRfWLHPalzlxt1MQm7osCEqV55bVdh
+0FH/l2oHASFA2HpMpQxJKwyGHscaAH6OuMLp2Z1BOrLOgm//CtJNUsgj9VUIHlFlh2Sy7i9z8uQ
uXGco7hyRIvOw9tV/DMH4EJTKUyf8nzkfXgEWExIlmPr2AlDJ8JjnqsP5iYCFlI2mA3tmmtb3GiR
G/K54CLcV5s+IrP/L9yQxcb7Jumeho8OBGZjHXpaefROVKuhPkC9HYgMBwUbzoTvk9ZSoAF8vDsk
P8Cdt99QlkV44iRnVMrtaOCMaQNtrn0m3Yv0c4vEJfoa9SJcJVt5uKnFPv0vE3B5HTmOmSrQ7hHC
r9wWLzEKb6MGJN4mB/Qy2Bjp2y7/m1habnzyDjGuZcccjD/K0v+QfCjUKO4Gt6posUjoJztbgc07
H1pzc4kFLXJ4N/CgEahoSqEuO4f74/5PJ+3YrwmOcdsb5fD4hMReIbFZuVupdkpvdfjPnQkyaq6o
H7+CrI2kk/lZ6zYw5YVFUD2QxkR0NzWBWckH5M+E733x81z6TFYQxkGbUPAjYlSZZW29151mCzk1
jw/iS7PnhLArrnT9ZRGcndxzVRUqGSzyuJ8CQLO5H+zsaF8ElJb3vNq09FjD0hSev8dZrZWnCkwA
eBq8VfZ2LLVXetwbtOfo3vr1XiOAvH/RQiDqq3hy0ZLzutCP9FuDdkb1beVEKDC4EIOo1P30p3fo
CygSNkL0gSZxSE5s9EYglp2LJG6ENxzvxIqb7I4qaWAb7de8io9ltWs+FcfS28wbme5x9eSTnTTh
/wfEQSR1B87AAgFS70SzF6Vcz1b9Cg0cBUrtPnYeeAZuEH9UKyMZG4ITwxFW034NfPthlZnxnMVP
ehn7TS6fsMRdTCGiHmwYeJlTpRATXlnlMmQiqOV72lJpXqBoHK1okUkUrpPrtnacio/tZsY9KLz5
ze9KLNfM8G+7WUuRtUFpkySTgvrr9oCCTxxdrnBvrh066i2sVIqVENRsA2Sssf9p18zsZDIeaY9a
YuB83img8yPqSY6lJ1CQx/g6/7kbak8IckaZJxttxyBjJoqk72Y2trLE/NZf024zOJlbsc1l01Rw
sDHGPcOk5YpvNSIBOpCRqHsOWKZMHobqk0ttjM6SJuRRKz2yqJcp0HXFBtc2zRS8djeWAE4xHRyC
GkU9/QJJzUl3NWjgVxXBPd+Etn3z97BbI9JTuGeYAvaemgOqwwF9UGOqEgxqDWuupHdFhREQN2nT
nHnIQ0yCLUKo/vkKSR1mvMZ4sg5vsJee5f/rPlPff3kTOkanUq7bjQD0Gr0bQVWnfklDXvwDL5mU
YpuM7bsZbBmXNpN8t6c2mOKriMB7Ll4aUAQ09n6u5Xpp2xiDH7Q+vdjpbZb3evVapf74PK2zmNuL
Q6E04cYx6tcZ6YYI2as0e2lWrpIkBzhsbOH9SJJfQJrJMGb6ezycZJuN+4YoT7kfX3SuJeE+z4bf
GOy+mOO354aDz+Fybxpvm5+fyztwYjz9H4u35ZeHbUUzbbPt7Kn6+oLeb3RjdTFvQdS20T9VJGcT
9JSBYtDYnAIA1tCALZuNgx6UeOocW7hec3F5NbEu7Qr9lZEE/Vxx9LShtNLxanA6shAVygSNpRBe
Hna9f4ijCaoAENpKTaHJ1pGP/cf6p2BzZD6DZEuIM2TzO309rdqBYpQ3CgSiPq+JFHWHucNgO8uv
51NnLxTShC6oUmsytnjozTx+Gea1h8cxe8U2GUNEcUQLuPfjh30CYtOav9zVLUx2hv8N/EW6I1mI
yeeY6QEEu+Xg5D7VEYo+mOWtTqz/Md7n0RByFFXHDr0Li2TXLo+q9tQlpRXbb/QsioKDu2ejrWGs
CuoBQvqVb7G0xWWnx1JblgvmoRoje5TDhxu0K4PfkzIRq9MTPufhSJ9Q+iBKyejvBs+6XmL6qgsN
XadUszBTYvL+UIKEaVj81QrWfxgeT1KxQSdtDMc9Kn1jdURLEDeqGSU8dZtGYOwqy5/r4QSkzNgt
z71/aF4dXXdR9k5hJgMcmnTS7LiMWnmMH6+jeSBUlOQQX4378pe5dnkO8cDPdes9WPChvSS9PaYt
0Fg2wca8c68O+kTLLpsy98npvn1GpkS0Z/4qczszquDtDKeV1sgs1YOGejJNHGerriLEJIVLm7c1
ojTU1WFVwmSKv4dPalFt5Pwb739rKE5BheFY9kDCdHg8wUnRpZajIZ1TeH1DoFlHhmetI+TNRqi5
+HgJmG2L3D6CqRdCHTfP9graBZv1IIw6OKFLlNnFRBE6qIEDmDUykFXV/Ac+XpNGnNR9180vQAVx
rItw3CeQdbomrldqFx2fDz/IcwoAiPpYj52gl9C19UGNktNVAeUWK5sbyphXouysp6uPswNupffs
6NbZGR40pYJpO7UkyavlC5H6AVn4trZ8EatR1Jyq698z5qYpJBIo8T6lvGai7brmnJUUdu2ZpMwi
TEbR8REN6B0GBw1mVz7qCMxm1cLbHIB8V1DBCKVjxjrhhdpRGg1oAxRVw0VXUazujAB634Om4n4l
7+VG7H9lAGwRNtiBOjZ//cW9A5ZGoCefiLOBVx/6gtzSN8wKtxHZhhm/Z4pnPkeOvhR64p2ZpDOD
0MBHGvc9TzGHLJ59h6tbFpQPTt0TzpTF6SMHV1vj/Kln3pasjc2CGVitjOa+mIx15E2SP86k+Vl0
7vnZYMfEWBVrFWpGNT3TJXAuxvYKZ0oReXUMjI0EtE2Z9I4H+Zh/gsJfnc8FIJA818LW+f7E34IP
dnR0fsh5lsIPy3IgBvCrFXA/iHrCA+lkoNqwyRQVpZJcUgGEVQOKivIbbrkErjpfNIGPXc2xz2HC
g5Pf9s3bwbGckD6xlBINphW5pb+IGuJNcxFVGSGzezXVmde1ZxrEt2v6Yw9VLV+8XahcpDy7xfp3
yQLQTHDGS0MbwUrfkvqCTOtamPk3/lxBlL9rjTWTxTAiAFEgeOV67jzYJ303Ra2iEqhdnRwrq0Dz
ZkHNJwneH0RRdkX5Uhkq6Swj0CX+YlJkuJ27j+Dqy4Tyw0B0x40B7yUWSBlPaQ0WxHnn12SGzgGk
kvTryF+qQ/9q4Ahzr0vWyNVTFsoSSwVod78VqxrIo69ju6stfdKvohXQ+K5HQN8JF0ghOxicYkK3
I50hZ+u0bM9RoW2N7SLkQTBltxr6J91QZLnZqIhwCn2dgwBiB/pCLIJzHOISBmi42SkxnxNnJrPi
cMNWJy69vahJYlYyjls0kcsKSf5dQF/l8hvmuJJH01l1zfrKaGnuJIAAXfAvynBKRa4lCoBpe/M7
gf4c/a/G1DrI4uVOzJ09mB4BVtuJSJ3SIF/wdFR3CIzCBsD3K0AaDnC34mKe5OY5lmwhgip9DNZy
IiL62Hm4NU5pUGWcXWUJP5d3suKXsROPdaPV5rDzqhcnYhKHTHahgvOur20S9epWQ6ibiE48avB7
krKzN/q/sXM3mH25Msn8gSRLJFpYUYX3Qjb4LF58E5oiQnmo6NLwt0e7Og3AkYjLQd7ajI94fcdN
iKwrh0cCjxT0GKCS6sVJPo8aZJik2pDck0r4kFPg8tkyxcbzLBHCr5EzsuPbVgVo7+LjbSJ0eWOm
LuzNLDYUS2IQVpMqv25pCkYtH2Lc2NDiFk4LcMyg4Wgr8sPW1N7FBRxif+bueCKlaVmOgoeppUra
oAOlxxL8cUs0EZsm4ojRMrXVewK15zz10OAx/rbSV3s88IutoRHe7JeV9d4P6nuhcDE1tzVGwMqY
LIOJV8UT8RPDcCDfGZq28YWugQh83gEGP/iQZGwlFH8t5LaAp4b2AdnfLoR7TQz7fLPEVrfHG6Q8
YB4iguF0LoNFaDbdy3PwoTwduCWcF/lhc4X01CKf73hNd4yS2UMCUiLuTOCXnrXox0m1pYP6LJpN
SAyARB/yEQgz/O12fpoYU39Me+5GVm+Pzo8rF8gfo1unZyENnawB9LTx3+lzS2V1EVzegk/DCsHd
rsHr5+gif/s6VOazUSRFUnRxl0V0r9mNwUYQf8Wgz0oiGAzFg3FxzvrtefJzfUvItqgPCyb97pdD
TExQxBVZglPMyVEsQZ7H4/XhldzspDBoVXjKaf9JXnzTHm7mUDVzq/H/g9//99KXzzFDUrj7wxh6
L+gzA5/xyv7YUZsO0XAuzPMUB6yP/5TKl8u/AHPDon/oUayIVtAqa2OMzD+hSRuQYt2F2hnLuP6a
IUvGjtDeGewhFE4CpKpwSVYVetvfpHTq/LUXFFHA381lUeNlJraPIE4K9ZyZh63kZQcBOlCDYBcn
OpkjyKq4FaugbnIqSJ+AzakoMV33r5b7wL4ZOuV+LPqQ0RAnvHxblEFYbIvaKxwezWxZnb4rvfL3
6QQjli6b1Fn/TiSCLfgIBrngQG2DJE5rAtNPXJZRCcBu/KIXfwDPmi3mAcq7hSK0ORIccL1iYoHj
neSCbQOcdoaiVu9HnzHa3RGxiakVO6+77lxjdtHYVtT2+u+ljtMTin14lGB5AXJQJTkJxtlSoLwH
4OIbDFcMZI4Xgire0XxsAJLoRXF7TPjy6b2wytunIEanqdiTlYr0hMyYrX5GlXSyWQ8G+kxMwGB5
bgXoClI4gB/3ChqizWDIF0gVj298D3fcOvm+JWFaR1ad9dEdhfxm7zENyO9Rm5UYpvgIutlqmiPC
Q3mHuBKGBO6TaIc44TcBGujgDcMRtlu4mW4LT9iALEfQJDxrdC0/obXy/JkSp0HPQIhqaSj4HvKw
yRGD9Mm3GeApOI2mF7aMM4YWYWU/1tgwPsfdvt4eK4c79FwP7t8ACVnYXJgwxRa3nBXVF4+AoB1t
3x/bkIM1vUN+ZD/gSStwu+83h5NW2c4T5i6nWYM1qNATwq4rowaXXsrj/MJQwLtXELRgKETwVn7B
+ctP6jQwwwpwlaPI/jpGIkggqlDQxJl5xrW7Sjxyd0IJwX3QyfUNsMDl01eQF1llyiRZu4PiQk6w
EobLFt/4oBegzoOoOtSUvzxLb5r07qtrayI121+ExsdNZ2zJzsl87pzK+fSJav9ZcEklm/LNoXFE
9u3bqwfGBU3EwaKIf0qVBMV441PdJTW0TD+ZfO2UcwNJsi7DeEof1fa7UCXamMbLCkB/JUYyU0AC
HhPjsujoEHKZEMNOY6ncXEIH13b0i5Jjv4BJievaJezthuPePiN44yn6mcAByaVSbE3K8De51Cnh
BHULbuIe8AonAl3hiJ6roebTMcHLUx22csXgJWaW4Rg5pvwEPWfcGBNij5z4+mVOvAWLBbwhBkSR
YjzXk50yU4FZIedWzIa4cYbFiMtSiARLkG/57u7OgvXUMCZ5bPmwNszMK4oWW0OgYkWJY1Cfa/e0
xlNOHavfk2NdDJ+N37XInYYxHpb/6pTj5hL1S8AeJohOG2F+JxvJ6pKuAJUaDww8h7X6cjtCRHkA
nyuXLYsOk6fiXcpBDSVOj9Aul3WLz4u2fMDGExFCrm2/8c6myl2KPxk754JQ4e0qo1LJoJy9vUgw
b5iU1IPMifk1tFUQBYpRcshZhVw3FVBV1dgPvbFKxO7kfjlMrM5NeBxfkMlxyQHR+XFecfOEqbTa
PGkjTZSYcDA28bLMhFwxFQe925YyVkf8cHRNdu3tkBZxDQdV6v56Gb5RmeiacbO80P2CqrDO88+S
dVFDvsUCAAgXqHJQ8hOBEjI1/QgAoyVU7aaXmkv9nlgaEqS8+yjjbXjD/Nj0y60AKHRskjQ7bISv
UehqVCH/dUpTpvkvR9D+9YjAori7uHFrTqS7FwOCXfiBBfeiab3UGVrI/Y8asJgYHDDGqFQxJgfB
oBa/gXWunmWcRbA89jD5fbc0kPbWjYr3U/2/aKL4aPD44vUfs1qQkH7oo/3HeB495JrUqcV/10nS
+vBnPgxnXhTTR1Noyl5nwpHXPv5/Y85liIztr//sBjh7rziaglpSo70mz4J5g6k+/wI/xjQF7Gmi
R8LzFg1Dsm+c21iQCbrh7lc2oSg5+BkSqsv8lJXKLbuo1hmL1tRQmXJ8sgkvrBnnoAV3O+od/TPU
3s41E8abYUVF/LK6lB8B/R/QG2z6Bv0YRV5s4ZxmcKWF7zexeVpabWOlLdaRVeK489rWpi69DaP6
8qLhd5K9IE48kIyUS8tROAzAnzWRT+5BNzJAYA5SEGYLwV3RYk8Pu+geFxEs1jNSZ6nUA/UIwifs
29nSElqMT2GdQJf68EpIqyOom7DJAUBm3EILppuF3JVv5iBbYDAHQbCfDcy86AmHIiQuFhmR67kz
piQtovEEVntzTj1qiZZkLk/7vyBGbf1xzAoApEr7UcJu/SzO5NYDbKmy+W/Q414ooODndD8gzZuX
lyHW7mi7ZbeUZQkoTSY87jlBYvsEaTVDkzxPm9s40u2rjW8rwiXCwptO9SbxUrLxBtVXUA6mc52Y
Z4vEu6Dh17uJKPBKmh06Uw2iO7dJr/CRmyUtIryxSwlCVAGyzv5GBgxzRoO4NFR1tLDxL0huJiod
WcwWwZjHAQ8ox0F/m6tjgAmipONw1L95weJAC20Tds+oyFIrfO19IQVfnpulurGq6Qd2e7iGZf8r
I9HiCBbNtx71lbsOf/DKNE0DtWOWl8oEhgdsLg4Ou5czERYTXjyemz1dU4nW8qQmVSXpNhhy2+UF
y3BbQpdldn/y5jrDSuhUFT5Fbw6+gUwX1aO9332kECkI5b/bR3A49OjtYwE1dmi6zBJb8QUyiW6q
ATtCHcp8YO8Xinl6h0fuad78+v56fgHnd9qUj6iVfqhDESy+8/7ofhL2ic1gkFRdKCI4a0kMSbwz
xTv6esdxp+yG3jzGMm4sXA5SEaHkuIgUrdmh9zEWB656BqdzFYbZ28GnF00tBpuM8fLr8krkoY8J
JUwu+jWvoRW7bIwXSZ5VgT0iFQEg/D54P5OXg7OHUOkuDqrFydMWNiKsZT6aHqfeaRaVOmIc6+kc
KLjHXNIgqyPpnL4SlJbQog58xsH7G6Ty2S7rnQxylEWYtQxmUdXcQEiafa7LAshFLCj9ynADjVUB
PY3zIe40D2lO8Th8wRwd24iv6sNm2dRyqe9jTFrLJvboU5UQM4gEbHv5XG8Yex6bbPCZsYTZIb2Y
Ta+ElWjz/s3PQffrq+Je4X3V/6pPnkKeTSAE4UZ6Hg2uE5G+c9ZxbUhnnFEaIAusmvXhXSoMOuqX
fJ0kJzlHL0nsYuBP28GTaORXxMlosGcUxmhtiV/Vkeeo923ajxOhRwmafty8VfK9lRFhDm3xIEOR
ZVq6DwmhTHfznQWK8uGNTnKg+NoE7kHpKJSWzxMtsj+sVoN0fggYcxbpvrukClm5RM9g9ADlv89Q
C6Lf0vy7O5gcdgpMT5ufX5p0kpgFkofEah3w6jtpdmIVOPho7WLZGOSQoyvKu+YXuy00bmx1qKM6
QebgaT78IvEXW8+oAYRBsr4TFTjVNDrsAXFd6j01IefyWjgyFv3BOvQj+3psbxc/7UU13+z4pGVe
vHyv20lFNGY68Yvs8GfwllchkxY8GYIzUV+d+hg2bK71SMDfZJirYb3Jgzb+TaB3PN9tdbKFnKRc
N+keAHLrtB3SqJaJG9b+07Ziiyf7gVw6YPVPNQBB5NzvN6vZBzfeh03YgB260ll26gCUAI10bONh
0MbBXcCayE/wLyCSWWQ1P4EYj0Y+hk3D23HQxPz/bbJWNDovxn30wS3sGIgXgNZI8SglJnDXZPWT
U1c41m8wnpt/qJlpcG6ALCq1DR0ulr2SRMRontlAxBxjDkwMMlvBj1RdFLEfjJ2zn3D9KJw/lNRd
MjyK2YFGy2sgaNQbKxP5nVPoDgXpEbkp6Z8YJOJpRT2z5yPmZeS9joElpbxFEbKPjfkbpYSWR7UU
dOGqOIQW4jkeghwFAW61AMfVZ/Pu0SuQI1zetaQM4oZ8i6eOIzN9dPHBzZms2Dg3VkdNG1J7Hblx
FIP8vD6anxm4ACzDGCc1vAoHfEtcks+/87GZOnxOd8Q5kWhHTv+KroYh+beAmQU6IG/VchQz5hd3
AQ/YTwiInpiXyg1AjRURfBACpoiW5FV5jBJfmXvPVtRWXMScMxQmkaenJy/UbUrmh5ZGhogQ05+C
3BQccGPG2qVFzoaYxSzPcd0ozN5R0TnBtC1MzrM2QujfbqpLWtbOvXqFUrQbs1epoBaERrUiMUJ2
q6xjvhRptSt3/oK9WZJ4KoDqrA8Vjf28J6RKm9fFZlYeiIUm9vSmIC09kiF9JH9Vq54KkVfNNyD6
46nyNG0QWErpj5dw0LH2iOD1tNtxZL7eeNhWwaTap9ZuEv8ZY5UHJS1zuD8O0CvdEMvjaEEjri0j
p04L7X/+99mti9GMZ1n+uLpQTIn/N25PGOYEXoo4KrfOYYO6IVzLqqCp2hP+UdLZSwenDTjiYSdF
vma6I40dSsXLXDB5mLwERoQHAaTmZ2Mab9GDsKKhDZ+em1Flam3m9am0vBmDd0Q8MKo/pEcoFk5D
z/ERRpdGlADgyZpie9rguACVYUifdOIwxT07+r8NFRp+R9Y/yC0L8fcBgd0xmOIdj2eMZyCmBfgx
DDYzEqsH/hlvi08Ri9utxlRuW+e/p3l9+Zy3zaRAmMtEpDMQHDnc1Y9ilGzK1V5SWZxKaZwYI1E1
jx3vWJ6urHBG3UQOTvQ4mQyRj+si+dn2ae7I84Kfe96e+OLfotvrSlSoarzP14F60FtBhMKmXpqF
Ej739E46gNUgeBnFOziJ/i0osphQwAppg8YcKqnPBUGdcGTQEDytzIAz9fUADhufCuhRADWkLA+2
0HzAoOSs/U3FuqLnRY+nvK9qApSj028X6lfac6Zg2Zagtz+cBkGxLqU+0GX6J0kOb+Ult4Q5Uff2
jiAepwgL7rfFJdlO/UFIIHFn9fQ7oEcFkkH3WEB8pOWLhCnkNfZQiqOHn7RHs9sAcAqrTKMCghR7
aS9bW2zaYd1iZJLw9ScgHA26PL6nlStNynSokUnKS9x6TIboJk+yB9SBU/46uDNe9jkowIAA0MLs
UFfrakwVPWStWpkbW3y1kaUDLiO6FL/1Qhg3zfeUxjONNYYJxdKNQZJfEFIFD7Ge+4YE2Ibt+nJR
FX/JxtAz/dGbDtDawarsEmvd1dUcihH8HAPAaLC2/VxGY/Q/JXUct9Y9rmRvrZhFqv6YJJkL1vW5
f7ga8hyjtNf0HNIwamhr0PtH7yFnvK13Vupn77NrF9cJaDlwX1dn0PQkSCa+T7VrfgdY2Pu/bI9k
eRcCD9G0hmPgPNgC7TubJxfqW8FAfetyiezwn+CfiAaj8cNK0c7cxOCWdV+4FBCXl0I9mXDpNTsZ
YCtDT4NmDbPe00pLC5RIgZ8Xi0X+H4Q42YpnEPTuB8qrdLRk2pTlRKFJQAmcAWR/u6f9MHfsUhna
MZpiCOXatST4EsNq2QxBt4Yuyv0ZmfBJOuPQLiVLnpgLkEL07UIqoI3xxztcK4lyWQNqbdV3Mfja
id+GXrl1a3YKDkmYEoSRXp443cnf1+5kBb89oF3iL7HEj3FEtkPj4cjZvigHjm9rSqN7Du2+agDO
K2jjqf5PF31ZWvq7/7PcpUA2gKWus1IpwQkbBTaZbEsRgMzlHez5XrfQLXqWGcOGxY+dExbWPsg5
u1GXFQsIVtU03wJ4VA5kPrRXsZncbo8YFOhcA8YXQ7FGNHPqHp9j0FmufsJDbEBc9esyfO4VGlAF
KgNujWsAv/8SgB0BgStPcygAgv2rwo3VId/tK7K6rXi7DJlNvNBMLGOFxPGhtawWEeUIEuOygCyz
EctLmfhpV4BdPMZers3s4lrLqyEC91gKFhADhqilRbnNjBFYAOgxsu6NmKl/KhzWlYCUbmv5o/ad
o2v4K/HLfkumLiqQpLMQXR8P1gVEqcTWFc56Ev0S4odi8t46dM+775uU6KF4QAoUebzW4IL0fDz9
5b1fGa62sO1+EpfdeZPqd+ya+cAbnyKq6HcgQ1ujmvCR/aqPtR/3iINIvVS80Ht1ZNOdb6FSTOMZ
TJVsjW31GmSVXpbTdDooYoad2RPOfn4eM++w5hAgTiNsNae6BYjHA7XP+E9SfZ3lo+xZ4HZgvnPc
1W3lCMcMKN9xFPydDArVT9oeXUp6lhhBQGRVQpk7lbBkNpYsnv4TX7AXVijL3JCQ0RffDbHTvgAt
yKCYIP8Gg/o3QBqez4QXNA0UCNdLBjN6Fju/zRd3UPumnuG1ulUsm8dOpUv8hYSszOkmmvPG7Zgz
ATqLij6B9UF5MldkZ21QBJdCvaIQGkgHgbvSGMWMuQ6z6LLqScIF15IvA8KYVkkW912bsRlVSHGL
2MVwR+8kjJ3dX4recRjEq6w6AmZwYzhno+oPhS7VwwnVwpSeqaQUbAdBfvoswfVEtxwzWaXP8RyZ
vOYbv4TLc2fItE99x6XIg//Vd2WDUwnCqRpMIq7L+GD1+3U6oVFxCbAb2dw3PMRcbK+gvINZM196
YiLYaDHbFLKXalrxSdQwilIazBzZ/1tSECfemxKspJrvcKW2Cfvo0ZvwZX6YomDv75JknEoEBIBS
YCXPUTHas2593naFZqBODvFlxam20evV/xN1OltQ3EibbnL6oywaCSe2u+P0/D9fE4Bcq7BxsCIK
Lycax0t5Ic0r23HHxBC2TudWOHU8AeVvkIj76F8wuOyec60DQDewXZ/nYfV4Avb8hGRRxsAESB5u
anN0vK+Gmwlj/6rSf/P5eOQnNDiRrOWwwaVX92K4T9IVP6utaRvhjjA47Ms9kN9UGUn9+dhk4s5+
LygdZDMnmkZYcR6Tw2BY257pc9PkeETlcr420iAoPCqHU4+BmP7SQspDh4MHhdmmnF2TaOt+hcQc
L66yjXnnSs8/H6mlmYnsmDucwahcsx2LxlX+1cNUgTykiQFYQsZ8++n4MG2D9AIQPrHevidmkmbj
bmVw9nTZAJSQAHJTbLZh/GMsOLyNRAOhc3bULkZ32F2QZRdckzp3qSJ2ttK07o2/3EFw8kr0zsMz
AcSfV7dSpa8DhtAt3pMZ1xShN9m/CgPHHxPl8XMb4rhlTX8yc2VPCSjBa8xzWBr5qE1mMGjMBPLf
XA0Qian1kOz3RGCuBcRLuyRrzOR6jS8Q0DRn/48uoFOkpfGWBbSvjhg/o4xcAfpAkpcjxoykMB82
yaVKxevinvQl80gXOlZWlRELl5ysDT2b8hE8YMBWQ8FXpFcRm3JsqsQJWdYV4+2Iab1r7mPrRoZb
TTA2QsuMZrqKrCl06GKf1YxABCFDM/6XR0ZOWC7fE/Ta/YOPaY20eHe+dkCyM/qxn4oOgEzcqSY+
+uSlQew00bYy36M5RTU38c33ei68XvSXl/W42l8snvUxOd+4VhAO0xlP3A9zm3+r+wEq2Pu/WVSm
LNVtxbBPemhwSM0coQM/SjYXZg/Ff3iMmn8xy166QVG1v4SvFaXe/L1XxDHIEmox9n6VkHzuMt/m
1Pg33iIelT2TiF9l6K0b95hHbdSfGzEsebOx4AdOFDHScnt+lgvVx2xmD+e2zuIpUx2x+pfkaW4q
StW76DsrDjedVW9x/Xohbj0ekaStffZH/BcWzVYUnfgaS2fjTV80rH/3tF+PMB6x+jeVkmaDA4Sm
fLSfDrifNEVI0Z7o0ZbtIn7truHbSldIB7dMHASjP0gLsfHXcih9NwRfYsF2I2SBpciy49haiaWd
BW9iWNUkf2I8KkjtvS1JXd+SDhp47nT4eZCeQWGNrle9ZnSLG4ppdO//1auE50RXhIF8/cZDIoqm
paqKa8eGXa0LGIxAHeWynLYTsnlET+bBaOJkMy5U5yRzt+WS4jztnz5reo+SvpP5Qe+KiJ0NXo+A
k6lnasyrtxD6iUs2FYVHp2Zsxiz2egoLLZ+mLPW2SCDlT7QSX3FJioKNEprxqfyOyrxYqj2CRTqk
pqI0+qasBDKRfWLm2TN/L+kfa+U+AdGIoowcgJFpMsjxwFDEzOso7cIN3HkWzlcjgxK/1gjtt+Av
B9xlGwePu1QxasnNb+eHlTd0aVJXBzNTHBI4yypo7M10HMviaJ9b5JdhZh25SLKEU9hlm8DCAAmf
i76RyakC80SUU4woxpBqB5lxjpP+Uh09kdYSYghNmQr75x+rudwYTjKj9cFWjv0Jwc2eALzxaHBk
XczsizKp72LoQdFT/LQGUV7opP4sG9PtwFhOjL82m4qJ3rbQToyeM4ELRcbbGWTVv/RF5ry/rRYg
EYaOKG2Yjsr070fSv3MYycC04gVirQzQEdJCC1vykDJi+kNK9INDKRDfz53E2yJIjYRq9qFYKgQX
vom4bk7tuTmv3epn5z4rsu0pwdw8EXRxi5P2m/MX1apvrbU/qKrxZ6d+xAgxzn0gd09o8Txh9EL5
fqv5tcnyC0NIb+YUBKJHZuN3cd5383Bu+WiytPnuo4zD2LbRVKRqAYNekxFtrlD14FA+ftNQzyu3
JdfG/l3OXtBtXS4TXFumcrG2qX6Ljg8W0Qwowb9o3DvvZkGx6yPSWSdUuAQu5xpNyy5iCQMw7MPX
AlFaj0RyBlmLgxstLhTsSiJQlFM/uReX/Ds+0mfxT3F7XdsAN+tYKBkuPDjE7zWYt8cW7ITH3t1S
weOZ6rb/qYfPHEYnBiEI0bF2t5CcJCxemjIlY+EsdTlkAZ8RSRQRtXIm1WvlHnIapZOyhP7I6vLQ
eoqWrUQEZse/FbgwRuW/5941GApOOio5FOfawHz0oXkF5be6qi6sEo2a2i8ERBPMQNYIw1zy8cWH
PJ+5HkOJR3VcA0MycNYR0du6TlDjidsWJb6NQk4HfLro6TheXTmAmgbAC3BrJX313OxohA52FaAP
2bQ//a3iYFG0MtRDjuSLgIdRFrBolMFned5YQbghM886sL2QFSMCgNI9fRIX5zbBUefJY2owwMaV
5viyudiw3mkIvlzrKWKQjTXP+T50QRj7+FSprDauMm2zQjJWMU8rnW0q1729mrBofdTs6VYWMyZp
QFfuZhQ+VgQcYdRzAtxfe4rXdv5XrYreTON3w4LAlduPl550f9dGQBh26fAIxH7vINBctA6PN89G
5KDr/LM6EwnDW0/vlYldAHQd0zbuKz/41dO5cd3nlocdA0LPwONYUI8O6Z5D1uUM9PgvomXpENR9
71+m7RMJMp33JFGewKmPdbiO3FTTxbO4yQlwvcKXyUiwLoWdhikRKDdzUum+59u4Bnt3Fu6W94fv
JruTn6f/Gnw4fgOp1Z555FkfjzO5rgxFrSXHHaJrkueIyWEUC8gjaKbFhKxrcnIII2/lQ+AHj7fl
40gAn/1kL9NqUzg2NJRoAabPZnMeAxR9ovbVMLwvgAEPE8cOxK/O0s+EcMGi0zcog5tCUtyYl8dS
4Q6ffudoC6gN0RyeR3U28/uksJJ2PbMES3YeuKof/cQBw+JUPEOmpVWh0j+BKsI6vNGRrdaqHMaw
T2ACSxNW9CmPU7mmZKBAYQAl+j1YOZYmbL83mtL77DcyNPr14x5+1QmEsYfGeadASDFfirqJNfRj
s+HkzhjOV+12y+rFlBbHYN32dlrf9QtGd0l5cPyE4cVllYdNXNDU6wnih74b4V6p4O3Sr5hC3UZK
EY+sk4xPBcVdnDUXXY+EWYP5xDqvzIvAJtZ1S0rI2LyzuCD0H03sqe6HilDT1qoGXWqQT+orbDJY
6w+fWMV3gsqZGvanzMGy182gHfeNPVAf7il13I3y1e7g6YJwfhF6cRQ/S1Rp+tYtyIi8+Yt1Ea40
fRBklIMuZjdcTrngi55zKmLUcH5VJgtANq/MAcJw0Zwm6n4W34vWXPqwpmpQwoOkyhO08vJIn2Mm
nbkdFXOgoVGE4KQTMms+j2AXUBBMQUi0xj6PV5t6VEDa/74S2lEMLyVs/yPbt1mvn7Eghkz+o8TE
wmaStgha9Sq8Yed9vy+pndYDOmO9nTnkI1qFofIWobdnsPUsXF4x0+aJRBBOiiQmluEZqVHoN6HL
qznUYOcG2cAVbS7UPYajPzHt8KWAN9uB8k2c7Gd4GKkVN9a2NaEqE20rRxF8kML/2ipVH6TnqaVi
zRdUA6gBnpL4FFOl3izvyxHcWTtsZc/k/vGu7s9cU9NRLPOofl6xhV42Lfk0ucWQBIbwbu1HAbou
eHDq4CbRogJDGSC/zB9ttxBCopmmxRFspPmQk24xWChNiUm2WC14HdKBb1GbuBzaryeZczmindvw
12DjJCUWOiRqGSeLV7IkkPanKO7x0s1xfEpJN8OB0dBiRTFBhZXz1YA5Cju+UH0op06xdlShM/jk
7+He0rjzPsVwdFyMTbJXj5RoVEnyhf3fArtV3Yfx/lfRGPrYjHnM8A8yR5KDb0IMTDx8+IT+46r7
wKUKQDRYFf/4rMcEymrOq2kOkcAetqzq/pIeGTAP4VEe39T8kb6mxXV1cGufZRQ0qVsKxJf9ykXx
XA4oSyVHCTgi6IMFB9PGzHUywUfZJGtMEgKb9q5IapA68sZtwfYtQJsUSnj07bvjbDmWYSUSVSgg
7Eh1mvkM+83kmFeihhCNaeR63Z7qY7t5F5cGjWEL/Ca1Lj+HrjArO8kuIWITSt3utJkLprdmhXb/
zOGhms55xniClyvgnnbva0oj+aeD32I0ABbU08MD9OseRTMJMlbZX5V7eTW85ERd7WLjF0HTTIqs
s1kJ/f/713DSyva0wqxKw2VzfY3Yy23GJvgqR2j1V1B3dkJLA47mrnfT5p+dqeH82Op2H1rMe1yJ
uKiq3LD4oKUM/sNKRr/zcVHAALLRZBQd8OSkjuxaAJ5L8ciAMF+h1dyLaKAlTueZ0vT+jpIww8cb
PnsZXsJNKfPl20CNUmcx8teKLZ3wMZ4vDuEj52Xk34mTqY5qyj8wWOU3f+Zl1MLTzXIbqQvfItdR
OAPPDmyTlV+fJvjrDpbDJQlm8PlldK8IUBP+YAQdNsFxbDex+dXoTmkMYUYGTP0ERb36qdsmOuUR
viDPlYoDyiX8FRKnYMa5bJlH+ewLcgMWvcqMP60lym7VKibo+KtcAUKfNzn4vEGomoAh4VP6pRtU
6gXVtJsYhrC7zJhJJH1IkxAXe+gb67EqO9bZNSn3KRTOwjjuvxCz2ceh44mCBc3OdITw1KWu2Abo
KS+xyYG7MYUZsExq4AL3hzwHtOTV9XlllrOmBUSKGmMOJ0oJ27xSWKJE3Whw95qqcLqwshLORdDW
m2emwhhdw8Uc+2A0neiqAdLSYdvKjel0VPBsUIfh6xrmGiBm2gEXlcEb7cERO2xr/XETLe2OxUgS
/rYJ/CZ1Hx2hcYvtz89Gy5XytvGY1bYbOE8mpcdy9Qop78OyE55hsMUsYhrcKq35kYLoRfoZFwSb
lyT4txr4udKjyaKzBlZVEgfQtIiXRcDnpmRJt7MM8RpzoLRvQw4Jv+ICkhFDVOIhXtoR5kMp0+d5
vZBBbwD9QXD8xvYA9t9ELI3Y7RSMImglA9lELoMHqocjmRbjjgFNYZKmPp4onHhkcAjWL8xmNzGA
DO//i0Q8bx5CO4jxPyY5XYwsblKDd5qoUC8SP87VH3/e3AIO9K3nRpGkUzs4TjwZmb28lVriLMMc
GzBrc3TGxOzw7Gbj2aBXU3mu2uVjJ/YdCpjrTTwIXa8Ga27kTeCIKNnTSsYOx0ZXyH2He+meQeSq
7A4L3ox0oBZcdLws8KjXTBmDl7jsZ+drt/DYA2ZB5O157R15UvtRrUEb4Tt33zNh2xC4In/aCmG0
/10psrJjF5jVqNLZSdvjNXT1FzHTm3yuhK7q09MJM5c221xkCN/3jLHKxkUhAoRRJy+r7DKGg4F9
xsXgf39GZG8VC0x1YSb+7VaVb1Im57c4YF9qHww/WBQcQkhADi4PJtE8h+Ugy/Mhjq7uhwdqcFsD
WheGUDZMrpo8CbXZcmcahZwt4stC49NXBziLIf4idB9loq8NoZTI/JFuWYfUBIZfq/SHUbZGahqo
0d9bdXNkFJ98eW28/2sp7/O3EcVAnJq8/RFf+4llSlOyOLDe3FhdIOPV0WTaiJ/UgXcxBIAdMUGh
evfnfzbaN7QaIOaIkYJ55GWEzVXmkZvqeQSCzOJpOXgF/0xmLgj6FGrJ4MpcSkbpZcCqII17T5Ky
dhPs7F0j7Bpvv7v8zk6n/V8ZILCfzUx26LD3GIrIDIhD20GS5o2D/6f+tbfT4VO2T56xY1FQTRso
VcV7z8dEuz2aAOM3KEjfjwRoO4zA0+5HQQ0DLo4w7jpuZ65MUWgIldEDuwTIZxeil6TM7b8E4Xl5
+/vnsYVdlx5c1/ZFlywMB4LV9YT9sc+AfRtmXW6V28NN5nv1KJvXr38vNbW9qMaJZ62xbtY/OgWm
1TV254MMTwLqyBZna9wiWaYZ6k3TqyB2QUapYj/GqVKz3292eisThC6u0L+lUKzaNoPblovPfcax
R6+avMS4oFQVuCJlyR9DY+S5aEonOQmCKzDkh/8iuzJW5BLMY94+NPIP/BWh1QgIbtvkWP8g9FFT
+fwao3aAa5ZwVvjmJLLWOOQiM8ntp4MzhJ3PE37dfzUyau7UmuW0xFjhqzYgXmwyeSuU9avQOU66
Ed8sigcrjasZCHP6mmn0EPVShBpKNF5VpGrw6Vi5r8XrIo2dE/rz41HgElbbhSnmn/5EUaMpkaTH
0xJCxpHqgD9CgLUeFtUaFLhgaR1+oJUp6uW1e2ejTPsQTbiQZuU26NycfvRvRXnEOq2pZIeJr2T2
1hp4cChWuiadJf6MnyR2PS7Xx2za4/NLjIKpyk+JcOmwP4Z+rpYST6IrxgWm8ZHFHXJg4y8GLvaa
vZAzIjZsykJSE8+PKVaB6A27kgUELoxWN56OCgLbCtLksC3F1bRVBNN1aBwSLGSp90jbm5zm1mbt
VZ1+iPmwuQV9PVCoG73gbzVsmrYOt845N3ZxfqI5COcyRnRjfBeK7M7w4Lq7BzJUZoI8OM4+pcZy
Bx4LJ/VpaepIrRjC1XOVajquARzLV7oBPrfKqIbW/evgpndlXNPdw60uqNEeXyJwRWswMzrk+XBf
PjHKhCzW2Xr4XQe9kgCBqDQeZJ+/v0P22ZaVYQhunnLQmi2dz8ZKfMzejfA44zMKHNQpj4mH20sB
1esMiu4s1vRQWHMEXJmKQsJ53Zapux/cQbLkfBcCj+t/ST4rZ714KZ6/Pmu6dApVJlhzpeK8WAcS
VQepHFPRPmIDgzNMS7Hfb7FEC4eWT71loFza37gWaLFoa3AbO+OK5a/32Q9cnDZO8QmESPeqcDsW
GvWkTXCrAH8f+BShxlunEljjVfAuNBxxvYTb7KAOKJM98jgA+9Fp95+mAQ62s8FOTPuXvt5SHhSk
w8ZhmnEGEknNO1RiTKO4qNv1sgzLkwB9l2MHs0nNuuekqW38tPy9MBW4vAU5MucIUh7wf49tpHdH
uiqR8pFxGgghMknUWAA2N9TBSIJZnAj7My81JJXFkwcbPwGFhLYBc73guNgxD06EX7t4WSCweaUa
NDftuWxX5ywtNOvulN9bgwRgvVqq3go5AgrXVxoQOEbIdh6rtcBieMoJfN6Iz8LUILMA4T0+20Bo
dEuGrXDTcYWt6ao+hXY8PucQ0hYTiVMwZ1uxoieKFYmWjtGro2s64O2VoX6MoPKCewuG2AGi/fi2
rwq30JQhhkoUIWkTfTP8fDuqSSyk0F75BzTER6Ogq59jjreXQYIhoKoPc6YzW6Q2XCI4G6Gw3M36
MF1cjzaIG3CwQPLjLtpJvI8oAwI1aHb2vf712DFCuv8kZJHZYzwhjMbYdh1PE6IHMgTHsDNfTDgk
aNCtoK7MEMc+5XOrIc/oWND+QCxkrgXq78vc6F0lRsDBrKKWtVPt9hFByyKUsWw2PdTIO2VpiV84
p8u0J5rAja87qes5d58JRV6uyJQSqJvlK1xCWb4DMcYMdgdx5LnjonzHrEdWjaGrOAHJF9HgfxIl
f3OWKXZroYSNPvM2NqR5tAUT8tpT74x7ZkMCB/UAFqlzsq5z0+7ijJY3fGUvKQPG0WBFVo14T5s+
C0b/d1luHQnryYarFi8VUpFiZnekLbNlw08Z26POU+tLmwQQPyxl4ER/9FN+cN/TD4E9mrP7mqRM
azY9DmnY6oWVsfiA1r00Ze6R6VF8XhVNeVqbE+vw/00K/Z7LfXaamT2DeYIhMi5m2uBXBRpHBzVN
ggCs+ctyeLOUahFOlrPlFHL1lI1DIBedLi+5C2hCpVxhAGtIUM0Bq2P4KQqXxNKL84SeEAUHevsW
L5YyLysxUqlVn8wKKJmmq/uZLJfiudOeSzLadkUBhQ56jrmtSBHqLWj2YrovN4r/YAHwzue0YNUY
NkwIXn4s7rZlBqbyLEZDxeUZspOPFx80AXW97lF6JbUYiC7hrttOwOPDTyvbe8PoFBckJMFTJZuD
DiQy7zGH8F0saI4O4fNiF96P92wxCEyYzXRbC/AOdVVOGIiilyrRyk2MwPhUr2rKmoeHUy2v5BHR
f6oFZRiWmqZdfBplWw8F3MHPOrsvAi6PygEXsfRfa3VL5Qmq7IG/Ze3t7eBhggoZ3UCvU90FvYwY
9PRY7NEukQvcRW6wiHMx2a+hlPNsUpAn4EviTRnjosoW+bToL+L2MkvAv5V+qLptzeNqceEjbIcK
KCe/1jxWAKqY+JtxfVciH6kLPfZ8CMBvxDcnaWvvCqFNh3x5o/FfxnKuuwA5WkAUyWVdNop0aZcN
gv92vOcX40Zvul0RzxNuRBqn3f8rpVXKIoHHL1Qc+MBT05/UjShkmXFSlGxQNaJgYE33VQcfrRqa
bshN8yYA2nPlj8I/CHfEX0PeEWQ4x8GNEg8iPpiRtaqde9qcIhkEnOi1iQdXCRSCWy5GHUThlSu2
vcVXxQe7nleqPwACOJxTPuyd+NKbCUq0sPJMUAwHM4gUsae/ZI+Jzei8/iFtx0yNZPum0RXucJIp
0NtqHQRbado+2KDnO9FccS0q7tfC8eUVNC6I3K1KaLHlXpHLYvuL9taxRnbFVB9VGivt8ZPt+xiS
GM/HlXHKE/iViFs3hHgKnVMfm60Xu7HVWi0qLUKyQslo3/v2Nx9rrigImormALoOBw+TP6trGI67
tenVgmU2J64N+37f7D4p4KZ/tF67WiLwJ4KX/mAxs9WrwopLfUyhnMHT0E3FOQ1aJaPkCevAff4A
42klSHqUjeZVBlldbJqW+EpVQnuO9X1N0Htfo7ZeHbeV91PTxXGrgVq4oZbgT49m5DNsBpCkc7TA
uIH4Al1s7ZDtoExJKY+1SdcBLLxeQ5+fqTRW974ZqcEIEMovEBRIzH4+RbcItxduM5lV8vwrYMbC
aKttWgr/bUEX3pQoRgGYDUt/4YKP+bNfH012yO1ENNB5+vNO5pT6hux+XAsgD7m/52uDDc4vcdx2
h0wuFSqdte9X+ip6h27tTesz2EJqfuVOgqzvH6m1pwmQj+qDjvEL58CcOEvqijPs/Jn0DSm3QsgZ
1ro7MXswnGK3Gc0RMNs/s0OQcFyDt55mlkSMf+XyB7PlwKKt/H/16EcxSCkSjoCcUl8YhrgLnUEk
XjzXLX9qhnoSMU1z4QoeOUEdNGNY+1FtYc3/6bClI8EiOp/1wIBqbbVitJS4EUhdSreA8rCMGpXq
gLgmzJ79wDdH4Zb+mRr1jcx8Tac4LFymAI9UOw6J0wH/pu8QRvS3YIgjUIGq8qdia0G58C/uXxOM
JLdHS7MmNxt6KXkFiqeFn46nbFDiP3w2QN1aqkz7n7hSq7o3168U6a6t4wyFCAjCwjOBkmSWFw3D
O7hqEou2KTfwG96Tumju5rjOxnlwg6N39C12GCE92YxyQ006dTdvGvVXH12Q8y/SsX8gklE8Qp9T
rgERQXipYvPyvwOn++HnQWNIYdnQ0cMjHSEhp7inrLMvabLYt37POyEjKzz16BmK/mNHmpcbK0p6
e/LSlT4Sq9ad/NW5lW9GwU3lD+5BhmqZE7cNOZyVat8l3iVpHH51YWfPHHgIkk5BEMj2ytKugea/
3Xbc+34gapXDnfThCdxrvM99SQll2ia0KbFQlvMtQqTfRl5SG/CEwHRsK/gZP5MKrOd+3Fe1eTgj
NA4yzv1/kgCbJZ4Bd7DM9gZ1fX/CAJSnSIhmXfgRYYDIkpVI50a/NUEhUbf2Zf7qKEa8xQK6wvR6
In24b4aOhPByq+vEt7l9xMfdPqP3jjoKrhztqcxAAcSaPZFJqlFm83sivPu1pL7zaqc3jyiP6QUF
EZ4N7lbmDvRLzWDzGYZPpLpZQZZF8RlIbUxLNsDi151KAsfog7yD6iCES5TQYr8KXG1nYnpJligO
cdRBudz7ah5+FCi/OP8DtzWqAI16FH4C699BLr4CAmsGpF+KrtVJfo4cWYQGWDGfy+2aVrSGRM1w
PjWipTr+m/P9Z8HvOz8+RVW7QKkasW3jcmS7r9eC789HbKJJpxZqmN3Fz5pTjAtxRcWybivymnK9
/LFXA50zqxHbpWYdtfSxVKoFjITB/+gceVQ2eTRQWfHt/T63EEOFWC8bRyXLeS0d3Bj/YQm/xopG
X+advxZJUJErZ0JvG7AZzWU6J6KZqWHCIGLIYg6x9QAEKGGLeY+0TEwpch+9e3EypYJW7UjwHcQR
NprGDtzbShz7IvCnZoT/NaIUDxuholHSpyHanUjvhIMgNH30mBwqgI7QCUw+Nn6a5Ifd3JwcjfHF
UQaxQNN0NcRwLDDFZI43vPlZLHoiurPjkxxuJQkfdcPURJmv4Tv1nZnreVYfmgeS0s/m2DnfSy1a
5Je85NYRZFdAmPyqI9XWmJRlyjWY6/zfTQkMrVBoQGQDiNhTlnWZdIvy+pu/PbBnmKAW3YTtPq3b
8Hn4cHltqMcGu6KpPDWBI5E3WqHQQ/tjzyGiADPfzOjgJ97Mtnsxl1BVVj2myGJTVzgHCH+AllKO
72VVkye+SmXE6+0zXCZkySrUd8/MQll8dQYkHr0mEDRBCRi6u3dNUh3CPUD8ny7E3vfNfaLrJeMc
/CfdeRb5shR2GupVLX8IQhs87aNylN7ELksJJa+H6+Wg/sZahasuUtWVxdixy9/6U9n1oXBj0j8v
kuhomCVRL02RNzkd5tBaDa9tOjx5kZ0SZkmLaDI2Y7mZjtJSwmnkyfB3EsN33cKy1IQCVNPd4Icq
8PODd9+A+QPVOCyvZxj1Bk3EwLagUFTj+db+zRIXWxbpEnDw5aJ4lwHhfrxXfXvjIIMJCnueu2mc
O5wbsIe5mpnbF1BBDQafRdaXBlcV5M37nhmf3pzCVQ6aJk9DHqryX5euekC1EPRi4u0pf5t9ACYi
AK+sRA/6fKtB4Ms7hCfvulgOF7dNIAo+jt4xxl4mEfdn0PTGUCr5BoEWRcxq5W4GdIneZCAJHbti
6mrbVifOYNzz/PXf8mBfZQw/mj4paI+bDEIudU4bDSdkFEi4ND9wsL3xnwx5a9Dv8K4rEuDQYZ00
BU2tLsmGuLdgep7b+W2ssSIBgpkGLO0arbip87kp6x9bfE89s0Y0NWV+6VZ5xR4vTUGpKa6fd2Bn
WneahIbZpOawWAXIc5G4uZ99np40VTMDxi6Oo7BC1P4ck7NaEea66ZbPfB6XON+U8cslXCYuumbm
hcMUlxqgeLOzUaom+ACbvs0+6vYlANGeVjFymCPiLb8NN7r/zhUjv54UcIm+lHavO37x5ROY+rDq
chugOtBf9cge2brsO364h2xVGfXuTEyFuFbsSWlz3pw6ImKl7YHG8VyeI5w4WFdR8G8EYHHBijsA
cUBp3BcIgrrq3SzXR6v77QCy6yTugXwhQPO0VWTwNcx3kGwxkb/5++C7it3FYvb2a8kIaX//Jruc
WCDmVxL/EHOwJjC32l2nvQC53PHhiI4G1YHrQ6qnVlhu3jy9EmTZATVSDcUGSYNMILMnstzsP9kd
hI4Rhc6X60jcYwRHnHhSEqqvN2ysvx7z7kY1XEH3Z0Q3uurjHnjYZb8u36j2EFPQpGRPK+deMi8x
A3eFWlm7Avw2Y1wW6TvAuqKNSriWfS5mm+XsjwBO4CcV66FjGLRmeB1C29//skHhVfWr+8sQV/Q1
7QVDUicOtn9NhnQT3WN5fbHNshWiv7i7zXPxDK6GDgK6MGrIAr98maWGJq9dxsDF9Y9jBHFrNDmN
XZ57YyS/XSyM1KnjlHX6Q7dURsh9ZMDevel54kjoU8NjFCDgMztcbJw9gXgGm70vYeZs6pj3bF4I
Saw97Vu7PBXoomskPFW9Av+uDKCbxdY8tYM0X0CLuL4IvaxG9eLlxy5P/1wVM1mqa3Xvnju9weL5
mrOjno68nXDmGdKeZ/N+IddmBC9oXE9ZgR03HihHUirq7Mm3tk11l9KzRY9Hpoq0lGv03Uz0S3yk
K2S0oOX0nAhftOT4+zvoYK/zSWQmGgE84z82+cYYx3ccPsWuZbwBbpjYbvYe4TEXBx40PV9rSUw9
Ea6CsebM2nzT2I4EsSdzIpRKQIPCsubnUUc/6bV/QWJDi0OymFFwOW4ZnwkTEmG34vy1tp8GE9cw
wBnvBHHN34paOKDuZ3ct2m8pg+9sMBXwQmJSuUF2WFvG2B7ozCsrY52q3v4Tg8Y8Uk9S4l+bVa5M
WEklovejNoqeEEwMKTrMG6ToGfLhOuPyVD2vwE9VwN7afKPMKJm9mrrZ+rcPvIR37np2fYk6g6DX
l33UQIXvQbfqijiASbYWZQzPMCrYV5akiCPr0YO0U80bh7l/BQEdd7D+jDhJ0DNCWPYgB00WeBr3
oMQM5qRLC1kp+JYHzRljflYOyTk8PszPgcAphTRgvPWSXg+R/AyeAvDR3MGHWKCvDz3ZmBCQ0Vl8
5weBWWvOYKdyUneeUM6Y4kFePGJWGws2mZUN4l70ASiuul6XXoXIv76G699BH6G+pUoLOWt6Divq
P9XPPW4PNwZQMpmGXCZULWjlTsMJdlwSE6VPnW7hYvtTkx1/w1ibglSJTN+gImBfpVAf84bVxlvp
8mdT7tfDTqguNd89StmOkrOjnAb+QkwDfFflxLAXd7C2grJMTc+HpVR6ubnpuzlSweTGDnVEEg+z
TPMYMLZfyKEfn6B9LOooulOpY6vzqv5q6BEqBk8+y3dQ3ejxtYxOnXZWPZMmtsS2UN0H/89MxN1z
R99acjwCE9xssUZ1koM3eW0n0lJHUPxnWjSB8oLev/sUJ23iJ2t/Yxp+zZdqwZ8/o+gj1sGjOLfg
E9i9whUBGGl7tPu7OgPMy2q+mSerMza1Rj556utoGQy/6c0YpxMuj6qMwTIVbF5Sv5r2vhv/fVOa
JSRjVG8cO01kLSIZqGakxvNGiZGNP7VYGx4yezdW1nuZQXS6PQz406tmsJEImNBHsQatTA1UJuhv
YB5EfvBWhZceZ556jRvny/k319jptYhefRag4zbN7qfZzqhgCzDajTaJ0K3vJ33XfG9CyQ2919gq
xp3a1SKxgl3+oqC2A56UiFrRAYIHU2h6kAVOo+/05TmlDkSDDnA/ABtc0o1qTRQSUORC/Bht6P7K
AB6UKKBTe768KBIEX21CcGdC/TEJOQ3W6D97ELP0eHC5vovdVd3oeTPkneVtJQAssbczOxMqBg2w
Nv0g+Jz9bJAB8jZramVVSWKxBq61sBRSFUgo6+W6hXOyJZq2eSG5AhOXHVQZhRRjyu4B0lrQEgO8
wN0/pqe04oYeWnfPHL3QMwoyYoPwX3xVo0ZOLO27bEyrLxvvU111E5bLyPutFmqR8sPbxiVGfq2Y
n15f4B/cLFL7m0fpibCAzHDjJPNTfKIGU/eqEcnQ7Akfn2FuXGOIXK+cPXuN+oIk3TBpAU4UmYq7
lhMI+Npx4Q+i44v0wKai3RSnUa40FwDxOoT6Fx/5o24hBZqCFcPmDdlUUJ52J2KoAZObmpfTCH7l
oLjrQUHN5WZwtQnaNCZ/18Af4m4y53K7ZtLeIQs4V07RKV/MDdrLx0yyiPn8/0bjKb6TLykKY4Si
nO7mBJn5FfT8XCRrUjxuP6nu5L1jyjUP6CXVfuTdrK1xSBBY5Xvht9SqNppxeklQxt+n/jsYmbiP
UfHzsRM+54AlCaZVBr5OTUVDU2yqiL8/SDb9huu/VaVe/oHh7x/CyXWr2xGQbYPrsKikXjdDoyat
83bJgXRLNs2/1be5Jilem/xJV8hOF9xY1tAkzhIOnsqso5hM8fqHXpn/oye6t/+7HCgeyRg2FgXZ
YClplCNoXXiQJ4DuM2FEGEVagyT4Zm5XYjcuJ/XTxhxU/aMQYwyjQisbgWDhuxn6xxlN9630/01F
HMa9p1vNL+q4kfvyNM5D7hDr/IM/jKiajPLcG8nZOpuVsh68x67GYZopQc2hKJHH8mC7ne4jc5ia
RGDhx7nPPKm+iuUQ4yQIfMBdZtApyvtMX7COQD68EDwY6gvNQA+tcc8NqTUw3i18WdFH4R08v32S
LCNlmEdIWaqMzMyaqAqOnc+/3YkH0ZuR7QvjOXKBCJibiiBElPH4sRpzK3mzWtD2QttmS+jJ9SlX
I5j8VFdrb0r2R5QBcLbXfBhbVCLO5HhweFIP4AmILB7HHXM1ZoIdbGt9Wq98jB4YY+jz/1YNzshQ
yXbcZcZgMla2k39OkwyOALS/FCDc1Lwr05jGyWmZwdVvqyFnb3El20t6lcvbnczA6QQpL7UU1QAN
5q8BLXEttjMuPpbhrWpB3ttxeVUhrCydIoQu7JAT3MviXoWVf+F32UmeM2RwlT8mrT/T4RkeuZf4
iUk0FKDdva3rUCVsAVKELN5z0WNkFXniC4I+AvL076wR1EHDTeTUmHYmGQZPwpG2owcj+reCpejF
X9hSkhn8nRdKbt7CTMsijx2a8zytc99lIU1C2tcFYx/c0wBhe0McMeXyNteiNUODhIDhgqsoiWBx
8Bdt7O68gsZyoveRiOPGmu44zHK0hCNogfHdVw+T5SobRVaBd1/ehS3RG8DjhMmE6O/GpWVQd44i
2prCjcSpLZ4PZCBjcfwOV/oMej74OXLBR3kE27/7wdEWtn4aqAh016uJxmI0YNevwJBqKu1aYTYI
vr8oM5ka55F5LNtgWEDR8l/NF4zCM0mGtDIWr4+dMHvBTAMlhgzr6YzdDQjD0t6CgYIccilcCcff
fvSs3x2OcEFi7x+Ivy2FntCEbpHNgPC1gIb0Plno2xmk0Ju1CH1VJORtBDe8yOjtCPoT+j/11Xxv
ar6T26G6ZVTUm5gRrcu4zzdN7isgC1UOZR+nVvWefBjjRN9iU4qgX0mTF+MIC4a2DEQaIu//cmia
QHemYaHaQSAUDcY6yeZHu/fDl3aDB6cWhsy5pCEfeSXJwvgThFVF9hQ1lQ3LPmgPGSo75fqR2Thq
aIJ5hVi7GBqUHVRL3LevrHDhwu/WeVSL8z0wakphn/U98Q+tMpvjXD3H1xkdGW4N4WtLScFMYD08
tw2BZc3OCrVSL2n/IRyQHueSPPZLD8peoLJEjPMyKxwdTkbAm8hjzMadQDtsPqr5dYFjp2+T6Kb+
8nGfUNixZOrKSrAzr70zlZjRlkdNMfKiE1yDe5KLy7COvcmmAK45PWcgCVj8GKxYcRsmW5OtdXQK
POdf25bWjXpZ2ND9Pl2086NWAA8Bax1r4k+fGTTEB0sM3z9HPXvPKTMKqM2sqy80IPJ+YStcDvvk
N1AXboY0b9HjvLlmMKTVG0sKqCHSR+9TWMRno5UVxdQMP7YgEdxTChvpX8mWLP5mCDklEU2xpWrK
znbgmCJuWAkT3OwDryru1Bs4TcHxtE2wnvS0xBg2OW0dgDV1whaOOuuLcD6Dkg5Qn9NOiz+N4mph
ZOVw0P+zowJ7zDWwQqBNVg6DttUr1eO4Ae4AnyPupufHWJmtn3YI6U+kxwV94jhl02Wp9k8C3Kih
U4kM7vWS49We3CCjh4kblPnU3bLqodX4xKYmgBNZQj6npJWz+BSG7ixEmOjzS9XE9djHIle2vAdh
Aru4qBi1JgIfnld4PyCDXNdFWXeOkspN8eOSy2xu3UQLAqwQ05UsEGNc1QMsDufHaUaABFp0kH9a
kgR9ngg0la201ZYXBBo+8ySfgmQcdLraMEaDTnmmwuh2NYVa/OMYfCQ/PGTUJfF/0ndTKluMW3Al
rYQH1Oo9UUq4G++whV41FE8eLz4MZ4y3T2JDhaMyu7UwtgQ8CDjPpsD8nt2JFxbuWW+xG4FLan1l
M883JDM1peIre1/5Cofw5PuCsx01Y9un770bA0BFzm4Y9dFHVE1XP4D9tqTU4yg2WsWHWFL6R5FY
K7aPM5mVPVgSZE2NBAchRFPatLyC+uPbHV/SFIs5AEMbWlIAQY3RbgYFyQQ5WZm3GYNbVogNp5+4
MhfoRITS77jMLbxR1Vy9Hjw7XDdgkdSAHK2lC07b/Xm86CbIQ/lzMv3lCUO3Yf8Bt3HNsoKcqvEt
BXP9q65yx6zg5edrnT7f6+aPTGsA+25L5qrIG3ymtTX792OH0rTkbCvOqI4pgM9vqB3AIZuEV3OA
/UIzIRfOs+YYn5mcQrWnjEF+Gp4Cr/+W7hW6KoTapRlJ6XOimQfh1sfJ8IIfRxgsiw2tDhtsQQMT
bVdnYJztNpMXPFx1e1wyxbaTfvdRwg/rM/9qWORbj59YQxQ+z+NzpKpX/zwPnEIeRzFb5O2fo5PX
okcwHYmAcpgEVsgy6g1NxEvpDrhhf42VbynJPmuIgB5q6ixg0CAWjI27IkqivXK7V1og4khvB5pg
T9yo87Fo/zYqaWjNv7hRIR/72s1PW6yhjS241tJR+wa/XXGML84NMr6PRcF/vQbKY3aq1SOzhJnN
QueA9k/HkNUy7pJHcPwbISlU5wSvJ4IbdKnVZPcWYkRJgJVdGl2jVpFsIxr9ymZ8tu1LNZWlKTvr
4Q1pT0mEu0bzcZ6R6UzfSM6HpNMzSU26AFwDGIGwMh2jsKh25hbHql9uRIVdGy8b0KS3kpUkhGfC
Bn4PZ8qF8GBJX71OKZOfPA9AKIZtb2Udl9XBqlyMYPrkFmcap3Y+fHfU71EKybMmI4eTto1EAnCC
/r/ROBKpRJ+Z2sKMkd1ElCpJrDd2dBPAioTJI2ZzRinSjVRoTnT3mu59Y8HLq311y7dGIF+5T6A9
N8/kcasmNenwiZVRsBRMl3y/jajkPFoi1m77xr9nqaPFfciYNzB7TwBaXh8nudn0JE9b5IcNu/Lz
n1tJg1IUxLB8Q5x8bfDrm4zt237g3RVS9Od6y33oXGaPQAhc8HijbiUUxRvjPkYMYIO6kqhwuFra
xkFt5VKaRmLvUOqzY06P4667BlXajsCWKqUWQp8Fh90i2KXK4fGjWyu+9xr4+Xj6KGZB30TTCQHR
7QI1/vROF/NhBIPUdvQFjjY/ORMOvS9LgT7lg98my9x7ZRwbrDuo5E/6HCopyFcidyEuLoYy4Jxw
N4FcDnXmbCaiiLCVZ6RrKE7COQb1Z7TLj9m+dahSMDRBG19ZU/n8Nd66f8cYRGORNPLoTt3vHVbO
FJIQ+5vTKmHaEjmUr6S2S1YJ94iaLnqMUbhPbj7OuZ7CsouMU9oioNNKUcviJEgtemRKaYL8bRbC
M6o1PVY9ayKVf7IWIRs7aJjfr2bq62DcZbYFF/prohHQvJ8qfa8gKxh5olCexgS8ANK/DEJuIVGU
HlpKqJswc14BMNn3d1Y+n6y8Qs3z0w8xRtwcbdZBzlNwuR3f2bB4Kuf1cby11DDXO6bTlE6vdmMd
fegtl34Q+gfnYd+EE6dkI63eK+ZTlQz0GZrh1WPoMVTdTo8Tp6nUGogv68VbitAkw/I0v2hg2r0S
ESRUlHR3+PDYBwgahRTDsGtvnnESij/DcMeVX1z1BKxfUMIydXuuer///NI8mDZUZCPVumJW4gp2
/1ccdMNBGSayW4LEHOJXLqhHYQ6DGrHX9b1WdGiVSGN4ojzO9DOYO+8FdIH/dgnZhPzxGESs5g6l
hOYL5crRnJgE/tRzh/JorVyaVLGU7Heh6ktY2tk7ZNvKZjA4k14+a/qhH0t9dEREe48PWIYGoSrO
WxHnZe9nF0jdlVfmxftoitRexjFycFh1NsiBV7J89npXiXyntcQfSOl/JRpINj3mpSiAz4ZLu4wi
99wNvbCeY+4k9JiLUITYTPrAUuPVieUuxIVE660c/d2AGVw6UYAXNyuUZE0QSYpE9KHK4CZAjsVK
YbP/s7uzwPIqyfuU7icgED/qc2LP9VcfsZ43IO8mKJIMXdfDsIpFq5/Ndp3AW/f6qEpsfih6C8xd
1QC+1j2OYVx2Eygs+HNqvL/PSbvka72v+4gVFZmdUf42PgzMMsx7+131lQYthqFp19PAVXD3nsuO
5nc7RMISnqA1LPSiuXLSNae695sIFje1r0WaKV4I9cZwORyrwg+et4Tg9N8M6f18Vnz8GQmtL8Qg
2TJ0vx8XyXcs2bMoicpPg4k0Z7d8gbXCoq39IDUdRDBJKEb7kybEeUvXyNZ6A5Wd7T/pMKXdIPzL
wMvML4yBe6y7NLKZYASmMflAdaq7qSCFKgobIXd7zqKot5KNN7BJdeMQpyufTnnDyCtYMP990zX9
udJSqwg2MH/9/mvmkjPK/p6k0mM/Moel0mCbJU5LcU82C8JohUjgmWtih6rMGQyFPZMs6mW1xw7N
IBzFYiBIQoZO3zPogiqPsR66/lmpFSuQESYERVn4vOYKEb4tso17b9FoVDGqVYTMXY/vpVE9uM2T
CLs/FULUDfl4dbgDprLisnSJmc1zPi4REKaWZGGPtV2wKOD+2rTI+1WyThDcWx+B3//AkaIVSLaH
vmWyZR4NzlqKcW4d1+Ef8FkMUKQKP6cWGrH+c65DhGHAOCdAVTlCD4dkud7rH6AOD8rxXgSmQ5uA
is2BKvzoEud1gCGVYjMpH4ILtXK5eenys4AizFMRS2ofnSu+9ALbMPoKvOVCHy8pcNcDEbwVU/yb
nhzh/wtm6q1KLBOSYOeIkT5zt6IDzlWgrdsmEy4JiFwInxEotvqlVDtarODget6NlQtvN9trJkm0
gAfScCZLiaaMe1WQL4uICz+D3iJ8LMMJJ5y6xuh3hQZRm/iKXp9cifeyz2p6+2TUqrAKRfWKhdQI
RRUHxmYpBB8OVN9P3kpEB28G8dj//qLiVhCAoOxc+a/etKXx8A0TAPwc3W7TQwekoBb3cocyeIW5
OrcjPDHbpO5iU+H70R1SqYdvUaup6JTSQgeb0RwfiuzsCihJqXkZS9O5RQ9bEdJAVUf4OOAWSdV6
QnzMQjFPkrAs8ZzEyP7XiZXSX3TUeVPuVTZtdcTidyZ6bFwghola8q+lnNhjN3SpVXbceKhyxc/j
hznmJpvYEg6ZIZ/hWhNspbbjSoHLw/L/OaTo7rWJiZ7algWF1oBPY1fpewarU/LUiS9ZHC3mgX/F
a4Rjs7fthQedl4dfxOZWqxSWi/7wblM5vQwNeOyMv9Sw0yfpXnYOJrzQININJsZBkWNTMZ0G3aP/
zYDbLhAa58TEHLdipba0/hw3ZdfVfqJSPoSPkWN0p8nHcD8vhhAxkYT/kkCf2xMak88qZYvfYzPK
WQ8xcp6d1aB6HXkNvTJ1eZ8M1dbt5+dDsSf+CrPZk91m1hYTZnRTjuPlxJcAvSyNEB2IyGdsONcZ
emI4bIqaMHh8GnKaWBoQfqwWKErPii77hKTAGAvW2xWV2JXtWPLowXLcBSs8s2n93cgCGY/SIqPy
YrlO443KHIW/HKl+NlQUM/yZISIwt8M/hSzIUXFmujESzt0wwdaIygCThV58/wwS2OTC/ZVHvD0q
tqFBb2Son020r7z2H7Fl+jFwgBLb/UdscHRU18kSJRm3T7lYSTxvO1MsIGhlqagqq8s2jg+uJJf2
HQDcUfpdYTnJuEwQ7NvTMUCxjJKk2QIgkzpGN8ATIK3LhFdr3cPdTkYQKUk5D4+HmE5PkMnnvHkC
8LzhrcR5fq1WQmdwZBVVBcJiXgW1lk9aQK8T3UYOrbF13okseSiYvvyTQBuSb9QSxouQgfUi6gJx
qMRttWoSVWhOo07ey+yIcpzZGVkmXJqfCQ46NbYTd97NBcgUVZ4ciDl1r9qU2bXP/JfYD7Y7jUdp
t0xmerBe/r0AINHpLsIk37+nP28r6AZ81cPFtd2mJXKaAlP02KUQgAXzSAAqcE1OIcm0G2f9xCBQ
vH4Ek7Z9crFU6qdgruFtbQU+dMC9JdW9QBx2Az8UL0qlsNKcJ6V5tZReRRCRkKMOAqsnujXp7OqU
PTLVGZ5sTWNkCLLmJ/BUgF3yfJ1F8eODBUkHJwXcBzz+aoQ9NnH6RkDUgZk/oxN0vCRzXgW3+3E/
/WDMqDrXwbyDfzbzaKKJe3KY1JbQl5vON7D/h1U8qmFWRC/kzOjlDlI/ul1kGHMCanzXwXM61/Yn
Nj9Pq8W9jU64ElxtJJ5qeY9Dd3NJVkiyofFYFwaqMlz2SChnAp34B1zIDID4mbYFhtAkSazhTEJl
pHNXqdRNJGTy4+3CDn4NNFXJqNTTlEBLL3R2Ym0W0+GTeZy9q5d8ONEOTHNJYdCEnIbSfLhuLk/0
IHsrzzcIa07r3K97CGF9MOYQX2gqoS6sRUpkHikZ46le021T8vyK/G15doiLWWFRdrcnLaPLf/CF
5y149TzdkvpX9WbI3+Vgk/BR0nNPqXzL8/56riKsXG7NYhHwCAMNEjDFPCwmG5fCYdYUpYfER7I2
p/T8xrgUg4MmffhiKvxGZAeNZbggcMYYuaSBMZ776aamcivFMXnzwG+C1Nwrrzuk6G/txmiV1GyE
iY/bNFD2FN1xFJHF1jWXEgynanNZEaAuGQl8/gx3KcWkuJwe0ojFOSG5LjbEZvkaIsRU4aKzvA7P
koCasbJ/c9r1z51/FuFgHrllO6hCw7ueiKQ6gn08jDbaehG3pFa5PJPBhkHx73QhgYZyQIvVlSck
tXYLhTYT4aLeB5q3GbI4iD6w0CzDW+hQpaKam415sHTPEIJ6c2rLlUoa7U58JM4t60uhiYfGxLUp
3A7UVFsk+i9JLayTpNYNktIfu7nA/n3jUXBbg/PTUTTQ1QmjviSEXkdDFJe0tl5b0GRa8PWoE+Jg
4RxJ0ed5Jx5jjAdq2xjYr9UTt2Fr36h0/DLrCQC0/A8QsaD/Xz5OZqOnzURp9Eb8Uf66kT27UlgK
Ct79t7j4fitJtRh7cCOzQHHpTYOptZ00yNeMuLG+Pc+Q8IZfEMOpYPyAGKdKUB8aBvmOMZzcZlH3
+BndCwahVDbzfDqv1VNCG4NgsmuYZjes3EQ0z6V8Khli1Jatsa0IZCC4VhqBreOcuAke3VIVGMfF
dfmKLccoIgQ3OzlHTDqWXhwAvE8hT3Y8F8nulmjJxXhMgJUyg6f9YAsoynW4OMxNx19+/UB4fMEj
OiWeWGKjdhnxsdvV4HskSeUc9ge5rG1Rh6lrYtW/cu/tvCZSwg96JhFomntO1YWKko8iwBhRZW2I
QP2lJpzAhUtx381oLkuiWwpH7hbdnj5YNZ2a2YszVjfsVs5qT5SlFgUAothxGEMTC+RnRL7a0zzM
LQK1ytypCp77BwSAGty8arhgjA7UHON89pNf/Xe5K7FQwq4O7jWCK/4EpdLFgXyHigIs5xjnEK7G
JLKvKf8qgxuZq+NInJe1WJLD1yxmIGAJUbh/GfiI4MydwQaukbnXMS5gUPXXO+EX+IHTzqFmNUA4
UVq5PLg4KTvxDCgVAaT+gcxTuTI74wZ2we1y27/RgjHDfQxmOmwTf9IbgagUsFxAV9cXj0iO7hpW
1UeryZ9aVVrGwT+SqKXLR6AXFKi2/asfs87sPcRmx/9neplm0QrNejuNSYLC1It47shf1MxP7bLE
H0w0wSOPVp5gDwucmKaLvZVySkaRl2j4SHRKs0U42s6JK6YjGjV5WjH7McikJMh15HaVjPKPADo5
HsKhOquMUhjwuTrCEknyIQkyNlFru2ZMlq/FHGdw3bNDHx3VvysT+f3njXas7F4AfMRdyzyjWLoF
W1AgdbCKfK4f894Ubs7qbgy6BCbgCT2CDeI1W+wNUrITh5b1tXrsYtFLVSujTH8mBVUYDSDyh+bt
XDteX/taqz4J7qJYe1xESQl5Z3TEwkidrtTVfULzfAUGUivY8t2Br5YPUDOIa2rvV8agBHA0L/A5
5tuJ+CU0so4Wry9ZR5Ltnri3dEplSU4VDKaVFAtnd1YJAe+YNrau/36uR1tFE6kQGrqdtPwYagL/
dUg0gKbOpEKDXlv4kcFWEBmQE+/1yzbtTTYHL3zcVB4BvXDKR7JFC2p3NuaHyEK9NKY/7y2i6ECy
MiELHBILipUCGTjZW83J9102m6hOepw1FAkIXk3FLThMWjR/qCwU33qGmjXHR++a2x1UVlK5QMVV
ZzwzzsiJtqun8YDjAswhq/RR6+TSaNM7AXV9CKHxD5pKT3nTcOQ4coMDoF6wCc7f6TYZ56sqqEaq
v5SsOQwPCIhnJBbbw8aWGhQ+vdVgoXiTy0NWOQngGKBaKYibH7aaDsvqPrbLC4wH8RxsWOV+pFTt
jb9Qi8A4AniuLLaATtDnxncWaBWSRbX3Gm1o3WSaavnpfkycUUK76lh3uetI4W/zDCTQQvomA9xm
cfoCcb+T8jRLsxV4woi6QQ+GnJlYhAyupaFxiL3EYM1gV85spBci/DYDvRnMdimvhuOqohZLJ3sh
rP1n1coxKI+XjZiqv5W35926BPgtbEMu0UAZ1seAOVekyiYk4mLiBbeqvXv7bZdssR3af+4H2oTL
9CoF/PYpcj6f6e3KknWZvmLxJ3j7CWd043dq1IHrG90FnU36hfNRFCzzvLsuYpJhGRHl6XKF4oYp
ZfZ1oI/FQXXuziqqnAWkk+aPfBiMqwxRyk2aPaQrGVY8nPNBL+e9eFuKaz1O2My/FSTQm1M4O6ru
jPMw0V3ToG+jBgbK2pPUpxnSQTdMKl9+IX3V2Q1jW3I0K1HpRP1W5WXdE9AQNYDcE4GqAcoxZpqT
ukeGXkRe6SpXT39CLDGjk2DsQxjRfObmg2AAGvuWSXIqkAeXlvarnMPpdq38bYkR+R2IBeieN3XX
TsElyO11/LSJF3dLIgCRjgdBuZfAPzSdVFmfUyZLG193ReAxWHG+VfVrHnx2uA73V6Gz2CZYaABQ
TWHJe84UopfT9AaXJO4n23m1+q+v4mP1tT8Fl1x1HV+3TfUDMYQRpvz49FPLW2DiYT6yYi+D3ApA
sjnY3o3PmsKjbgxvoDg/c1NJeIPATN9oOwPhfbv24EdLNcTGhBpT8pbRMy4Ixo9h+He7hew/Z2Hv
xfehRe3nI+QfbBOhFfs33/FoKcKbTJIeqbiCRFf/+q4sxFxqAr2syY8oKnJ09sBK8cU/grFPQb7t
K7nF4MX0gSLR8KL20rBN6mzYPun90noPLL9MBbEdYocMgMZCkz7K7Eur7nmp6hG6k9VkQxHox6Oc
S4eGGpERYeuj3vFZDEWnEUfNWdcjXy/OFsf7sXokJTfXCUJ0i8v3gUnYYNZJoX8U+++BMwESmvIX
CXmQob5mmD+oT1uw+R4M+zLzV2iNxKdZ8/f1KZmqCNFLKGdYYr9JqXZFVkgRLysK8PbhyFE02KiY
gx99yPNsLOgAw9v4M1xdaq9GRicS9eSO9r0blfLHQiClsgRJqw/fVZdGe7E0kUIrIb/FshPspeRz
0BK4aGSrF8BA36JAbYjQPWtt+ix61sKODFtivGAZHRl3iVbLKhk6RXUUcvibUeX0LtabCGrVEL6T
u3rQaZFq09R4JVLrMtnbynBmp6lnrMjuihVkSA2T8av5/2qoaboqarSbCENb1ckkEyfCpWG+8mVD
9WkHnendLa4zNi6ZdYoHIkvj9nZku3wzzCcREnfhwWDMMHZtsf+rnb2bl6Q/7YGBiaFCLPyVai79
MlC0VQrZeNz7Y60bPULnT9bQ3ObOD6HPaoLZKX4i4VkM//ltEvtJ01A02GU3v/Xv0CzIK+7dIBrv
gZddehUu1Q8S5cQPqKEOK6UA1pBKXgLa8V0hfB35viMaQJpD0atLuXYx5XmB3hBgC7/7XXEbpziT
yOWZg1tXl3P+lF3Z+Hagik7QcSA7gyaxQ5V0RalmmBOzRva5siMXZFe0UYPRhcgcj8PAfpU40bMP
5qU7aBnkUs+j6wReHJzCPtVY3bLBxlGkTc1OPlg8Z0Q9U/Av7LOY7rCo4IHyn1N25Q5VnZRxxk/I
Jh2wzxo9mff+2A1KifDI0mRo9eydlsZMAjIlCFQsY+Pg2fdRyERh6UdtbNn1zrGsMFwt+b0+aH/j
NJY+GcZKEgQswn9JvKIDIagChhgVC5N+yWnOHNPDYyj0IcapSHhpCKC3WVklLaBFwhF9vWoxEo12
dDQhRPoHsjDT/6dU7Igtdew2gYDFyxXQR58H6qF8A4NzkLYqczGuaYQAZf51q9SimK+5xjdMgEEu
hRAK+xWP3PNdnRJCJvYEKsw5g0yK17YM63EfemnReAklsECu64/olm/ILV81nxzzywkYnY6k3dxV
ydrlv8zXResYEBgv9zr7UOyu5i6FNAOXXpJ4MvKHYBk3eHvInwhsS7Jqc/yFmP5UtUYn0OiMkzQI
O0Kb2H5Nsy+30yZjIlSIfCz5sfwefwX8fb7CyNiRkYVi25RDskly2LFdsody5zQJ0Z7WwSXdavr3
Mh+iYTiJtLUISU46u8YrAtbzkKZZpO8PFs8Xxc2MEOkHlvtkAqUZ03bl6E1qKV2uARxNd8EP7zXZ
aOXAB9roSn1O6YjCj7O5GszYOrmfqoNOjJ2/ZWvYGAsMOJ+KDZ9t1cIN/bzNxCbO5JrZO2iYKgkB
NYWvqAHN2n9RBP04S3xbtwI/xa3ZPN805xEaD5FAHuERTFpLn8rOLfKVAmVvT3QDUmg+YFlr0lUE
BD109g5VC5c41uTb1a08r2fGwzKXRuQeSs7fQbDODGMQvh0n7uA1trjGTo48TYnvvZ3yGOb2ykai
Rw2rJ6SEwQOynhw96hmSn74konmPKTEwsHsFj+IPF2eFuCoeZNZMoaZoG4mjEjNb5fzzVVsrhaQT
9aT3dmhPdkRVq2XpqzoLNx+c+GrimoEY2lj0y/RkUjG81yVwFLJ8Sl/S12xTAwnq/HarruFCbT03
ENCZ+twDvjCL1IsT1SY3xnHeX01ZWI568BL7FSGlOELn8OnJ5Q0jBy6O1lGfxEq5nHStWsZg2DOg
auVvs+UlLCxNPtqNZVr+AEM+lQ0qA0KZCoei6OE9oegHCIMAKM2s0k5L3tWW1r6jLBUOq/x8Royu
0iDtPBdVBrZx2v1fRQaLfummg8lIUXXb3NHADoTG6v20si+1GpEMToxqzGEeSkyRdlB9plHcJQXO
os0wzrezDIeZa8hSNzDOvGpgLNB50aiqpV5/iXNBrpURSCLekoC5TZFvgNyJvZpEKw4JCRd8Cd4G
ELM+uzP1Tmjlzd//cdF8tp0EEwjTzg1Jiqhycdb9yBbZJrBeR6OyBW115Dk+yBTYOOhwDLnzTq4y
swE5qJJ7jEZ2clp3Ypynf0b8UQz4af9rc1LI7PjgtAwz3c3fCiFV5k4UDscb5xOyvVouW5PGzj2S
Di20M1sk5hcn6Coe/4sUOiwARaZHVyM63ADc4Zn88KQuKJFeQ8CMojn5a0O+tUrlWSi/1cF8CJcF
PH8eDGJa8Yfmju8yEosyrd4vRCLWIfS+Kglho0QcYHTnkPkeq1aOlHrO7z9lxYkkKlWxYAXb8nCv
OePUEtT6PXju7BGIVbh6kZKs3gzU77AgAw9XMfe6BWvxL2DouJdZrgLKIE5rBUtPbRlGjBHhZjeC
G9OCaN8Hj9b4H6HCLNpx4twLDrtWFn+H4A639CHBEHscITjdq5lQD3HAhBNjJSB8TrSrsv2cw88c
oAaKKMf9JiuQbQr3ycoZyQo76e+fkrVnW97mVdd4+F63JsyChP3F4xdLm891bVwJVAQl6xSpVFuS
Vd0x+yJes93vQYjfp5JbmICx8WUN69BwNk4OfkFjlsM/0IGLTDbLkK+TTA6Bqi9fHbIY6KiYkwAP
rwGrMlc6MG+haSl+7ecxQ92jtOIQ+K1NS76UhgIqtR+uO2zqkx2W8A2ertdXKnLbQsFiLwu0nmn8
ICL+MSprnXBgm56L3b5gaCiDyDPKJdWOsJW+Ld7vb50QsYa0Evc3amzvIwSzSUP57n503TWTIWp5
QW+j5fGzVi8Bha+KNStSmkdcSnlbl/p854YaGnvfg+MA1vDQDbY9jHAdiZsWjtW4AznbiSfmbtj9
H3cq2wxyP5f0HzTGyd93lM9BTqnm8EzoOgmBOt1GK9XWVH2DsOlRAl2tdmitnGQDx6t5mKQqoGCr
NRUMTVowcTtwJrZkvxtVPS/ywAvarWZBC58I+nI42198UlibPZjOxS39vMH7V8EKHVnTs2XDDi4D
kFZu3orSzmbKIFeUtUaeWvJiXs+2qQVr1S8Ol4lRQKgTT35KoEXCwpvp+aH9CV8CWAjUkV1DcJU3
w1GV53WOBDta8H3YGhS56uWWgf1/BATbm/7s8SGHHlqa2LNgXEWZaJVbJlP2W1UfWWUXswbB/HH4
CRPtuG/84i2ZqGkhC9B/QkuhfGGrmQm+TNirbfpN8GmalZ8vSav8NffoK14sVXwD16uRzpB/Ku4+
ljnyLyccsjdzcNxR4n6UvPczhxsInm8l3BW7k8CZ8EBT0i4aTW7aqQFWaRaWgVM6nPBnfZ6XEpR3
cPTlUMfUPxztGxTNnaDEk3hAy93uFbHW9FVWOpkEwdl6ZQqGgOwloudkQJZTD6+qdDvxFcKUBxrz
czJ5bDDNGzmfdCMIraGmDjZihzQpEF9SErYCxDX6BLNKMYotlXsO1TIYCQCELy/5Dhm12vMrPjWi
GimRFy1yF6qAWquTUrXz5o+RTgAu0WgGCHqc5x34lmdwnvM2CpmdbHbogE0CpRDM3fbysmufnYz3
eeOPFDubRoKo6RsZry7Pp79bxSf3i3DgTq/q61sjDo/MEzNwCWZilc5nrHFi5lQ2nscDyIME8S9V
/WNm7ITG4rRB/w2Nx+iyQIrapCjH3DCvNotfeeinyvjafbbykRJdv66esmGnORS6mFWdp/8e58Xt
1oMb1s6rf+RlRnojHqZR4fxGUvwLGGMh07vIJa+iqrdXGlSxGemYUpFVu88MKwlPbxYs5g7TsSpU
/VZKU1s70HiE/wqDXrKaYUTPgrE+pHmZOjiH6rbD++mUb66V1sh4npIsMYSeBB04YX79fMbac83x
zNMkRw5D6KEGkIiOura7f96rkIiGwTqq7NA+kXbti6JcpPiHlYmd1PNJF6LO2VpOrhT4bcCHT5od
6HoVgl4XaENSCejf1n4caY1ByJXnzKSjoxLO42/aS8RrE2ghEt4l3OENAuMzUB1lgVh2qt01Labg
ZErfRCoqXjp28FY9gJ2J++xLcqnDOw+3Bi3AsrCLUvYIvE63kDGjDgK20fS9G9HoDFHpnYPT5JKK
FNb7eiHQya5J6SLfcfd45uhghM6/DvkyD5TDruJpVqlVOVY6hDZlKgPc7rUbIXJYiHODyvhPwx7I
hbOTy8tXH/CeQOOUbIS7vOfy+hZE5rPdNAWOVjEIlQp6MpvTseiJubVaH0DZXwaayhG3QZ1jaR0D
jYqhcO0uuGy3R6So8yXTVb2fZvYgydTRvsitKr0VvqyEqFOSGbuEyoa0lDzb7njo4hWBci1ws1pS
IYuBzLR4BmuISxg9kPe+SHks3uF4cW7iO2HevwRXEMfLCnZtbrX1rQPc1eQ/9dxzZ7X/O9I681mV
tpB/bRIOelZCBdfST6PIr9hlDE8SMr21vSgzJhnV1qxn+lxBCH777ZahOmXmAcp+YqxewWQNHEmp
dJHGrONb41EBDRwRvywX+dv6TINK3+OenclIlEbypGoADExuoGOz98cNLx5lc4hAyLbMkWnFaqGw
hVNTSnM3zB46Joh9kfJ7OSn3wztZnea4AwNbajoEsC4IveTndzkiH93Tk3HCjOKxyoyTDm6nRqtK
8pDDSKQT0n/0waUfPNp+Dj7uHxoseVxIE5kvUFEZopQYMe2CLlrsVBlBHjskahse7A05jK5lbErH
8AcO8l9ezqvg6MfDpK7wZLC2oy4l/X+H2IDl4vQqGai9wwpD0a6bVIL3jHmR1M463rS1NuUtiY/L
mb3rPd8TV5lG2mds/oClieoB8vG4wV6L9/I8JvLXCtLdczYAGsx2FkjLILGjkTqzFIF21PUUFA8n
Uh0Soi8WOhd74YMXiNs5LdrPandI0ZO9GZTRKa7U9qT5/RXQeL9tsumIytTHqDdq4srfeuGU8LqK
9TlGxNeCSISGCIWpYqArqWWLla0n2SbiOvDd83snRQFCkoKb1Q53rvz4zsNPx3HI+ieW5bz0y5cA
UDNk5oDiIhMoDB/enLED8jQ5/zaQ7oej3rKJw1zqw6kcNxXr0o1FXyTam0x8BqjciOXlzfw5G1UB
yC0z5VKcPqX095I9NpZb+bl1WCZkZaibWWNq8Uju75Cf6c3hxlBkMGXTUfMJdllC8Qt99OrGSZuV
AeVUZFibxHGNioAZFgZpWwd+T92KbmQDj8ycOpiU/ppxTkhrTWjEu+mfOXH/4b7kmYgIoNDCmLyL
lseb6i1IIY9deA3OFT9eg4Cc0AuHY0saCsGXoANhidG0D5XS/HW0Z9+9bUKupm+QNyYpcOUayoeO
NiZrmPmJRwJxF8BRpkXssrqHAaIO/f1v3BIJA+2ble3CYqcv3TPsKKUNCCd94FoKyJ/3bIm5giLh
4kTWDs53N8Pp7DKyquyIuahDzxqif4BYEmzOqBm8hLjG5VeeFvuYStBM2ENlAXovFZlDUTvxvlxU
2DUPZWh8DLA1mGmK3ESDScQn63o5v6I7f7ietRm/jtM6ZGhu6m3Mo/kV08ShM8Fk6UsK4K0Y48yE
peees4vkh/5SA6d6fgUL0ExGdV4dxCPsGETWGB+OkWxf3Y5D8mGsFTXCgjZttbTXoICn3Bdg2nLa
GeJO50kUrIR7h7+VhUBdmpQu57aHTp2tl35D15/jhhkgRQkZ26QcbMPfMf6zjQTzaIBBGZXW0+bm
3CcQUcVRP7qBubzPkPQo6qRXrtBAAafh9+iZh+UHiXeeeYOtAK9TZwKhpA9S25z5HAOlU38Z5pp3
40MLKk7UEt7x9RcOKmmhmvY9aVaAy3oXUEv4YIkKVrsyZ4qUWprkxIZM6jq4dn4E5PY1ae0GrM/t
s5XfYyujcWHz9wcIoYMfpMOoxkHFpktkELlPelikFcTbvvovzBt+rlWsdUZ4wABA9myN3AiA7HkR
Eo0Ho6NmTB7g/qOmxH759BkwQlkYxQhatx0XK6KR8mikGk1lXADRZARkA8h3yv6FZmYX+S+WeTUn
EjHaHLlfSEF8ise8czRiPbpQPrs0eoY6/fsWMj8VlUMKt0zqsLN082rOpZKlvSQznFvbAzwsi12T
8rtkQ3MAJd+Oe9avc8CBrS2mdk3KK62pS1hWquBRsT4yEWlqPUrIu3IlO74QBPm6CfKNGxiV3iz3
oY6+zP5Fo7LIgi0Eb1QC1Zjn13+ZZ5cxbtTGyX0TQsPMJjrkhlSpZgjEf4mRfV9tKbAfChn0pN6f
mxEc6whlMdvHcR4EE9W8jflod83+frIeMl0DNJzpfiE7ntu1xHLLNp74ahNqsJnwulxvwjEv0JEy
kRW36gTyFUD2nromjraOgB2Gp2K+ToogzFn219wXWofR/PE6GpR8IGBrQW6sTr1+d3YvXqZreRfC
HPe6BSkI7ktNUSVeP95PHGmkKJSAaHllUMFA5pBIahV6sXmFM0dXxLOTLnjWrAeDA7XHF8XLnZ2Z
8JbffoBI1S+2inREBa9wcm748SmJS9fiyZJkQfIIH73CkduJJXuJnIWkVQpl6rqUldHm5S2yNpLS
qBMFR22KuFzp4YgSjZBQWNkRdZ73Tvwixr+QOPy0kE33Xx7NOPc3CCmPoSM7Q6QyzwEq0oMClc84
A9xKSjn75yLbhnmS932wZkGN8M+kptn2CuQ1UQ23v3V61kJwnMBoSgc+esvKXJiUEh8RlpkGD385
APFuo1F+K7Tvfdkt1dlz6+KN+vlSq/uCfRHPXwJxmKTs68buweeG1wzfNtkfMYM93l72f4uDPWVV
n24e4BfV6sWVA7LfN8eD323Jj0iznl/4q9owykIOnA0qXgA765HbR6nYEoPgHGwigggdAXPRrczC
gXI9ciheghnnaQiVt20lIJ1dJTXBPLHt0HeCnL8JvjVDJblO4YO8VQbKyfdH/GZlrHmTO5q+raEl
dqsQIHZM1vre3vdffbT1w77AnnSY9Zy7jMBapAVPJuC/gqj9cGSuTxPmjaV8fpLOyQcCR2PHnOjd
eff4ue0yP9Q4tMmfbd6T9TeT8JGv9ixovCpY/cUSz/R+ietujzyXOaucITjja61HJnHLDqsvIcq1
AIZbXfrHV/CEgyAAK0bc+LHGJ/4dKRaHmLy8byh9qoUe/ljDeUGKvWRWuuo4LS+9Gb+JM5pn3+Zl
waNlR2r5UfqpsvkkwEujTZEZc/+WjFey/TCbcUt2qrNWRGZOUTX+cH4FGvfB9xfRF/D4ef4+slxy
YvrNR4FH2HkmncLrNwH5mO8wE+u1Vok2Gtpkpoh7hjy/d5IfQzGBu5QpNixHHdtoI+LTedK8QoYk
F4aKRIJM6xVDWMf507rZf4t08Ok/0B6jBnAUdy1GTx0+8CSoXVG9tWneavNAMqkow04OJZ8i8JAY
cvDAgRTk/Qd6oB9WCWMhMNEa7K1UpnPg85/G2ok0Upc2XXbrcainfgBu33mSdxc7H5XYC70eZ9iJ
QrxsE4TVmdQKUoboxEAURt0VMXv5w26jaJA3pUuur3soZGX0r75NohaT6b9GOvLV5XodnQUa9Ck3
9KGRP8kXPw1Pcs67vD1XTonpLPMyjRbl/lUniYnntgSS5wmV+XHuWDU1b7uI4GHu2ZynIriFOWzP
TjLcBRD7zoOSERuBb2p++XmvPRFrESxUVNGYLzI2GKX8qJ1iQqanIyqywTFQoZTB4HL5YkX4L2dM
vRr+YlY1TUtlIOmRXPMTq9RgwS7Uax3mPq5yfkWgGM4JXx41NKPpsX83CrdQdAbETvTQkzcBVC6e
eSoS4D3ux2I35+47EM23GDFReKL/zrHF8GLPujuI2a6lLIGSVxBbzbkk3TRdLZnyE4hdGUaUGMPC
LEq1kLpcdDEVQhiUi5U0AawuHZXAgEYWIoCn5BBWCiURvfs1mgJU/yMqBpHYldQfipAr9kALnthu
LIdUAAR6xrlMvFGdWhe4hjjhu4kVO/6MT5daS+j09lwkuX6pHEBUDPdL3+runogv5Bajj2VjCQx1
m2LocSHHsTuZMFTnkAITP23BdKOlEogKNmNohJPYa3tFlpsS4y7RC05x7iTu6Y6+QE34DIalowUA
T+Oh2pk4Sp5qEADYq5sFbpRjIPfi6wBbhP+3H1CmBly1vW62QuA9K7R2D/oSocGP8dQfe2wVAMNT
tV7Ys+oFIz4HKi+VoNSGwsbTIlhnLR2wmb+78QW/GxNfxvAmqFEItdPiUdX6/+aM4xE6hcOSejgy
9qz58+pqT1gVXLJ45DUouBBkxxKj9yYxgujy6bc9AsZJ1svWgTsXftQQgAau6ow4On6I1cfooHdv
i9kRU5dViK6r0GhvzrTMQDkpRlgiNfQx8I1DmT4Lnr4I78Jyg6JmPV0y2WgV7jHFCA0aU3h5dKii
GNRoOVeXy6vJnf0GhY0jp1vGBndaVIHSZn5GO7f9azfLv5cwtphmpc02BbhJDCd7O+xLUI7zhz9x
DBJSL/mPCV/LvZ2ChNRqsVvbWz63fBDjhcpBFfczmZZfdPrTcSPwpDSJ5hvd84sHDTun6V05JkEc
3Jp1gleWji05CF2Y0EnNvLreQLdZR5O38qEXZo/jQzRTS2EygWsVm53RBTo2ullniFluu/AtKvQD
tgPx2vM8+xnVS/RqhC5moaSGzko13gSsymvHMjIzjFMGCDSfxCZUs7FVBy7brEtAIPbs/xyLL2A6
XjYbMmgWOvG15FG9pEyFsN7tRsLqAcWhDiFB3FiJ0CPPJ712HwI8DyR4y75zeBT1dN3jPb23PMcx
j1sO9youl9uK/2HL6Vo6RH/0EawayC2qTWzI6CQF1XphDRARX0kd1umkmudQ8lcThXRmq0xog8sv
sF9LV18jTr7mzKHQC+nfQxb5lutjUDCmLzyUnYPSH5Ckoy2pNS8TS1dAG0kn9ycHPFVFtPLBo85q
rYako1YTduKMMlPDN/IN+tcklwfeAcg7yXKdFL6Qt8WMT6AyNQZLtmNKsNPQ7/+vtVGsyMAVtXvy
lEHm70pfnxfynCwlu+zzUuNPqspimn0subWO+moo+X9KAtBV32uLF0WZTtkh+rICfnaCDRWdI6TG
7SdOiZwCz1pFSB2J0ErsPnRFjCjAfEcnaMJHGsOhdY2MD42fsYCe+h0o7oRFGtQcvnMzUrco+k/I
qfN8+yNrBoLgHMbMsunZVlznflwK75HEKNtTy3kEguj0EK26qgGvn4TDYrX/9dMm8wch45Wlr51I
65ww69jdmdKoxndSqXLkTq5DqOAr4I74cmEAYvBA1K7lGDQUunrQsff4CYy69lpAPeolD4djfgHo
VZpXZ/bt8HXRnTBjZC1jvN0yH9rRMSR0H5AQyVs48yXre104+//zoD39gIulTQzRuBcinUHRHgWL
2iXF0jgyqsib+prXwWBdu5pWdEvl181Qjti4G3sDH1EBEyFZovo6bpSxF68ZCE0RA8YNLei3YU09
0DyQ1vMmucB9KEQdqlXljdLWxlo2qFZjuiWKau8il5RaCKOIiQJSp1Nw4pzdRX7qf/7DdkEsKeaa
MC7C7DkiLSDoLlcWPrvVf6tZvtug5ftVclCA6FWwegYNeaWMQgkjarghC2udxeFWJdecp21aNsXg
2DJncuj2UM/JwtdIgCz86IzI0quQfWDSW61Au6A8Dimh5BHkrnUMRZDoxLY2AacaCRXBNwa9487j
PAjVkyzQi65Qr/MMwhyK6eQL4PXD2cqRXuXZO6zr4hjg+iOr1n0AZrsE/inpLMCgYvdUqj0qu2HY
PszXDlCjWPVjOg5Z/DElG3LgTmfN6eWCUzrioaaGtaZv9ywXvh0sq1DW9TLcQNo+M7sdbo2ts/xL
3R8PkSngY1VHv7IjodL7KLEfoLaWfdSm09BzHb1duRnCY2pwPLJZpTLUKk2TxcK48apfhx4Bdeeg
h/2uggXsVWYDiGYnGuptfBeAosW4S4aiPg3HMLoFPoTRxY9sboFKQjf9XJcfbxJvXCXJ12uWrdtv
jKv1R8AGjq+MawLCCXa1TJCJwWLIhou9u5Uq3+mD1vgRNYlD5f8j0rET8LqjxGkXMJOfOxqU3aMz
Ku60TjvZoZXCKi6Wt0GdC6jKnpXU/vU4mi3EUG8Ts6YED2/Ks8mGVeyslO7Ng9R2heYnj1hoA9bc
d4gXB1azTHOS1REXZF2yx1NCOzuCIz12D+2WxvIANd8glIRJ4rSXcbvMdPdLcCCEwoAwylMYqlDM
g1EQWYvaL0e2Bm4MEP8s17okRR40fVYmaHCtnhtKbnnh3NIoDDnoIfZf7GA2ewBRC0K8GIO24bbO
QZR99qySU9Bn9qs/TGax5gvXoExLFVqvi/P+oWXF5aoZCc4CgHcAsKxf/DjrmU1v1aeDf91MTQSi
phqGZZb+8ZrXwqVHaTbk36DhNqWgl5VEUOcaHE5Fe00ASuKU2Yis1Xh7LZigiEYsgdzW0lLNoCU2
LaeOP4bEAQvlkgopE5KPZXj6N33iMuCrbmNSv6demq8J+VTSG6jGxuMmcp+VSvNBcoVT4lwQTC+x
fC3I0sd4P8m+zQ4ebOpiEmpo8wCJVoogDXhIJ3TcEDvfXxTieq7ngeCzhkf9T35fg976T5rQRktu
eUvHVKMM8BJSKaDf9+ERxnfflVpN7qJEtpENuo1hOFH2KuDyyw+5pYB1mVZU4VNlIKRCGIKD2zSc
OtmDOXjRaI7ViOfGbyQDhVwKFZ98JN8tKa2tqyKVrlMS3L1/aEWH6MwcwBSRcSDdBvsPUNnZYgz5
T6zkyHOnBo2Te4BlMzEmlRs0eFJdF0IK5jeENo2HQZS4LmfDYPdWHpa87iX64WMPVhoKZJxkitZu
JLkENbMF2bezC0lbj4+LllfSbvuATVsdHScVk1kLUH+iVhUbGBN84xno2mCui4RlIfVm0Leadx51
ebMlP4Mk6teVdh7nVol1L4Uu5Iip6QbEq+m5Kisr6GBUfZktqgiGjDXcRaWoJO6d+2f3CQx4cvC3
RDdW6115iegDjhpO1AHCFSOmnLbW0jvFrjiHBypE0cfMBPafE3hLN7J+qhvD3N6TCAUo9jS8N+/5
vFFOmJA+03Ozz/i1KqfvfhC0o8MKd9kBrF5b/sTgaDUpdEyFPRHk8Q7bb2F1YZxvyhKIJKqVg8Bc
rvb+jrAA2Bvg0zGbeqKXMp8Pc5Abh5NdBiKNzsCtVkHXKZ5/KeoxfhgP0ZPVBzhJ0wZFJsIsbbYC
Sg7TdIZbn7Ii+NX6zlEZust3W+2rbhTz+voQGdBBdCW2lPPuE1+Q1MOQZ3W7gEPP34uvLiTewXD7
PnfAn2g7r/SoMRenCDS4vCvp9tRwKNSzGL8npMrLTBXBeA77dh5xFb5dGnDBn2m1CEakc3ZoNRWD
CO9lU73X5OrpQV2KtASIi41kvWjLBV4tFhLhN3KMGGHhMua30M8pVkF3ET09ku+jx8AaOJnvebfL
VG+YBrmk7ix0HSSK+cOwm6wU1CskdLEF0Zk4E5cBnV2K63n79KNC50jXK31ilmvquplu4MH+c+X6
X+CmAjcktjsPn0u2YWnQ5GiEjovCGeX8ieaChyF89utsDiCqhFHols6vpfhoUa2a4dowAB5h5jmk
LXPPHsKfPA835Oh1dTby1dzpwv2lZcDUHj+R6Foy8C3P9MO8bN6OSfjCi8JrwQMB0zYTN5fgCyOz
7x7ZlqAXjFNN42VZhFPVMbrOv2Z+vh2xmfT4+HRMtGeTpQSdEIK++k9g56Bb+b99mimLw90IsPhB
uigSuJSIv/om65MWkXNfl7z17iwr+XXzbbAJnvwUDY2lxbUCEzwS0YK1wfbl9h32+w/pKp2YfDw7
3lw1V50WWf9LSsaTEaezzPH+mCu75og0/EOFaKL5h05Kh0zOH1vxzJxsjnE1EntlAk66E0UA6YJE
aazuAsZh8Iqe0ftNG5UgjQl6ZmAWI0Tt+MLKUVokQKXLHV6XZEGMs2YZb9qymuzZGhkejrO8pDVk
3dI9ajtYpfLH7TZawYrMkrfHAtIQiEjBs/97ZjRkAKd0cZHvmF/GZMkc6cLZzibyMC+PTQ2VPIw2
0X3yitiSTx8MymHOWuozDJ50ZYPx/pt+iNU8wCFhu4k8331DMM8MZFmfyAmnCUdPGY1vW1YHYuUX
J9p+6WrDI3zQ/fzyVAZ2YoO3vFtD+rfHI4+Gz9TaY1IWSrk6OWI69YyJfSDtqKY6Ve0k97b4ceAV
uw5XIWROknLlqOb2cLL7bG+c0BOLCcsNMBd4bEiHoOE8ti5SprfLFQDFOACdyDp++Hht2UZ3BlAi
0gDRkvQFFq5D6Y/CpIjk1WVQpUiVj/zn+WO9Oz1vSzIGa88yWjBmNsWqQ8fgfz8MIZGbkaX1aL99
vKr343vnYBlWVbSYcpstVdkJMk0zrtmHULwLC3vpIwF8CRH93aUPJuSyJU17eevfRLlvxDqqMcbU
jMCj4Cm0e2ri0n/xGHWki+ZbYaqGcEiPVH2dT0wbdEIflI7kzGBU91METgHGkk3tdiBn6T1w1pbK
XaZvqGkbFIn4B9CioC4owl9O5688NliJR2iZ0KEEtngK3ew5cwhbo8FSKJM0U1zO2uP9/s9mNlDM
Y3awcaWdZwh+5ojib4s+X8ddVqpvGWn+FHXV2bXiZh5iFbTfn7Bb4QZl61l8HnB5c+C+KqvpISAn
lIMEHMMueJJHusoWYjM+zd67bhVXL/SZZ0509kFa5fFghyAynDouSMu3NRutZTrRdbFT6V7P29e0
+6lvwOivAwNdF4S0Juw8yhFACrddQWrxjqpwSrsazb9Z5uwttCqLKxsBijTZ2btdAFYfR92p1YoA
P/GqTh9F+p/Z/PKLcw6igxHwxEIa8F/D9dCAyZtJHKHMrAfEJ5SuaSAilW/O0d54ziKDKtu54vCO
qUdpXmI23Gcvu91bzF3LJYKCenSOnZjVzY5zqLKX3yKhiRW64ACV9wdZFEqK27TLNQ99lx8vujwe
NpCEmNNW7ExEGrS+Kulls/ezL1kRjgaTxcFRX5HwEi7P0/A/bRG6l/QNrz0nNDmcv80GqzjweLVv
vO+OULUeu+GncxijeYUzY6Hwvs6PsONzB5mHZ0dVFUewsDfQ5Sldj1koREUjbO7vxIi5lKxwwNFB
vttIFLePQwAeN4sgXfEpqxS0LzmveBFqofgbmeoZNQYlOXd60nLmu69HDsww/Kg+NHpKLNaf4hAs
FsJopyaY6W7fbxoNCy9AkiLlPy1MqXHDvQtIbpILn1lPnpYJN5YRWFxOZXNc8AlPk+njF7uLxr0N
zC2bGO7Jv2iii8a9USqBiYCUjUvVwNUCh8rF2KSfBxh4yYoYgCJ1z8ndcCi4R/o1zWmWij75w2u9
L58b+ExDLy6IdwIoqrR253hrA8XWi/UJxbm+YYbhKEILq/89CgaLD3keB2mxXzaWb9na8xlgnrjJ
etpbk50UZm3EkgPqDLhZZDtD1JX3v9jg8NQc2yfIH/MQZbgja9IYenHANb1sJ7rQHAn4N1HskfAa
26ni4343zicT9+9xBBWNBX2LJuvpF7qjKqdHeugi7pKqVOhdK+OMxYQotl89siiUuWkSGoR1rSIp
NAdif3qIOVwEjGkwJ8l3VggRojnSMsRtn9y3ef6S33ZqNJQXJrywwsNL6Rr86Fb4OyfJdmqP5XLS
Z0jZP2+UONxQx6DlpeBBrxsOk/3tl8WduYc842EVDFef8FEH9kQqzChmlsw4v11401XJP1oEJV15
QQGuWs8uY1naigxzJ1Zzse5cNUqPMGQ1nklJmTWab+WVYqVJfizNmuCVDOmh+fkuTOiOh3cNOXj+
EnklOc1pagzhVi5nmxac6txkfRZhMU+FxUFUQutlU6fSZMQI4aSZ57Gt6k0L5SqOODd8s6cJm15m
P8VpDwJ8ovAJU5Y6HBckII6zDC06TyCZMackY8KIP1AP6+ZFvox+gEoIYjAfHkXLr5nsvX4+xH9t
byKhorMxFis9lm6vNbK0qk+FnPi3W57nkGfRmF/0LxjKT3l+Ke8hLKpEXqjaI7ye2ztt10ECuCcF
VEBdwlKQ+erfuNY2QO2HG/bB4bGSy6Z09aCdRsfuGSdIhZrN/zS6ieuDZAwrqy2knH4AdY5SJjxP
vp+daEL5p/ZqQ1IJ4LymOHJEOuZWvF/IA6NZi0NOi7Opb5+nraTV3DJ65Cb7Y822+fRzNdMl/uCw
je/Ze+ww2ok+PRjqVDC1Fljs3NKfdqGWZGKCLVDcnb9VcO3QWRVrFTx9qTc9xcJVeOrWdW+91cdl
Tjir4VXiXhcUrqN+T1JoEC/OnXoEO094oYdOW8Cjh4WTxTZE2IxSrLPuFaN4JDJS17sr4WwQN95V
6XTKuzpUPdVp3zVBGRu3o8SftJWEcyslGRQz3pRZ0lxCeB1koh5pt+rT5pqPU9DB2F7pdQUEak7H
uV/DMt/Yi0JxZ6faFypynHTR9A8m/cEtOfUQPVl14onapvff/rY9dvfZHSHQ2X2HsZRLUDsB+UyP
CSu9TuX/wLdYTA0MwMieyKOpQoIKyr6xuLYbkW3TIw68qVypT6oaXzwegVE9Dxx99md37Qc6H2Lv
4c070Q33O03Vpa99UqcGyj4LcHiKfp3s+jCgvgsKAeNcd4BMVo9B5cR9gxYy5IoQE1NcB/VKmI/r
mv3CFVa21bvTJF1oP1gIkY4OzU3tFcLRI5SlA/d81Et/tvf901dVhaEk4bmuNUi1mo2F+iOMg63F
8veG3KrYCKBRQ8rVgMlcS5AT2zs7aVAa5p1AA0XNxwBVdhvDGZWvDwUwgetzrb8gSPZkJzZZJp7e
ZGbZRfOyJ7zsC4+kwUpakhSZXcXLJ8d5J6UEPUrsTQ4NqBGOOSr8YLCoeIKAl9t6YcT3dQdGbA7A
2cqIcqfTeakIq1agu0CNbrtG8PR6FYaWyg31AiPlzFUPq0Gr8jPImsVPWVmqaF1iF81MR92rIxAP
onyYa8IwMXfl9JE7bMj4c0AVWh04pClCQbrqn7ZUVQGssh7in4+9/47yQdgS1LxFbuL4wiwxDGYc
QKF1FCmcSRxhH7E4zYI1MXro0QqpTgNbKGOI1/bAlCsnz1A2iHtnwggiWGsV5iisLMq5ak2Wk5Yc
lraQvRfgJ1tqKf7Au2PI4DHERlUMX8zdEYKCGfZbk3QFydRim10z1TBaICcm8O35Kjfa+Qz7ek1S
yOWGpQVTsjw2u8ZMk1nZneEQSvOy5W0acovqLJHXvRVYy7auOSbo9XGkt3uyJwNAmpNAMUcG060M
x3mmCr+21G5y71umHfrGqnmmKNP8BWHu92akm/0hG/71KBlp8sFzI/qSGiSSUV8VeYY1sq/BVIzh
rh/cG4rCWuu6AsZACBAqtT2G0MKq4wHM7nBc2oBn/h0Fy3VkhxENSp1+iQOZVyyhLAyiWADKrSkp
2K4CdVf2v23+OGVxHOcLU3rZZo3bgOYPdDvRC4PiRyVqAR+tLWEr1VNNrlCAwH6oMnzptl8iQrJL
LuuXjXeu0+Zg0WlirWsZgWL+VtX00B1rnjidRjfwjjY4kE+4hZefnIHWMUJlzcDBZhFp3OAYBewa
Fd6RnxTlgNNJ6iUIOLcaflAoRwMXnhUymFZ01nEU1MqlQszA0p1STTUdDgWYAI4hgqRROd4UEPOh
j/daoCd3UXKNbG+gqSYKvGGpgWcPzcBFKdoEpSMitYNqs1mAKjhlO8RNfgHrUU4XydH+Oxscvlih
Uvp2sRbamSNOTIoyqM0C5lnvBP5x/b+IC3N5VcSZNr07gMAcEBhAdiLhInoe6uivyA+yiOlqmZKU
HYp2Qt2vorl1u8fpM8OTEoyxJ+dnNG3AJrcNp7A1SGQS7aYA6Nz+V4G1+Kg+/RQ27osvZPiZziF1
qgio7W9WiUlMWjXxPZszivH/YftrQ3pxlZWEsQeG3OWC6k9PDolveDGozt6FZBRCW1Aca6FCgpkq
C4x5ffc2PNrwoPOX2RtDEdNd33D/Jjfp5qz3Nrg/JjGM7O9Pmlo+zeIM7T/sQnWz8fdCFconiQVZ
+uCM22lW7tUBHQVnt4A5CDfrqlrcz62b9Ro4hVO2dmgsZjr867eVDn3sZ73KHyd0d3/s3aGExZvC
zDQDVTJNO0+bB1NwQVl5KURaRo7LaSW0zXKtF+yxDMzmK41daD7HFNnBOGsoXyid3dMZPVS0PdqH
YBVQsiI2VgoW7vSGfxqnhYd/khu0RuNVqyVTHF+1/maiwcFXC/ZYweLPd4aY9ttfOtNtFrEbVurH
Qg0B1R9PXxy1iRhOy6JGfnd8iNVRYGz2lufT+TBpLmKoWelN8IYirD40V9mLI4sxZVTi9deqbkL+
xiZ8H0PAGuYfW2ZlZ6XXxnlvzQBzV5ccCjHzY1Pn7IXAkZG2m9EUWNKkeaY50WTpeopHLmk7yTyQ
y/+aa1mq54dKgi/yKOQgB0JgsqQ1+bEJvmXOlU34OSeiopBnuXsrstuzaIiZtXUuUtH2+V+oLXzz
Xn0vTsV9C6R5OrPCJ0DleJ933LaihgMbPlbFxVtKPm/diSdtKozAuMbSM/UvITkWfDFbGts0mmdd
8+6+H2l9if8EEKhEOqvKBqfD8HbRU6BkllxasHVenqLjiWRTY8GFUErng6Wlk0Ws8oznNghwFc7B
LZtZm8H3FLdMxjVgVY6tCNE6H1x1bnObyZ0fcfqYhZh22BFeH0u1BqruLFFSqoTLz+w5udvkoQFI
8nFJk0zKAPzuZTpvpvPUMdc/YIwiFF/rbRzOvBcIOU3iPX7Cmq8j4X+gozenaOd7pJk4hgvkEwMb
cDZQb+0t8NdEB+nk2eOrhVu+PhKE5MFAuzZBDvCr7HesdYtUO5KIjY4WGlOKC/I4ti70Of9yUu3U
JpjTLvOKv5pLLA9xcpyqtp/d5gkvhqNtP7Meh86lW1VgzHQocK8Q5AM65Xvwr5+grwIOkigDNk/j
bnpUFeWBBC59AlDjdTADGCC8Le4jNtYqxHOa13K6hViA0czHzk1mCl5r2pjVKOWIOjMFPgKOhVTk
GOmGPnu53B6OEyKZB4yXXbcTQzzTDYP3X3U1MgDo0SLF2Ndmuzxh+Q3Ae8z0mOYi32Jvd6n/jHYw
xkGBNeMLu7LCAQiCUMV0RCFpckIOVRKhvmeydwnHQgz0S9RA5nkW0pDSqpXRnkdewT/R2OqSf8oG
sNtZrr3XLWeDK22V0jjLHQUUvfB6l5dTySehvnOWLakozBQKbN0fqYbM0WdTJAWGCCN5Q2rvIKse
EB2RGkne/Dlt8dr8PyKCv1ErJm9+pIWtJvT5Iffw6VYzgzyHtgycpYR/4aItspFbjxQHhWIZ4Kc/
vb1vuoV5DmGlKVexs8x0FJF1xKdg4ggg25pwpm/oNtgONL9/txMZGojRjtsCwMe2ThKy19OXxOTd
pgp3BAxFkX0xuxBAP1KNNiJvO+9txpcOPw5CQYqwBc69cTcG01pRCeSd/E1huC/Zq/n0JXHS6zxj
fzOcJT+1cIuP0uOxuKj8sk9D0unBCAUyTXAflwnvSB1pVayKmsJWakk/dXELr6SOTHgmmReLX96b
eLMkebHEbMjCRDnRi7sQvfkksIzR14pK4QgH105og1fFItpaCjJ673h7Feek/XPw/ft9axvI06Bi
vm8AClZOF/kvgDYMvesKjNH63k7Y+ds8rGCCdf5uP/oVJ7lrRQMXRZ6ZOrtDGDaswlMF7kUukr+/
/hSfuHXHXvjSZI1C5DNPDlJmkxx398NsCPFhWUcVFXOiC8yntngLZf1wLDQNmxvORwKg9rxJRlJW
Y4E9Y1OC7Q3zKjY8jXMT3cflgr6YYtYORVXe6Lfs1UiE7AaVRH+OfdgjyNQ2dWmHJAUpjc41wKOO
9B5wjT//vGQTjkyvz3FAt1h0erdmtaCeP/X/+PNunCuCmy5yPUMiwSrjw1utZzlGqCTUTs2CpO5o
Ey6JyoVrPGP38BvHrs09WQKpthZzORCxBhMEy80vxLmWkmWjS/4QtzEZmYiadX0JGa9JI4LQStuE
OHnWPELKVkUJiXCSPZsYPrpIA24X5uvAxcLapusCk5BltI/SXuRDB6IWvALkCOLw/0qNQDsul247
plHEOCov2fPgIANAuTYUn0RfMccN3jrNdlepKKRuqOUTgxEtEseCC5l/ZVohVK/Xokz/WJoKFDpw
HX0UXogzwiDoL9pE3ZSsaM1X+ndJwYP4HORzMpV9zSOa9EIUJlEQSaSHMR/91lNrIkeOgVUpnMie
6cdX+E7z1ppGt/a7y0T4A1u+xNiLbJmSPzXXgU9ugZST4c3UqC2uWstPs//H62LIPTa9g/3LIqP8
FU9d2YRAzEtHj+y82q8avWdb72YnjZ8Gq2QRGv0eT1Og3HDNsdDXXPR+cdaor4U7XPihcpl7aUqq
k7m9EyCKW3lviBFbXioLymboAHpAD+ZUR4PiazHacaXuk3FrkMkMPR4rHD0vrkZPh6Uunxu04G1A
ypR19QRyN0lrnAi1ilavYecUP8i944zU4qFkp5y14A8lwZwjxiAAcoO3DcLjTloSWht+ELKIbYo3
vPUUWx3uj26QMN2yrwYBYjaS2WztxmgeN1SNHZFTbIOlZAo0PMPM9/T2vnqAL+hZ+OK2WVm8HyKn
O7724zk6tlSvT5S4l+P9LdQo7SUlc/8kmqCRFngjGUPb6A8nfgde92N3yEsRwnHL2PI7GRndmhfj
2XADzW7INdFL1f7nJgQhszKXUM8gWJi3x7n8sXf4KSODt4VH/OuTS7q1JgPLFFbHmR+hrqBdcD96
dil+OvvCQYw5TI/WTTqaMhpGYIrEszgvPdnThVJaySizjiYjJfnuhLb9egmjIRDI9M1da/R1498a
lGKCZrMoM1gxDZj7Ia/P0RZlhNgXsoPoCFhUm3krDogrllIXI5bS3TcLLXCKGc8WS/LepPpzDmp9
GpdlwhpJASMv8USiwGkrruaSTzXSunZWTieJIhfv+s7N67lcfv6Q7RLClIyPFgJ+m2YOylXPBGBG
r2OCKd/1hMgighQ5/NZ3loA0nkHT+XGlOOA1tOfmaGJj/Mi182CxEPNK0W9Ac4DhDr8ZJw2Upu0r
n8fn11FM/XK2/rx5pGohOWX0301uv+h8pqS4zWvLyj8sXt851SBjdqSKKE+RTYZZKY2FVEMvOmeA
sb3SPFLjlxLwwc4jjJJ97YsTMIS+7O97zdysQ426rYBov1WtR/wgW+1K0U78FvS+IKxPpmjOFlQ3
xKTQp1+bNaHSsNHDZPvYa0Hmy40K3kO6CZERFiXxoM/t44klVUsgWv84A/hguAzxQi/twIIG1A+p
c8Gy/BxJ28hqQ6IF9hZ/m7+DM1ZXCxrbSPjG+thnfOQndRaEACZhre7XjsZGxWCpnMzJvTWj06mr
A0+pN6Sw7RR1enjOvPb3+yj1moKGqgjMSAgG20xUcQ6RcAAB4vFUfAT31aGeSHy5ki8pt46YxfMl
Orvu+V07kAO63O+2S9ApyennXRYyx794XrTMUQtviGJ6/nC1bhNC68MRnkyBGFYDYCTF4SlHsJ8U
/45IvuPefG59bvL71iRqCzjjUeoPc+8lug58hFBHUFyPRjjJjdV+PBLDX1pc8fLRzu7n7c73Oxx6
h/7c7Uxc50jorWwfDG3weK17SXQsF/zYcaT3dJD1VxZ7W+PKo/4VOumGNB4l2iZNPFEVFxNDvgE6
cupUABA2g8HyWY3Ck/q46MfCl5JFqEquyXx35iB7EMUxiurHgeEWAkWpPVJG/6tFMPgxw1dOMj7V
oVRNtSF8atHxD1yiDr+09G/koDuB/HpxqJMGLlgB3e97dypzQ+WgXKTBkoqYGHn1c3mR6IzvIC91
jR0fxKY/2XRG6EKprFjpouHdoO8wZwVUIP3HeqxpbV3vbuCdSnlHvXeC43aQOlM6aPxGcTd+99cN
aFHTvEenfsKPGJwRPymLvSASIV9s72tbpLPNp1XjdbF6LpAZXAs1fVoVxKKKhxeWLlC9917PuRXj
1sGhAv8kHScnBwe+EHbAGBGCEx5wZ4dhSj4LRpXxQd0oZzyWZufo8bGv6HDJ8LZvkVpIzKopKrfa
3GSo99eCK+5Rz/4kJRgGP5F/MnVB+Jyfa1mAS4vWVI3R8vp8jK51qwIDZBUWXocjMMCAmlPHrF97
DnRsT/G/HoJVkYSinmpEaZOidCoXTaV5KebFInXmdmbo0wFMbEAyg6Lgi0U0pA9NlKCiDDeHbbje
hww/9kwMfgFrShALJGng0GauATUPKxSkQK8HxQdpp97G/Q1In/3VmStDNYEyEX7k11Y88jDXgLMb
iyEzC9NYZEGx1bmQdnnxrisBZhQ8ZVkr7O9IiqVCxDHnstZ7t4rysGI/tVF8WL7aRXSdhMLQRoE7
fKs0+Y/XcLlkkTX8xHcMiv3tu6bwlTUdMosZoQtKTYcd7nndrUR6GWIxf4OGvmg3jlItsQfFPM/a
F2vHcRQoPVvG8/dbTuTst80HVZdDtCHLx+IiggiTcmJBnargBNXqSUUQkEpR9001qZU+rasIfju/
gwiRJmJP5HbJJyxi+OHwMX4a7XB70gcMhstk3ak22opZJ2Ev7G01wdwXZ+JwP85wyUKW8wvIvf9V
qPMw30vUxUX9sHZTCZhsYrMDHpjrM5hXOl51j5OgF5wPiMZpHjP9Iov2q4PjyL2UyPLtf6/T7cX2
Xtnkdh6GSUzmlP57qGJYNZwALG4jVovM+Z6LpVgePga9uYoRJmckX44GTpbigNq7XqWF1Wlsq+dj
MfTP9LW95tcVORD6n5Xtw1UEXAfTH5sYjxoOaitUwabYjGkAGXnDft9L+EdTB0yO1gxNOYEi8tRP
7b+qT+weOs1g72DaC0Jjdo1Jst/n9Xo8FZ6Ms/KRZ33YRo7WDWlOYBBKgLxP98z24U5VYhT28fJZ
TGkFs7zhlOSKuWEMdSXz/1n+vw51n2XI+SiQ2UUjrMqg0uN5++Dtr77F6MMKOIAp4NvG/p3pqn8p
jX4UMR01++hkjAcPQLcj9jP+LShfklBq4Ub0JUXigKmaZ3yu/y9ACQlisleMUapaYNBLaG8L3BvY
Aj32FkKy6pp+7y9eC8qq5NJARK+l7aW2gTPX6k+PZav1xoLb0sLTIyScd88vbMusGeQgs3GuTKGi
GvQBBLaJwnyRw8JkAwwNh3lHRTOXBr9MdlyC9gaiSL4gaKjCpmNLJVm0yllodKdOneOwmz4btqv6
ZLlC+5f6kvKVQkYtIi99ujK1RaqsapLKv2qsfa2QxL6TrpGo5knu9nO/p7hUO9MhY2S1DenEPcE0
XgWpqH9lcL82VrnMHPiDC+qhh2XaGa/GPXFJClu8vTcYKrIogKLo12p96hCAq2DJpArldwswATqo
mE5Ngh/Ypwe9EsNvKAUWUislL2nLIewN73X85xY+xCrDQtiY7u4PIgtaW7jKlZu1Q0DxKH8o3gmi
vhWoPBJBHrHespJte9wRjhgbkPp+9tCsTbmBl8Tu2GV0zaPTuTtpTs/enrnQFAUgLx7fJYLbo/Dl
uqbPBBOF6LSPjjBPJhN8Mk4gPEyuY7YB/XdyB1PQQJgKpin3v8Vmh/FLwCtMb8PcjJtBz7BwGLRB
1ZjleOYJaoISyJXDhS4Vc/XDnzW+PFh7JznVypHvgn+IvygoXegnoerhVErBtps/mzsrBp+Dumw+
A86Hrec41Ad6/XP8KKwPaJCY/fAemhFaYMAhpikgXOEKpe89jUOgNqr6Q2TxbC5gkhCo9zcn0Q1E
Q1tNCF3HpFneIwGU+73yOvZNatkE9w6UDqJjWj/n9muASBMosPz6echwiKNc/30Qfm6XxMMdvFjq
fN07LaYWAhBG/O8Vt8d51FXHCr1m/xjXtRsaMdIinhaJSW10DDqMpjIr0S7AS2JaAyPNFF3zqMnS
G4mXNsDbFLUoayt/UrHSLpGmGOn7xjUXM96hhtlRK6HevessC5GGZGItmiA/aq9+UQT7A5Y4xd1E
l2hmbvvXWVtb5ZnkblHIjbS5IOGjgQXWV3k765cU+9qLcrDaK4+swl7hgJE23Aq2J4Cb7AkON+Ta
cLoMLQaO1HCoo2B4IuQXBgERr0emaE0MDXUUU9B8LKeiB1ltel6N4pdzJHcC/4ub2DA7GrWM+12k
CWsMT+Kz+BzO3p7YILobs+MvIpdO1+0Jy2JAfJ3PaSf5tmKlg9lLJ0sVgnunVUbXR0Ub06IlOpSF
ugit9WbGtGCIFRPwiG9D5VY51aEK4oH3WWGaQcy0s1F2oeSwLD4rq8IVU9mlUmd3e01yv2ficOxq
llj9/MdDl1VzJ4m6vHpDOloXvLaxy9yDGU0WpnWA3iMY2Da0HjIUBmTm3w3tl8mLiYhn+o2Dcml2
ZyS1K5Uh13MduQsMnHC9VyPVRvKP+OTNcLW88M9p7gyeZof2hN9dxY60yJSzmiuxoLJyvhYsAz/6
PcRTjMEiCfhoa2sFVStzhhYUCXy3a4Yjkqz/BRiJGI2cyKa6GeeZLVh1c8dMDhFRn0FYmtwZQQEs
7TE4nD4WPdfC9ZVoldtOA6/Ay5quIlz8Pmcl3UA6kvS1K8ajbBzcFDVoLabxfGGK/ScQFauFmQ2l
Nqg+Fo7gv5L6q2VOwRfWoTmEQYgdtdNxu1xdx+LdpmDXH+syYLZVAn0TarFVim+yCtoWLxbrEE5n
sQe2RxjmpTy8efsh9N25O68VJOuVrysgXoSSPkSFxGjTKtmolqiDDK/1hHFzGe7J5MoL7VLa5oVY
/tjTPjhFcp8x9m8+zPa+uOc/O/LfTo3RjjwUWMcqR48QfU3Mm7GZXW6uwQHtbVKA/k3+xLHYcA/Q
rk2e91eNm6lelxEcB0dok+AKLmWXay4b+XPQ70+UF892P27NJgIFFNG4UlVScMss74vQL2ssYq++
jHN+BoVynbrI4SjYvEle5qTHT8LkNnHoK5T5hB324ywURAvEypcm+Swq35qLdWeP96dbU/Tyyekj
P8XIgbVihZuykdB6TiU6uLVUwWHcfApx01PYJVLEZrqYtA7pfO8xWzEdxQCeq7VCSb22mTxnKtop
vC4bhRxKGIalf5TAhJNU/zIqzLkAnKZdZypG8RoVYPWMeX9yjKVAoRIMMMx4srW3OpSh7sA6AC20
9B7/yRmUm5NtvfhnzaG69wnCj6oqbJSJ1PbiSOb25IC2OXgfSx0l937pqkTaEP83dgfW3bXHv4Pd
VBSVqrSEwWvZxNuNoION1wNZBDAuyVLN+983CNKwCArjRYfQKeo/C6GprS5KtLBeoTu0icDY7qeK
gHpYguWkEpYP3DMrv5fVYPKke8jUxjQJJ0JO7c0oj9Bu3cyy/A2SSTy+gSy/4tfTI55oGcUpwEwb
Sskj9A2qF7lMaVfJwGiNrGTTPsZg10EXE/cUlxZYc3G7yP7MuWUpXG1G/7zsXit9xYbN3Nm1N/PO
okzY3nM4OuabhwH0NFq0l7cnb667e1qPEUoejuobjDDBCQEV9cQrfrf+MTGXvhYJiyT9FsCGHGEY
qqFSiQbbg4dEegkP7J0k1uGeqe0r+OohfktK4ufFJ1tD7Tal7xGT6aji7EjEfPxuJ9nSnieqyE7x
6dGKY/fm6UghuQ0X5VIu8k2FvNKFAvfveqChOJs98EGDEJWWJ7rJEI0q9yMiSShWoqVeX943t6kC
OJlzFEdYMAmSthwGcvs8KV7jVFXfvUgpG1MoeWg5ejKzN0JJplXp5DCycI1GPjaCb0shbog+k1XK
gfEzJLGNJ981HFH3SPtQjXAfC+1IeA7YnOkimffGLEz9WOrPU6OZvr0TvwmU2HpjgL0rx2/LD/96
4TER4ZEebSmwdoJE4W0+oilR0RtEoN3d4zlTFcRSCIvk9MerOWTW5pfsF+1SlGOPXC254W0meBCS
59NXMurAqqhEVmgjgEoRLHvn/fTPpqA8xDek9GeWMABPaXqjc3JvytqOrc28hDk/lvl0OFLRFIrE
knC41J6rh+34A/atqOKCPDL+657+/blYj2GjkCCbVNk8jYaM5pJTlBe7EW7OD2qePrg0d8i8BZqG
L5iaQw1j9HFfkLsRDQTiisrZVm23tvgIwH4j94P1/bjcBcOmEUl3SEigos7WvWfhfWduWVOAAAXB
nKuuHyAQR5ig7cJsKLc3uWzF9wM/8xdKfe1aboBF6MbiYoql/+jtlX6fswxfn0DMQr/7LF62XRvA
mOGVMBwLZbf4SCw4tXDMLTTaCHbsn8Qjxkz8gMymC0qt68rpFdwCjI3MmuAnqRkpKQaob6Y5EfnU
s7KqiyFbM+xi7G3SINn2MZObghD3w0Ll7LKKsd7p/I9RHwX4Rt1Joy9hhTNFXg7NFOK8AzhX5kGR
ajrdqTBaIFR6DmhjQwz5pC+DV0AtZ2C8BQv9XWLpnjtOnhx1SsDxPTF2vApGYgE0GPWBb4IrSWpW
WoD0aew4BI0cnZRpPA7ttCZEN3Ef8b2iDZWxEr2dHSbQG9IoKYtFZnY6kOzRAIa9uo8/AEkliE65
0KE4U7uqSwLiNs0kxOPwPVFt1OVQIpTDTfPB0O5NJPFRyxBpMbqqR4s6kB+0dSQNS/XYcJ8mMgoy
co699GZstDh4CQIR3xYTSMkNXbJw1wiqkxIKz1Jj2U3Cj92yuzRf7nH3wsgaGwG1PQjNzcTXwM82
7Uv1pvS5vfthmDJ9n3Modn1bc7sOHvBoODa4J8eHGvAT202Z3sxqYykk0PNfvuNbgGswhhCifzoC
FmcxRi3tJfSNz2XDAFvzfSqtwyT9Fg3bU2fHHMU+CPLx1K8UEIoCwMRakbbSAUykQONPyqhVSA3l
+lnqQZVL37wb/48jppPKc4wYKWCYU8rpwxnSwZ0JU4NEa7gVLiup/HNTF4Ko6XnlNnTvpoYyV7/I
tUPM+Xysw0bGxVUmkF2pNELdV1KgSM/944WlSBT1n0/h0G+9ru8KkBs5N6l1J8UCuBUc4LBHVCMP
oryTgJ2fzDdpHDzTrcvBMpImJCRCRPE8m5/Nb6wwR0RaBm1vkBmzWKTVq/Q6z9VLkOzu2g3vTgQb
gOy37si7dm3qo4gvbgyYHRCxgmiNo0wnAcO4XKNr9xpCSmsxAB2tz+GBuhMQw1axpnk0NUIBfZLN
RPE9T4B8nDvoVEIGcLXNYhsT3Gq2htQ+xtyxP8SX+4zEC5SeOhD2AnMfcXjncNv0fYyuWq7Fp5rK
Gor8m34Md5ok+LdNSNxs73aHgLT/l1vP/YooQBx/fGq22ZP4vcLEgrydQMK12wD97ZD+vsZWto+/
gOZjfgzdOz1f8DijZAOWpr1W/JyQ7H6MmAU3wV+jlyFY1OhEuF+ghJ7riLK4dnUVXbkmNmTvVldc
JWKRM2idLiusDBT4FONLx3ySe+RwhaoB7kM91rK2j38gcx3pF5qedtbCbX2k48m4lBqMOvddDqwH
Xs/GTZs2Zdjee4rM5bTrQ/J86CrygQesosQdkfOmU6DM+OUCq1n+Ke/CveV8bMEKki852RA6FEC0
YPHfJstHWj2qxGyEXozbz0HHHmsHrAq8Tumqv81QCiMf7hZ8P4QYEBFc1TS/Q4YgqoF7gLt0/PMS
tUURPyRbG9yKhkHj9UOXaE9fIVgwOWFRwmggwpW/s8Bji3xy023KfShC2LTa9VQ0Pm8MT6MAtM5Q
y/FxjiLd9WdzRrx7y0YEXfS76v/X60SaMWqcbUzgsobP5nO4330af7Gu68yl7LRj62JfUIswkbIE
aeXxLxhYy+b+45Br46vLuIRSbjDvow0ZKqlhK1xVXw9AR7BpXNR9jjvdUZjh1Yy8+eXSxltntcVY
eHQGxvylSDMK3BZVJ8TWz1yH9nX8yMWXFdx8KSedxUqH24W5UKRDspgwL5X0a15pRi646268c85p
PyGQfkpxx1WeMhm8+NjfGT3JZqaQCdMcPBms+0LTgxTWyseQK7bAZ0kK1G1epOJpHXJAqKXe3W3b
v6Tx39O2buUCLC4d4mbg/THYZXt0ftxeEQKz1/tMyl7NHcluMp6so7luAL+NBCJAwgS8AFwBdVOF
VrdFeRFOmUZdTOAC0CH9bzyIbwDTGq3dohDIygcDNrTTbx9/ExZjNE8shfN/WhZG4hVLpjzxyxd1
kyC9aN/gSU4LxNFbfFk6Y+JyMNMiTKffq+V/YfdMDOEo7F5yVXTwTgjzMBlOa2Y+2x/zjAAoUgQK
QxylBxJ/QvW18s/Iwhv4UtDW7yeZqU1dkp2GoTVg1ZqqZEK1QZ52Nqw0V4Cf9lVmDscOIcZxEjF3
9y3Z9vWp/wZzCSVvu8qVVw4aVba1i9eOpRc4JKtNSaD7gimjWyEXuVXj/K0GvkmSdf7vsLNFISTb
6MjFtV0p3jxsy2TO2DERP0V5jFPKO+kK3BHK7VLGgBgZJD7s4UVHjVxmf70XIdrjgUvf1F/pQ9Zh
1/5nkPXnXEwqA+9ryQXbCSxZQGB4omsKNowAK3v6dos8d771DQUbR3VdXn8K5hxy0OXJDBhikeI/
UGqwtUnNOX4OnX2L3X2QqsrzkMewFxJxbfAsspX/q2XeF/bSK6/ww1hMxeGUiKbECbdoUfoCRtt3
0N/437KDIPSXP2E/jQ+nc1OYGVwfNi3Aw3pUDAyR7MaKiTs8j4fEordZdBHp+o6LuB38jm5WJoXY
QXrCaAp40n/AN8A8uZ1bInCWgKkK7K9ebz82PC7r9sHpqSPrl212Wl263s6m8F/gyICQLVyLS7Q9
DahvKRerWQpInpJApYybh0HJO1JtwArw4eW0YKO6PS7nr9tYXxQav2s8ZevNiudppSPLPVLNxKNy
ZaCVkzpXHgf+dmkmX45Cfl5SE8Y7OOxYGSMdN2aZBJFH5/a2L9X/IJlx3L4WBgn5si8OMiUVGcjZ
IPe8Ye4oJoyN1yU6bcsQ0Eqp/ENkDKyHPBjs0+XtVh8+8QCRC84Pqsl/xu+xQ1HcmMee9a0Fms9/
N9jgGb1q6fEIEUlHsz2T3+xAECS3699BvbeMSWlvm+skdYxVtdw1/9QCujWBMtvWeXr51sp2c5e+
unI/hiaWpww3hVy4zXU5QCZROkd3UFK51NcPPGGC5Qt15W4PFL7ZVPd11ie0IlcxN7bv8sT8+OKB
m+tHDcyr3VX40F13Qq2lbO5mi/unBaXdxpcg3jEv8NaCRzQXzbZiBezJOy9/2c6RWSAVmxFV+EqU
5SZs8ELWPhdPU2jsC8ukwwGw9fCWj8MB3B6e3UBnvCCAc2U6bWLUXIrS7GG3sX4iW7H+Ns4Gil5O
z96Cl2c0mLn8H28j8zjf7lGIChG5dYr5FVIHCw6rGVOuY95K0ihlCrCtVCAHxpckpgMjGE1Sv73A
oNiZiMLZ7+2jgczrSOsNYvxkbPHd3UGAIL+d+nSTKUlqFdTVd99E0AafFq4iSAv+iuRlUHl4iU5e
Vdo7PMn8jfhVfwlzNl6xu1hgg+/7nJ34/c5xVGgR8FAUJwcCDs747jFovVomtRz8EblAdnbn3pnR
QOCxLlheGsNMFHizqHb0xij2anZMh7unsa8r+cJf+jVm3MTt4zJoFRUkb0uUM/6Mi1XLtDZlWHbi
t56xYAPx52p8H0icL1hFoVb8tc6F7ByvcYMjeRI8TFb4OWiBkw5oab8pECF3r2HiylUzPeSucw3s
bzo3gMicMWwaRqFU5mMuvDoQ7ziJC9R5vWbvv4uaPHS/OGBYGKA/rD6DzIehcs0U90LD/lUcAW9f
nBqBVj2b2HO8ZfXbtf2D0LOPDW81pOpQDzk9HxhrrOxp/fKCbUdFkYdJVpnpLp/RP58WdIJbYzlN
0RsuNNahvzSlRpesLdnbeIExemiZ6UevTuYerFGs80TURwl/fJoNi5k/4CWYJR0FcUopoFpLRDgJ
SKhKMgKGzOVaASoWslb6cg4BRxSPRTl/aLdqRpvhowoMpud9vjBqNmM0l2WXGc/xu/PvsX7Grd+m
Xk0Kva9COu0kPBgXBs85mJzrvtJiSfQyNSLDjjZKYhCOnbl84xn+B0Av2Ql/mB1OFB+B51S25/n0
SDV8QXrDvVZhIDGlDG6zkoWv+Ygmz9TZ+mv4zCch0yNonkD9Th+kCsHksd43W2cs19Lm1kWfSAOy
OB0hNEJLh60gcYMtX3WDRJ7mXUdxzERmdBUXcWa6/ECbhro/5jVei/wq23GETdkL5XXS/sRlkGui
LkBckTibUwTG6lUqEkuOrcumYJCjjKkXpM3AS00AB7Xe1o1zwTQklfF15gs+TVDvCyRW/QCMIbHk
GWOqLp20f4E+o1GhkqPv2iIiAH7sFatrQzfDQ+3N7kd9gQmJRvXG5dBHOwp0h1AAj8LrT6jz2itb
jcJhjIsFMYUz6/80DMNsL4pnJ+YnBgRtS0IRYeJka3x8Xe2PJ0VKe3dO/i1psOxIGiCbpFmtH3SE
zZaJITetsYOJQvrQ5ZbfunbzVPF6Z6s78i69Afua+VkwFyX4n+lSf2/bKMIncKQhUube+dpuUCCT
vsy1QyesV5/iOOqUfj8gUY2HLA5iivGbR3jYjq0Z74kILwmwe99NOxVgE5/LTON4GZfFq5fS7r0s
GsjtFz3kv+GZ5AaW/vpQHPj5zgiHYHpQdXoSOBQ8BSJbW4AnXBZaZZcPrgyOPFSzIltpfwoZtkoH
aLArD/jb05F6nt0a/Fnr+vGc4zgf3pIZMN52eAQdudt1pC5IObl8cZonMZ9bo/Xj7pzfXn1d7P4v
GpUsUIIjLR+y77NFpElNI25mNQYFdLZP1BRHMiKnCHWGMHGMrj6ggwLr4CfXg7r+ijEtrSfxCLtm
W2eEq6V82SdjXUUPQ0LmHRquxqpw1ragRtj+JFu1q+yd4q3QqNpR1EUokMkKum6sJSwDi7T4fVin
ijJaM+R4b3dIEtmdX3n8hC7yrkBt6kkQTy1lZY6ol5RdzvwkCdl8OnS/fKRvw7SZltNNYew7XjsR
n7t1MLxkQAEquzx8AXs/EYfYjbOgDMuiKBvaW8NJzsF4Y20i7NbnsAtwqNwrCcDrFahwjWHHREut
1A/tde282WtFt+dx1UTv517/Lbql92MNROeCauVV0xuZ4+1Qd0v6MiyLXHXKh2o2r8pwNW9ehctv
nKXNg41c5EnJ7/m3D+p0a0/Opi96sin4b+zwTSm0JJdAqo4o0D0bqREBbxUjHBnd8WGl9lwz/lc/
NoyougZxFlY1l5ZNeHbcZ7xIkJH8bs2Y5ht4Lah/HMqFv8UnV0XqU8oYHsK6Fmy8GUJ3P5i1XtCv
FXvel5QpEGzHM9TwNS42ke+pTd47bmHAojN8qWWKnHj2wPItv00mMW+j+EpyN2O8c6zaKBmmStcJ
Ks3jawDvEJ5r5qvNhhtUBF6UJQWfqXGYWzlLSsrGqXEO/Cg05+aUWdSGM0nWAvGYq9Y7TbAWgqed
b/kwYRhHfuGlhW13J8K1OR9p8+yj+5/7ALtSL+WJ1uijyS2RzSl2Or22wTFtoCqRQmts9mMmAEDJ
Atsb9q4FIQ48lLRBJSO9TomVxGv+lpZuT+VeDvHFVLDKi/+sugmHyqhoJZbYPkqNEXImOVEy7/NP
k4hv0jYrUK+ZUBzw4JgDSy4HMvoH8hb1yrokzq3eLmasoVdEgLnVp8tf5WIHyMaT7mn0EJLPusj3
mrSQ2tm5y4igrNF8DV88eSQa3MC3wG9xIpWPNOQCiPvVOWH8ZVCdZR6E1v4bziz7BhPawCHrFnKg
8oyFaDf2ze9+btMglAJT0WPB41UccJcbL5VcWIBGXTZ3nrb3+F80MkxG2DZ3DM0XzX05dZ+8+6tZ
A1srZ82zhnZsof2lFGZTATXFMB0ti4HtuHu9l749hBeSEol7tHleu6G4LmffOTN1Od6DH3IR/nY/
NV0V3u1KMZXsD7539rI1OB2SBN7AVFbhHGpLhYJLl8RJOyCmcoabFqWXiraEymSgMdav0mgEQRJm
zyrpXvAdw2GoLBy3fcOg89/hDAhPKY88RzCiYHkAPHXj7VsGSXfL5urCQr5SOMUCkhKgpYJLs+4z
vIOIcle+ZhbhGBSxGwsoGMJb+QFPKumjXTqF7qYUGAK337I5UjgACdCQHuIWRjR6SxzIOBC96HFK
rD0eijjOuucAPlAL/u5Gc/IWQRyIF0yrJZNuO77AFVPaE5giEulFd5aYPFqYb40qX5yV16NTHuzO
bAG0xcPnXURarRcP881c50nFLTPM6gtziYIGaOBrkH71ATNDFSr/EgkLat/GfZtmHbbWLLL+/VjW
rxSeQpFRimQWbcijxS1hAp9lSSDkYnPXbU1edZdQE/Z6fKv1wES5GfxdWSfkAGApiagzxsKI6Ojr
mFfQxfQ6ajN2rtak47PgNpkV4Y9ELf79kyY9h62u64JnZLVoSVBG0w7oQcaPiN5iOadmIZUDs6XM
c1J5DHoXBTgFHLuqoITH3pegNSmmB1Cedb1u98yOodPW93ZweePMOhHFV65U12SW5MK6T/OZqlt/
/oAIz5dsztFVZi2AKQ8Gfj0J3qyRdje07d4DRw4+53ZlkERpW4bDhu2XZwnY7P4IozywNoqUI+lh
GSlbimbIg756nuD4OD5smYlKQ/akEzPQ3WoZ+4RUYEmeKEhFKbHhNoJ6kIBzawMMylYVDbcWSAFl
BmfEmT1/dihQ0mQO4/vj9CZk30ZLQfZpogU77yy8seEqj+hudepOGj+d2uvggojf4qKEXcM3V3uk
OunpQOJF6osFYhSOc0+ISJL2YKqFMfNqJcd22Zdyd7BDLHq22BmapxEsXCudCPyYvacYjhq0H6y5
wvYsJySPx2kNzlSVom7s9zBAYmTCaBgM73ce7iOKK3OrquBcobcvrKKaMOBY2F5EAiHIC8yc998v
9mv/ljASyiMbJfCVdBkzds3iN+3sMi7yf/BSPbVmweWdesjFa1Z0+phoZPfperUtJCtCzJJAZM+r
YhipoFTKRHcrZZQ40+5m3tb161d5SYodI6zg5VcnIzQc2ZlxN96kvNhtHuhqleWsL3R8Kmq83l1B
qWaR+y7nfhHaycx4tSb70frTTKDtmu4oWl+8rWr4UBPyrEuKyUG1Io7LWj+8OaoekfULj02lIF/Q
NIr7GLF3NCV77bopQ1l5LfDRl9VLf41YfzlbRjBdFvD6Vw2UI9AXnd8+3lpqB90vNhsQKehv1QZd
oQVDzPbjOpUW2cBjTiNQaYL+6dlIZ1ImwVM5b1X+fKX4fF2zi5ssTKkbZxSu3Q/+0P0gWnnBghs+
1RgxsiPTE7bUll8buO0174ZFCKpSK/tf385fINlvAdWfUSWo7zBlfdNRewflanmMywiK9QFzm+Q+
eEx+z+xIql29En/ZSgbDrTC81ycN112G7CJ1AwPM8CKp87oBlQcjduTWTEWgL/znkf/9LTf9kVsR
OvNDe+Xy98mDCwx7xt90HX/WETbH/DU8cqsw1MbGc9TP7q609JlyD1Q+YO26mCcnaLcnVFhEIXGl
8e0FLRrx7fkBG2CJgBPnIeGkl5jzSA5E20xxxCpusWr6esTrMNTla3bjjVGxzhRc0AYIaWV+Fwhd
erfYhf248KPI3S6bvC05c+TKiRB/6qlbk7iCuUIZsPl70ksTkAcvRRTH/Op4iJbxOaDiud73B6W5
GmIJgezhxN+70c09KxyKGGHROA0+OK56rPhE2w6Ipjx5mMdVt8JViajqnVXGK17kmCPtINHkThIb
u1+L7y7/cZK+PY2tVEWMO+FTq0lgechOW3kz7P3q9rYUEVHudwC1Srrw0bdv5ADmll5+DNhGuyA4
X1ALPqhciUJKHXFL3TTawm9GBfkdlWZmARU9Gut6TRDetClvpLW0sEDGwAbi7CP4lZ+FQIJ3NBLE
Z0QQquChYJkPM4tGSAh4U41y7hhoNTZDB5n6sN+I3gMVx3+aNHd5AbWLjTmWCaJ0pLf5z+DJztyG
3MNJY/KkE0O/8POfbcxntYoVHKldhXFimdpVGVdaVjX2xxIDGz2N9ERuP6Zd0HanfO5WxLnrGzlB
jakjlKUH/60F7hfRBMkiKaadVDVzPsDuJvAbX/kik3rWXdTu/pvdbk8b/jt3r3xscplbyWyWug4K
bjI6dkKeH5LkHeIzGb2Rr6NGhVKHj/oasSlLo94U/nN2ecpPbse7CBXjDCGxwP6+jV0ZAJ92UIOG
ZYfHyP5AlddVeRf8UtCW6+OnBIpfm9SBnCr7GUB/caiLxeHrRvHvV6X24somdFzMFU2jczFnmxjo
29v6Mhf6BESeVgwyUSpweWRjPcMzsc7H3JrD/cLnU1x/81xJ3Pp4D/dxsflHPcF/mBNYI/RtR4C3
AUQOS3B/Ci26Gux8qa3Ww4tIWGardwPUZoHRXR6mtQ51DFwQiKsXgkxPqMvdjAhkcRQoSj8yRlHN
Rn5BA70hUJfjksi2r3EoTP5gWEFmwgajwOMBoSwDUU3w0VUkKuDQK9BvY7gNj43WF1fhhHNCWGcV
4sV18ng/IdLpRY6FdQIl1296XY3Sg5PrUZ1KJGJoTbgXmv3ogVetHhjLT5W7U045qi+TeqGjs8C1
3PRuR4Mjbek9i9lkq68VG4LMzV//lTA2rqvOxSRP1IYRpJDdUWdo99VC42fVn+/jhnYNKkf6vX/w
iEpnwyCs4DZoeZTFCLmoOmwf4WHE/NNb5oWO+p4eLIuNWA/CCad4ceXsGGLK27iridT/KoTZEhMx
k8BZrMzhWZFbRzsuX7XsozbLeXWpnrFC5OWe2kUcRVRF7kvOhuEm9DyA5o8A3mENT4N2i37Nm9Vi
TDm3fweYTU99YmagH9ktqpxFw88QrhKbAFUZDXJK2er5Uq5O4HJ/yLm/DLK89Shj2nYWiB1JYhbu
nDvzGSRlAcXMgddMWfPexQbRYJYPb/9wiL/NeQD7EcWQOtezk6nq9vpaCazYzpBei6RYWHVCOvVc
se3lQ1cft0mpES1lHKSCVRsDT5dIob4Jzt2q8Ubii9uRHQcuVa/krhMX6me6Cf2qZp8VL9X2nPTX
+usX8YVeKx8jWLA2edu3sJps+eUojfom7Tnt4qVIRD2affAovtMispAPvRCSaOP1oAKlZ/rDn6uc
qVvdrKC8AfUCHRV2SNY16MsMFxhiAbdK2RwZ7buXl0fGQHu6efCQsxasqCtRVu6Qwlm9gRAh19ce
f8BJ8KbCxG7rX1DdhAdplX/W0R856p+JAn9nbvofu8uQfngTCyjVUloAeJ70P49gNUYIXbBXpaiq
rvzaeZrvTJHmn/9RfE7U6vlvNx458xW2D+v7ud7+94LqiarPckcowF+dtDqb5JEOtquGFTJtdrMB
oke5zctDv8O8f8x+8xUrzzLSphi4PDSUn1RpuWAR4xY8koshRvQb19UI8Meag/E8/plEs0ggvoYn
TCikaqNipoApvkkHFcfy9Jy6JOo62l/JDe3lhTmAnvbMp+L+5pgY1G8U4TfpFnKKIH0PAYc0v1PC
t0HjoGIQk4N2oumag8cZ3tcNDzY+gray7DhlqOYAmcl6xeSfusJh97j8gIrECQzcjhdHjS3uGfac
LdOuUp+ZNU+HUlbxT044VVZuv2dN6lVvL+tiCYzwM3VcrTnmHOyoxjbNKHhh5YMNRkBV5IyiGK37
XuBHzOaT9a7NpOzcsfutRkLnIwiTfveiXmk/3f10ZTHP3kXStwTei9t+T7EwWvoCpmtVT/LUh/0f
CFzIgYRnOEFoSUkLTteM8A5/AZwWydjWm0Ypk55pu6SuoLMlS6a5VAqE+qmwSgkOKEO2Pz1VMiPw
Ab/r8XNOrK4NQw5Z84zxZiK/RR1z39Pj17nchUGq80AIGQw7xZSeKM41OcqfvA9kIMgdoFJweyoX
BcVkva7KI8a5DaJ++wa0lneRiHWbJSUdE25Qmq+dg8kbdSHnrvOkok17fMTuAXgB0wHqHCcXUqHE
cFcjK0ATV0VRB0M762aJ2P8CAgbwQD5sgyiR8NVGAWRQWejC4kdrbn80nkswXq6yypEucd9MshF3
MfZPj2Frqs9J7Zpln5mkmJPY4tKZbM2xBDFvXNYBtJNGIzE7AvZ+suyIUfGzrOFDY/5rsARyG5Pn
mO26KuXMj/iA/HhmnIAJsTLz563GPRSU7s6G60tUoq3fXL+mvbMjqqdN2hz937kg85n88CFe4jy+
xRMlVO4A/hIpopCb1vJdt77VV/bm5R5C7x4IA8dSOIxuS/J4uUqVQDy9CRTSO3NI7STjTHujd/Ar
IG0NIyJtO8NcpgLmk8YiCK3ldvYrklB+2cGcrzZDAQZM3iMJxuuunA5psPo+r1BfpmEEj4WLBs35
04LpvXDKyg/LaPSyznW0p+OL3rn4NeFrvrVu6sWSmcWdZSljTvHtDat6n+tIWAvtmmmdcWsYmL2z
v7cW4ks8rWA3VQMzhMuI4ixoavpdNc6B0nbOIFsoummLppmGmwUr55pfsmsRW7UsaFgJy8hUKBfj
UHS2HQxEjf0BSatKP1M06mfVeNErEI9hMS7WlMKvYZuMHxxAbDb1kQSXDmY8Mn/MNTcgY4Iijd31
2U9BsrGrRByhwUo2S2ACWe1BYAb6qYALuALRUwG3zmGFDdLg1uNJS11WwL0376oKTJyUaFYgmsy3
NqMp8P4/SstzrOOs+Abrs2Ki0EH6cBi6V//W5JT7J74iH+DKn9RGjrf2g8Vc+vyKad+WR0rt8OAZ
iHz4tKZCRbYOM10iFoVAIN4xMpGhH1I0U/PBzo+UNUxsT4b45YfVLF1eBxyTwMghSzg1r4dKTOzQ
+oygD+klbeUzQSyKuoBzaEi4Do8MTHCqpsPvxLJxb9CuuKvvrKQKnCyN3obyQ/7nPME5pIehwu0H
Loky5wj4yu5C746v9ZsScIsfnYIc/OBREwGes29tZyboLu4t7a7rnCGyI9J1EbKC5Q6P8Apns9gq
DtzJc4nRfE+jjnmxMlxk2VOx/0F3D/J0Iew3mjVeV5rasZlElVmo2QXaQVQcVaz4iqO7CVR6ZMol
MP20lMjKv+XyRA5rwmHOyjteuOSecma0bWtYwFKW9UqwYvhl6zCqIr485DJerh0l59po9g2rllkq
mE4/LZ+F2VvJeek01l1Mw3P9rmq515yiGCawl9zhy2TaiJiDdLfDmCFy/jWhsZmlKJTMrjTFtI+m
/sKBoFeTWYnrV22T4nDuXh/Gf/rluPd3Bp3aeIkdAIItCLFPBoz3WHT+JAYcP6nZnlL0LUd9TWAY
igMrs1w30FXrXmuRuO87YchLa/53YKxpHne3JQzIB36QJTwOyve649p9kA0xASLzo5MpjwyJ/OwZ
8VXhgJtS+khiezdsValU7HlZ7Jc4uEK2lIRN0V+ZSwvSTSsXj7d7oita6O0LLlgjCMVbSGUoPNls
MxO9oUfNzu+3uPspH/cyBStdDahCiV155b/Sb9PoJOrsF6nzqRMkyjtkVeKehkMdje3ncHWaroUY
Swy0Vjc71CJLFg338A5j6K311IlYg1Uk2EsgtmaZI3IQ7L2yc97O4+H/MOA++ZXmUvFdAce4TFkI
F92AOOD0UpfglWymye9GTD8V/B4Df4KXNTlKaM26eM3/kqsXHhtfLp4dbF1KwX4sdMI0FLB9Lwn4
4apl1dG7V+XHh6vDYUJfDDoO1HKvUUCKE5v2To8XAh+NB/9jYQ1hos0CXiTRwa0awfK+dPRKnKni
bexdC/bpDn273m3D/1gnnKgEuDHt464FZ3AbSpxO9zPf3WYiqW5qhMhSJQqY7+9ttJV00B7Hpq9p
sO/ENTanRMPPemVTZqjL2sOTiHimqU7KKX92siGz65okOMndcL45CWkffusDORmIoX2R35WZJGNk
EW012GwCiXoBlksGGmxgIv+9vhAEXWWajLavJgcLRInzZXVgJVnBRkFG7mkOnQMRV4kZAnZTMgmd
G6UImocELNk8A7oY/7VXQ17QBxsYza3BJ+Xe84OPAOu2oivI4dmaeJ0dJdKZ+vjzIwBywfh1/RCa
6dnngQihk5H7u34D0NJ49RTknA7MWihkKw/96EbDi66qcbA4TOhWT9RuOBGyQe345Ju/iX8djpzM
nC4eP+EhPiZT2lw78c17JdiTau4NBzjdvo65Q+tdZC06bycUTT7RELzg6ijdSvG+k0s4iXZCYt1J
LeQL590JFSb7cuZ0Kr64WcWuCAp4L0QQDqdCuBlzPgKNGBl8ikQQxpCijh6W9PA1P63LSDYL+XGe
6hmXJnMqm7HVnL9dtWRSkw74JhwZwZdxOVzIMozTYXRBkgkedZPOsuPCH9W/hAl8pGj/hk6FVqKi
z3EJRsMKW9DGE2SCgakFcLF86vCZIV91I+TUGoJ+94L4iqCO/blyeV1doGeRLLSuaHQivoDGDYg5
KlVkcsiLgS8y+GjBwbyjtmhPdBxQvhtMbDsGFU/XxivwKTaY3FRaooh4Yqj6o2isByP7f22w79it
P9Bm/pR9oUFF2DCIfZuUXSdWJaUX2E7VWsWN4IcxJLu1aT8m6TOC0aTCng4+q6YftStCqr7tSAOv
uYDmxi+I4bRwx6dtXrW4x1r0HaWm3KoE9CqFESTewZlyMeiRlHRSQ792ghWGtwYeWvNh6dp+B3fP
fVRsoA0VF7UXfS7mA9XdOe1RA0TzSLp02v9+65ofqRRjWYrelT2FFAfZNk6QEmup/qWMsAkOzxsD
pfq3FmRZrg3JM6n5LwqJU4xERgp83D5ev5BgI51aQ9Sal1KpS5eCsLIQgU2MhKGTy5scb8brkQB4
5hJgM3cfe9AMN3Plzz3d4WnvckmdPXtlXDSO5z112XoT03bzmXt/VPosj/XneVarZnTmpidUYd9Z
01szzxqTMskTC3xiWABwx7vbJ2AqA4t+HHqEjaGK9vAFDEEvESFUtRXuE9zp9olsTInxxwh7MVFf
Ex6HnFi3XQLchus0V0+X9FDOsHiAIrt5ItE9rg2CwV/t5eZGsIgBVbT//lNyjLwkF8uax272CJNo
eER/zK7rk5pEPo0akgpvjPskzlBFDGu9m5x0nZzcOA0dJEue/CQwxnytZDc1zs6qqJUi12UA6atu
ohlOMDxl8WRRKB3HIWXr2ggeTgAs4xcwWZh0f6bV3NVbyWbtbup44rDuJ64P7aV35F1onKrubmZh
KvWWd0Os2r366yHmKzQVhSA3SW1IoBFrCA5zBsBqN77O1vOYBp5JqHBcMeRBI+2+vslWc+uBUppo
yycNLx+F78UTlTfy4oHLigvlO1VLOWk7W1WzGUGNkhfKPjVit1Abg12s3sZ2iROh10nC5F7Sid0p
8Lidzh9ubyPOQsC02cTnP+0fvCG4efgJlDYnhRaCtn2Me6TDZbub/QeXDtePCVvz7FPgXhUH54BU
ALrNlj5WVsnKYaOLxJNVdj1LhHwB/yosS/aQSSODkZuum+aW9u0iK7MNCqD2R72zdYzQOfVDAuCw
Lho0p10OFpGxRX/CMNyeoKYuQKc+I0uLcXrAYKi0Xh2+UpGra3WCIhAwMZGuepSIiCBge7lGCTNZ
ZbqJ30Nd1EPa7ZvlI/7HxYM8sXhigQvtnG8vW/4STWtDzLx6OV5o1uHrwZsasUJ1Do7R3z8gywrz
j8vLhe5sJZnoIICHgVVPwTQtLVj/v+oqh7fanHScBUCIUsasUqqgfwWJrZwF4oChnyvFe+m31zx/
6LC9vFuGnIy8jMV6wlDQsOWBjrMC/5pUMQ17DmomcyRFHUwmhLlRCiKoqZbWyNiUpzCOtMH1Ydmp
F2GOjwIq8luYGACj00/GvAMWqJqIej9+SOWlSvOwEH1CpB4IqgdAlNBj33JnSYJF6qm+KnJ5gvY+
Vy22bPhLJoeOQA8QqY2Ip3948ZmL1ArUgxpl4IHDukHYsA75BQaoURcYGKzsVTV3BaEjSZ9IO0we
2yPPoqK9VaqhvuaYyNdyvzielS+89fznpcMTbBpqs7wvSXl5F9SdFBxitPTcE12Z7WWFhqIe2YmY
nhH89rK++kA16WI3EGA7sWNidhB3Dtnpv2lMOp5rxpCCqQ1+S/EXzN7nmUk8R7CT2TdlH0fJdeST
D8NgLp5lU1FvS6uF8IbPMRcIz19zG07nYRlmvAkLVMIfwZmE9kOh8pazIaLlV8qAhuogw0q4n2iA
R4acE9WJVmsYYlZKmxcb2duiby1OStmjy39REc/absCKv/lypxxstz6Xdkx2EnbvhXj91Y63KmMa
LLF+mtnLAzbk6UJ8DxCCxec2PApI4Ma/RSGFpZVQcldm32WKTXPeyxysWPSJ0JWXJ+LmD3mHuA6o
uKaDjcUVLBqN1q6BC7VXRo3TKVk1XPqgQ8bo86qgpMEnqxJ0jlxtgeAPbUpkyKSD8oCp1fRY1zBW
I/CBv/M7OUuA5PWFjyFVxgFK4TK56nhovesFDHR+dTZnYZpThKA98YcED0+zlhJxJvDnn9NuRbeC
Tep6Sbbnv+6DgNI6pYC+UND9MKoL/HUkuGGq0GAabWI2tm5FKzAg1NvLTY/elYKOIyJqICLv73n5
S0muKD1IfwFZtns/6WEcs7ozDI3OvyRyQoQxv9hGkdHjkZYSRvqPiiRulajuD+Hxl0m2yVkl0cOO
OAOB5k5o54+yz6QRb8ZoQjYZ2bcHYNMOUsnZIj3XVmwhPzgtwH2anH9/Vj3eTJrLVwl2fLn48j/B
XQZxkamsUyj9/ulnreJ+CJID5LwislTCHOFSKv/0NkT6lkTP4pOFl4sdyC1eCktX/xVphihXMoiD
tAWWXSVpvBZIbV/+Am+Sm/f5m29rxbrR17LTFt4l1Pm1DnHMxe8VDkMY43As1RgqI8CdeC70KDvN
CyQdsZSBzdku3ZyFifQix1Y/ZSwbGjUvBQzjVKHDhWh8EA/vAdNIzlZSj6PUG3ZcSthOLrojwYz8
eGIRSXrfECu65YjttpJyKe/utEskQlG9lg3kDcnoZ14yGNv/En6X9KOsOb44Iiit05kZWvnP8cqu
MahqcUiXXvoa80oPTfgEWVDH5AuvQeOjmC2VZ1WenVXOX0T3OwSXu/UtHcFC1dz5alJT2qeAhGz+
/c77e8rB6vJVfgrVmHe/feO2HDlGqPHxq+S1CATPV0g+2wPunPqFP1OBu8dRHv6KVo/JUG26LPVE
jptykV4R90iQf7IDoaRPHcd4nML48qQ2RkdNfHS8Q1iSBVCLQ+sABu0hO0TaZn06ePn508EWy1UD
cujPJ2TQ85e4D6Ps1Z3UdmbTNplMLhJ+XykwT5WHxR+wmYkkusecsOPoDcThZLY6Kuj0/xQlJvMu
/aAbltOCiDj9qzn+92dCvSQ87p8zoAPtuggssKrnV/xgzoSuGMlEGVhaWbCDg4roo1bm1CgelNaf
ykyIdP1FuKOhgeOew0mk59rrJR4zT1bpLheXHG+FKpUVZStMqdHetYSYwNruGUnjVRDn6Ul23Bdx
NpKfLclMSjwDUi2YOWlh2sCMtcTB08lOSQf6EFtirkjfxKrThlO/xgsXDXRIjQOQn8ki8tZ4/JpE
DAvaGuA3xi3J09DwqazHYsgWtez2FQH/rAMieTELJAH5oWkG17x905vFOu6fxIPzsD8zeBy1KXX9
gEb5rqSTPEWLQoD4RdzvfJ8xiyZDlPTcBM/eppbhO0iXpbu282veePw+8gLnWIoJC0euKFgcaV6r
fDXnbjX/4ThcrShGhw89IIhS67GAmVeXYvTiCLvYLPGpXTK6ItmG8MdK/1dRlBdYdcVp9/Uqvgz+
IHP2C8Mi6LKPUAXWaFipV5+uPAd5xm37JYlm0dzu3lVH8eaLPIxSFXurcohmgjrbR9FcK8310mPF
eixCkP4R5pJ3I0N1pkNjHAz7Jz8ReUWBt8eoFP8G+2p8yCdtwmOPsIO9+6kW0oB0Fqdyu7Yw4w9C
Hi5ZZak6qbvcFRKFZWK6C9gqUa37Pnnd94BVDUGiJmTMR9yYIe7eTFsEDJSvwnOZIplU/Agk8axw
0BA04WKnxGSvM4EebtAGMXxEIAyLtn0L4THtOH28k0D70giBFge+9/G4IbRGqOQYDRuyqkA9MyYh
aS80E0G9wZC99OIoZWRZ0SV63wZVht+I0Nsk9JgqHfHvjhlXTqb7ecIKo8tKf81bTHmLVygJhNgX
5OqKZz6rsgk426G67VX1QmzDidtFRa5tA5If8TeKqRnWC7ysNSkdHFDW0JLlf2WHGmkZHhWtx/1y
C/IYOqrDarbWRbHkCX53XAQB+yVNJFv8GcqmcbFHqD+vyMTsEc+qhIjC1OEpsJyhAQYWCiAuxdn4
ttwlGE3mtvQcJRfG86Z4YLtS0Rwl1vWQMEUduYfYCcUeIedR0t6vTvsdK2JaNAciI7upSEIE1FXO
ZEDUC+GOmjcI71y/e4fmqyEZrtU/nPCpxaXd/r7UMe3V9JHQJRQ+Aa0oggt/n8A9nMRQRguO3FfZ
fVBhuoCkl1S6tmE6WNV6YEWc3V7C552xJlM6wP2Z1w6pSzlw0zA3ShxpD/PpnQHTEWhTvgHcVY6H
KdF8+v1XAu8wr84rEFka7p8aLuLJM8sxBfL3BGPRavW80KKzFURp4HwYM/Uz45LZqhOOCCZJww1q
Gjxa2SANO+7gUO4/cFT1vRy7gtDDbOKcfzkrieCBvJko52Y6iHjjrj3BwQ8AW6YC+dl+DMkclYq1
Kur7RHyRSlVQIaqmoJE74kB0YqdYEcesEQkI4MHzyWjC1CTtBPwf+A/rMqfE/qUV2HbhtJvdcjdW
op09XH8u03P7vEkYkWhBTWVIloQ76EXR8yfWW2NUToDFU2orUiVvx+1xecu6aKUKZ8LyO3Eme2ut
Mh7bn9arVpP0lF0lDSjdNM+a8sxQW9p6x8Rvpuzy40beJA3R7P4Ou/XRFkI1IwOlNXZ3q/rr+PRv
rxQyi4s6+PCN33ThUZ99LhQAIpWTg4kzn8Fj31BuIDBf5ZxL0PW+FkicOrTErtOz5tySU4jmeYuD
9rWMBroUDwH3wagGgrI5G1GS8b1fMdFbtEgzPXLOg6jiej1xus5F71PukLm7rGlBh+0euIhftX6M
1Go7G8UwLcwf1TpgQEzX3zuFF2hiqoSdngSEl2qO0GgysIRHQzEZjyNzHgo+INwDuEazzBTJcLfs
hc6v2D0fzGKen1SmL6d6dAwyQG+lwYQRdKke9TC7EgCgH9qG0GA0nLsWwGdEHe6uCLRzDHfufBL5
9zw4gu8GU3TKSAbx8PLty1GhfsFycAp6SEGk8WYgr1TqbKwT+ad9jUC4h2ffqOVBcQ296Cz8Mvzx
RTGwf2aTpObq7pzAaUksbL8vhnL6uxCPfgpXgY5YaCab2kCjPNJQC0AvR9ZWY47pHIEDXR9NHYQ0
BntYAhkPhaRKdx4y/vFu0M42DKlfsdAFFUGdDOCVzDctLBt1On+0uxezv8iQcKQijsx1EzNOmycy
EIHojM1tdtx98/+tYIXy2+TXVIR76abngbE3MoAiItpKc/scz0isrFA8JeVORDuYNImocmsmBCEw
jf4WtBhskjBfWRidc0mx96zklofFew2sNGDzqQOqLnjLlsy7HDAAoOSQPUu/UbYbONK6SFUSVQto
e72wRwVkZDM2qy4RJVMOlgBwdmvwJuHjrBo32Bc+s3b3hGiMZiQOwM5nWnPxaFdryojNxcc3PhGr
/HCeZqw+uhhEJYu8UPULz6B5VC5VYb7b97TW8uICm2anef1Xc/uF6bGISfbZFPM+c2qidyBL6FxM
JwXpRMehGIxqwmxlbYpPzj4yF1FV4UTtgVUzwmHdHBr+ZU62EKm3hmyKy02vWHnebXwOTDprD+o+
tJmxlg5vmcZ1TAhqG3xY6hN45/9FXMGQWCDERjcOsEVoU3rvziLaRYuRqACVgB/SzjwuzHNQt+HO
v7zR124V3D9vOtMPA1Ottlrldo4+mxFveOm1tsHUjzhL6+kCAbmgIi/XJbN/HwC4fAWXZ4Y3+hGS
MIMFxU46DUUQJmRTbjPckLHZUYUVWRN7ncHO4bNn94gELoYVAIo8lT1fwxdfwl5YkC041j5QXGgc
+13KqYuAbMoj7A5ELDmiSBjwz397ywKWFF8QO5WajazPGWEgDVqCpMCMojSE3iiHz4iT1aa4AwFc
2y3cPJ5vZCW4BG0DdDgvalY/O+fShTlc6Hdo7GMZozPJzwxo75tIVXfMRaPoAdR2FlNwDKOrJOfs
PmNKL9j3CYUxXGhQeTyUbgcbqSXx0zX8wvwSRkl7d3c8jwD6FpsSb9cEo4qIcDULVZR3irw10uq6
LlyKRK0jwd/Yf6plr7OByo0XXYnZiIkrH5ViLZNtlj8UmfJPuJT918WsEKVi9s+FaoZwucmXrCVO
61ocdbqGyvTqOR81h+CJE/XxTisfxKeIM9TqIZRIXZfY0/jOMWCOMZmjToFDNd49wZSwD4stMsjv
SqTaR6k2DO+Jvo4ENpi/ruYGygke5d7af+ukKDT0A67IsoIr66n4jfd1OysH1LN9TnAy0iPfXBtu
qiqcqHJkLzouY6q4+YKtU4U0c/I4P1ruFQPnV/KoioMMJPKv5eW30MZJORVHFL8X+83A83Ims9DM
1FdpESLP9Kd64SLn8D2dmg7DhcKYrgXwV9D0adpTk6/UEC7EdM0oDhYh2xOtgUOnGMFKwnRj7puJ
3VRr8MJ9mZKnKKZEgtFFoI/zzhDu2QrKlrdYAx8ReBSpIlHyOV4nHQyrdzkdvzxtK70eZ6+59DZA
CL8D89n/WMwwuTBwHPZyO2DHRAoBZHP78U105U3MQOuGCSbN4LZDtg0vttbBJJAXGIEXLbodpSl9
Uit9MZjQtHtk6dAnvizdnLfcvlCVkbfHqDt/9L5GSu4dCd1oIoq1iNNiQGF4WcEKjUcDexviiVxF
9cFes3VoOaZ0S8RvpMBhO1MnG3rvssKHnrPKbcXgqa26sPyTsJesXTcBIK/f/9rIe1+9l4n8Wexz
SnkP2DKMkq+fRGSHm9gPURrobW+e1kDIaOaR2rFysVcwWIadeWG7aRYEC/2nrTpxvhghrpd7gRaO
QKoUliemSErDw4reqVe0Jc8PuQDwzmeVMPz2Mn5KjNiH63dPd0xg2UMCIGLLKCmGssd7m7ELlZAn
vpvUKl2XkwOIE0b5dOAbLOCgGyfmEV20NdL2R5ndLGMu0pKBXoytV/fj7o3OEY48fsZ2Ds+tQaBw
8zJy+IQ2w+RP5l6tr/Lkf0VG/ebQtfthFbn1OUEEwEG1TbgSWbiLdeRW/kexPDPjcimNy1UELqoC
7hlbK/qPeHr5DAgrydKGXwRpuUAM8A/Poj3pbZN76HbxFyqocdh/ZIkNMyIBTVCdxgwtPjaSdt/6
LoyTg6o5OLKrIWr1CEm2GcJYOt52F1zpmUe++lz6UiF9ayXVZcCPzEPqN6kLjDOxaasb48PcYpim
rlEdE6Jw4au3P+V53MQccLOp7+C+BYEJ+qIC+2f55HIWhtNwlQc11S0756ZdaVMwIssTjBsNjNdo
Pb1GQYeyWke2pArZmLQzFlQcd/BTdLdML9NXe5uJzjFDG5iitDf1Qw8g7JsGkKGOJ+6IdKRj/E3M
TQYJ6Ckg7YcIhazLyTsKjTLDjIPea4zlTfL7Sivt1O5a0zn3KS32boM6tVBoJzTnfxnpu/6ccUT+
PhMzJsHCzOucziHvgs/fcnlXArTKKX0auu/1PBxFuARgxvQ8VKem7SbZ4A8kiwibIwd8eT7NuDQM
5iOUln3j0WfNyaxSTz5i1ti/v75catnudlMZ4qh7syTowiVRKU6drVbXDBsmPzAkb/4ljHeOwjNw
VdJe2GImQ7Mzr2rpW5Lzy8lFYNta9k5skDUUQV3brOwIx/Rz/1zZKy6FaHPOtTbNkp7Lh4/V7EgK
eMoEKMnZ/AVRrOAgAV53LoMySibwf4BhWZ4lW5oMJz1p/dOhgzHLT9yegqSce6vSlH5JmbA2iyHG
Wp4uidCub16eQCgW409C2WFP2I7bxqhNvhtVKeXBDyIT4urOrnoMSow0mKmSvTHBDomsm4i5iIDE
1Ykfyho6SEXwvJkjwZDPKhEJjraJ8s9RCoi+puBvgOZVRpsFGZpHtpSXHMY15yJkPVrJuWK+OSSV
M0iAv3n5cHPWY4IxYoS9vQEWh+9fm0GnLP5Mmx33BhtU1Hs+cuGVH9GxQitC+7LngNO2YbOncLhV
bzvfGtwwiP1yeHyfpwgl4F3q3gu6s+6naeMN1LiBv8uvLg75bFRpK9/PqZGbVJli/91s+dUgkfx/
LyhexGKRa4VcLgV9mqEL3rI7bTcLHNUmRSBesywXV25XfjubH9xpjzhk/jztqi2uCm/iB/+/0Yc/
Nf+6hP9r4cViramEPIjRWEQ5/eAicXaQEHD9C4H8a15TDXgEhSpVUE0MjeTAeE+s8JyYj5NaH6L8
kullJpJqNjSafOxOCrHRMNLaUIR/TU2Ef4kxdrJ0ZEgltq+moGsAA4MI0/Bd4mJWT3qCybdB38TI
Kd7Nx8IO03KlOEZSvZpOnupr2T6rvZR7EWvCAYXc5iLRntkq+Gfapm/iYfaGFhYn9Q2c8Tpm4VWF
1eM3UnlLuDKVz4jXk/Xup891P5PptKzzkNnm/9t53tjeR3NUkig0fzaunap3C+elK2pRKQfvUuF9
LLDK6/Vs/GAYzrNc80jCVY/gHmHuQUgCc98qYresJ6CyGVVIwmC2jEBkWsjipobZQCZci7oZ5jJX
18X08lL66Vg9yIXvKG21hqKNSDu59+tccNe/qVQ47FUBUuYC4RPVWEPv37WEl23r6b8Ag/OSJr6h
qoqaJVFOFYlt1+sQNu2/5z5uWBfGiQCgrR3yDZiSOi1SxXrECXjREfafKAS3xUYBZq4Z7xU2MqBH
GA2veSCWbNSFMcZqapOLCVxtQe7ZWig92oob7bogldMkB6sYgzFlyrR6awv88hNu2yo5we1yGyE+
mWUNMQ9St9ROgpZt4H4mBnk1EkMmo14Rhf8noq7GOt8ErZCaVkT240BBekSed1upDspI2UE0s6Bm
YBYHfSRZkc686od89NpUF3TebLarA76yRBkROkkuIATIzrk24elWYQzvplJAOQtzd2xYa6mtN6ZF
G3qMgOdxhGnd371fMK3lrvEjmstGs9LQVY5U6gODEgsIpYkh2Nt2j9BMA4HQm9dXD4eFgbjbILNC
5yDtyQKdcgGl6dLK4FB0fhtrFr3gs+Tr2/uuRSa0lk8Zj36eZwqc06MiCrTPiwLlcywhv43M2PoC
5Mo56DjncaRpHYQFTA+c8/dNz/EBmxIpHmXZKQF03eAoToEfsG5ujqi6BsDbLCGU6ms4xTqbvUAP
kNMZIP1mLDXzfQEfGyyHVqaWxf7hGi90RiXxP6qDVYUNaZZm3Ligl/jgl3q3nYG7/5dur3jwJvEW
EqFiUzM/vPlJXlJC7T7UjK8x+KScwsuB7ukJSrtVMBLEUt5PqHZVKUYRo58EhXyre65OSNomBh5j
llxOnayTLB3i16V659Ia5f6ZkS+aEWza+opouFayjR1W49YANutSO975qDOz5KfRBSFlPbFb/3Q/
vsZZs7Qde51VTCMatixEdv+XbwNqp7BJdF0srH5A6AfKLkb19+8C3WUYH9MnnmYB6P79giCPbqob
EzXo/6pjPzuwICJJSLsvg6WseCXmP4YLKNX9Rad0riozx6PSGjUowgWklmF2p47r7zWQBd4Qlm2R
5ZOteO0VmhsNXA1vGmUBpOFeK433VxBq33cu2P54hBRrDe567YfY8KUTbd6m45fvPCibdA/Biarm
/KhIFXWZLdZCy520mrDhOARJ/SAFk8tti7LI36fL6CWecwrDvrLJeZ2R5rEAKSOhdw6e9JrsS09e
UXwOsIl4jVd7qjm8cMcUmwY6kEej++UbxlOl6njk4BW4GlkSB1veBi/5TxhkthEWzGtY6N0IdWJk
D4Emb2han3oKPgaz/fiPcMbUUl9B275N/JjcUdOXuRcOJ2oB2xOIceTcpNypIhFXLEcIwCSeuYQP
wTqKLyKKhvwfEMYHrMCtmGja9hAJCXwJWy0Txz3mUKzux2+nHx8fwni1nXkTeQ7mGMQnSgmnc2c2
bMAcXQUIk+ePOgobbK7259vBVxoSaORPak1gXMj2AoqFcYzacBNK2mYoKaSJDfUsLW931DBSgcP2
2uRqYv4M/i8IhIgWjH8HnHV3d8SWAhWJG3Ak+rMsBIuBgU4jrKvmXPk5fKthhencrHyZpD4s363D
D/pht3qRBhxRxISFKuAv1eE/bsK2CmlkXOHqfppDdrQPPMJKR07bnRFaD0ZdqBiQvxr8UrEQ35Bs
WRX1KLRoAPsJUijHT73t0vTj50s8VuKb9hoFsJ41go2YD04Rqw2rr4dCpJsVSHQ1ibsUtAnWQxJt
tW19C2KuETr/sty7CbhFvx1xZyLnNavUKpvxs+fyxVU20nfxwdhjHuSgMeMYzi9CoqYbPUs0E4x3
HUTEUs1GbeRKkRWjXfFprsuvHDEV55c2jCrurF4MLGOHV5ikSJRA6ef04kihW3y9oGAAmE+2bXcN
MxXfyTitMKSfa8Pb4KEUyVNDnZGx/Q7wlP1CGny2tc3Xx53FTw9m118K09DqB6eu5sIgQNQzYMmD
2rUGGokywjJ/+IMlG6EFpwY2zL14V7943hrnLQQlSCPOGuaWoAYyR5RvXrd89AHNzG0OrGk2CvB4
9z9YxEPRzrAYZvqHcB0IxgNyzwEKL4kpn3JcWvSRyEys/jtB2xDsrfdMh6QaAUMWuxsmeE8Is5j3
eo2MVqxQOPcF9Nny3L0tx5UXlJbaQ//WffqqnoNBbwNZm/1A/0//ut8SFNaqHTOsith5PDAqlv/4
jtAe5hOYHaL3r2Bl3LGho6tNiJ2GgHyPfryzaLA3bO7iM3sZBUD4pm4v9NM+/V/rWRlmzUEma0om
UHpNEhuc6cx+8N/HifFpNJdELOnGHlRNlKn2kUEcuDctx7eYeJMGz36qIngFJCibkKBVMTtveoVH
YhVI+WivJAqPBJh/Wl34s4T6ozGePf8j/P+Uwi+EkHqbRd89zCQb3dod1qMvWYmUfs2QF8BCeNgd
144VoUmPLMlNJO6lb71dS1dja6XDpRjP0ktXTCoYVd0a4Y61jd0Ej1g8hMg5USje+F8YfH9J8vhM
TiedA6qttb79GQUPEI6Z6xkwuuGjRljWH85BPYCELC1/7J93t3zwQycXYPajVJWuaP3YfIgv8hEq
B0QkPeJ9c8Xj7SzObjuKM6wCuIuzsIiWz0OJxc6oKSvdUWeDJUydT+N095c4U/Kq2xWl1LsyMoFu
pzXPKCJx7FHZ20gqJZd5aRh9E5LHEFDTkxk0ACE84m9zRgRkBVpOm6ryCZr/09LkTECnE/Qa6krD
HrLGpZraNoIgcfuSa7055PzLFDHmZ4x8oUmtjAro5LqFAtcAfn9uGLJ9hQd7XnN/Q2kXd8rXlyya
WJnMRCgvzG/16VAR/U+WJfbL2HcM3uRzAkJJzi3shlCaHIWHBxGQo0NT9v+PCGWRT/Ns9q/KRhmS
mSD4g83QVvwo8xDkVUW6yRHIk6hFFYCAK27oI4bAT0XkO6yevC9PyB1EhGJCJ7R4krAEW/Gt2xhV
+k7/se2n3KlzuMPtnvxr86bhR5n/Vx6NeqFVG7+hxEH3JGbgxhID/+zlvlskSlUZYQ/h3ofmP4I1
i3pbMFFM+aMfNiBtA0rZZyPQqJxaJdARDJM1rnvku/aeO+s8y6v16k4pGqGcdrtyqqPymlT6Zug7
sekfhXJrTHH1v/P8+EEYo0q/naaA5PF/E08Rh8gZXR4QGziYO+t8inr/xMC6IEZD9g7cLe/OHGjw
yMyVF1DqsJXQzF/cf13NxXjiHBD2jfUqWxrEeNwTcX1WYc6nguBaql52p3P1CV9JN6I4L8NrcaO1
TfqW+AQ1/TMyCeOGQfvzPJRyE5zSn4hvg075KGC7OktPq51P2KK831nT4a6IpLZRBVSa+tJPXzmv
sMR0SUpdyhn41o2Bg/7XiMB8iXUk/egV3F82xciRnYiqAvB2pHZqUQlvZfpSJ8d68y1Hvh81/jMp
kP6Wq6ascExstN5jUFAxiK0i9gXFhZNEuM86FjYGwg7W1X3T70jDSRz3r3JQiG1fWLMz2FAJIOUa
pk4E5xIC/xLcyYk9JImOg7LSfZOhGlD3jiPYhqvkP0cCzEQ60KXKNp2k/7rcAr7JUtzcxL5yV7t6
KSCo0rtdlHfzdMIMxftDGFZVTsAwCDCJCniJDXhuJ/FlMX6XFsvpeUCe0yXsN71iYEvILePQVGGo
K7Rvw2BGFYQgHb3fRURXHWDLqeE325mJ+JTjStLEDD6Gw5vm/QeGBSXEfuzVEfOGOXuv562DC9Bu
XUrSx8hk71QPtcreWR7vJ5JxUoQpxKAAfHO3hnuq95PcGmJAF4jF5NEZ0QLMw+AeOjIkaAtFFopQ
Akllr8ZOy6AZM+5Rw7n+9EsnKScAQ5y50zOAJWmuFT10d75qfWA6TktO/bZAptY6NUe1zHB2/KYD
FzUcuzMsxTxEAxcNa5og3mi9V7WgWFnCJkxO2XNTh2di0Esy5NgGAc309OosIggdQd/FA6P5qqZo
yoc6G2KPrFEd1qKcnEBF2Bpo5LdBhPs2m5hZodTkapYPoFXaM/ngveYHtaeLOCnubcXDV9YkIuSN
X6rpQv47qUDXykcqZqew7lTiDnh0ank/oOSXevQVU7u2QKlTh6rRPUmN60HKrjFI1++16sKVIPrY
ee9vlk8Pm4EEUAgmQsGj1LAKsn7qf/sK40mO1AE7keg9bUmze5BbPA6Qz7NiqssOZRIWNzI0hNpy
1hSK5MKiLYo55VyjBjN7BqeM/CSg4iGObJHJE/jrS/qYwrAtpo1btm9X6CLsZkCYLNjPhLv0nmQA
HtpYTsnEiMW5vVBRUaBQ0vzApESrU1XYNOlKmRp9/9qcPXnjr+nPWEeUNhdD4IVe/l/miVH5qa9Q
II24Rr9ollobFTWLjECIgG3iCVvlpshiq1teUHsVwSkLCU6m0HxyNj5mBxdHViZWsN6nJr5TgHY0
HdPN3u/235xeVmz5IBU7uKm0PQP3VfkK5NfOTaj7BIVnq+Tux2B5gWdrfvoFZNttOGGU2IGqYJuD
hMbAP9zUZiHrFoAtm+C5fbWWeND+/xbsEg9KW2QzTYmiuz5JjjTaZrEzYxvLAZvBuFPmzVPmndVv
5Niv5WPsY6Bkw37XrVb1/LLjVU/zA/DnjloXouSp59E/zo19IDY3ZkncaXoUG1jQBEZ1EA/ldOMl
3njz0knySmC3WawL6YEtV7igXY3MgqVsxdo2hl4N2sppYq+TvE9EnLg1Yg5BjFYNZlVlM7lSWZzo
WmodFjLU84uTPPDyTd95KzUJAm4MgpWb/kXON6yOpAZh/3lx4aLQEH0KsCxOZAn6ZzcCgp+bdn3J
ztQyzlLITxOjNCO84t7Av0e4JRoxvFLu2hnxnbGzevwPtd0EelQ3u2OXhPHt90318iiazU+WjXWN
Gz/W0/fV1OuPv6gurN6KsNMXc6xw5UYEwi+hWedfsQYCZOUVm64PbbDjqRm7j0LoVGYCjxFbkI5+
df24vROhzAaryvZsoLzpY/FwBJwhCH4mks4FI6fLEeVUzmoEbtgvaKxiESUeNJ2azhtOAapwF4D9
UxLVvHLM3RaBb1iI+LweyURNYDQxXwY9imhRidEXDa3xWCHgsDrc8Fphc0PQ66J0yrAg7f3/T81w
KlZSgCZuE7CMtaFMtlTA5wQB5l22fvoEUtuwqk5TE9o2tDP0lZUFqA4ZagapL5xMpOfI1G6afvn2
h5n6eJgaBOoD9AYYNeCg+7bliRa2xXEGrkiByRjlF7si6MmH2KpEIEPUz62HQHyiBlZgNAI0lfi6
rLrTV1daZFrlpHDaKVzV4YO4c4bKQKjMhrYIY8Pyd+51PJ/814WmgQNDIoC+q/sqkXLUe9+cAPTC
QfRZ7g85m3siIG21Hs+T4FHUzTz3dhHzJdpKUDxiCYJziEfmGYfrLxfd3rp0NIP6J7hqno7bXwZn
Sh4VRFQoiyS2yonP4xu38q5GAJAXSyT4ihAwjLDIXiW9fc6sw1xZ9CAG2ezGMcgyY4M3+w6Rbb6Z
BjdR5W2wp26FvqoGsQkvE5R1lCK9kXgZEQhf5pi//KkbYPQqreZWJE+8/apvxuQnxLelDYvYpHRr
3+9gR23XQSqK2Og6eGsGqy7b7+eEuPHWorXoaE2A1vGC2ebbNOYjkb5WsdL0fZs7/tGSMpOBZbIQ
ehV/ERY7bvJG90z4G/4G60xWI66bxi7PE0mx80urmgWVfu5c/DAFEnzU+w0DTRGyQKG1wzF86fNi
d3tcDfSXgZaUQlDShSbn7wZQYj7cfETKsD192eYBkIvL+aUE6wakSRh79Dr66WugiWS+lU9MDOcf
NoZNL8zqVI9fIU0e0BQyniWKXCFMpae73LsdTFCg0D70yxgUpZPcK1GnSDyC/zInoyNmCLgi/2PN
PoQC/ATwLNSLEfTD9MpAB8ctia+vUZZ2HQq8XzteW9byfWp814LRePR4HplE9iyDqeB0Ul1uVmEJ
4XOG5HGpvSD2lpx3a2blGxnIcQmdkXVRthLj1/ZUZP4FbNuruG0HMV4FkxGpQ39Bhlm1Ewq4IQSU
1wTmaB9VzUSvynYy5uU+eAQ3KFVMG2LuEes1MceaT9SckGqk8i/ja0/cQ1QXYVMNO+bEAUq3RkLd
zGcs4jASm4Q+DxzcBu4tV4WYvlFOl+sqBpYiYLkntYgltFXhEzhiAGh+EuBemM3NKRey9jD/H6Sa
7R6bisyjJEIyX3LMO1YmpFe8fmijx7MjmcvwVeI5Q7vjeL/4mJ91Ivj55KNQYW92APhPI/Sbs4PX
Mn048YGfQ6rf1KMq7wWeL61/N+WyfOBctqY7C8QkbdQcOkmNEQG33YOBKEvi6E19MEB6auL2v7rU
jMhN4h86g/srV+qqelyM21mfg/j83HIjWqc4JX61xavuWIlL+clUu4aR5/cyTQcerE0RFhPfMc/G
t1tN8qU68BCnMYxKYF8QPri5HXUcjxT7ah+3yMZ6IlPIFEMfvB7Hvi1NciiFHu1dvrU8bp6srh+r
nFjsa9cHa+e/vfTUPUQWMg9tO6tQl4c0zX23yZTkZIpGhypuEAMzxuy/aYK0ztusgiaLwC7IGI32
h5/Jvf4eTtNO8QKmxXQhzWxx0gakQCMCtbn/IHStlo2kUqw574vDEx00/QvumIgvmTpNkxOsu3cl
Y1lR9xm94UWLBVHQeCBGGA7akLr9ycv9oGc/6ErJqWJ0JoUoUQh9sgzDyKn0OsGtmzuauSsLr00F
Kctxh0ZG3lGJQnz80fo+kAplL7fkBbpqvzDnjyqphARVZju3wS2OQR6Fj17liaBmCsgBi0ZWAGiO
O2Cn2U9VSIlTGwMEh2d8TRNdrvC16lREIN60tAQEJzqIwORmSEQjevpYagaklP6vHkTFsBrDdYiW
bM0YZC2qb7J9dPuLVEfBT0V4Lnuywh5qKfm98t18mkxs/w562JcoZOmkZ3VYrif39p7uix1lvAN7
jaexhVNaD+9qwkdlIcm5D2QXdvaufFnQK1s0XTPWhIM6e9d5TxPypDxeiZ8WqWD15cBpboys+UE7
uXU0M0v9pG5JZ4OmmeAqtPIPxU1+kgyTw9LdFv14A2eOgALpM6xeTQ3dZDdPXVPcIGo2MQNEaZ+T
sacsIR7ghha4eWHPGIOBOU2iyh9jgcpx5+frCSPgR1x8Ssg9PtmHnOGWgaE0nCETJ/kA/lhA4GLq
JUUBw4QwduPBzGOsndLVRYTBowtLduRqTStvD3VbecL/Ch8ExNEUQ3pmhlE+rdh/2nPoSNplI7dp
VTJBttdozalFZttj73q1aPRBsn67NevqKExGe6BkiYa8kvIA4QlmBIrERulNh3qfHO+t9eK1ZFo2
Az5cvW0sbV19sTtdX+3LqSg4XmXW8k+k0srvoBLVwM7s/BgOl7Yk9JwmZXUXqQBxTdqL1EeBtMqa
lLaFoZ3hZCsMwUdgjg6SMErdSpR3fh9jVwPVmGpL+p0GWrj7ilHuDKA23iAPorzsCQ2bbYt0gWcV
GoEr9WzfrbzfDf0YhZs/Kxrqjt8C9HMGcWRtTT9lLPDNiwWP8nbptq2j7Z3sAFwa+9xAC4zo7X5X
1i/islMX2o0JtQAwFdUzYThB3f2YxGl8xTxPuzslXc6N9JWPMuNfm/fmJhk6gIttCyP1v2+Ocq15
WNVg6Y0heylhY5qEdKczG/7V7ueHs0EdSgZBsTVsmRvHfu27mXRB/Cw403xgEodFHrsZFBymkyNH
ke2dhGUXRQIiTfq0g7jhbHaCfCoPmGW8KL+MnwzU+efrufpN1tXCdWlFqOqA6BTdYDNIMm5aV8U8
Pe1gWFzV0v/xbWHzs4Q5XZjFbt16q83i8EoeythS3GQuqb2jpHFAIekIv14Ps0QWrgeCefxAboN8
6txIIgyXGKNIgQBn6w8sIabhEJy5fyDo7tD9Aop7I+mAHf+7r8bX868V0BML079OBfnLvBKvnOqG
CdrdVw54T57xdLA/676Aq4qMwLiwLBxbOtwZqADMqDPbb6DirKmVo0+LgoIpuL2856rbQZ9BcN9m
+UyEaKSICfGNB2RDS4nVTnVBm29pWSEF3ufQZss5GLVRnQo8+zNyZtXKeD0QhQjtGHfbXXxcx/Ax
o/fF9Oa97ZiUy2SapvJH86sppNcQxQPQAO7TPcY4OKRBdCnW45vAACwPfDYrLyPcP1/Lnv3ke0gd
FDnHV0O8t5Lrn0Ndl4OR1Fac3jprD+7F70zGrkAgXZ3jwlCbtmcJ1XY92Ig9WJ1l9gT0OFemBCuI
L2ZfPPomqFx3i1XKP1IJ6JWqV2O9GsDCLNFFOeXSYYVJjlKAVQmGLbEu97bnmOELzDctxjLC9wHX
fzZuB+vey271UOwF00Rh/KpeGakPzXn1WUWHf1DGuz6yYhHVvFnLANxUGS8ONXrk9QqEPHKKhOhV
RJRl8oCenCucVfjGXtjP7WiXu6ys7Px2bmtSwAkdyAPwb1UQaWvk7HsonoM6DDSqFUV3FhFOIhDw
Sy1mL938uOkSXEs1EO4KtmaNRvFpSAtd0P1BECDVkoWt1fesmsLMmYcrnfbsc1DgvlGAlh0tqlCr
kD/v4CTBiSauV8vbsmJaE+72biig1FG0vDjRx8lhwNrrdfQSHK63UyTTi0xQq+2Ax67PZEToAlMa
ve746zI33IRJpeUfNv1sMsFaCL5VD2a9/C5YOwWU8XTwCY0GAwtlAA6Jz//zGFen/bYvgwQEzcPl
jfOceagDKBqMXCIwePK0co4jb+7uY0wIKBqGlBOZKAaZBkt8mapfHrDzYEM5mnx2TM7yPYKxiBUE
azdCarDsAtBgmD3q916pMf/oqvArO6hB1RDINrTfkrEj09FQCo28fHVQkGwHoH6s8fCEEmP0hFlU
AtNPa1LfUUZ4k9RMJnLwj3u+fphWMX5U6AGdYxTJmOVjiqLdUR5ULtiAGSeN5hJ4NQG5HZUyCYHB
iWJea/s38hryRBN2K82ezup+Ann4VoTjCjSpT9bK8NVS12Dzqbx+Qd7CyumQjnPj3hODgNkbiv4U
vfBo5/JUAxgdf56EPASEda1dUp9Y7BPGbNTa975DN7PBWpwyjt+PzJxT+JJqZUyO6O20yw7Q7M+r
37BeRmhs2s7m3xb1X+rRM394CgTnHmL36x3dnhNIqSHpu6uO8glbi4mgVwPOR0j/yDR2kaeorliR
7HEKgD2wBgU3bhZw6mswKjb+Q0SyWgJ4lgqUO594Jp0QOVgGNbFy8K4/NCJyqTaopz0ijZ4AFJuu
j1cRpwKa7qOViUtGZtZzJrxahhxy51V58W3KIYh5bXl8N2e7vbBJBv9PUilNhwBGI6o6iMaTTBbd
pRvAWyh6Q7BYgGLfwPPI5NWfbYStYOjTOpG438L3z2TaFcWAxzoDoATFFPiCxahK8wVRbsto71Ud
ec48cC1XiUc7Aj7dwnCmMBNTalfkcqzRc0cjaVBzNEhvVvpl0raI7qvy3TN3qHldU0ox3FNZn4iX
G64h7y2yoaXkHUE3+6p6d0ecXgwjFgh1zss0oO64yfak3uzlJC1N7KfT70TyGsCBoneAXalpdcDt
3RaQcZB86B4dxSkBhyo4yZSDg1cjfzmukV/GHTqDmH4+8DVVgNcGfYNzt2TAd9m9YaflO6JkTMNO
wGV4lNY4oz/SRUmCvvj0UsHBxvrZ3uem/mhLWShkl8Q20/8URtmlhwqlj977D1rprpvc5P5LrU8G
j5b1g/q+Gew8cV4GfFn8nLU71qr05dLxbnGh/DzbwmbxwOiqcToC/Xb2beY2D88qY6AMktSE81s7
2oOBFikIq0BIQO9ucja8y8mzbTHhEA8ayn60Z65Uz8B13vieSMFSsrJHYWPN0PEB04if73dsOHeN
GnkAuHXrwqSfV37EhNHhedxP2Sus/rOXqorYEKbx3mcK8q1QIj0iFzMCXwE8VJjVsCW0a5Qz4zYL
qiogne1wrG+2adKSU2eWIAni3uvf9lW7tcXM+0oWIby96YfUbH5DlH8EZuvn//SCrpXPA239Es6l
e6ME4Kin9LU4LUIAsBmrQLSUIWgpSxjYHxC7YpVf0SUfPWiwpTAgffctQongplWWnG68FZpZoKsW
osXb6D3KxLZoKEPkOqfsiSSMO/ty8WQFN2/AEJqvceD1qcNRym1M5w8LQ9FdYTZ9vDE02Ts6o+gE
CDK7HLbhIVIHL6iDA41g6WYnR+9SgZ7+7XqMMNCU7AbnpiKNjo68LWTgO4luQI4D937NuhOyPvVv
25BQr0//ktp3dqVWBfhjuM63QUJXi2U4ahFmDPef6lO2Phs4FL+8iKdz/y3zdR1fw6YWzE7gODdq
ystmKulEmeW21jlfaK1ApfUD9GbdwN1grZALzom0aHTklYcY5dFODHGoJ04wcShsE18yMqoQuObL
8MIa8JF/0eo6GPCmLm/lJ4V8xVnxgTH+nlq4L4ZejXPAz0Rw/gclq4FYRXpBWGDhD3a3MZczYFLp
hI7BwbqX14oQmt9+HdyNJeZc8rR7PmL529/OgTyn8lIqG1lxDV58frPU6jkp0xOONiT39ySqF2Sr
KawqNQT3aHCQiVRRzeDAFMWsKQgIGJaJLV4z8BVTttgVJC2CShrQWmAGXeBh9AbiOJGIn/p3bTf0
QYwIWUkt9wpvbV0ifYMruC8XCCLyup+WZ40L8hODXIv/x9SFfhEiIPZkUEZDFcoty1GxWI+soeSm
RZZ7jQLDDpNtbHcP2KMWyqkszXt4aBCrlj6BfiZSmYbPoRUiN0O+2bhC7PNLPiddQkun5lQ7udhI
PiD8qHyj0xpu6qvXmdFMa3L/44bBLH70vVm4v99uX/Ge/SlZnE/JSpFzWNgo6nPdw4t7YIhJXZGb
+flWyUj3Kh9k0x+SDtSrkeXcAapkjL8rJ6XlukmjJCOCO75RmvGjG94KTIP9iVqk6/QNtAAKUQP5
nAD8MuN7S8XdXuDuQRUWBHh6ScoCw3RgcvZQ4bKQqj2yGKTJVOp0ZgV7W3l7uyUpHjSXhcmkEuLL
u7Xf+iNV3yIGTNahyf71eLMqZ4XZM/ncg+7MRfNW1NRJgB7aj61+qjF4tgLN+gIpIHU/LG7v+JTL
l7NsIav1olZWOOZEjAeVkPXvFupgm+sFdMejPok3HibE7U5maP0KewUN8JfDguJYwsaJ+SS7Xagx
7mwd2oQ9Iy7SzrCm7GTl/XfMXq1WkrE3kletbCnvRONCC6JlMt5LyqA8oZEiPe1SHVxjM43nX3MO
VLlZ8pWJBVchq3k/s4wuNFhbfQePUCCLj/liNreACJYBpy3oUy808qjxFy7/XOULd+JBXRVgjW9H
2Gcw0Wx1hYGblxPeo+jneuhRtCgciMogIC72n+LthD4mDKAWLI3aZsFM3WepbkMDtB6usWm5QBOO
mm0X9EEYMuaa/gMb0QmA777PgOBMbxyUz+v41KgE70m64hNNj9p8T7Cxhg0ggfthUrmtrnhmXbRb
09qHs67bTrdQij5HzA1Fv1gHxtyMd09FlcHG90KdEp6oOQgHWeVjrBvfu2X/VIERdkyueicQxrZl
jld2Hvt6XVsmhyhRMfwbCQfG84fsTAZZh3XE6/WQjib65oYzKtwm2kOkmfe7ptmNacs+vgKLDX76
P1D0ZAs1uvwhZLS7uhVmrp12yGODrdp/XdWP0SnR//qsx7pxblFZgZ/r4lfyknVuAAqA1USqo93S
roIFz8bpIY2iV5DjY+u7D5a9iiJPvqJd387oWI/8t1YtYzoD6zyn49toDyElDVcjfqySqzOzWyXg
P0tDcHYkjanuz11i41LrRHkj7/ocYNweJQB01FDS2HHplNwFxU5Xe9LqQNDEwunfhLeAhlu1UE8g
BHtQLDF238nQ8SBa5NZ3eE5HCZ3GrqAEx8vdVoPWsYWXRovZ/dOlRRBnPVP/Vs6LkkQVdq6df4pK
70ow/SUxa1nwlrjr6A/sLEG5l7Uajx/6cOeBpxA+EmMhcpUJo5Ik6QuK3Un4cNTli+Ur8zlzGTR/
Wd4XL4PXXpmVd0qS2MpPxV5Fx3BL0mBixFFhd3K36Q3+d81Jc/gHlnUwHzKgurCLoylhddCrAysX
ww7spf9NKKAI474lxggQcLfj4yORjTJhi8gQjqVi8MgYyPTQhWJ6m+I76+ltCkftQAGDnJSnid0F
R/wcRfPL25nmZCDc8Buqc57r4XBsWetGXROPnkCf7W0FDAtl5Y9G5DBVRj17+7gd6kkhmNzfhNFd
wTPleSvfAas+INCNUuSpLPbJ17JQAaVntAoDrHpYuepSRqqxK2wJE8xYy0eCUMLQdB1TossffmYy
k6um0a57xl9gBrjxwDjfkmo1AE4uqUJ2U85gE4eI+fOA9dT9XrVN7ShZv3Do57iYlpZ2qts7xYg1
wVUH8r7Hi39CkIH+3aylteQiJDzpGY9GZWBgLuch2owFWjUO/duj2zX0dap/s8iVCe28/8hUM8la
t1oD6Iu6cTR5lFMU1fBr9BXLxr8XyGpDOCqdjuCSGuDzLX+Ybs/0ph52EW5QCqwFDGwU+0gcj8jH
eF44NYFuN9rGXVTw2qPfaJtnT5EQukoQLqKRR+OKdcwHj5/mkvEexs8SvWDmQLH/pc6lsyL1QvKp
zSCNYw8CpSh0kXXKdEqSw+b0Wugu1dUncJxCPrQcVZdXyz28lbMvGKb8C+M8dYYv67oQ32ekmEBD
L9wGtKdyn7R3b2YtOf1Ll62jLVRBCpm7ifmzXSwORuslJiYUulvF1k10Zk+0WohwvvZolZXuyYwx
Z6J3W5CGjofaVOVhTQbvhQfE60veBPpTWJ5aE1V7VaImye5xbWj7+/iq8arkENrK94API5he6cLN
dLRMRtDZQgm7Ah3SpMViWuVMRRsVXzzNU1DaWy5HAXH0HaShc9UZ6OFRAiHYcPifZWecl+fGduZz
JpLF2bfSDKA8zTVwaq4gQStDDonpWuAy5MDY6pJhlpM22AdZHoCDB8PsBOFpd30avGeZmozaU2jr
WWskrP7Z50i2s/cSanJiNVar5iWSo7WvkCBAWs+YQX1yyxzdcpyywpq2i52EKOckAqiVygPfNRM7
wrMGGERy2NCOjxC3ht69U/1Y8cfilLKfAFYmD9xC0+EcICX1ADwxhVaZdfqg+Q7mGiDwavOHdMY0
QxClZpRDIlT7wO8Jco1lRyeAg+wU+1rj+u0OAYe6D0m+WPSd4WaKS0hc+WwZvDf34777hGh0tpyR
WHfvZsMHBpSVtDhcNz3y+z8z3B1okMwUWhpEQIWrPvSLAwYarygEMra7wNGBmsiKSBgfu5lFVDK/
UeABc7blxPzbUmhWHSlP6LIqwmTUmrkIy31nXgHPKTglZR+4u5UTyJjwGFkZzu0Ja/sSK5I/fw4v
vlsmkeDvWVRWGdPsJvnTAB8GniUswEWyvUAG+CdOpxt+yWd14eveUkujthHVEM2yFwv8nLRKYl6x
CYz/d3N/oNrMI69HyFhUO4KR4D00hCHxyFoajoNJFFpLAV0IChDNWGWK5m5UDryrWkooTzyC5/fY
Asb5daxkAN75LGa0imL5hV27BP58lIYVdCURgtoxjp+kjVRdOwtC514s/x/cSnF0Yr8tefiQ0ys9
DrqvjAwxjP1gUraSmCqthZwrXsC3RlN967ldLuZNVmuBkEt6g/N/1YRSYwDW06P6B559Z27E408t
OVJzp7XvjjvnwHiU/9I9GqDiiipqqZiCM3b3JN/U2k65A2vdSyuzjWBA0ns3ipwV8uywr2fVbQLt
sQKUR4Rg6HNeAh9DgixQJvusUlE0aZa4TTVBLn2fJTZZv//mpf938Gj6lgBeDitqA1OeCA7vt8Rt
45fOMkn8wRD12VwbCV5j/9aGYJWPA8abp8UN/1ja7XEhvjug6yuqI6O4sSeefuT3uyd1PGwKWQu4
P90N2ZlmuJ9+VqDPJqKKA5sN9fSXmIL8DOa7zMHqBeWK+TYe1T6agRwPb56uXIJCzWXgMmLUUn9K
X/LP2fo56YoaMNyWcfVk2TMcYccMm1xHKPvRIEvtqhJquyZq98fOx6b9pedjWrnmW7YJWprO5fwD
SUVkFO6SEZibzXaUY6eXw7XngRY6wYwRGwR4Hi7AGXY4aDG3pTqbl0JJm+BNoQm+EIAJMxSmcXGU
z1d9ZK7tYvE4kxAVOLzut0G4xhwWyHeWQZ1S9up5anM30PbDHV4AASdcY6wfiHh9NHjpPdtLfKLw
sOk14LeY5MihO/fC+cS4/5nwnfjElYj9Ner1HOSRsceYvzc/6qYCsRFyTm7ISAY0wx9cQyIW2cE/
hl5jAnxogEY9Sc3GKYoHdgeAQ/BIlnkhHTQmQe9O2cAwlDpfpnCW7kfWZU8Fku5XUPcwG3ntNa/H
aCFWtHHETNtlWq1WS/62/BxLy6AAbZDfmqlm4Ud/8Nc7rEaj9y4McOWr9RdSX7Gnfl2K/bX8N1jy
swfg0dsgyQpv9dAo9RrFAbzw4ZLrvo8vh59somBGXTdBXjBgKgnBBiVTxKYyVHMxxhHSa2BaW+EZ
UHYE/T+6GINkO4+ODtFIJroDB7+cM7xppRIonPlciAR7CIyTOW6MhZoDeXP49uagpZEYVamK0F3A
4VgfRpdP3k0KSrz9Qg9gB2aBMDEpUU9aUGO629N+PdO09YBITJEd/+PrYiTHngcS1soiafZhcoXN
kyd1wPGpP09Au6Xjsyo56nebyilSLgzvU/BadwInryung7HLVcJDzARE1g947tGoJubGUDAC6Oxn
Rj4hCFxVUlPIYRWI24CeXUGSSuo1l5pmtCUVXm5BRMWQzvaDIdWsXeavK+3nQVxZtxGYeGd8zPpB
03LuMHbgVTpoMZeDIxY4/j6mMy72bvZzyGrOfZxbyyFsZ/aVf68rAoSBcDX7sObKPjSYux/tLqGo
fQjoMjtSgrv78er1uKDyXMX1qQdYuENwfeWTCHE2WuDdETEeVwUUwu2De8cwA1vES1XM8Py47Fkq
OmumAfe7gi9lk6yoK6P8LdXEj287Dsiz1v0VRwd5i4MQ59fJi6BKfw/hCS3FPcavfT9LZuzBJBzp
OKfDOnAAxInyLTrPBv7POlGiZQN/3J4UJLUGOOVIrBMhs5fZM1+T2BLmj1nQsnmM9zpy19DebN3c
lq1CpXWtfepSrCoRc73gBmVIuOjjeY1sAhfBu6nQb0aNlPwMsPOX0kpZDBwGsAZ3UXxDQY633tni
ir2puK89lXMCk+B0Zu0Wbu1oSa9pfaCV7UEsbLYOlArG4wVO2R1K6BlYrGbxl/5QWXqsT8lDzJRW
C1HGAID1Qs6l0qjFoljRe+XBsPOGFsnxH/2theeCYZRY3T82vDo4Xh70RfkDDbvMBmQasQtXxkR6
7MVj7mN+Ez4+HQqX/loKIXtK4apaGeG479ToXU2nL9wKILE6/wkLnOPIaWdSW7qUd7ZEsEtCZHxk
htKvOCcyprS+eqiujPDZeUv+pdYD8I2HZ7SuoYZEcZ/J0K4KAOTFTbk/J3C+IhC5jRBggtjBx+Kk
I+jdtypKw3kgVSb7p4qyJ3MAns6w0QbykKpWkTZ7P1j2pxh8mogmvqTCDyWyMp4puIEAGqxM9Nur
WSrRbyiitLy6I9L4IaZ28aKhKuTHifrKD3YHNx1ZqVBimf2qkYk5pkRj1Wl2TH0jpcMJkmwFWaVI
qQEONFxVcr8A5vk+mELIRszacyiOUtRXgiezWZ7w+wLZ4rH6+zJm1QYKKlRdRRS8Q+mafAiPbdUQ
2M/NKE7+1ugpwBkdnRK9kSMy9Bwf6eJnI3koWLfnf7F/1ByvU2iPEJpNKgHzM4Len218Jclfxos4
6vYTBKtJ9mktmFx42NTj36P/EAH0LupdhG+3c3iQpvC9LI6OM20aJ38LVTqBwDjs62rOuLQ1EIEt
MAN5kEMjvqoE7bsmWRtA3mYw8oY7riZyyfhhq9NKzpWwTAYBaxjMUbfrMDQq4Wf575HTcZg8/Vj6
mJirR/qgW7MZa4yGwXfuKtSdl6H70ETSpF+dbIuGUedx8si1vpZbQhT/m10AMio0QkbTLvvDMkgq
RM/VRQjFqtGeZKqO4hr2aWQNzAtc+ScCom12e0ukxGI24F0CXfOmZYYXxf6CEWwevRG8tvmZrpTM
eDBFaSuyIDq4slupuyCxmB+tbU7MJR7Donlghj9u4Z2dlmHqdm6nHYUBE2ZnSqw/Z7Gv6N5oJiPz
N6FAZRHcLwEwaowxkjiY8sYxImVMSZzCG0e3jt7xSHrgbjrNjZx5EfVT18E3FCnU3ZonILuumJmt
AIfgAZzxSvvgJUiX2fvlumA9LLzyUP0f5prMSlLIgjUer5COTsRCoxyW8rxbWV/T3lk6d9P7+USt
lBQlbq/6I81Et5qnnQUdIHi65dWqAF6a1Q7zz+wj0WLEjimlmtLI949BcaBMpKLL99nhBzbSzsQ7
Y3Vo4qPxyEnVa8WczhhEmZGZAbVaYp/HLi1sEEtds/D7OOAVFDndNkuHIHP6YYcbPZJ+r7pNF9Y9
jwa42uwxyCUd2uJGUKi0ybJwMT/mvhNAk0xcVA/bmx2JP9Obb379Yx8E8PVyOTp4m7zMYUHQNx8f
QBbHE0f33ExoU6adaNJZSDH4h3YaiNnzW8EMo8bvPQ4WejqY2UtyfLz5+3H5R8wlwm2theMLScCO
JXsS4nmnhu4ZNNfYWVhfwdcpS8vHGtU+u3r02iXmhHCtQTg37tAVygwtzhNQ62wHIuW4t9iRLVOG
hdEUYI/HXSWAG9NR0PN/CMeQqRXh9pd80rUrWniYIvRbO5jLlvhmA8NyJPjU4nzaI8CjXrq2X0n2
IoGPIPxQp9td9vmAX+J0SKM2/8fhudMkeRoD4cJZp2JnjpScsK9DItqIlwBZeBxP59aLMRIU+jDG
PmWl8Xr1mNuazgmbhOQQHKO+S2q5s7AutoPYhRkyDEbfyfdasWWH9H70foKY5tdG72bHTZqoJk/J
x0FPjP8flCBRRPWuYM9SKHqQDtyUq9LF+qSQZXeYMAhG1O4DyTz2idsSyH1raTqSbHQgjlrzuUjq
lRwNJs/UsGYiBr0lVwxQffeTDca5Nrla7lT832lGWoeNDs6gddIIe4l9DU3w6Ii+GHePOtEPFQN6
Xt5GpyzXhRyiYUul8c7mX24F7Ob+lDvh0EiGYdeymqewu6UxU1Iy7GRSrPuamB1ktX0tZULwzUYN
YI9EdPKu7du/qKPTAFzBXzghbobzhwoxFJ+IAXzYzJlyw1Xo+pzdZ8GvMrowbqLWLpKtn9JhCP1W
KHo2onNSTub5Ohwkgll8C4gk9dcy+c/E2UfFB25ApKZMQfBmATcgdr6N2vvxAmjT8dZBPJvoiC+J
PTL4+IxASnQh9jxWWz/IkJ32XSuW9mSWTMcfGggouGniJ5uHXZFqNiLXIPA9hRF/Pn90j+HyyOIJ
Ip9m0EzhuvfCiX/uvqyjYksvRt10zUoiCiAw0hnbjrN5PDnsL96eNM6Y6tQ+IXX++eSBxMdWbo1I
fnJonZKDy6DiFtvq2SvttmI/Uk1gZ+0Flp3B1JIO0+UKyVk0zcmOkmTKx5WTWuN4pjw92LX2vJyr
i1kJsWC3LtUQ4xn27qxONV21OI9r4BdONVKL9TfLjTfKYeVmEZC40yGjguITm9Sez7OSMelH43V4
woZY0O5xY21mYxyEZT1BUDan2IArpdRDV2m1p3CWcSh2u+vZf7V58nSsij+27dbsjsyL7ov0MQQf
E+o6j5xAb666/KBTtDesRgfNedbsU6U3sKUl8PEHQ88KHNBplw0qHoH67bfqV5Je3m0b3wc+fNhS
pA/21M57c8eK12jWcT2wU5Mk2+DTXhNtH48lNxnvYSZTrJAaoWtVq4nbIuPslXHnpr7vI0gvkZJP
z9lAFTH7UT/Ep091H2KChI/hIDlVAVm0RpbbbEdhm3cgZ9aDgfym2XRov+tMOBFJ2Km4QnbK0gwB
EhrMZv30cYfT5gS40wK9s4ubyu2auEUhMXZofQzTaF2jYiQYLNkazzPlJGZno+tHiBTvH7bWXjhN
vsDuVkXSzMFMDAPhCagx/n0uHljJR0uczmbfAnrZioX8m6Pcm3KNv1rASze03oxJ24Aanz15zAbn
aw5oFHqoJ/3VWBfSs5ZoTr7sIMNPbuYAYuIuqXS6jcJZ3/lsJ4Dly/UNl1t+BjEDuV4m51bi4K8T
faCG6OtIoatKEV/3Sh91UWpN4GlAI0VLLKBfgx+VpxZ0yoMBKvnyJZ3+pk4Din0g9axQEGTMV2hD
6xif8VC/uHZc/LwuDHe/U0dCaHOgEW0XTfNUU9FqqhKbVOvl8q66IZqEErIezqNOpFTLf9dJtSG3
QToi/WeUjmRwFang1e+FicvKD7OZGgjkeOEAIRL6dMr4adV/BGehNKd/7A7uUY2B/zYjP7yu3bGx
p2S4wmHHksdkRdLyqNV/AHIIyoy/fs5QTY3IfdnMMjZabTmoILCb3UW7mKiuihpQsucPAmJ27jqC
thDxddHkKSZSh1Nyy1dM4xGY5b/J760CjZQiDSQ9Yvi7y5Hv4RTNmovL7S3rtIP2hkOG3PmJzlPk
s6IuZefQmFQa7QAfWUFI9JGCtOd/Go5bN7QoTIGe4VajtiQAd4k6N9ynOjDqIfPy4Mq0q3sKCj/1
bDRnIpDfvdaoYjtqDreJB2Yr/cXG9ebK42a5GgCslDSFE9GwixZ+W5jNGyH8fE/5uVO0EuckQ793
yQP2zxfunHD1qkRA40f2Vo/CO+VVMYmzxbeZsN0ApLxbCNGg3gmo5XhWUH8vz/EQN96yu6DBYUuZ
XfNgbQhS6hg/5kT23ldygsAQ41VBr3iKDxBqATHsmM0oIQgLvGt/ON48gpwIZWOoTGDSyW2UF9KH
Hv2/3t3vV0M9XTncyWbZELDQ5eXd2aKlC59vjCdkJ+uggzgf775IYDCIKWQXz7xqxRRVgkIWFyga
OKoxPfCAosnQSJxELvWytsh+MEXXTuRS4CdRdBDndLwpA80pveI8r98YIptcaCa+4Clc151+Bz0B
eDmd3kNBFEf3l8DmbOwJXvN0KEp+/32NEUXCN6rZLgypbXygG7vrOUA5nvMKwAPG/+Ni77FqQKlf
mpIP0kaWqhLJeyTHLb0l67ooVbkd+FVOyPPiRIu9EbyWk1Wr4acJ0G8+14xG1FFHeo3tCxVKpc+S
c7kiWP64Gj4vdkhO9opxfo95XsPk0aoWLIkg/YNKczhPMNuOnciXjAbD14TP+n9lfgTZ77WHxSZK
+D/+ohEcjtySIdTizxfqlAkmhh44jg23b2dysj8te7v7LLKv0fdwQOtcAypsF36JM+j8aP87J+eH
fAeU6o5+UBDtqCL0BQpgYEKAHgW27ORjSa2jMC25S4LVe4cM7D1hIIsU3Tqcayh0N4np3kgOmZ95
EImJZea09N/ofq8AjfLqNN7wSt77AkgYTYfmQ7fLwQKvy5BS41ycMRK+GFs1zv/gm48cqwHedWO0
xihxkQJphMOIcOi9JlMEw1GZhz06seJgeuZJxZJ9a3p4vCdZVyLOSlD3En1MLDnJGx6xWLYFqhDM
bhzZUH2seC7VXhV4S9XjzwDu8BxKeH9Y+ot41xdXunl2CN6yQur0uHZMGmf5G1pv7V2CrE81aFaq
wbl2rE0ZFPCaVtTo6xrsY/N4TKdYYxvrsIVdb2W7ps3o1FOczPdLY+e0slyEXmSRXr8vx7H0jnLR
Qn5sl6SI/+hr+mBV9O8rQUUqUeYXtTwrj+Ba4n89A31P9Y/GIpq19uzdWSCYhq4x1DxfxnhStc8z
EdouaxpQ1JvpSCSnfka8u5LiLADiNUCzA5R70/7rnPTmYyr/dB8ugjA8gqaTD8CvHbNG2SPlwkui
cddWlk8iWb0f8GGi2OAcppzvnjfuB55LV7wQG1vvt6RQX5SB9MbtJsi+ssoNzqwJp2oUfaGSusU5
95urAFFttJchh3pty861zlQ0fF1NQTVXIpqeHQG7eujvhAEdh6v4GyZZms9dtZKw8YLpEb1PQoFt
CFuvehluPtevmLY7sLWPDctktg28/cea7PSU+4xgW9cywJLy6YMf8RJS8Px8x3oOQGQ7ggHze3bE
O2qni/6X2p/gNJsaQvbhyDS1cB/q2LxAW9ABtH8VcU3wmQGO26HRAL29Y8FaUKaIz2lRBpR+/8jI
SybqXrk4aCl/9jPS6anov0tKr3s7mDdITNdIKehwfyVBPAvnG04hu0fouzxlXJ+37YHpglLQC4MS
uzX8HHLRZz/H9SNtk/MTJwtitWZYcW7fXoGf/ggBTmVYBBqlS/fJfZQ64dTLndmov3/nsuUlmBss
B8wKnCWX17DoW5vVbZ/GELeA8BuxrRC98e9cHO1NRyfTR+ONOEGY6frcoiZdAhhpuA4jqCnxbbCW
0YOd6JnhHcxMEjH9eCQ7gKmabT50mGNXjebaIWmuPPsGptZLjfK3gZ4m4ncDFKrOKoGcuITOgcim
Mr2hg9Y2ojgJunqTNQKnP72Utxe8cCMV2zfxEamsfQ4H32eIcy7p80LlQIEFyexOdbA/KPS+dp0E
qTXpIqAmBJTrWeacV/jzQUrzTf7DBcMPOUcOGSXueq3p5vNUmSaY/JcovZC883AwBJ8zDbYUN23y
wsaKSUKiNIM7bwGLUalFBqe01xTB+udCvgwwsVNC6a6+gNEUlUFYWBIeUiaZpx+m2tQVgCBpLKPc
lEFImKjSayewPP44RHoIadW5TcECI4poPso/vCu1zjaE+09CHLRRk10CHId8ZR4h1jmsRl4L7vLu
U/p/XxQTzJ7Iuk10Zd8OG+khNULgPY7aJKrJnnVITGsLM0vV8ddXHbm7Oqjh5A6u/TCcW/0WLmPS
6ooF+kTCMAzHLsLK0IS9+NSfglCHcIhbdckSQJuWJzrs8w5m0EpwkkDhzFKgZmuEiyiWqiyMt2fC
VHIX3foSY/kI1SibqFfv3C224yLxacHxBK+vZhycaYERHsttXLKq+HCrh4XKAP5ZzT6c2Yo9cDia
xniDDbi/BjPM8padA1AdN49/iGvw1TdjBaVEjHqItaC4rzs674ENRNbVsiHjt6rb0PW+Q/1YTrTp
qj+NCOq/bTmHkw3b6pgFf4i9gaHhcZcbnXvKAuZYz3K3v2mtaeZmB650Eq6mhhs0vSiBFjpNrqHP
uLHJOgAPNj8WYhbiBCgwwaOKT4XGNiskvtMn5BzVKV8oJrfKG6gFa/mSljXdIIKeTvQ04ex7d7qW
/DPYMt7nejmZ122Deq0JlF8l7WNptBla8AYK5EYGrkMmUfaqrhzsWWYXbEZwRCX4FXKA17DiBp72
veFmdO0hcugbCWa+girZuMuVVumDziiczCgnwlpNyljXdfv6NEf+Gw6WWO5fOd4qHVIe4iLBEjBh
BPlqPKdEPL8DqbxB6+hs/FiI3mM8N8HPRL9+uacAO8fIJ46mIm4f2yo9vofCLhDVkVbs5ZR6dUJ6
dH9OPnxX6apExqJBd3KOlVVTBEiVTdyUhbw/C/KxjkAcl9j8YS+zOisrOQb51X6gRq43DoW8fux/
VjiFqvSQxZ2LfqYizWECO3nvwRGj8SaLFJFY1XlG+ERludvu9Ab/OCC0WZUafXagTsNhYeX+oSHG
YdIo3/oF+pxyLoenKkr3ueSxzM4JkJBH4yuJ6gxoLdVgIE/dWjyGZv6V6neOmQ2utghzn9jNBX1b
Qyc5BMe36JNv3veYeT48Nx0ozWFZ5sqY8mkh92zPInfG4uQJKzjqV5cRgbr/F6GO1nvFZdEN3+cp
QIEluYQHV/skmHmqpHVJsqru31TSxXjQr9QSnlOfLRJOEdGBlPIOuNpmozx7Y0h/8HEKfu3zZYCM
q3HIp4xoKFkhg3kEh3uXTKtapwyCAvpL8K47miHJEy36esMa8bfnuQ4j+s/Wj5BKp7rNEmV1XWMC
ZxaaoMk9hUgrTk3FWkV8cuv1FppGRZThrZ9CYM/QuGL4X1QdwKGmIduN+LZ9WhvKSBG8A/OhXL6r
xGz/EYDHs+EbT+4m6ra/DqtaX718klllkVVMcYSuBK0OM3+7cceXdgwg00dOrsrdXbbjiP63gRay
IAkPvE4X99pea2GAuS73aS16uzCHNv/JsTwfDfk4TpGi/z4194v+V6M+AU4S4p5yt6PpzFikNycE
PdEKsMUYvYI0K6soTcxEjuxKjE8vhGVbENVxRWaLaaOMTLXl9v5X0zB5iWhO/2AUIq9o2og744Eq
QHmPqtiYrx2a03ImZM6w4eVu3rnUBJNCGlXoIj2v0MXp7NB5minY+woBu0PGG1K2fbifsSQKjxxi
OQ7aEaA4oyi7xtwelKwax800z7tepfOOUqGmOphitB9s3ekYVlE9PPgNTpAvI6PgztrNK1p3glTR
mRR+3Vp1Ljz6NvJlvuabGhIzj1d6Fapa7dYdwuwaBUXcczaKnYgsKKtmfF1HaGjtpT/jTLgIy6Ce
Hqt7DM7G864FbL0UB3wkttyhSlampr55Rx0ntxXolBVm6qdis0tOpeWtofHoYSe0sVKSc7Uy/+rQ
oKWvIHhIs898rH8UEI4dxiG+oOtlrSFetw4EBAuBUgOR9uBywwfQYhnZPPRrLU9W/qkQb+kdzLSF
LSyuRWL5Lag840vc3CTh4R/r9+6VOktTjil1cJW7ub0Sxmbl7hkXD+hyQvcfm/DajMOn6c5HSoL3
uaChHK3HwRnmRWagmCwFiuQTcNYQJYUdKSBTWt7SwHcv24j2NLUQSqa+ZmbVUgr/tpB8FtCggA7k
HD9i6M6ftcfT9+bxFu1g32EgS4o3B4yug/rFrjLF/lveJfoTQPz1IuHDSUb4xJv4IPB/hsIDpn9w
1Hji04m7YJUTX7xzkjvymK6YVO7Ws5ILwsERHAW2DkS3YlEtdkoR3i4iffTyhS6bx/eUXwcxRZMs
HmUy98YcQFUVHkwurOuR4hh1xSHWsMCO24TvEeVcRf41M5wmIgW1+52r2heMBEckFZFLYEg4V/ip
16AisrN2w/WpHCu0KqT+NiLlUY8ShDeioU2so16YEUFCeHlWKF7+3e6/1DysTde9/7AtSbPopu+s
6b0z5YU6+jOcTkYCu8agGLhalJXPr1zcBS9+z5MO9y9JkaT6dcmHwijDPvFk1vLOUF2tLPMQDrRi
mLGPf7ForlfHS6QOvcyc4odvX2UIksGvZnLZ2tusgPZ/lgdApLhtfcd/Es9/Nc8/tChlH8g25T85
xQWs6CtfRiLUJHLwX7IJbaLj0HL/IufdYogwIwH+KpXJZ4IsC75bbkyr/KywvOa+a4dIvNJ07SAs
TMgInJ4dOukjt74NAlhcs8ErI3zUZNl2f1cCCUgE+kKVdjsWPjxvMvL4q0jlYsLq/o48sDQmWNiI
Z2YqsWsMWupzvZNi9ec9PWwXeGxehDUmuOF90IPM0rTY0jeZXuZO3e2QYkaV8SJDida4RakaK+j+
sbijEsFrXQILSzxEfi/0NEprE6fQNpxBa17h3snlOFI3C5N0EdPgXH9gmYqrDja8d3DIT93MGRaF
4EKLry6ZGTznyiX7b8AZJmIjWUS+FOumq2E4PA3XgrXNEDy/40P93Jb6qhxh3qmXCKiFWGf4/Crg
kF8w8gXX4Ns4rY95VBwmPG/BXshyw6HglMEzAw0EIWeYw2TtDc6IaxbBF/k3iFqkMjP9J+AuQSq6
VnS7wQmSrXR25wbKsTa7kEeFQunU/GklnLr01yLmbUAmU4asoWYYiY5uw1gw+c4v78Wy95qIC8u2
om2AuRhF3qLOCv8Sw3S7NsLzkYyk2s0yA55pmaI2VxbxMyfxQ8rIdepSLpdkcwK/sWBf1DPAY9xl
BHnfZj3KudsYvt7cv+SNK4S1AKtUM6z8HktoyaRf2Hw1R9LpdY/3RBvQjv7wvVhqrPXBteUunpmi
4de14JJAFi0+f2TxU0c+yormJjY1IhSK0gJbLXina9Gd+D0acF3ZrTePxFtlZToN0uG9ouywP1B7
lRopODyYJf2l5LBCeVe+LOXODGIxDtmIzw0DQY9xaK3/+g1oWm86M2HbPi26oHL8ZZqhV4mLV0Mi
UcFqBVrEu6eud/OhyRhsb/M9CN3GP4vXhKXefeiefSJr84QP8px16Y9tdt2xva9qj8sz8uUV0am6
uvj+1609xfN76ajIRfIKYti5Lm+FLqvuERxw1tGmBUuy4+FA6PH+BCpAtXdDs3AsPVCBGcXyjQVR
sJA387+QNZfCf9LVTQUjFgGsrYxj3HfBGOxQWx0VAVrCCB9C1az8lgDBeNQ0evsMlRqdUhs6RePr
y2OW9MPNqUPKNH+nGXv4rsYaRYlpcEI3YXRFqVn5CH5cIrsUi2hvS81iiPbUAf3jlRJYigB8tq/h
I4zPk+FAcJHV68gjT6M/GIDSYmW4wUUURkqI3mLAufcFeoUiRGdY7euTG2u4+Y8X5gb4vnPBiZPJ
7nfk83yrbrC9sCHTkke7NebnaYaM+qT0SfDZyhx+MxadVbvVtDjW+nVjV6teSBGNFIVM3k95gVSm
4q64YgDNK2rmP1Bp5hQJ1NVzMNLXZqhGb8inPpE65GAC9ykYoWOuMMD3kceD47lbO6aMewCug2n9
FfIFSCk5dfXEwe7nm8QAdNAzMebeLI8LmZ3W6NIgZJXyIxfPiujUS1JOXmWeO1K1zelUUtJu2aQp
sxBkq6K+hXJLSx5IGdqxGAh/G82GPKwt6yTIE6q0LKko5GwS9VipaArxiNbrGESqaSkHmkkkugcV
RteD+akeqEOrscRFULcoyqDNqmCFx2LScGmeI/71VldwXQVGquQf3PRC9qcnvhMVHUnFvTuge6cp
GJwFb4xJb+iU2Tf4+8AqPHowx2nvpA4QwwDJ3zO1VGnms4A0YnEEF2ySMPg/vlvEoJoFDhSXmfJy
tZ8QoFJjjZKIK4TSytI/A+V9GkxWjpUNCsgVrlEqT089C4LDEGxoHjb1ajF6WiwN5BPTEDaj4K6m
N9Os20LEOC0fb2RkPj4NaeoFhMBfqSWUR7q2QV1RU72pZmZbe+DPx+gZFRzH5pQVIuaZ9nb+bUm+
Xd/rBpNIGfipY0+DH6GzWmTG8ZX9DneWiQRru/jaGvh5gzFvdTBJ79fnOi0Ms6YnGr6mB8FUiMed
FXPE2w8APEV8YZQDi76fU7/UgnGvk9WJVrnSD4uf2PQl4CnL7XZk7LY6H8Re37DPqXbMg5bYXDZb
pgDVhGGienGEfQRRa6mbsWIQ7H0DxU97S8F5g7ktyqDjSvsYxzy0dO/KWQmKiYhfnGqsxptV0fLE
iezLJVi+wyvedoXvaM2CFUBm3E35OPRCsz/ng1yV89fiAiNUOI3mSGobWTtoe6tWuYwkRHSJDyD+
/3V1VyuF93b50lCw5FgSUeHMiTueYt0Tnw1yMxEYXgvNw53yCQFpcedCe90ZmPllRK0vTw5g0wNs
YanLO3PmKRG7wU2ZlJWWa9BGdgGdw9z1ErqWfdJHEorhwiyJhIm35Hch54bmTDN/4aCuRsrKFhvB
6zG9Zuxv9Fb2FUUVC5xKErMiLE8mn3+NtldXX49oO4xgBMRABa4ZGHWA7qtha3VfGeXLxkrTYZOT
0fi5j5qzRkrcHFqSMDsv6TnISZHMeDNYQPN4QubN3WsE9BbtceVW4zwZkxuftaL444U8jC4Jyga8
akLImcrJqxjgoR2qkFacQUqQpxIldyEpI69gOfpiEIyAYta2jYd6qRRXg4ITDQSndSfISjuWWLlS
6kKd/MzG80lGsiEtVITRuFMzqkQ1OS6AGDnz8Rn/9Im9eMb1Mk3PdW52Pw3L2krnX9xbtN/3GHUD
I8dkkE/lPYEuE/XwQ1QP8cKY/9f366fEy6FTR8MBi1k3N5NR69W1/WHOeuEMt3w7UrfJ1qUincWb
E0p9zFPKZFuScjSezO3gW0DU6SPDEMsuz0uUm/VtZcqlRARhUWLjHWxjQqg04B9oIpvg8PPURneU
KaETreHbW8z7auqLv8+qeS+w3j8AWufxYRdzCXBlqOpvx14rJucc3MMlOrB//Jfo2nPCK8JWmQ3f
z+foCPmTrD8ye1UcfrM3wiinCU6KOqk/HYU3zCt2P8uxjdAIJuxaUt1NcfhgNtS6X8E612nXcSE/
zVXyMwDKMLUOXsVDXFZREg5/S6jBAP6OHIoBUIgRyWxBkP0O4at2uB2mHxuyXDaD7q0wp85ycZLw
gIJEvXROY/qBCVCMfZrigP8ih9luJbOJp8rDuH0SkJSuXXYgtfdaV2yx3bNUDGVPD1X4Xs+Gc3Gf
wLvnIwajfK5t8fWL+YFTu7KlEfw7rq4lE/3JoBibHBRAh6+uN1zsma3kgSBqZjvRaXoCBSoxQZbj
x2cISTnlAaesd1/U6aEHklQ2lysxiA2wV0odukUQpUqsJvyzdqFojEM3zxijYQDGj6Oh4Z5mWMYG
Y/pMPhzq5xRsKM5loJ/ooUa6U5gFLwhuSlDrQXuRMyMssNVgoWw8x0bCAg2Do4NGidjjhNm0Fjxh
d66/LmdF9q9Ke3cQjk32KQH1GWEPGoJI9/mqq9/N365yzPOFZFukw3H/e4f8KBRWl4KsMoucfdJ4
m8gbdkwVI92wXGl3Ms4IqyRCIYz6vEUAULBT0gzk0uejynSC7j1pZYMeg6Py+s3ZUeLLrciUk+B5
DAvKQZQKB2ZdX11Ci2MHmrf/lD3/SeWv95mAtKZPmhIbxHNMFWDjQJz+hsp2iZ0ZSu8rgLKy/qU4
9RLTc1V4fF9AR8Qp7XPiZFiVRXp1R7pYg0iqLF4ufHTyxYReuI554/cgdMo30gLODbPy5BXV96Gd
IdTiZhGVO7btLaWxT80zRAp4dihmFCk8fOXkZmPxUunIzXV7004e/YmwK7jn43cujobeO/fNjWMC
qJ4ndW3aNo7Xxc4BHw5VWyJF8LYOg2knHKgPVCgG9zy//qN5B03w7XX6O6ffoz6+3KpIT30FvVB7
VXxwXBAyRA5rNAFd3bExCKLX8GK9+E/zIBjfguI2AvOXi10hBsPWPCzYDZp42eSPDPBhB6WtC+V3
HKeE1kK08YQRyNnTVNDP4VVH+Zz0VwqiJ28+EIQuK/ftZwka1RxKZBovqG9AuK2RxasTdjWap8cK
U77xcS39mO2ZB37RpUMGFL6a6AC7RaYk+DgUkj8ikvokC5cT9cbMQpxTlxTzajyvRhf1UolHolSu
7o4M+P3jMahNt1DaPCBhhikI/y23rVgXFY/UwNUD6yXkRCYBc287E7fsL4WuvSfdnlnf2GLkPdGD
MaLkCzODEyNTOcAANueqATr2Lfe0VvHOZO/p7mkqSeZolvzjo6sgrK3Bs4XVkEOJ+lSJ8O5kST9U
gzidB+ACd3siLLGnoeBX5+q0RikD8DjZnvA56aZlPbcYCBueRYmhSvxwlOB+hRhfWZlHxmhILviJ
8hhVFeTOIGAtjrsxsON2EoyEG6mwX5Q1GfO1aLKwtQLz3xs+Q4fJlOC2jcVd22g+VBrEzdcPlttW
BDCGGxucB40vE1tgKjlfyBaC7CP8OlWk7j91+UIujAADPguk41E/e5IPZxL2bF1Zh+JrvKqVDGGs
gRf0pTRn6oP14hJkw03ieHVZ8lPmWsPkuZ9OmjXkL+QXB7lYVr8pi17sXnJ/9EF5jVPLJZ2ymTwb
0UWNBD8CFEVbUQvoQ64Rsevi/kMAxWvfeWafA6xVfeMD4AiR9UiwTcWdMad31GijqOq7mszTICO7
eiSJmYSOKzZAKoH21jRgyQZLtxJRIrg04S8QSi84PW9/Oz9aHHQ8rxEXOkDZvidVloTCiq5YeX/e
cdzooWOg1zqUE+NfOZ/mLLPp8n3ljxoPagffa139Xcjgh3LV0SH5yr7HaGxUzxyTCNS5VOLbCxKs
z/bSyzYAS/d21EPv4gmY4ZHbWc4l36KWqhGQEFyG5vezK8xCLgEoSiV22xoWsIBeiD72lf5n+Cyd
WKh+GOPi3WYoBzEssaFG63WIDxOjWGJ7Jd6J9bp+CMmi4kfcJJ33EqdmPDvPZjJ9nzN1Ba33YO7r
SollrKSrbbT2qANUKjkWnNxh/Pnz/w3PVoMtvwjxKLBbocxbZIyWuDI5S8uP7zoOZiO5orIRyvj3
vijRt0OJedEvvvSMPOrBxDohi67ug1jmxlXo4Ne7Y3cNItKJ36LugjtG8BYsAFByeOP2I7mp8V0t
bHHbaWlDACe6VGZYomTvuHDGPBVThqSkzWC2eNyXfuImkpXtaybRF6EQLSvr3k0HxwtdIsrXSe0g
q5VIPqb4TUD7clOnm5w3yJmPGzbT2x1H8W2sgagZaWrGtl4RpT1tRqWfQjHO1+EToHwpjt4cG6Cs
1N09nEiB5+Yv+oFkspT0Npg6zm4jy0HGPK+c42h8bny0o7kBEg/ro/hyypOlvsKKHxCe0xj6dyCU
HANUXBCMzzEdR4qCl55tMMxus882FAgV1Su9L0Qe8yn5ZP/OsLSigHcz/yXohbLzzBl7drnCHdeF
HOFDyWeN+AptOQMM91SUXYJObg83Z774ErTOhjUM2D1ouZSpIW66BBZHxILpOSf1RkGNqHowXfE3
ZE+7FNRFGCf84EEE55hNMHllUQFD1FkgAUbxraGxyisSNjdQLkyli5TRngmUsIWsyVwaJ8KD3ZHp
awWLwlsqd6xpHc3LSFCDaskNvgRUmgkktzAJcYE2xVPhoBHpK1yXTwHOy8opHvYToY7i5Fl8awHZ
f6xD6RpuUzphct698bXLJqVv0FNOqInpvRMfwXngqZOtIt58ieP0JiGPe8ZhZmzyIIs/b6ExtJHH
OBBiyVHZ2cGGVK/eDdcFtevbIY8lSKPBH8hYg3+xRLHdkurotvjtiSqUsy1LTUtt7m9gk+LM0m7l
kTMd8cNowHGl4VXQiTCwpC4PYjgfgv5KKTtVCRn05Z8T8mT3g55upY4hHm+/eNaXqvU0MD+tUdoi
FnlHiHVUpuDGXPCUmntq3HKFdxXDbYCprDz4mIvebIP6IM3mUcRMJp1ZOEu5oaTvBNRsiKqXcU+6
ihq2+JMJgTn+Ie7FLHN3LI8n9srf/cKSOSAmaCnkrmeaiRoFWWEy4ilCxI43m1O8YOO2hJlRgf3J
iIoA993SLdk0Z2+g+ai9FOsaklCZOLpKlgazM3oyReR84bcOmyD+POAnjMmdUfziGhHEdrlk953W
CKXWrsSiA91cWWWWGdtUcE2H3GucUNw/zFFPmRYgP88BYbmJkIpprKVMq9CrJbBmFSpL5uDgh/fI
VYUfO4jpIst/dDAEK10Gi3fTidpWB2Ch9sG6rgPIbT7M3OMMBE5JgbCnvAWqfaBOMUEicOW7fmJO
kmCoZv3OmtSlSLMIgfzRSV1BtV12V8zdB33aAI+HjuHSM8UISN5nkZVtMM5YIxgGiAFTChGAW7ZO
Cb1fstN2DJUafX/xOd7AuMWsDNChaf70X9r49wmZrAhFxQ+JF1KPfKqTGi9RJmf4gS26FGD8ZLda
s8mUsyKE2EbCAAK1FvBnhzXwssv3RRYJrVGWWL2ta7iZXC3HRLC94/RNhCtAHJKIo/IpdIXgK3j0
8u3omYF3gu1BJpgoVrXBvvklKOm0MWKWE+k4hbpH0QrBgJHSZc1moUYaoGSZR0qQHNUhJPfO7h7/
lzzgSqnBgqnoXStt/bF9Oz6mKNk94KHEwPbero4uV7wTJVWPFpM2hRpJTGx02Ba25QPGPvIUewuM
XStfHOdvnJ4KTwXiKTDVIOM4xD5lVW73uGZvOl0m1GizitgEpJW7Nwp0dJEuH/xEnQ3Tk28lAGww
ai0NET+n40hFcbO08UlyqGxYNw5X84hB9q3fsxYINh+GQ1alQDvuaICQRmIbE7aUnHg5mzoIG0tq
EviTJvkLQXl7thmWIWZQwJ9QlVoKqiyFOoaJlql4iJzlBMg/E0rzn+g8/JozWOOxaRkgQj/yyk4E
zQ6f06Kt4IHRYCfxsu9JZRG750LIL5SXa4KxkOVCIyING5Qty9jKiERK/0Qoy52lFQ5vR5APx24q
wSFVkihAxkaRQwIElOx7cR9x2EtVsIjFEG+1VCMLX7F8UsgFJgxu621ZG11flZ9XtBRtMNDttOOD
Zz59pIZNsxChipjdtebQePCMUmrJ/SeiDqQLJpT1BEWjOHophMfOKRA3Dtcob0I+9jU3+d8c/LoT
2lo3UexfaKbHsNHzXsHsfkFPL+gWEaHrWnqtGz887oGnwYaLMnuJ0uPHc8vzWshDh1sWw3yh+xNo
o2B7Zht9NLyDHUA5QEYLhTzRaxmOXPQOxcC/UsJ6nOiI/tdKo3+uyQF7xPZWVIuqe2fqKVEhK8l9
bfqPscCJMPSr6a62g4Z7BKR9fUiULIFjDkAhLfPIq1dN2yJRU/OKHV7xtgOy/NAYeyOSRVHaWvbD
zuNzc8SbWWNXV5TDnTOaeOnABsMVS2XabtemgoguJG2J5DksiAINl+ztvrIpWuZ0rTAisbduaMMb
mGYjLEhFWUtbZ1N1OSvBg0d4KbdjeVpLUSS9JaERfB7zO4wKBwWhIwjA2mJ9ct3r5VZN/jsn+s7b
77Rribe90TbrxZ7nu34eNaAuNwmKZf5rvo+DHjpHnhmPFc/xXsa+NIJ9PcV/1v++slmAOsUThmcn
xiLsM40/XJBPdgO18IMehw6rZK4Ls64xAuCAesnDoOEXmoJUiumiZm+4jG/ztyutro22E9BMwu+a
+iD8+dkKxEQEtPrLuliB5ntabNRSwhwiRk6wleI+sNa0iOQMCbpHtZ3SMkW0WqGaJkEvzofqqtdw
HvDYR7CNQ1zxC87m3PSmT/ysMufRZk4es9UPspHu6oxgx/cII5c4oxbpv9a1hSFFAcmlCbRPcwKd
GIDEf1pKLem1QBnAkKFLH2XD5dlJt47yULAiRnBSsAU5InuQEBe0Ha82tYRuVTdUFnTura/s+mPx
jchlHSB4oBNO52tmANKN1xyee5RQpq9acEAsCAesqF3lmPvqs123eIAwEHGSMl4Rbx16F+1qGcF5
fxZ1gxrvZGqp2eCML16Dl+olRSAHDsDljgdIQqmGSEfBiVi1xPKHJpwgz+acJy7x8qBa4C91Vn03
sbuaT67U7LgnCzfDRk5Uhec9/5qLMlM7CBARWeA0nxwGb10Eu2ATKzmhQzJiq3LLu/xURagmbHNy
96S9fgs5RTWFS52lJv0CDO2VbBqVmREIJf5dpd9av9rRCpJviyqpwMhR9b15FUMFkuLlAt61WIox
l10JN9xZ87Cbf9Uu2Qx5Mlb/JML8JgQ/wXPVT1gKoFUUSxVZgf3woGXzDd4m33tmFEUExsgv+DEb
oLyWdOny2OwoBXZuQuyLxRYYh2hbCM3doK4tMPOVkBspTa2p6kdN8DOTOt7zhVcl3B3FCpJD3+Q0
rU2P7zRVGsDupe7JdhIM3gHUD5Mn3cfqzyJu+KLwJheTme7pKFd2gNTnYwWBtDT5OvDCvjDxjnRX
nzss3o0TrrygMRr0PyRp6Q8aIgJNl5yaKD9qBpLSmfEAHuE7/hdE7l9nPLYRPbzC7/3gZS6NLK00
kJWY2jttYPhz6D1GGDLIlGvD+ogdnSTL11LH9QEDh3IdncYBaKwHFMYppzN9rR+fnpQfhbIqp7mX
t1jlHqe2O1epckQX8l9ef9t00jCDuHQips5ZVwm0Fl5WnwBpZnhyvdE5P7wCe8ZG0NSHX4Yyxpvf
4PRVfafxPagcBq5B0Cym/FEHLOWKmtdbIDT5dxhgZlHIKnsSO77cb9ML8nytWbh+3iH4QVQX/GWd
HHPllta9QrobjYQ1T9Lg9zqOichNU6Ex6oppwx7ensV8wVfAl5S5uofJPjVBC9TT3frt4Vhv6pey
++00GcxxGrF40YK6A13+cScwj/fRHAM6k0rVeCItLdiCOXjaYEJugjlpJ4eyWB3dY7mi7VqWssFr
9Vrv/yALHPUDC7KUt3A3rzqpljY3IbCpqEOlQ/I775ztAXzG3if5yBjrLgjKdW+q5dhLgjfHSqmR
GzfZVmkB+FNaHaK/TTh3asnkl+S/VQU/xQ2yqncNo5UPuLZ27h1pzRUwMU2ABN/7wzbxA7FVYiy2
GzK0uNCCM2NKAQ5kn8RmNUGnZFi3qqJaSd3ZB/eofZkgQcuO7jnX5E9kol3dJV9CVd1mibRklXlo
qMx6SrcrERENY3n8DS7J55XY165ks38NZJQHxtE3HufjU6vsFzE+GzhfVkyM1NumLk4MJ3fPR3UG
MuXrrrzpSaVUAxU7Po8D2Rp7hAercp6Niz3h0hw083a6yD3ZK/3ZbD45TsaRjt922SAUiKoUBdW4
sjB+GKzALh2AJxVSAYIXNf9m9uR+7RAVIwZYOkcQWOYXvPR+qp+XkgOrhBzQ++cpGbDKvuYTq+wh
hwbPSKSmTsGX3J2Pp//0/BQndLl3ezjK0HhrX8b8y4QI9ZLbb+9UpZfARK7l5vaxk/mMUHX+kTlJ
LTfxKqVOxrQyEWNF4Qsnuz5KZA5Mdw37RAvi91MgoAoSPUxvpAFbf6vrkHvofCgcd4fiBw7TnG9k
n+SwaDmgvxZn3yioa1OyHG2c3F14Lxtn5sivuL111TfvcAkKWedSAF5JqqgOKkuEU1PdZcHGNpPG
GbwgewPCErVzlP7PXPzOLTvkPpIzAqxPJmjfscuAGMTg6HZQNYFWGapmxwKvuILUNreyD9wuLN3m
/ZpZlBflsd10yS5PoWpYq5QYQdTqsGx0tAynwtNNbGHk8LPqIz52NXGki89j3GSUmrC5k9Od3kpq
cNsGx6k0vKw12eyo7hTf4X91ngzkEXey2IZVKmK2LR0Fmx+VVld37L+7bEwgMI1PXWGtkqpdZfBE
7YicUBPchNdRBBL6SG/dhSWbmkBtfhsY5WJN9EXdtsP7/y/8X62rTHyWOW971jcEnfFoOw/Y+sCr
qAhEVnwUX/Y2XGuwH/0bo2K3H1SsfmNMtaczcHpce9YaY9/SJBWjp5AxP6JMLe4WdVCTnT90jSFU
Qocf29EEY7kiNaDaZjuhLPex5ok3nkjWvCJv3dF7/HwI2kt8LPrUFgvcleXmnCr1qOiJdpDwS177
zdhJziFhaBwBaE3laFnV0L8yNRhrWw57am9rZ9Vv0vVV1KYNq9FQ6ONUl/qXhWSiNJhHEwKE3rIc
5ELO55xLuSF6s+9ztN1FWkkEZvRd3WBSg1axo88AVKUKUuqXCfv7PIEHOPO/wM+bMcIdIoBg2Iqr
tEBBfbC8F1k2foSTw3LV/MwoVWks+tMXKwVGpZkhqNCqS0SlecRyLfKY5LB1hDv+69WBZLdQvdt3
cptFbXICQ51F6z2JoR6WJJADHnchOKyZp59oObxsELXgUR8UXC/EHTfoR+kOq7wYKEOgOjcXkWaW
cAj9NXJzKFi4CNZYACClh4p4jTWDQEoGtONOPRFcKBQwOTKdhYjsUsTfXsxL7+amuqoqHKIb/jfU
qmYP6Ba+nvwd5pCEaI6pcE3P45r2ZmoH/VU2PD64xKAiLWuQM1tEvX4WuT1lt8Yf8P3m5TTB4ZF9
sIOl4/NY0OC1BFJTh/hKcKtz9WIXloBssG0ig61wYYwzzPK8V1jtwcETQ1vex69YDmkrWNZIqSVO
XPPqn0MFP5ZGN8HLP5bW3zOwc48S4QREwa14uh/g16S0hQ3cBwI61xKtstuQhC3GvYkm+2/36/ar
2qQJUyR0dvXfL9mMPAvQqQdln64wV1Lor7M82bn73nELgqqLO++/Izu2TOKCa0uQVVdJfWl1zL68
L5xtTHEnOKKUpvHnMbeOByrbRwyHve9VsBPfIdbBN/k4Uk09wgFhuAdYxQoMWd76+PEah9fm8cYF
gHRKX/8JANJ//jbQndA7xalT1Wbq9Wmwm4HryLcg0WBgWChLaRYqz71PUtTtRBv0sfQRqzTgsx2G
MWNmoxGdY+SGLn8lugcbi9VmrJCvzTbl3pas0Io2JHU4GO5cw60YGudMtf36vIrwkc4fQOIi77WJ
sd3YkVssZJ6eadat/W7ZkikJoxFcvDlIscBUseZ5PdedqfMmHsQBK76/cmzaVh/mbegWHzxwO8/u
7d0APkG8vX0i+qjoO/XbOKZeXxtDxvdUl4RpedRx7qtl5ICZ0p4VD/vJ1zejJ/JHDubSoZN0r1cO
xbZZzYCuHNg+2iC4vx2K5j+X9UeAyw+IhvGtsbMdOsX7jBVhvdDFX0X2DWz97fukvh9yaUHV4ioM
jCg2oFn85svI+/FBfwBaTg5F/EgL2d0EAn9gxqO3q/Kd12aUk4ix/6kl60c+qctO3Rruk8PGOwts
0s7dFywDpAGUYX9O/oAKiLvu23QPmhUpAUpo3Nsbxt0reKtsldblcv8VVxg9BdKT8VtsVqeezeah
GszodU84HPrpUaE1IYzC1+iKSEJzwblrE09H0XhZ58Z+Icw+OqvRh5a3brNe5tpvSivAEHsqV1Jg
NB55yTuBLN5YNjQF0Hiw4KwPnbC23BiL0HwON/Tmy6sdwRbzJuJ9j4jUladovl8+0aNc/M1B9aJj
jCxoNjB1HcyQ/rHjUxRtTslUkLiKheWKMGdohWoMzCPpoyrYA2mVmRDiRyOpeSUBYs9ieSgOacdt
mW049406el+V87oCzJ25Pxih3LNbcRveFCHivGrwIT6HJCINtH8TJ5MKJWz/jgFIpWkNAp53eO4O
JLzlAWSMdCVO1JYXEXXCB7q7+1Y7SjAct104+JHhKXY+bsttgtQ64cOn7NkUkK5AJPgwEJ+8gSzr
JNwbnhjhiw8VECEdCH7dQNEcOSy1HZjt+XBJmDwwO931S07tPgtXG5GwmKTDkRspnsWsM2pF5220
ceJosTtsLXLlz8bR/6mcEUezGjR+Gx0xceVuqat1m3Atl6dvLW1S0Ve19Nf4POTyjIVRLM4sL/3A
bP70JbLEdpYrRH1acUNw+qTr9C7ha26Viz+8ljsZ8wRaGoDL1bVT+GbmRIiBUvJgXYNT3I3QzykM
/kJ2dHqclNm5P4kuw8oXfl5MTdMpZvIj4WG5czLuAH/y+n/koff6yjahajai+4HadNv8XPUnWY9M
TmF0WPqRTk5VrVOJeQmgrU3EH7QM++xMz+Sli5taGcvT+M9w/QH4QQGw4L/hX61GQy7xEZ2SaFK9
2Sh3gsxgNpDV3IZQw52epJeWVbuIs/Ow3MiBqBIsCDU4VhpSh9dpabGto1fMLUuqMS1Tg1wT/SMV
I2q/yi6Kws9yR+bZKOQl7oLJECHIdZHDGRsY445lIZrokuBrnxkFwnUpT6j6e7uXPzAdednjhUYV
h15fpfUgiAVrrsUTZQvltsadiLHkipJD9OyvGUNzvF5zWSf6KBxfunC2hHZ9PXqPlcY6WP8uxsoq
030d5uPE888uzFgYhVUfSmix/TzMLVmVyDCB2HRjXEh7qM11AP1mebx26hiQTLOnjp87shH3RMFd
LntjwP4nAWhz321g1LmyzgLth3nlGBW2IqJXjcouG2hFt+cg/aGtmmEGB2jBu5BbRzxdZkvtBzbC
I3ybnFIAOLgL6eoIkmzMEY6zpF8Rz7zkxrbcKCXuDRdAnqfpmzFbRY2Empw2FbrXTcqYj5tOQFFT
lZhWJut+f2PTpC/UO/DV73QvS4d7i2UwrE3qq7bBXuD/0uNMbh6jY+oG4tMTTTh95B8y1KoiQjLK
SOqe3hmAIYRsK+HL8DI6Mb4OI/55CXHKkrUXFZZan5snZF49QqYWrcW3GXmE9h2ZO3GZiNUzY2cF
cynbYXwRYSBtKX56yyCpDRlXJX+HkaZ6Xwc9cH/r8whEhbL/ZWGtfOz5iOv0DDouKVdXw2f63GQs
cIZW3bVt5y+GXEDprI7Lpg2sBp67KVMCGQwbC0YdTa6pmbV62VGQk0IJ5vuz5mp12YsaX8m3ttSa
Seq3MXp72WaN32SLNscGIMjLIfAQqgfgG3LvR0/OaW/mB1mO4htL5Wcjzm4rq/otNrX7TM8YviUa
VUdFXJLX1s5AEVJz6sxzHuYq/+hpF0dVG9Ok7tflfWgQWRVJ5+iZRVpwLpgQ21s7LDZ4nXcYyYNk
p6pAIX4zHINgfN5fEdZuxQd+ejc33p2bYNR7kTKw313CZcxnlA3HEXXQ/I89QtqWIZ5xPHh2n2kP
7ClBfQgb8FSizpXkG9CzOfjgZIgynREixEYdoPCintkjijbn3TwkJlv6yMIb0UBx7u8+8KzAq738
aJOCFAozY58cPuNl7+UZ+U8xLLyeNUCki185c7J3P8HMOSyD8wJyhbJNlxAfIQJ+24glcoZDuWC7
dzajEAhFOKcCFoYNTprCSh2+Z05UQrFKp7u46NkWrfKbzNbqScDv1cKn9bc+NJJAaA6kImQq4NqG
HuiFw8qQBg+7iH8z/4gXiIzEH44BXg24U6YVD/CenZoxI+XCPN2G+TGOPvcWAQT2V7/uYJMjIbMZ
HA32lCMw6QOoMnL1/Bze2CUjdcU6Yw+ZlBjVtTcYbkWTHo+QnQgeD8tVI85cTSFdNOKBg5ghmDWt
KuEEj+Z0bZxPisOuRogekSa5qvfeSyGkIQLfy2BmlPOBeWYJk1ItG0DNApPZr8xpMg8vrNJjVCUn
f25P4cxDJBkmgqbBME7xcqD+XsI5GmMGC/jgcIpdLR/FzQ9Jkpj7QCXal6bQYIxmyWq4+cZ8NrcG
MNOoD633cvtoJG2MDQaQvf3Do0IHlmt1w9bT7NP+Jty90Y0DkYMl8pZJmVm/k1p3jNkaz07bHR+y
Hw3IVpqMbFDNkqv7kNyeEbS3FC9HBX0A7aPOUsTMQqJ4uRVlu6mNAkPhnwy43Jz56vxU3BJHV0Wq
z/5XMhnKoDa1UbOxEqQ6Y0t8I8ajxa/+m1TMn35NPthwAopGteMu6LhA6PScjzxiOB245SEFPggl
aC2nYvkqZ4B/YDOE14kAG0LExee1gtAf/McTt4j1sDAWDn1m0IuTILphJEJ6ZgMT13eqJMCF9r1l
12XGZ6Iff/51svXFROlPidrPBow5GZwa0ORi3JKsSmJ4cjmCWFlvvOo2KEdrsFFjViSc4ZlDt3PK
30GXhdXQadTeCPxh9kyGQrsQcR2SwR0D4Szn7NfCUxrSLzdDEa3p1ZEo1qDYSHZ//cA14CKlveMn
wHedSfq1bH1fEW6edfHyCFRlxjpynu6VmC3K2O0qnffO8+wYwpJ1oRpE8O9BY0JzakLxq/z/fpBl
1Ug87uIy4tWYjbTO1PnA0AGs/dqiobFO8lju9vwli/y1P9+Twm1r3TU1YpWg23asBD607VMKFpPX
G3tjZj0b/lsoKS1gXykB/Hokl5dBcRe33q6pqeh1Em4thIhUqMYsbFtDF9TEc4Y5RSSFUgKEEMGO
N/n+sDJdIPKM3QaAPQdP5WForNn+5rGpQ0Ly5+xZMxPJ45m5dMv3Z8RF15Y+bzf73nwvP4P8NzBW
UTWz7nmocw1RHq2lIN/t3fRX5+8VXxmE7Z7+xYwvW+XlQlg155KPfEX8mc+I/NNSuxgZcgf4gpRR
tC96V3lRvCnX/xdeWW1Ii/8aLHUQRC54VKVLjPzttdtE/5YJ72hQpXqic0P/CTOhOU9boGn8rWPd
YEsz891GB4CIKczpfTv5Dxk1w6hmx9BQrRu3HO5qz1+7zKWqeo77vGcyGuuHAL98l6hSk6Q2DrV7
OdSmohMOVU8nEQJpvekDyFBPhXNKXSL6DwRtyYsa0hgYnRdzhRO4n8Nz7o6TBB4HguZ8FaUkNyat
kGmFAcPUeXxDvFXlTA0qhHZjSy92Zb+AftfVmf54ETNG7GaL6rBtU9Y6YXdnX1WzdEB9jX7i/SAr
5Y/ECIT8d1xtWWI4UqVgpREXCKD31DcO3YlZbKUU6Ii+LbDBuYyu8B+WsujETK0L1BQf/xo2CJWF
jhw1I+UC56Ycq2hWW7n1AMGQMEL+M54Kp55QK9tcGmGeSKxk59Litpb4I2S/XSXj0vsDGbY55B77
o4Qv+fLPCVQx0psP1y5Ia2iugywa/Havrjbdxu6AwpeY/75+0qg/N+y7XaBfxe+bNDwUYQEeUDAU
tZKyYKz5pBBnvM147j+LJYKYB6Zsp40F9V44XzAfSzRCAK0/pZ4KHPs2gFqVxvOsu3Cvebv4Xvud
enpDr3nBbsCvRp4eX+d3BFMwG4Zc2w8JIIIkEzltwCRyjoEeAmz4C4TpZidCVgK26ibXWxF6QslP
BVnL/8qgcx6ZcqP11P8+CkGPr0txvIPrxZPxYl6s4U21HwjCkKiMSu6lcVmgv7C8qloh/UQKo3YS
ZUmBTlYUZOgwsstPiJfF/xlD99pTBzMLOJ/l0Olu6NSpu9JNaVSk49AkOwhu4ED9LbEpweDe0l4z
6K9+bLvbYF3nZmsZzvzqQD/McPQp2eFPW4iNu0ZzwrgAlJQ3b/aDLA2mpGQUpfLG2/ImpOX8cGY2
mCBgILFs/VvmjDw6WQqb3PosHtelpsLWW3L05RMWlGfSmCfbrSlTJAhQlPmV/Rf/6/ViWKD0T2e9
mdKTT5SgVY1ztpEmTzO1AXMDBB1jI3Z6UCAAl2Tavugk72MvjvrgWNeonM0I8duHCWKCDXyzrMv/
KWGGE5WNgLgYS1LirqpbFAbwbYd5meZegGr7ahH8qS61BF1i2PbUpYn4T2fOizB7/P6rYJat/dL7
5ub0Ap9eWIL/NvcqC2wQKybkepukhhy1GgbgVuw6MDY4piWXosyxDe+v8EFLi7JxJoZ6xUcPgC03
87/HKpm0+tiBZjQ6cVFkzcadL1Qphv5Vrcz0zH182xB49M8oCtRYfACbQYbGLZVprAuqZoczIpzy
YU4Fa3quIuPdt+oH+m4QxVeiqtk8zT00DqS1MAP/WrpJaKe+v2bMMLWYFOHBkrK8dox5PGEm/qqm
sCzlan1kwnzVRv5gBNbIu3VlQ4Ezz4ayEJihmLuEnTR3QDiYsdbhdZ7m6rAbI5/SqAMo2FVB9zZM
ndHEJVKoIz8aCm2vd094MSaRkpB9Aw7Kehp3xsdp7JDgeLRVaz+jS04CXtH1IKMyC2xrW1/qGzTg
MdmfAIidprx7uWHV2J408odnM+qvrj+459+HA/RGGHWXypW82MAqi81Yd75JfIu48deSnJBHJXVi
X/LVsDWVRn/kLBBiZtkaXH5TZvTfruhm2nfQjkK30BfNmVzxJlpXoe3PyHFbmDtLldOX+6wzXyfA
NZAmDY3vHUDvFiWjuxFnu0XU8u30ua6EYuVJpn6WBMfoB/OAMWfrUeCLATcgppDR8gMHTPDcK5VK
9aAQ2+5Z1V7VAs6S37e8cInPpdRebMuZH/Vq/yU7CD39nP4MpBQiu7DjjK0V6zuSE5xTrQl8Inwl
huPuX8XOkhInCJpguW4oh4b1QglanzDXRmSH4Z4ACPMV46y5ZFImX4Lb0+AxP2hSlahYfQLZZCCS
RKvjm5iq05wyJWTCRyEoUgcGwmQmUdU2qMqUeeGCJEB0eaNkTw0N0tIaXxXgUinSuyAIDNxoS7dW
kM/O1QcJBlcjtvDUBqyRX3LXO4KfWupBFoo5rKtm01/oXpI4Wkc4xhOqOp7xVJNtbvb1NwRLHnCH
TyqppF/Qjmw/gL40c47y1gferNWNuJOcBgkGwzJQcxHYpmFSLeh7X23+frA0C83nIz4WRsqZ47JF
B2abmI0VUEZFVzAB8DIGvMF4ktUdnC8Nl7YiI18e/o5COJIj9XvodPKIgl8fFMYpIWEKkSJJw21o
Nvts9+7g+f3SnvllyvCqqSvg7BfKs1qIMf2ixsbJ/KSkTo5wJuBGm4J0sJ9r8bTM0BLy0PVqc9gb
no7jqpkaACHzdaBuZ46hGhtH9H1hXmQuoFUwa5+sff86H3mDP7Vi4VVGiJMaVJ9qBRre+B71PhpK
+ihV8okY3RJc1MiwhjyXzu01uD72n/+6ae/6vxaAu5SSWIZfhHzvedLcdMNazpe9ZK89HKqNc4U+
6RpUI2VKP5hKXTVByQIlKkERlBBE2njsRvUIQU7eMeqWQpdQ9aNzHl+LEFQAGWHf3U2bNMMg2L5T
fKHMiuNwnQuX3VZrEThHltJQKOiSvSOQkKUnp1IACsAJtUHICTs0KMEUaGksVocDqNC8powNAJj3
2wAWDcq/gpnjKORSBZdprYmFcnxGpyEzKUKvFj7aNEkUzbtuKlQdujartOW+d2z+4onCfz3Qd4MM
AxT4IQBSXXDZAjOCBGkm0PKYNj9MOZvtIhcOMxxLZ8kfUpxK8V9MVg7h1OZzGu77UhpqwuuNQcAR
+Lma/Mz32E14doaNuN+R6j+RHVBADEzecEWaZXfSvarK4qg4i31rDCteFONtv6Q/P53tKHiaQRl3
gA8HisZ008pwduTzvosmd6MW4++amTubh0CuxL+vC4bYkCIU/3tjF6k0soQz3IaYrt0THrMdN6ZA
HG7ziSwb++4+UXODRJavxE3+8xRLF1IHfG6LqwX5xYzPo7k4dxukwWfOiHQvoUz3CUjjTHhqNZ9H
ffT3U3hrh5RtWmWiaXraxKzpR8EPTI2pWbKd2ej0DSgaudvl/bf2Jg2Wxgw7iISn2RK+CJNKcwMl
pP8tWMmxcZ8xMJ2dNbv3vwNXuArfFMyW8aaO3kMYLNPidNiaSGENwzBtJhRjRtTKnLSN0lmiYrp9
dD0+q8AJyXGNt9wHGujix0EajNG/rExJKBtA1rGckaoyfF60nfa2+iiqMz98JXRiOrjGR2/LRU46
hc1aMH4kLIbSnrjB1oMc6sPceeOALxtMuDFAyxSTkKhO2c9QAS50/R3XkozyhfoEXHm22OdNQwkH
QpEkRXmTfQvhlpKCB1HJ3gOJjWXOjDAGWSXAD4hlDqyE9Pi1Ms6vA5Er+Av/zvfnRvke5Q7fBGFF
UODNjsTDNTvgsIs6Wm4/dEum0EFIgnaK6c/Ip2wZRs1cx/V1xsEMCrNcUn0aU7fHGz8xK1kYxU8k
B4Ra48NUB2PQo6TcFyE9yO99Vs8NrZnyyc3vNW7Xj7hH2QPCNvNbRsG0NBlSQZ1NEcKm3KxLhFKf
hQ2PcwhFY8j00vcXbzNPHTy2JUN/ao8uBil1tPPIyJ7Fu6j9vmgRNpSRviZwXwHHTpEeAORtpOd6
wRaYz0dC5BDf/jMgRwCsc0X1PcfcIjfYSOwsZae/IqAyZrvoCld2AOzLOTtlln/VtWKAvlITIJo8
wwa8EFpK5rjz1UGBKT/3Dc/zT4YLqejw7e9E+W2XpwteZuYy1BFfd9dw0XHn8JfpgubTZgtYnlYF
7u9KFCetRLi0gCpO1jUI/INNm/MmxI8Vq5KRyfiS6yVuv6ogiCWC9R2sjDCSkYcZELytQpxqAoUs
LRQpNk4xbm0GxcvmkJKmBtYqTlyJhZjeWZW+h9i3DuBZG3F+t+1OTprS63FPw3AFgSDReVJk5Rmu
ciBDfZ+38pZmGozI5W3nxhmCZb6vBf+ekWnjTl4LzOT8j5HY9po1naUjSklOdsIrVhAcYC2LI6ST
Ol2Q49jmjRLcx70gT+TEf6wfMCynufSm92yb6sd6Ntu/ucELDK3lXZw7Bu2Df9tWQpp1i5RXnK7Q
OQ3vTFcMs9Fhn1prKUbHJOiheCstJq0KUtFgGw7xvVzgdvIIem4MFYO1xkad+9xJztCXT+snf/MV
O29JfJN1cUOlbgyN/h/7NzfZw2dFxY1I42xrFiZ3juOMuyzLPKZAWwyM9GRiRMjK0Ztwi6poAOLi
q6yTlnfIHzKwu2pD0/L6RfPsSbahrJZ4kai3WN2bnpDdv6YLg/BvnyrT5YKcfBIUzP90k2/mZQJ9
mQd2YF7ZVvRbCAJYT7uhcSwSYNG5JxWjn6iiudfmgItI9p3UMuu/MhzqZuR9ohjZcKEXI9xQ2YEV
M0UTOSJz7F28JI+5ObDeWIiAEnLzKCrLUs9FBwwxLLKFRFpqAZy0NfZIe9sK3hoAgFg2A4kpn0AG
fyIS9QRIzRPnrWPrGTxbGTM1j8L3yoWxnqvgOOzrUr9UYNymG33PxQoc8uED9LxbRy3MTocd4AmG
/O1k6+AtKZIXTvyJ7sLthaUfrgTCIemowcghEH8TH0A+a/VWaNZOBjSh54r25Ah/2+ddIOwjFB6h
b7aodpieJ+HaTtC5gKSIB1pO9ClfHZ1blvOHZiAhkSNE3kzHgryaMQHD+ZH0zWTPpVMzlqCy1NnV
cyWb3HGwskTOSWWHZ5obkFUhr/t1py7yDqotn61clXM/2zrq700w5Kxy0n7e31lcejKuDs8eiPkP
U0C8Eu7zRKY53NQzyxl+6XqeXCnvNT1aCY8QCC4UovS8U7VWDotP2cV7GP8Uwf/ZUGD9iBUyBDM6
Npe/wcQaH61qtp/1qNreMU6MXjWkk/ElV/sbsL4VFWLS6kGM9dkYfi0ANsXl9+eydMIsx9yqSqqR
lBnTMANWFAXvxnpU8nAKTjXWN7jzQqhV/ZdFHckTi06o2Xw4g/JNltXi0oedUv7uPSjPsIzB83bO
ANi5le952EIlT3slOU50ycQuiheIoRTImwSgWcuCpfUNTzEV4IM0xVQ7IrieZcj46KKDRuK+7Kjf
5vep6lU4ZRHMJjTSEacATMr7tFm0iBsW1sVvEHXRbfrg2iFGjjbxM0Zeg4ZAxfGV2Hd/yAP30Smj
gLMgiv0oY6WedR6cz4/z8FcbVvEJjjNoBpBzTbYwabNei7N7o8SfPC49G0VLsV2lvyEUBbpdrBVK
WB4nVBEFrAlqxB4MVscM2nafo7qHOSmEN/dQhxhiAbfb8VuLHDsmNoukk0HbnjPm9R5zqAo/Y45E
IW9OS9Ut+4cSCoJeo3bxHiSZlhbadtBRfdWy450G7VvGsYrnh9ErujXppgA+xA0a+d09LROHif+f
SHRGbos+41v+KSxCbj0PQnIAtdfSzDHtyKukNzgz6wDWWuTDYBSK0jN8d5gtB70ew+nvzpVuu+80
6QIdpKzraQuKTlVrSpKDQh2rCcV3ccJxLyG9ns//kovUJcJMu6aFICPe3LOkcCF805D0U2fG12JD
E158pMyhe1OJDL+qCIno5HFblsDl0DIh7IKq5pLDlbVTgEq9kBaqannSfOQXApLLWst0NP8hqSMc
o+CnCVBPXMVcALShaapNotdHc9nn4ZHBwiI+xb4fZpYzntXt7QZEOACRAVl4JUDWh2MKzEiTaPTq
4wQPtLAAzMzVruiXPw7VhsamTNcC31AVL5UWumD1g0a7420AVoHWb3ki7G2IFyb6WHO7CP5g1Sb1
7et44zaLJf47r0i+Ft1yQADXq77LF/3Pl46mzhsX8xq4M8vKKrznty66ppkKFKdSV0K4EiV6atIt
LxbwJMCxT30DlwgzxoABth8IApFBDh25eVPJIvnIjJ74suQhNMYdXEgFlqRgTaxdbSwiQppYFkrV
JLurRtKhYcwTrrRaB4wB7mDRn1qLGpQyNv+hupLfWuANBx5y7tY32Qj3Xy7WkMyjPu2qzuPTHOsd
Q7PyOlU/WnZHiR1dxysvaFxVWZJXTHyndgpizkn96IjYqMfpxFt2ARziQwLNVR7s4DG6PIw60rxX
lwvq6+j81biqHdWeBk1+9SJ+AECJcSn4nBEcKusjvvtEv/MHEd/5zJKjXyyjqFBP+OZVc4SuV3LD
rhsLKCgHM5ghZqq5NUUkNUjO0AHSWPDUPlFCW5840ebgq44fTPEikn/xq2vdIVqcvqDfHaczFCMT
iEc7DxW4LGbtqr6GfkU6MrD6skQ+Te9rGgMxXHqdkUKP49I8a4md0uLYfDxt9kuc7voLcYOGLB+C
GmxwE4Ykg470MRNrdC7E9cx9m9V7GbIThwkLMv/lR5iZo5hXXb28XZBA5ZnG0BSH5FBL5bWQgvUY
um2DUhv/HxBa26YCO7TxmiSR8Od2z+KeE1aVzcUIk4E2x1sqUaJhD3tB49HQWJT69eIrWDXFImxq
XGNJzme191Ag9VfIw5rCrOddzGoTZR5DNExdrsR10YGOwXFiQtOoHNB1gq9Ovj899P/fI19B6XkV
cZbemykVCQU/w/S+AJNxwrxBINsipc9Dy6feiSVaG4mutLd3YEP+ECrkNwLllHUIwRqqgst6/mgJ
Od07PvQMbtoEU7jz7Nce+SIrX9qKEQh6R18R/sDThYWIIhcN2o6ZisOOl2Ed9dXjXomAKYPhQNzj
fhXKWg3E1qH1rwB6PA0LA0keC1fGkPMn8pnrk42bKlQ5nllosG8mi74u8WeL3rHLRKluxRbokvpO
QIwjYZl9XhOHPSakRvNBnvq57mgPI5lJox5drzH0dBSBpDmXNqkrhQLMlc3CPX7LyafX97DrjVzc
FetMUFT5BeEBkDmALylvQXuWAeOFWj3WJarQG1vFO0b3kjaY/hSZtKQi2pQ4ZmkQKGBlI+6ECmTm
5zoKuQCVRYpV3ZEqGKWuoEWjUA9Rbdco6DkcPyc+nK6qdlZb22NSgia6SpYHlwhu9W6DljiFICUS
UovSsr+quizRFZ57gv2LGzEytvQ3LT0gK8wWy99GJyEqf3+NqIVdfug8AOQ4aCt/GPl0vT3iFO8L
v+AwUSA8x8k6hFi47B3Cpew9oSzuclwmZmP5tH4u+LofaOWsQaCHD3TtpZMYyxy090WihKwNx8lb
X4lxGHQKuy80G56iJJNfTqYWx5a246SwIt3+aWklWmjeA+FGdHSn+TAGP/aIfwDUp5Lea7jEkcA/
POXArMWMvj6ZmDn/QPevWq87MWAO6hZYRhWJ4k6V7MNqSEKyYe6f4hTsigJzoJ1R0TdITYVh+cMr
uoagAU0aVYN/8vWHsaEkD8mv3PUrb/qQHd0I66Nebb4JatKjCEkVR9EP+GjPfX89zVVbxL11nzEp
+aX7Cn2uIm3EPDFerg6BgB7RSIYTP0gGnQrocG2a45pddnJSOdRiWrxndIrnU19wJFl3JFtEWUBC
AnE+KMpRG39mu2xtMofh+kvuoWu2m4pslRwNmfOpnvO780/PIDtX3CDdx+mOA7Q0KegrtFGrE9r1
S6NNSO6Br7NhifWOJ3dhAY/KezWM1kj+6y+gZIK8TM3AFUFI1uCmoqREw2Rx0VQw2FLjOvVxtJmh
uOolD0vgOoxRFziiprhJcxUtjBM4+1VOJlROvIwGYP2pNjgXj1H5oYQan6h9ATAo7TFk6XcxRwfU
T/IglJ9QIVCckZx5JCUxvyO8/c6v49deKnqAzPwJHWHZEtHKcB1AtOnN+hBZmQ7OWDTeN6YDxHQ+
Mp8pBrZ9kN7QNsfilLb/h7xwxQGtoB6WqjPgcd7lL2cAOq8+hotdXdceV88swqqLOL/afTf6YfBa
h7CrLsQCI84la+LIV1d7i9uvrmWv0UIynrR0Ow9Y+2UJ8KxiEIi4J7LdL/b/ZVfao6re4x4MgN5T
zKIz6DUqrKuLt3P7trYdtTUBrTPGfhnsGL8lpSqvgdVRcHcmnxQ/G1baM4XIlz0hbC5kVALfLz1R
rax6KML4KhTihazQye9G+d09y6xCRfy+SyJWZDB2uucohRlVP7BPGbMhL41HZFe4VwpAhm7y6LRr
7nwI8Kk3vYQmk4/777wT3oswA0Wb8dSLouRvcRs5xLQxKsdPbbdkFZd09Lmu5I7Xgjdqs5eS8bRC
ML2S4UMLmPREj2CE9HHNllkH3njEalJByHcbPUJbJOO5uNdyR+CJ3r2RrvOX211Pg6JwMXEz0PS1
kKA4EOEIdJI8b/soXKBA50LrWqkMYIgJg1RYvlZJtf+mVzYP4Uqwc++tR7JndrmR+6uwMrI153wC
yalzfsBPgOjIQ7elPdWFtHaHlvozhiahk9rtqq1lvWSPTCfEnNcMlNEGAhMg+t0AvceaQLUwwp2B
m8+igjte/AoWDAW9DjuS9gRRmJImVv3djqSkq1OypLeAQevfTLyDjgMdzHjTnzQJe+lF7ay26gwo
A4myqCT6qVsQ3xemYBCqXN7pwFOGjr4QbCvzIyFXZJpqwYjyCWxtHKAJ7d7RbUcGRXrBEauHMDib
sEket1T5JJ1M5sW1WNq/EoD1qoEfIf1fq07vf93dpC2l7xKgFhU3reGuMuITMk5/Sh9KdQEkMkCW
zZ0x9XwR0EX3d7U7Rcz0EYzIyh5SZA9VLRGAlK0HWAxk0YnD2uW/cOeov8F9aCM2MyyhILvAX24N
Gm2yXh4lxI5CAmksMprUg8VA7MwdM385WZreR0oJCOiPM9hSw1TQJT4AUc+P3LjAU59x9EmsehcP
C8MAv81ZmSp7toLHzu5w4xaTFbHvG9IqNcUHWFdWuBkHcLh1ZIEdJ6pVLtfeNny+GZsgfUiz/4ku
e/tNUHS6d29J63QAWp9LdABbYxzgHC0dC9v1fOHQa5QmAzrA3wb4AauvkRb/9kyKqT2X84UoXoOH
V2HEgNtRAC04L5x02DCBpenydD3EwzR0Ido4XPbtcw+Qs4KyUYXTIzxx/kwem0TOYMjvRys9YzjG
Rw1RuELk3nhLEZC3vc9UD1VhDIsQs7P2G34fOnBhXMV14tXWhr8dDxktydIeV3Gbw73Mfg8PQWt2
ZGpcql3wCSFQQTYvXt//YQztEW7Qc8b9i9hwnGA2YqYT3mIzwJid2Gex079zSeYlbq1iT99GhxLm
kdfFbKbI+LBOgqbEpcT52xyT84YL14y6iMq7nDFNNKdsT+aylX60TSC1HyDXHOVtl6XEnIi3B6FA
05U3iu1RvXtoLt2GX4xhpqTEIJCfVrerHt62gSYzwytue4vJrRjnW5eqYfsP0uE1vLoH8UUCw8bt
1P5Cz4YrsWDb3QmOhiunc4H2bn20Vkdzysc+ha+KlHOV3mUM059I5vlKeLGtVUWCffrszl2y4X0T
79/KVu0SpIX9cMy7nVSMK7cdRNKcda4mzGAV0ZcNU3swMxfk8qqXhpM1gJxI8/3hgt8y5HiUH2+V
0xf0rM/OxS1yDBF8CprSIDXiZ/1J1PHl66H4XBwiPNRdB8mOsK6hILblx9zOJgDxVtb6wy/R3mMH
zmkbfUyTdpDDMfE/5dEYi2lgT5ewfKdadV8iWk7pxVti7HLZi3sTkTDQxbpTO88zOmcrWliA8OnH
PoDuY5QcsAIcAN4NCkcCz6tpAiRVisQLiH2+D8WxCmTPAy8Z8p0FVIdPOSDRfkyCM+JeIF+PQNe/
ZNVFCxYlgfnNYGuHgVdUJTi4Txya8Yu+A+vaWKPw4A1AAIy5g86uGg4QWDOnk76a5pJOkefHNg7O
/7nWdrt7cIzD6ZUOUQp5qzm1eNw9dJPreJGwWXDE9t3gTPBIbgT3JeDaXKcR4T583Pw4kqJTysd/
kuZ0WP3JwuuK+0H4mQhjh7F7l44HXpOmpVC1TxrgPkRbV29aZsXE4Eo6yxskfg1/am+F4VrQJ1fv
UBGyPkvvUJ16Lic6++rzTE9iTdDqUhZedTVeBat5Ez0eVtzTybNTBB2hcjd/t4ceW1Q/kWW5D/38
gCA/ukRo6r6zDLcAvjxkMWCvhrUF4gY70lz+VRZq/RqrICQ6ViqZRO7wiurlsXluxnuXTdQ1GXL+
k9IacaXK73BVhXApnSU9+8iBYIn3Uh1QJ0/8Qg0RvJUCMldVOjeNSJ+eeEt7u2SqfdegW+D1b1y6
iLhlRFbWAzB0s1aWsgF3AmRv2+3Q10QuGXBXt08GcK/RszTpAH59g+iuOmBZmlvAszB7gIX5/sTb
G2TktJ8HG5RuIZcQHMQelHfdiVuUELuUbS+rKljs0N+W0RHHc9SgWN2WXg5lXh+5hbxot0iGAxHj
7SUlfLz0cXKlfFVd9zONaPW0DVCOp8H0TR3EQsxr1m2QLSWY0sJqjy+jtuJxo7UoaIaoSEpyVkkl
LAGwX2xcaH7Q6RV7jvMniEnf2XSS9p35cEv/mMkg+EN27RWmxW/sOg6gFRuY+NrxzlJTvrwExiIy
22z3pMs63GcOTnis4w4bSqqDb3IoDXIqwETKXVTYoLB/3xvPs9HjpwFCWMd46vPTbOWKKXHN6Mln
QmHCtfvofk+/7hq8Jv+g7QYCutPdcdEEKZDBowOwmmXXnB5OgoepAhvzOUR1E6tHlvas7c/8p0CZ
Du0hCQKn5OR71vOl2jabeQcH0+wGMmi12budcdvwdALzujR1SzzvS0GlMPotvualJ7rm8Pu7XOho
lL5MMBTGIeHY6o2zVUqBGrDVosvn+9vJOxJJFi1rSoalEC987cDVXF/xq5wkwyA8TROI26kPuG1t
QcpFzgJIgYUwqq6bqy0rKl5an/qbyAnENyi5/CuHQVPtMMjCALm627+HFdUTPdCRvI4iJpEgKRYl
QKPv/MaQv8wSxHKqvoKmVGdfqZwBMOCVJkfWYh51r/1r2BY0s9mJBPwOUc0IAo/x4rPJNBYmVqnA
XNrYz1cW5saaspggYQqDdEqC+XAHc1dSF2sSg4tVxjijQd2M7z0B00mPFGeiirk4v1ARf8YXXNPg
QQXjZh0Js7PEzOxQ6fE/l/AzHop7VdRF1rYz6ehkOFA8lRDLnDf7VOQ2v8U4MOu8uiYmrGzdTFio
pAmAuNw0f1FU/9natqI0Sz/XVHLeaHfyeEmWMS+llPeq949oa61wchBZuCgi6gFj+4SJOFAu3O+j
8dfGeFMJRcS25AP8gCfDFGbKU9JHXV4mGHhzUnzgZpZaq1zgDMoSXwjIpzYyJbCltQmh5pOAxY0S
hyO3fsY7jxcWvZEd62vVHOFdvEv0eRY82lyDHIp2zGZ5e+Lx548P40zye38v4sMLB1LmRz47T99y
EjyHDPYbUoq8Jhw8IXxSvAu7P2JjDz9mXce62Q2798/Zb9mngiTGbdQs9DGoDhFDeoP3aGgtyNmZ
NUh0s3jEPyYnTFo5qu7Qg62HjWUCfRKmI1kT9+hf36anWsneV2AGUdBCKgBLd3lCwkOErn9HrqT6
k94tBp/YLvcqNA0W/rU+PoVTMUgfA5LB3BQCQnngVrn8Xmp8T+li5lxn0Fs1dg3p3cKU7z+pKweZ
cqMOoMt+jPRYzqtTq1HQVmcoT85hviix71gUKIj7NPZwvC2bq4cuAWOmFDMkkbehw7tUasIRqt7V
TNJL+vgd7o8Lcye4R8TssRUc43ihmp0aR09LLuPsEqbfEfCYChrto9yg/hh69ooG4bGeFtDCVXYH
V8MQYFOw102+dNs1iwqz+AXbRuvg27QNL8iVf+OVhiM8EkwgClTHVuVq63kZrPNQ1AAXDRSEvH/R
OI5vrmz46CouONS9XFzR8CShpiesqytBMTKF1fPntNRYykRpZAJBNM9iKLTfca7H0ep3dYGkWhu/
VvspBkLG8dB6R8QNnzvxILN5uKpnwuqpyzaXRSbFYg5pFVNgIA1UNaSaMfeKP9ELPRdNqA0JE44f
N3SztYIPSNhDx+cquc1F8k7epSPEjC2MguZXFK3cncfld/yqWJuUdUqPA3Gzb5PouDDS1CzuQgrc
r7ZVDCsq/kkxFesmXxsYVO52AacdilPWRrK5A1e2Lv20PmMiVIm+qxjHESBye7Lcw2LMlhLgnNca
UYrMDkuKh3mA9cLE5kgy37pRdteObgyib+qkhpEu7K0RXRL8Ei9bFZh0hqvGZiRydYAkaX64yLll
De9RY4FH/mGOx2CKejm/S2kN5yF8mJnuPXQmK7PqGB3xEo794fiWSQoj65nxkel/CCpmywOQYHEt
uNAEYaesNXDunwqdMd+LpoaaRRadfA6Sf1hDEr1BlsPrfQGvWP9Z89lClOe3eswBQJU84rvIkd+P
Wc49PRA4wHLaBwhV/etk0St1Kx1yQcxg6KcE6hIvlpMJXKV+fqDPIeEplxQVOBrBjKfKbCG5mvOW
C1sGRmv+2uKsg4mhfsKSKe6jQc3skWl2vnQk2HYZ0UfPrZ7nEVUM5v1qS/JpWYUqDd74nfSTzUfV
1SCtsICf1fOY9dLZRLjFz3dQwbyq29EAQAvhsj03xA3+4F7PR3uDpWDPFOoNB3VZCbCvRDvVW7CB
/z7o9VYyk99R1hiLBlJKpnH/S7AaAoRVPLCGbDH7AREzcjbe2DXyyafIIkhZrwGWvRraunMG6daS
/n1OUbv/YriM93eoXY+qtihCnL+Rm4XZucdbNL5D9wInuTCLsxnstnBclgHeRZn2a5mJMG/ErjnU
LJJ9pU69IlWktbSZfNQCDOFwQTjOGxzYCNJETChRrWkQgB4CumlMxo1ClKYUfQby5WbbkcjKKJ5+
EtxSeqxYljcXrsmN2tQlrHsqLn/p0BniMwKhR7VsFkwV6ju8Rp1SBn4BtbQ3qW+gryTj5L9AGcQD
ucvrAnKzvvGmweTDWgeHcBZJaFsF4eZkqVgPN3JRemENs++v+r6dsktuAp97/yaBuuvj/JO6AtS9
OnDBGkH8B0tL5ySuqnhVCRIA4FZTKnSOmM9CSHv1w7CnYiZJW9ubFPz4FTb3GMj+ovBN0ytW2Jlu
AVl0HrEtZZVbBKl8wvWg7PwgSXpv+5QobrML8L7CxGoC+4njJxhwf8cZciWps7LXALd/CIOoHh1y
Sq5ZK9fZACcIRwGdGQwtFV3yjnXClwEnPqdUVTDXNhj9UD4LZZxAy129UJAgOVsSo+4ZZQmtg0bj
EbgHH4pKSM5go8+XkBCWIZkb000n9tyJMs/bWQ9V6b0Gf0JANd6tGd3zd+FZIYhNrJDoZtdQCXy+
HSPoPx5ULqoREwhZ5/0pcL7SZSFQ+gNbGwdnVjI+ytktRDAr7yU5HXTv5uKYpdPiItz4W3Yaj3sN
o6L/dB1bDL51b2bKy8XtFisuwkwNjFmBMpdt+6nsx3X01UivdBm6HqyEhILz59Vypj8v8rGDEFW9
rSXlEV1iMDHj3m8/czT/m8q796XbwAqBw0C+ZG2v3PwF725GBSk9tmOKdb2RDaf+bD0xeHFRF2xT
9d9a2GXabhIb7VdHiWbNmMt8KAuLeGnOVKyx5cMcX0XJQcd8DDCe+cxtp/JhT9XOgb0GgvvJA0Z9
9Tq6ES0VO8TM2DXbvC+WLV639gRcpDWcQFoZ1/aQrbf2yzZp5VFAfR+exN1c1e7QCnkP+lMrGIxN
WPhkX6m5x7rV9fxkvF91G6ZWKTGnDleg88T7rgwmBBoQv3Xib/zJnAYj66G6gNh3+jk7Q5Wba+hk
7zhascZ+ONC7JRtdbbQGmnUsxA9ctqfZN0NmgB1juPY41w4/QnM79QN9iVN6wZrEuAFrtcsJBXTF
no/4Kc/y0b3vL5naualDGahW699UiQ894ROkE6OtlrnSpTyh17PaXkIz0JhjVRJRBo8+G/pdjZn1
krG2msJM2b5Qe+c39N/+6YtPBoBVypRhDxeLoXDOaBTVi4l+tW4h1w5Iv+ePII/kHUK0xoxdESme
8568ZL/4O2+ExB4tfVVZ+6nDX/NkWOcQKlCF+AjajYars6w1RYtVFwbFGjhknfR38TKM3O4gZQOD
lH6Ed4NQGicipEWNmp2Lbn0IGB5e5aohLsHskN6QLMg5MczJ6LoPc3tM3GEif2Y0laaMGlx5Yag0
aAOGmnzgQhE0FZCToU5jgx8AiIcHIWFaB6RZv/GN3RpUql1OCmglyFxIxtL2LWKI0ZCprYm3Slnv
GVBjhQsYeZLruQpwgcAMOmMR8ttewmZQ5k0JIhjdO3e8/1qTxFXCuhDQNT4K89aMfYsq7jsQOk9M
XRV0jfE5mslDARL4LBJJzjYTR4X1DUmjMZQcncJWsfMC81s2nxyBSy3YqTpvtlNLJdhzjZvgnULW
jPRhidG/kVdSokK83BrqLWhvdYz+Q0+D/ylw0Ps5a2h0CgAK+eXQDeTDGUeatXORGxXUnlCPCE5R
9VrvV8X5ii0Qaiu/DH4cqra6anZzfrUA4xYAOiblnZkyUjAHC0oc7wdEc1NXsKflrGSgtBZ5q8WF
ZrbSQW35y2etX8/YpFkfk7kgZuW+P7KLtEJw3UOQtBY/2hoAzDLYmlSrU4yu14YZI9MNZSLQX8Nh
M22Ayvw++SYICIgQH9ZAO4CSkqXLM0tH8dirihPh9y0vpE9vbSDJq87oXLlu8gE27KdMj6yun77E
SZF7V6YrIWc/kJjhkUH1bb9MvhEe9i3gm0aLvawPUrFUS+gJo/9Uk930yJ1fsc2Naj+WqtztWYYF
RrxDdQskgXRGQMfhEcuYnCEVQ1ZQIqWLKXLVd4C1IR6r96o9eAc5GbZBiSsnUCf4ZHroUFPfAkCO
R7r7PRW5TjyZwFe2AkneSyVyeiNpLi10YmxrmCt5C730qmDpYUc1O4AaqFek3ddcJ3SClo/W/pTN
qlfw1knu6Uts3xqNWfqtKYzRMaZ9lUcEw6DkQo/3NyH7vqmZ5PYork2KnxJ7FXP8oefyC+qabnQW
zZZIzKhUxo3JjvKGGZTzl1pz2dsXZaBYPjETLuZRdCwQNAUjktFpgbiejkx7wmtMCHCp4Yw8qu9T
3YmmsZbvXjAlkNDjTXScEhUR2ZVwvl3MkoKcMpeEIL3vx7E3SstIBNVTLEtPOhG5HRlvYrtSptm/
6a6em0jnKOe8cRdKNl0BEbFpR4pGCBfKMYZa+PbnCskuV9s1JNesirt6UcfARlvysTzHwmBJVfu4
L9ZhMJO86f0NmVIKc35iRS7QER3XosZiDbLZMXSxNNoNT/fPLGdHcaZjm20CxYxp3xfzjjxD2A2X
Pc/r6sESHxDpVGUPXROVheDIIxt0Cgi7KZWPRMSg6s2W5uiD0z/wBRaX2DVE8xX618jvzF+HrRgS
A+JpyQVPXovuB+fksI8mMLgHRpx+alqxaJi+4//3th6w6UJ52tuISUsUxze3e9pPGh+8722msUJG
HzJmU5/8CaShs7Uurno5oYKd6LrrBRX2OwtRO+4QInDWjFdvdN3ukpQSYVmqJ2ZVtUDh53JmCHtg
0k7Dv1dKO1+McDb8a/ImmNOsO8y8Ft3tqexz2RrNeL9KdDRE9XS9qaSKzP8rblF0pa/nWPKF0uh3
KOaos7cNJ98bx4wJjDkleTY3fn4Nfor4/jBVzgOcETZ3hpDCMW+GCqyn3clHjAeqrzn7bGIbvdCY
s0hZxajTWEOMNKUkRO/4e1BGOPRUfsHpjUd0g+3RAVk0LV4EopPDPTsamLgkIQjfXaZa3eW07GVg
AJNw7EcF+5RyjJAr0kyllmoPNnKTcT4QOR6MExdnFbOWv/X9YjDOyeMU5vUXiH9Bahic4dce46vH
a5VlrTxBBViVHLNLFKvTqHwuYEnDSctHYKLntR55x1vORI4Ad2YiV1FgjC/1gIek0QC3lUyhOWup
uR9wxEsNjXMCR3nskXgoiiQVi/GNp+n9PPS3IRUoOa3tACMs3c9wfXJR4Zn2Tn73+SBjUCPv8OaF
bHl25ucsBYao1KZX4JR0tlmah4jPHjrX2BwD2sVYS0U47H+oBaoAug6kB90OLkHfX8s3+Ca7jm9+
ImhehHamGZLuyOrO/sCnTFI7J1DWE2ZjgdBzeXn4I5oFasTxOSj98Dv+CtBn54juYelZ+m0i4CPY
/MxM+S3f3TvBqj8jujABR8f7UmuZx23O6cSzXoFMPffDyGowg4lR0Tl3a7V+RNggo4SQtxFRZQn3
0SkuPLxK98H4wWr8at40VgWdfps+n5m4U0fXF5vrsRif0J6Ahtzh53O1q8Hr3hJ97XLjEqU5U3Bx
9+kSQ/XLnypyOT6/MNC8TC19UdioKavkKzrIaxzlvLuut8I07p5jpnUL8j+OOypQm/7Mcqg24aeg
JMsruQ6Ysptb6kdXU4l4+zFPZfANMgsi5i5aaI4909oCRsSPDNm3ofZ05e6mdRTbMjs/wQwtE3eV
9j07Acd+SMNPmstKeHTwl8RLgBgAJSebWTPhcHiDIxQqjc3l7s+XewnhYksydtX6zOiZaBBNYJQ8
1S3Niahcz9lDVJs8WV03NDkYtZI2ln8ER380OLIE1E/BBlEcAOL6JFJk2U11BCLJKbvLnphzET1d
Axsm0+g70Y5/YXo2Zc5TWIuSC9rY0DqTXgmI/4KMpLS7iPBP1iAGrJlcK+PhzjOjwiqBxGIdMY6V
N4d769digFvJjid/OJRXPIrBPo8eDCgeDP8bvCzOdgr7CEbIvjvllfSeOXDpd3CUp+vnv+o5FM2k
wfGogkgVbJzWjwz4yMGZUdQtJxbc1C2JxXtghPFA4CamX+FO4767GXg5Okd9GzD8KrVBcSNl7kLS
7qPz3UKMpRnXma/68cyryj7sCQH/NFfnTAqsvZqTnBLmvTwsJ3th/DzvPxSpC6c3IVkAx5xePGLP
c0DOzUXPadqKmp08birRqued3c9StiohzlbWLNuUuuyLMqCJYpXUl1tubf3KPl9K0D9HFtjEKufW
kSTdaf9b2KhZKT1D7+e77z80hZhiQsxeBEXaCtOFgYgCGnS5w5L5hY1uQ3m2JFPN7rUVmzX4reBL
EcJsn+TuiVPLBesOHYOd0PAiC6AfJd/G0J/HiiFOOHp5piuvmnuB4QzkN4y9cdWABa+KgZm3DvCx
tmYjwBlDvWArSRsJ+ez5eTdwQE3oINwR9llMWBTchWuo4V5JRp5ldx94Gl9xLKLyflDVRETJ9sD0
UBR+8XvdCWC/j5YxvX/c1VxVYpNowUzntU2F9EMgjGMruFb4n8jebhLhfFyGkul5XsI/2x7AD01q
PXFxMKNiJroPRo+dr0F/4ZuRY9YMzied1pSVxWb+s5TXShSdIjaB30Hk/eKJsspeSC37w60oY33M
L0G7uQsE/VPakFeOsPFdd+K0rNja1lRA2/HsnQhwExDZ8m6R8nmrZmRTDB+ihTYDCaDiLrtHtCRy
maP6+77JHPfSGnHlg6Fn0xZ0kIhSom3s8MCwXW3STUwwAnU+akTirTH5pDBiXtwH97GkLCYVeW70
R4BMpe4nMXf7SrEpuCEpMox4nfl9/HWt6Y52ft8aDcADslTZ86u/XRV9b2RTmz/jhghLtQqczpYp
uEzPOYAOioEFUHJmn+7qn5rSUFLIvOpqCwoW+1puNcdUtAockDfOVQAa0UkVi0JqD52vTrvqIi4G
FUnyUqiqoYtQq/ShwvJwfnSSrHQlIAI7OBAU54IhtUSIEg/dbrEHs+duGV3+aSU1macByxoR8yft
8Ua9cgVNX/s/0c7xxioklSJIqEYAWiE7GLB3ebLC5/VkgfkBeu0nvhF2Den5dGZpT5g5JxhsqWdv
K34mYc/F5DH7JjoauS0nknxYWOcVQGwHTBWBPobDmiOXC+B5wRRR/TLhbJU3HKgI+fXdWho0NPLs
twz8TaKepESw5KbwM/zhYLxEaC2I5kl62ViW8A5Bca3DZLHTpwWqn3kgtQ0bIsfs2Xx6wWqtUE8I
FGmnDTGXzdTNspWeEEZmOFOntM5ac+Ic4XJmnH66R3suDPynuCmOp8fzJ2+xkmVKSp7PwHOg4Oo+
9ds8OgsVSWvHnKA7WIFd2I9tf/z1uT0Fq0i0NaDxznT4x2KYjDsBaKY4RUO3ytebQ4W5/sIxHFGs
VJXkDQ80utZ7Ou3yCTSPGsBr42w1YjPASgHq5EjS8G5ylbxLrQaA/zG5O1ANk+ddySPWOxsbRDVB
/SBLN4yuNV112tMtBIUsApCiM5FteuXPCsZ4WtoChJbV/3kL2kc6uoW0KMKvBXGtgxelp5dzdxt2
7Mz80CTR2Cbu+039tdzZsir+Lf7dnepUeiarkrg+LmcxW6bNg2YY47wMqFkqMRiFu6Jb7W/YdIKJ
StVLa7jc/9HRibCe9K7BqiaGG5tcH+CSd2E+DbvP8HOuRyAuyD5SD1AdhiotyvCqsTPKFrfSZRb4
ZMcoGTUOGeZKdD1sI5S2qTo7SUX3cnppMXFJEuuE/qsOVrEijak9hYZ3qL9oQUuVVrniXCOtujV5
eX0hfINW7/CCV7/IVtMTaLoem9hNl0jJyQf+8SUlpIzoY+TpOUtesmaHjNgbdYSK7RcVX9DZDqbh
cdy83ZEkoxx6jDNJBp8nWpPzznxHnO/GcmXfyfFAqSdxGamMbzhdnKC9Q829Uonnr7SkCV9HtD1I
P+Z9KdR55d9uRFCSHGEpwTKMtKY1aZHN6PpmCHUfO8ifhtNRSxe+E7swmMk/dzXGr8pfbx2lREgg
0EKsEXmVKUbkdUjdRhw5Bfn3K5M800I7vUDEK0tuaekB8Zug28E9yA4XtSVIHGWb2O1b40Hp5YDi
yKaf4fd3ykRJB7BYbw6DWUI+aQHa6giSfG3H1f206MZ5oty9RWgxdGXz6u35xh6bgDPBjqe0qGKY
0bs3O3X2wrIGd2fegjNltYrQhVjuOE36t7PRiJBhOKYMmJsWiPijwxZm5cr+ZIu6o8jNCBEB3Ica
Q+FYbI1ceQpooHKNpZRJTpQuKwwJYWOb9CWf68exLuecHlf3BaxAHDZZLbj9nb/URmxMoSewvnIH
YO7oiqR4LRA80bPB8vJUDyoxUuyFsQF81mATCSSvnVNGPIa2nBXzF1rroqvngBrsf7WQUcDwIQNY
6R9xtR5UABoKHO75kW3uvMzoLKF51VSr1wmZWnVFpdb+tKKK+lu6fJagIbxhY/hmsYpTqB4zHgpy
YWQl96TeXTz2a6Zd2lH91k1R+woOyJrl6I4qEMkMVkb09wDMKP6pohATttxCUpdjRMMOoEL7PgUe
NTtQdnFLlDxlrIizgOdg4aHZSwcQwd+Wf0ZudvlOMh7zMMh/DUhRbvcAOAJtGWoTuvAASRpKKN82
LOI5o+fWBe4dqd7naE7VmAb9AAH9yWmRIHFJKoMFNRQ83mUdIE4lmnOTEy/tQeJsT61lOxgvUSxU
JL7NhapuB97d0kzQJARqwsJBGHHidtUkk1oZsq24FY3UUMGAK2CaITNiPLCemsKxqZs84HBAU2UB
VP68LNw1xhJo8ZRbkjZLmJf4txMq9s/z5vWW436dscXq64//tav/Vd1u99ryuEMr5VJ+UvISlDyn
PktVy48Vo6aq8/SWYT+h8IrnLOEWUytZYEnMjvYWEUCg5m7GJGTR9fGdmGC5wq4gSbUMHV3tzOca
ZPgxFTIPfFhvM12u48XedgwLe8sFLysyfA4WZBU9ZrJsetBtJFcnqH+HqbgFEx5LdmJ3c5Fk0YHo
169D57/aTol6jcGNBN9IzvAD1OPVAhTD9V0rNkcyrhEIBfncBW6r23sKpp2E5OMXpwp//bdoHiWl
cjef80o36wqB3MhjQmHpCFNkhC4bv/VRtjWdQYEVt91OdMxXvex91sFd8PNtGYe6THQDXRL8ubT0
xH1s/4n4iR3/KNhvX7Mx5MFT8yJKKE+V2xFTmJMGIB4h8xe5Lmk7ihPE0DWcKOzUFNfbsQpsnX1J
OwFPJioilptlrRMs06eFaQHlrQ/5+OpOYZsO0/VeM4anoE9t4bFKmlKn60+7UFEwrPJDbwx3A+fS
lcGsUPUPscyDdqzUxRw6SKT+Q3mlHBc5Wu+4cSdCI139z8/pHnY8uriQ5psdYW9LiDTBJSmf7FbX
8lW+eaSzdHMG4KkVAiabUuoUUou3lIqIu42mHtIj8090EbDrvEYvl96VjV7wBpSIucWrT89DQSzC
m5BebAaC+BWDgVKJwus25H1fLERD8FHEUtr9yxw10CYuSy7+TD1RRXHgtiMGHwYf9FiYydEr1mug
XywoiDjhUnYq3s8xHkL1Cot689eNEqcO4BHuf3C9AogNhGIWxhnxaHoH3OJcofHQJdkh45DTFX8I
sqjtiie8N5+nF1m4kFV2+1KqR80fl/cWUtTeYoFUQRgqrRAK1baKviZ0mg1rNLehQgBzU3z6isXM
F64quCH47J8rFUANzpsBZ4dgkxiUyLDyyw/6sWtvKUkQKI9lGEvYVmE3Q4NQ+UNgcX1nZH1whBDs
NPSIpC2aI5t5eH3lO0Ru0sLR0A8Jy73F5qNOaa+UPU/dFf+eP1OJJBjgio6xN28FURSeSRrguwOA
7zt2BMbQFNvvjJWQIGOAzOb/wknva6rdsAdP4yxjYgyV2jgILoWB7b9gpdw9sdWxJAKsVHNVljmz
nkxPVZ/9aZfIe5BC3q7y/ueHi0NCyhjjaRpXolNbDTpFJd9aIBfAtey20g3UdFuAa8Bm1ygooyg4
nwfKrehMiBtn8YDTOTKD6BS4QIOhGHkku+8luEfw+Y40onFw4kytg7eOMNWsohKNGs8t3VRNjmQp
Pi+oPNEchEW1kLBMFi0F4cXje6H6mbwy2ThLp+sjUsCT9wUe06wGoX0R+pCaoQw+T9DBNT4s0I8Y
JbJvM/OwDFdSh6eue0xZKk1fwn0DAGogzRXhQNvzu78FpKybfbPZ/KpJNBHeHIoIypH2HeMRLouC
Cus0b6jPUKl/4uTMwUNV57Vuoy9+EYaSc0balZwvSCTRDhd1Zik08NoZYoVRhSKutBWl940cGJK8
CZTDlhDwhigiZXWlSMyAriPh7y7dp0G42akrZSRhgwKhR6cVmKck6zJIM4FKea3QtOQFchqyrnbE
gVknhj2nyrAecByCT/p2/6wUsNdmZa8T/PfbGZUNoryEyzMvVo/f8VKn0s5A/kTLsXo/lkP9vWOI
+LUp+w2bYL+PtM4T+ObHVn8bubhFLs19llPjK3kKKwT+1WeE9DVZoxlZvoUT51fLMKM8JxcBoMlZ
eI1mNfqWexq2gYKw/WrksjvMBuVfrnqOqjummJ2TbXo0wYObgXRrCaOWKSRTLlIaWgHNPOSSBiCX
jDb3Q1f3j/pVBvWXTXYXRfX+N4n728q6xoJ0lwfcgHvbw1nH0KhKZMlyHbONQPd6pH6WF1qI2VLg
LWmPBSAlW7e7RlDffjvdPAdBLp0w5+oht6FFMCuQDHuhAqXWWccuWiEOLeaZf153rkIrUcbTf6w/
kklKlgQmK9DRBX4+Xf1lXrrb28Wuc8zo13O1d5AUzMvvuVqPlqMU9mrNytJIodkvmdnTp37ebRDR
ty/NzntmS/Ws3vlxDCWiEsjKhSDiusbGD1gkhjuhK5+3ONLMhf3FCrnmkwphXRc+/B+Vs5DTc+pS
AoWUb3DSzaofYiIVx7FOXyGquoxaWmczHmnKzOEIkRgkVnG0ogTVmUwoG4OmQ6kfjLTSol98b0nm
7o5WTbIjzLqfhNDtp+ZAx92qg/ORJISMrynMv7Q6vaCJ9Qr76XdVByLVUx8d8O3rOjPmOCvSoIVd
QR4tsNUTe3ADRrZZ4IhHPWZwfd9o/7KzyDJvNmoslhrTVuQXhmN3pWSUuvY+sR7SxX1qpl5jvkmM
iTr2EDMvYrKyeZC46k0Tx8/l8UqvH4NSQkOl6F+1FqJBqBD4LSdWM0p+EyfzJnRK6NkUJhX5uBoY
qrQMDUBHmTTsbkKrK11rdv52h9VRvQ7vYlqoMtWj4UqIf+HyfAnkv17aVRvJIby5f1GkzBa6/KhW
SEhEXM4MrJOHSMkVtwIhL5dXYdgQBn4e9JRN86jbL5aQb/qC10TYUxuQLRMIIeYwOSb+/MoEULeL
/pV9aB3VVY/WLtfPPCxTMKL6ONgaXHfPjuxyQmTbPUTo0ZR6JQnW/ldMqpCG2TuJg+H6Zc7H9cKy
EJGmqiB7L/6usnDkg5wdpkT1qzIGtM7i+zEROXgRgV/ZSRjT/VPq8ZVknqK6S4S3eXwS/NO7MpNj
b/pYwpL68upCRvR9WobzD7VapamTexsXorufCA5XwC52s/gM2LBweVqDaAymyY4tL6/fxc0CHusN
yhRGdApyPOCSk64i27BOnMTQHTQXkLAY/WwEAJC7vjpLUWB3rSDItuk4VmpUlVZJ1+iu6po6XqAY
4iD1fCS2En9xowz+x7tPPMiIH2joxiYSf4MkVKbveHw/DpZRzhvKD5QyWtCxAK/T5gjeyQRQrbfz
7/nsb1W1j5lhmQdSfSp23o6wDf1C8GwvzO3UVb8LZnm1z0Uw5VS74YncGn5qYUSUHkBDAuTqlJuC
8S67HSiK/ZwYjjZJWcklvWzuTS+HEVGu1wwY4k0FaB3QOAuieqkmWQKO4BjwqEnvy8eVqF6NIXSM
FRnWla6/W7ZMhcrtRJM3e2n//1nXOuAi1PNInkEjB33CqY4z5JJRvQ3Ntxa0aK5/ddzWimZvoApk
UKqYhwc+W12izBp2OZgwS7yI9qVZdpoNhOzU2502cQ0Kht93niS8v7zg1PIMhEcDyIi4xPTctk+I
TQCHrSjuia8au65W/1mtlb3NmkX+8v5CHjEcWmW+kPy62gkoms4Fz4LMo540Xb5klseicIo/NdXh
jQW4f9+4SdB0fMH8a8gRaWRIh5YQ8J96V73xr1nvnwMvcjeGIiB3unoeTi2Uez2c82iD8eXF/IyX
qJCCIf/lo8SaphPcqs0k7DNOAeugffL08XgVKJGPTYPa//fV24YjuvECAOfGcISfCz5vjaRSkEDg
AMCh+jtK4gH6hw7cEhlH16GllMGKs8yy7zGNeL42b62v2Jc3M4NSqxxihcYvOalhS4JfPpExVi58
0qxu8x2zDsuujBhvLT/byGqtB/ImO0jl8rBqZT2L2o/9ankRQuJ90PbefMlB5FReZVbHbx+BDd/t
rOHmAnhIOlc+nHlPMZ4Y2lujUeZITRsfpSJp8L+TXtc3JJLdwwaUxrhV3xrtKK/zn+MFKfUBmabZ
r/mHlQLNZU1O2stDQyPdQvZZFY4gijmkxityoz0oUTW2LPAw0ldGRsbMoVFBnMjZNwYwVT4rEveX
4pAqwvD+0eE1b2KO/b0J57KaABTugjvYpp3JD+y5yo3Hh3hTHnjo1fmVkUbtBmH24t9DxP4PIqNz
h5YDzw0YpvVM5HBlKc13mA1vwtGzlzamlutRCToIWVQBvybEcFJQKcEiRhrv/PjyvKgdzvQpnnTd
DUDnuCdUpHwuchvPSszhmh7WF+UOiUY0up0Wy453pfhblWzUDYVAaIY4kvyLO/HB5vQZlinKwhLX
TofmGtKnyYfTq30tUAnLuJdO4w92D54wmk/Qkz4ZrJmwMktmYqXuHshC+p56YmjC3/g95yjBsgh2
4pXl/OrSPlnIpoxnVxXqcQ55Wqc1q82BQ+FGv7vD2mBmPosPBP77u1Ohe0Qj/0m0F8sGisbGPZD0
i7WzETofrNpviAZ0w3OaUvrmTGtXHR7HfsFyaWQHxnzfrjBabxDjnwVM96lKcntpuKY3L9AcJ0ja
AmfyPOUdZ12fFqWteXYLAqx6eSxRMjz+FB2t4Qod2h51wUQqJyOFj0R65n+ZCQGv2RcBwPY1It82
YbvWCjqf+C3VfGls98+dXIsJVUEb9IaO3ygMPHX0WDmyP9C7kZhyh/Z2arVZBmiP0iYitD9uLHSz
++gTRFu+XXlIuxX39f9FNDh/K/jCWKKVr+xtxkBNpuCMRMY6O6MFnGdXf+/GBxbe4BrpVWP9hvXg
HaMGnEAyThPoz394C7N7FcKfCGc44QttTqxaWhvMjc+mq8G5jXAl+zfiuEnRSG9U+is3IyUenKM2
aK54piMF94B4j1c7ag9egj+6e9mPG3ORPU5hYI6Us47A5F6D78J5PXsqsPPkzr5kMKI2x8vMM7Lu
IG+nYxs1ZdrB/c0yIeyw1AsdbRQ4IydHjoIkWWI3A1zqhr/1WVq/mXsAG0SwznKEcJLW8DkMqMZf
LgQb8Y8KD9vxRp9phhYVjLwRVr7lAAuhZjcnoGvzAjxFXHxzQRzD6V0HIBwL7dlBrMdFg9XWaOJM
rwbjvqpF0ixgcncCTA5vDMxg8+IakAC1XGGt6XXlm/yswQUVnnzQluLY2TktYT2lm/m774u5+Vfp
DxutVa5dpg2M3HMmDvPWnSXpu8IDndBjcQ8keSaDrUfHUlFy9T3I/07KVXiKdMXlP8DNjL4739XF
vI3TtFL4kQs4uiMsKVe0PRyiRoZMq85j9woKTQSLWItFiVpFvj+3T7d/3oILzW8kGGP+7n9sMuN+
ejXRWe5tImUU5IW+CfDKbDa1ToBy9AmzIlzx/i7sL9Sq1AJILaJGSxJElBSYphCOcVplKGLYfuvb
eHJ2FoQKTkbPfVK522yFrovJWyxOZZYUW9X3x157X9B8wyeyHtmlh4J2Fva6pazUQ4ytz3yCOMEN
76xlu9Jebtf6g+Dm3pH8+xGMDURZxSHWgg/9Bw3TS4pE+H+UZYaVMXzWPuLInajaBHu5jCOG66Ft
2yMKntu2OsqbNOk1AVxiQrq0CwJlcC4LXAUzR9SJ8+79dMfDGhVqV0rzNNeVSLx0+31R4hrM7Ffb
35YKPeCg0yIpYIYb7Uzho7MAPO5vJocrUUv5OXirLoWu+1krNMOtBWGSXZs47GuFxJ/NFZlcQNYG
pdg7La6EpcXyS5HwSqyaR6fmn9anf18px6J1O5JCWKzomANMDMFv5dmkRO/w9g1j1zBvKbf9opJk
tb0o0JCy1PJSY2MJDbNI84N59BfQLB45Uh17gFnv64WpLQQ+A8ftS3J0ACGfuYmFoUKsWDZ9hvdu
ylDLxtmXV7DF4oa0Zdkglk/nqoAuWQHGgC/nczA64rzR45MlLda36wG2/8RxaNIFaUr2fuaER+Q4
kznH8sI02o5yFX0Di7li2tyXTnti5r1oP8BgsEgEsHsIW0C4Wz8Yy2ju1ABS5cVY7u05Do64g3J2
vUPZqCOQCeZ5KukkEylsyKqQE++jTVg9l93LNb0omzmMbMy7RCfu1i00u94ql5y4iFjeiTqjHR1w
lOerftxB4oHJz1PGFCOol6nR8k8gizoaSpz9U7hHVcewMJsdhS5Wgj1I6CVnv4sEc9GWH2NtQxCs
MUHKBazDxZo24JVIPZHVfA42qdcZBBI/BRM/pD9ulmSaujT6Mz1r2nqLV9YuJrQMAYvbe3B6/GF8
suLJ51uJkBMPpTTtAQHe1R9jePRZCclhcn60E26onG70WCgIGCZZARbp8hBBwnU9HnZQLkNYH4m0
9u/PTDPJeX8y9BF6vyZ6uteCgfmDUT5+9yR4tpr4k6aMr/rlid1hYYNhFoEXP239LJs0O6aO7unR
4ARudhOu6mhZ16EVd01+xr19el3X9neGW3Mk+dqHoR/tv5Nn1eu6zhtsY3DlIVA/pk5I4v+rvZq6
BqNLnqaT/3AU1pie2z8Zhy9coQiDB5rhv3zsKQHnTNHFPopKpSM8AOGh54Ut7RHMpZVyf+hcbNNp
S0TfvaxuzuWmqUZLKoBPwRUlUfHTgW7l9uJznt2tfzhBgBWZw49elpHJ2Siao9b6C7Eb1SMBMPBk
a9dxxPE7o61AUHpX2IuY5DYlW9NNsNdeKpFgOkkcODdwJDkY6xMrDY5hCxk2egb8ye7UsGAvBI2s
zyK7ZxGGlt6TOLBwuo9fNJF+GIPXH3JWc7Pthc/+KU8410audpIfZlztu2rsr/H+0RuoHqDBu/sO
V/iYzMmWfLTstWF/su8aEoTL5FtuKHAtAvNBgvM8Hvg5dLYOU5cFhYW+VGAN11arWeEo9jwfjNH2
1OihPAg4CvGAYGfdyDZec1EYemFALyMo/ZUR5A10sCuYbdJ74PyCZPrA4dCwrS5RXITKIddavwmW
MS/TigBkK0ncQdbQEoN8ExGlHsmmg+Pp6Lof3TmZ+Fq6la5RTGBkQ8LBPn33VIlmoahGD079IIvQ
YUItviN6kVCOLDw6st4bdBPBJK3T22BvgknxBkxGfK0DViYb4KcDpsacrrqqLDccYkBFx6Ug35WS
WOlEME1nPuoCS+LAaCsE3iVoZJCsuyap7T8epCQ5c1hiLxOhCgaisK9RuiHLRC1KKu0A9JDMYOab
gHbdGTJGYFWjbQ0fTJNyoFfpzGcLpPz20UgviFTnluTTIEZBEENviIVvh1HMZGs5yP3zidbJqaue
SfayI+0EbX1Dll57FsPdZkd4SZdqIHXKtNeXFItpHoX8cFVZX36hXGD88E3WMTUBUewjUpLmRdAF
efun3qBiR/q0hMuucOVewIlSIu41hXqugcfjD6R4N2hzBqzD5oDomsb18FsZIur5G/EBzqGrCJCj
oapqK6l8HTVyE7HZ3ya3fM6bBM9o72TD7b7csyFCnTdvMvi8z7tq7g1JVa4FjkmwZKIG2Zxwl96V
EYjlN+hubQdghjdHCn6RUEpLXla+rpnPFjqNrSEiPc3AZHns72ZLBuMrRrh/2T1Kt2p5kiFT29uj
6qUx0hz3e0L0CRJgoYszTH3dyGZRWaieZ20/keUJnnQBVdkr/zr8KTEBe0iVmtCNtniM8EJ44Szc
AeXQSkiiSIRqp/KBpQmlQbZVJmFI2vVir26fg1cHqwpxJVKi5DjZyPACaYqVB5QOd3fGgp6rdvH+
g+Ap/KCLSSBTBRVY7GvpShoZGr1GDF44hQBzbJ/70C8wLd46Faucn3hBj+QaINxiiRwBJoNfWDx8
FThS6LBT0bM/QYmxhsrS3yIE9wKdsVP2MoFqF2rzbZobEldheXVrOss30cHwyAUl1g2nBTwfoTId
9ifRJo7An2j0Z88JU4LngMx0zyIUAn8HHxKYoLFjPgfQdLx8/KwTW+NBOPud0v4ys3WQHx6TF6xP
YtowZovqC8RLfTzdU8Oi5zHC8RWMGnYpvYLwmvDYk+IHu1yAUtO6S2LkWzHySzV6O55GUHiqlNEu
xNudo3ziCUS8k40IL34Mag+Orv3qFXxeJS82IE1MTvn9CyFFgRNkLpZJfN18+/zPjmZBCju5PsGB
AU9+YMR/w6+1NCkSispIITDGkAkkySGpWzllnzJC2bsrmI3uVwc2RTfMs3w32hGTB6rd73RyG4Rc
iOi6ViX4Kp/rhkCN8HHhZNdjHKcH+keIUJYPCSgJDS0+F6B5YF3pNybi8lAG80ZNHzE+00mAwQlT
KrNmzfZA1RI7XWrDWPXerIIO2CIp4G0JQi27xhFgBPOL+9omsdTNoGNXClmIBejvcwG9iQ9RXPac
WNjI6BkNazgmWcNhdw/GxKqpOHzPnXM3KqnreZ5qIvGRR+oqxwpYqauQTV+qDqVB8D+nMPj2TTq/
UubqqFT7HbB8uxelXDSvFUbqW64WmtcGcEhvyLm2q2wR62+VsPSRsfbTtT19ErhgMDmLLKksqO2P
SJZQC4QLz4j7AXNjvohHIJsqAvTZCiwFsxEaMT70rtMS3+vmwjnycSsctoeghLjMBanLUVSQX3dY
MimGIfSem2mzfijWS+LZmP7XxXnyq/UmRMFLeK/tTPppSHDlz0BOr3lxDJvbxk+SN8wzwhCqLqJ5
zUFGVmJtqxLl6csZIRofDg7o3soyll9diAYmyk8v0by1On3RDX/9xVoWH62xA6nradQFo7jX2aTH
FG1qZFjbX4Qs///V6HerIiVcyCIfEEID5L4qPEKfDar92/fSnj9XTAt10tH18bIVLEBo9pSC7FJh
ZLhqtD2JqFTMQcSlwQnuLx2sK3QYUhaiEtFwZSKhgGNYeYcouI6VFFm87g1M/yvkZsANmPxPzNBM
0tMv5bglQVwp2hDsMTxC4gVUZ7N9D+OVJLYi7mxDvXshth1hFJ9jYpw7EJa3boKGqblIysZUDj2i
Q2Du11kMxkxmqdrhRhqrNwzW9u/u3oJcsaQj36n4bDACr3es87C0y7Kt3uzDbIm4uUezsz8rQKSi
kDOQsqiRPikC9xccLMMjK7k7jCeuwK9rhkueH4dFR4/ONCAtN9nlpxxLCuMPhhR2dWL7ktl5RduO
rC1AZF8+zvdkjg2x/W27ELYlSA0/FgP4/nMK3Cn+M5fVJra1vK+sxcVOqNEulB08IKBIUjSK2UcI
/+Wp4dXCazYZio/BLkNF+NtgHv6U+YvigZ28VTXXKThA419+TB7IgF1pH7/PUnzpHIKMInC0KkJ5
u11FUF9pnsIAwjDr/Y6Daf8y9l8a9m/xaij61A1V5fl3RzXGuL9l76dzIkVwtmYFFnpec36FZena
PeWpom1CS6hmHtQyXnp7jDAcxCbTz8v9Tb/sf3bWMVlFtAVm97ji7tWoSai3vnOmjwcIv/a30MXl
dEJDHJl2/QLnjT/8NHjEfjwgSLgVW0O1hLDgBst1jct2JThWK/OdcJp3xD2cwkL5ZQqeW06g7izq
PLSB4IZI6w/pXRI4cZirgw/GsJxiKSyJzKSth16JexP8Hysca59qwkw+r1pTwTjzwyWwXmiceLZm
KwoKMVnAKoUICRBa0/I3suy6MAvgXVB7jwT9zXo9ybGmgOiBrwdf/XrMR7NHOuX5uG8BEXGOxdpp
3Zax5tZ0nsYcracWlctH1KOP6O+B+GUzxmod98KqlJzCrW+bZoG3fapTGrX9nLpV3xhCGeu1gySs
lLx86bZx74FiK6ME9aAg4Khqn6uQf1dLwMy98MlxEmFMQdJzcpnfXc72vRTHhFsIGO5nuyiGl3q3
40rPck8oPfppW15QPtci2C39TDh938xrNmzH+5RYWwFmgSbT8SFoTl/rfce7bP7Hp5Ql8tnTxXRK
toCLgtLN3aIU8mxXJ7WWmhM+OUDV1Rs+2i0regN06pGurZ8VBnW4fKNjquGJvqUqzRmwaZq9ze0O
C5ZnVqqEjQIjpYiqlVnL7nlzH0dyOh7BoiRvDhxdw6RFiztYbH81+pM65x8fBAGB5r0IUrtz+xBj
pJReF0gUXSMKcVCPbFE+nBwopVRb3aXHJ+I+Wk+EJqTrV+bZ5mFgdcv57cj6JVygaZg/L54MMP5G
1A02LL/CUq3YZ9ZF+i1HufdvN5lofU+XUtENPvG7GDbcCLHa5ccyeJv1Wqe+eAwRA6SMmRrzrMU2
cM5PcNsZHSSJ5lAl3WIuQkr8JCXk2zPidvkeO2CL8kx0g/cmQpfTMkQ9vdr6FIECW9/rWZlr8+qx
ldFd5AYVCPkSk3xIT6xUGGLH0dAUSGMS3SJYHSe74b2FaBYEijNZNuUDFcZkHms8oslWwbbRI1uQ
g5OfVhWySEOcKGGJp7sDz1lS8YKdxtSmW9xB3bFd4e+3VzmlLNfnCqs36eWlESwlL8Cx/Lg3hwDg
vKiovNFEOK3QOoBTed8uZksqZD5oHbqvNh4Czyh444UJXDzeWTVAiL5OUbUVcUUeeeo6HZCx7vYF
Ru3dedSAdDolOuB7z5CeRaishIZtEvoGeO82lbuiYKWkaYSkPK+KfLARmnC3RRt+JKNxTaW1fBlN
/4j2D8NXCfi6PzrZEk0vJAwk3tZiSZVfuUHOzjo9wTeqbXnDFIyhpQjOx4xeNqT82lHbiRuhZKGk
+zeoUDOobBRjONRZwl9rsIlgMgjfu2nzWhirF/l4bSE/CbHkSBc6CQR8rNhDfB549aNvr1+mgppD
MkYhgFIRQQC4G/a/fqRcsZYADAKIhqIpUo+lBSvQpsXe2ptpUz9bpQmCwUhrK2xH/ebu8mDyMvH+
Dx7YCeHAsT95hVnHICkOrf8d0CZEnEsKNo1Pgpg3uJl1L1ZFmfoXsGT6I39bdaKrdatSkP1RRbbC
MD/ds/ppLRw++3cwsTyZ66NaQE/5kDCPAFZCIXKY4E1WiXjh9Hadqh5Sy8Q4eGLgus4ZFpoxr7Hp
OpAMiivFNmsVQGs2VLEz0KVjvrAdqCrdt1JwiRIy8rZ6jvTb4I4wsqhKix8DZAnY9+n0jFZe0B0r
Gh35YNtwCuU7zVjOdO+TPGncwiehjsLTF60XhLDC0rYmM3uCuP6uuH/oc4p3go0RSl7Vpi2ZVoAq
6+bgPWnhGnWB3tfZ3dKe4/vlJ58C3AaDqitUj3tpJoAsgJ+1LKEI/pF7WqKGN6Hy/GmkvshBeR9I
PrMEsexCOgxyThfFyf0PtJ+hJO7QQSGg5DuZwL9BrK/ApYQiHlsp+KQumTuodFfVt3xi+vBPc/OJ
4mdd+139GwvXg/IOFQpVkYaNRaZC+0WF1v7gX9HJ6aVTDtZz+Hsju3bUMOFCHiNzYh8g6pWbzS5X
Stui+MkwLLB68h8q7hy40Hajisd6l3OI7cSPXgFpkugdG4o6ZmGLdvrX9SLbYNPY8f29zfreC9WW
FsybIhv9g6ODFGu3FpPkUDHxzRr4je+f2V13+48FNgJ6q0AYQIyrYnl83EgU8Mx/r9neXxsMtU8T
mgyJmIRcWKvdCUFFcWmFzVgrk690i/HR+SAfNTAP+D9Qb97QlgxJ650SYvf5FKaxXYrzW/dJ0o4s
Z9Y8qBfm5KUjMripZ3favHENE/E5OcJELHSZntA8OwfVYsIBl9DtKeLEP8AS/DOLI627cI3e+c5f
LHEyjRp493E48kd4U23ZHIRYE7ysSwdDwtnvJwoQ2VWVkHGBOMfsMQ9TN7cbXjGfvp8+0Kx8L2Mh
yDVGOaQeKmVVRImVKQpSDUVC/D0A2Y2qaZIAmTWorcso9k8o+Z7Uj8pq2U0A/HLtDFw7tGesBYpZ
37lK+KEFZf0ij3KFGxApdosGOv3/waZB3GYQOS+bjyUirESFXTD/Kh/xkdS6Z8ivXLGqRU9u6BFk
yYfceQPbwvrqdUp51PdOZNXRfwF7DfFG9Y+5/7atcLQ+w3pJJEao9K6FJsXqSr59Otx76WgmM0vH
ATQ9wQG9LVwAJc3cWEgW4emLuVZW3kyuJmU/E1pFwFDeBl/MUy9zaFRbMw2yJ4u3QP+cViLb5uJM
aF1yNNRPKij9nOTlT7DCVKU/LN4B0cfsqalgKPFPLWdyTbMAFl6nA8SyriyTu3UxUfePLLFawQXU
MM4RTU4DsLVLhNlR/Qcqz6WdCWdJVIGH7nGvygxrG/DgDqZMBoF0FbxSqeaaatDCuMV1k4cngWdP
34m3EElM3bHMgJRCdroIHfWN+jyHWoy3PDh4re9tEeYLRbMHIK0WIJ3Tx8lJHNRXpzYnJGQMcLZt
sZgT/Vgg9cD2IwPTWye1gt03b1AJ5PI4qwuvDiOj3PShUNEnNzKjS7wBMzrXc5pvf/yk//fkWo5g
71uELi89H9PWaGsNUaKunGB+7wqKUZPfKuO8yonkLAskG0AF1f6gWTqNiRaxsxVmxJoJKG3nGe7R
WC9k5gs3ZJe9g3NMCmTqJXf2awtloEW4g0xzn35TObO9Z43WO2vYTbs5UXH3lC7/Tx1xWL0NvCAQ
b6fAsTJizjP6RzeSISbDOyt4MWXKupsNLyE60g7MKgO0+zIfsLEARx2Fq9+oimuWc7Th49fsCD2A
rwtiwa+Ufs4+8HBD2Zqv8Mw0GWu6f3yBIB5XDcQ6kkvvG6l3M7EpHxb3MCeoMI4IWwaF7vpcFOpR
EyP2M3VsbxDGDTP4iSd2foZO8gDvVtNq8EUduuUujNFMd3Vds9FGNBFuj6aBgPnnS6xXBJ9+IDL2
LR3UXS9Go3rt+Q31pS4N6xDwuWrEuqojYG/mWuej9Yu+9xxx5d5SSSNmRISGmsqQIDmyhzMQPZSm
Jm+dOj0PSw2ogU83nyL5hQ3Rm7a0kIZLyq8ByBDrmuw7Q2Eo0PMYK+fFlTWyvBXYCIvoVCw+z11L
FiHg2OUsMITh0/I/AAkOnaEXSdoSReG0dwLm2znCBJfcx3XvHHwCt77yC1Zy8iHdxJhdXRFKE0V5
J7p76OkCe033JtqS29AvcPExupP0Uksj/jl6VyF0E0NXZTpxAUh6gpmTTckZ3olwbtcs6pSbJAK9
mYieScRrZ6fQQ2fWVSD5XeopI4NO61wln4qjKWDxAuI/T/hg2Qkh0BMKPWLp2yWU80Z25NQCoIsi
vvjlFGnXQlzxQ5snre6QKfQOIHlZctFL/E7GBxzY7HIVAZoPeAnyh8q3Xxu72ImBdXnqGmbILKrY
kZLfUmB7vMkdaPrXws7Flx35MjRAd3NQlm5pV4DDoZ6mgd12KjhxjFylxjLS9MRidgcbpZSqjOjU
NlOvrA2LBqOplIAnRK2AnZh6ItJFyRTdtOCAQ84vBieJwCXe8UqGu7GbCQoy0k4In5sPfpQ9EjWv
LhJI19Do8WVF2AXvrfsm+4Dx+C12+DgFAicX1BwPeMdaZLqFW64mH1nNghaS9wmGlm0poH8SfMln
z8anNFNmDYWgtgq4oNIs4jU0bDN2hphVTpmtOSwtN4wlgV7nXJ/ZhhbrjxMFJQdbDYqQ/RWuxty4
FffNtYK1IRCUva+uvK0IHa/S+tdJKl1xEy53KMmmWjqbAa5inF72aiVP10zY+TLZsUl56lMZBCQG
vtU5jdhsCql94TV0HsRqeQuODzyya+GmzCJ+QMg7Pjy58whBnNXvBderY3uxNogQ17T5FXJ3jd9W
ieyPjCXa4pizxZlGf7+gUWpNFvyj7dYyldEN+9m1viIwQrRIxWrSIh/MCtZeRvZdkqefunwAhZ+F
c+P6G4ywrOsj6BTB0bzzKJNuzUZ1dpQmJvOTBQb2DHy69pp0OY2YEySxmuFMY6jAGnv+x6M/4gho
84XxmuozWhEKRJtCXHD2YIgq/i9GLnc9ThZ+Ym07Q5T6C4QOEspRX+65F9CaVuntwUx6CF0NdZYX
nDhUMIuAz/+X9JSmn5ffKChJ/0EDMpG7CbZJyJrMCsy/oNCBmmKhHfpfKyoadVLyu+PUmsZcIFqE
eyRItxLaLmlyGeOsKPdulbtQ4vCkUAv1HHSTITCbkvGnglyrahroE+BW5Ick9AyLxpOTTrfM4qjY
dLA1SH8RKp7wFdzMEPAHyih75Q1cw9y4Hs9KVzDWHX/GcN8fQmDwyd8AKkMhO2GK8jY6IJH4gTYZ
pZfQH4zHZxR/kQsRtlMO5bdkdJ3W2zPgjDhyxqPbOdt2goLudqUD2KgN6YgDevynbTJiNbxEy0fu
RtxJXZLrhg2tzJ/cLz5bhQtz2eMsrWmgctMDfCXdC0rNiARHZYy+XmBHXFKcGW3R3DatGZNt7OZE
HacVXlKmuZ/l/xkbM9YhYzA0xdQxnKncDDVyOJlP8eF9sjKZoC4k9t48tcvdEBhmdf1g6MftrU1M
T+wkYSP0pVw1m4HR+Kb3+70mqT6YgXq9wjNySENDlXIHbFqUR22vecTzioO38pYvtofd8PS8dLiB
kdNc5QEhBnH4mCvQfThCGLJKG+QbqPwaIZkIpo7nslGXLZisoUFWQvVsYKjZl9gvix3aw1cnKWTp
T8bUd5kPmF3FbndccUiNp+ZqQA29g8+a0b88XhzTeU+IrTLrKc+HhYEyD/d8M6OemvqRHCJJ2Mul
BFp3UH6As/1Pe7d5lxjugp7q/baQ8rUbwhqaIdPUXORpvVry5Bp8fXXEXwKyPJQy+GV+QEcjHKO8
dzO29XW5u1ZJxY7042MOVIK6jetniUD3xdofNSqIAOnHYYrhDJCUMgaUOfP5TySRCFPqLrDkf3yr
Qblaor9ymtTBoSTWzV+CZXoC/0JBtRkpfTp38nUikZoHhQTvsc00VX7Ey4l4PvJVImu+iwfbQSDp
g9xgEXlMggQ6/8dXzZAnKbSJCrRSj9gt1BKKVTZGINYamXyTKFzByJUgrjBAPMMiekteRWzJ1mhr
6ZnxD+nkyN4AkCWe2D6VzMcjlz3JbAIBy494lxqwm4xUFKYGIUV/ZJX/WvKclbv5KJqgfawoLols
bb4gXoQMJonMe0JuAgbE9D0cbAXZwuWhJmp4Y/dk/IPUtmDYMxb7rsTpC5BCBVLBWiFzhozDtV0J
TIDxQirc0sVU+q/xy6l0kFRWP7As4u4GSTo8vYZT1DLtCBW030mR3jO7QThjEpUJ6z8Xf3cR9Rwb
P1dQyUxwUczRj+JCGYUOv5Iggrz3Dc0Xkc4fnLHc4DTB4v0+16Yyv8Gw4iyZEK8VAu+Wm6I2OZ9H
7Dxu4nee8/URgEhurlJCW346AAwAOTonlDwftomh2DLN6padKRpJAH+XXveRkDVJfeqmEjBav+OW
cmQ8DaOAjT+VArjvD6xd4/neRvQGZTmk4y3gZgrv9gpEHA42H8UEFbw24s3YKWAg61R5BlHf4L04
NUhqStGt1f4ndQ6DXCbHCWELgMZPrYyxPeE5lXfDAjGittwEdw+Ro5Zoa9DHD6mIK07thc6W7qZg
IdL1BkFM0214Vrlo7ujLQfAdXt+bgaN3IOk0k3IDDZnKLDINyd5R+0wESxBiIeNkoUE9BBgHFwxd
AeZi7KMfc8H8aeXZchm/RbbyQ1bqmgQ3IbqsprULc81og48MY/ZlEd8HC0DSyZg5hF0Paw6DhS7w
Ec5W+Njg5JENrJbIcR8/nFgHlWsS9VQCFUGLtNBTaX8M68hzssj3WmLfatl84xm3u1CJutZB7f26
5K3N6xGWO5oF7FBtOVxE2tmTBAaeXeueLLdQjMvwfaROQQjYwRzLBms+c/gYefD1dSUp2szn8vZV
dssTZlUSJ5P6fEp4kg0vkqhN/O4Y8eMq4v9se5BV4NChLH6jSVzeM3BLtrZLEGF862x1JktBB3vG
1DU4kDRMeXOd3oearO69Jj9vvw+3tkxkuzf2xbmkbi0EXvaXw9fJFaDO9HE1B3kFHQZoyymCMu5y
9XuraXeJq+nbaspAoWJX55fhoo2akGpJ6tS7lBgY/p+23dDtUfrFIbDeA7/KZ3sQfkIDsLwwXus0
LopoSwiwpFBzPP8VJg6u0yeponDZFql2wlJ/RyfWV5GsPtngtvYiRUEEgNJ7LFyGCU3+u64dG5Dr
hx9EynA+ESt/ZvVhsPmeYBsUJhpNELqOh2qv9f2A/4f3KeecqnQOkTp69xepnGrkWeXKOLeA3wqh
C00Yl1hv7f1mm4pGF1jAWUJz/OElwQeBmWOruxtwd0IlmARmsKvhLQEW0fdtaQ6IhNNHml4hPfpK
rZhqk9klVMPjF1P7PGn0V05q1dPEv4O1u4d43A0x5dxLTC/MXCj95eHKKnK+mpmbo50pXTwY4TDE
g2lL/CG/GFfYi6rNRuCjNODXa4FdITVMnJd8f9Ot8FnPx43Xr85jQt/uUrmHWTcrJNedV+x2hmts
9utYA3RDK67okt8Qr1pP7tjjQQg8LgfJlb+GmIasVaogK4lr/JI7igpppsi/2uY29qQlo7PdYptL
viuQNHBx7TmGFv6K5VDIu6K5qKKOCdqiKaBpTw6MPZLTxJgrX86aqp+uTUWEN2coX65edYuC+EiI
0nvLLGM6wOr7V3+3/pgsNCSI2memmYbOCibJ39/uv6V8PdskuIfepRCLUmDmioL3EZuun5tEvuxw
U4mOcQGqs79FAuPO3N/HlfL3qaFPRtTnQ+DM1wthUlTlfE1H34QfroXVNVdlR4ze00D3BIbx1xsW
GGoJyVLgSFENon7bPk+2eFR7M7BS4SYd8ZOD7bjbrQaBeGBqhcdwcX73yyA1hCnDCYpDQ7ZAeLEu
p0I8AczQa5D7mg0KjynV+1lGQoP+F1Ozz53tbbdqtKtRFkcVr47kOLwI5qHe6ki4ATLRx72TMLlr
OmYBMW2SQhbPdexcnG1oHZXt/9ZMhPiPTks8OZOuduKjE409E76rL1XdYiJkhQbluGN6UNDQunYh
eS5RvN2F+onKgHSBh+3+DzGzcoYG00qHW2CKKDs1yfx+KC67oM3qDuhr87XGiVBcfPAHy9EkxAq2
Xs3gl2iSHqv1oPAXznRSlHvKZ3lIa0w5PT51HN+bVQ9FNC3yWw3Mo7BB1Sx5UnFsfYL9gI68zj+v
KGsGm7KU0jEXkA5PKaURXnEn5ud6fCrVdQ22GJh+cw9C3qGhJaPn1vi9XDTF5KM/YzaodguX5shw
oG6HZpn1B2VGTvCquv+5U7AM/fAZjt9bR9vtDIMcVdlkXT8iNnr3SauDoPe+N1KMcHK1bspaq3v+
Kgd4ueq9ZbDYu7A3aKPxV01XkIkZOfkEJdsy3Tm1qsDQy+jct9pZSOJYrttg10OkkrmBeQRsX7f9
cSUpHG+H3rhd14u5Mh9Wv2rpBJ2iXq2GZFkQul6VWAh90RkvwmNF0TyKn5LSRIVLZriEr7gBwdG0
vd65cL/HGJ/SA7r71azwVQ5LqUgEoTAStaiA9PQGtnO35dpY2HtG70tVJt6FQtKHE3O5oGgS7Fix
Qop9xB8Nyl2W3opYIlmEoTbxK16WoI0r04H6Ab2xhZM9fJ+rBxX192KbFNmojxBwVJlk9t9Vsurw
oOJxR7EWZ2fL+i/bK86+9xSyqwmuQ1eiLWiTdLKEf0IC/crRQAbA07s5L5AjVIkx6rxjlvtTj6Th
dJGLNbT3kl+Pj4qbqBPMCqeIBSt4R0PzCwTwXE4lCB80T6//HZXqZkpKN8r0fH6sqeV4mD6r9RYJ
KMClzj7Fk9Bs4XgK55UjNCzR2Yos3ZoeYyVT2Frxk8r0wetaAZXknJcx7df8rrp8SVabmF4UQBdy
o5/lAc3STZqDnieE7oBiNyVcI3gmsmPxxvB1kQBXO+/9NcRai5jzMPKT23lx9CfL6dr8YR0BiN4m
Xom+zSfuuYfyVJRXDfxLudPKhjQF4J+RCjPHAB44BVcq4Pu4QKAwkm7Sw66QW5PBSSCZW84dTLe0
cqdffeUU8SH1cZviWh//BcObWgtaZa2IB/hhPM2OMBU1lLwGxXMl0OvRrvToEexMO2YA1eqKVDBo
iVkMlULmhZyDrVfjKQJAvyFrWpKaWi8zDugD1LVMwTG+bCdw3eapw3W/+yJqepG5Je9qSUweScVQ
8a7a0E06LJRqhQaErQeQNQ4z0ex6xnoyPvcO2ecFaFblSv4e2B+3Yw9EIkjc0oScLKc+BrZoqUoF
2w19bozRhpDq1Z39s0CAZkKDCnHCyo1z0+aptWF3PzrfvR4QG6mHNXu/wyW+Qc/eC7iQR9j5GFAN
RR+X6s144mHJ+F13IsI3M+y02H6WGjCVblTbRForlqpiWQ/e3PEwzgtwF7uYzvYCfqURlgZ9m58p
x9XrgiB2rbxWga6y5c52afWMOh8X/9+XT502oHHkLf3dMrkyRzecxH5kaGqCoEbSbtg4cPDMPEoL
0CyM6jwwudfdnUplIGSjrRfCrTG9T+oUKLnvOJASlpNfABUszAc1WMYdpxCD4F+Z2iPH2cjoef6z
FNszxl9pTYUyO/e+tHxV183oXpBJBd7Y+hvh+sDSH+mfJD7eurKE0hpGXPbkbZlsM6+CEDS5hOB5
L1f7YRTPrMXNYjuAz0jlybVKOHk4I8dJ3rWbRaTz5P9aL8Ylt111/9Z1yVBnNeUlDfCUJt9Nz7nG
iUjV9GPUHx2JAjeBvQWYM3ftMW2Z3x4TvpcTPPTgGoS5jeKuK3h9sgoVzG8Du2mIUsK98Mht1/aj
glrLNsojLSlW54oDU2PnEGxT294j329KI7ZoCc3q5DB79T+2kIg3WhzA+fjRcxmo+jP3l3CtpLj9
iWZ8tINda2WPONHtiyMAKDu+ZSedT827k4kzjS8IbSRz9T2tbkaL8imrmdjf1qS1ymyRBOJMR7KD
MBxvQfAgVeOp36HMZZlCBfoSdnj+cZ+klpJ7TPiOVRJbZ6isAi4kwtKaryKp4u9CPYDVX4L97fvJ
CVSdwvhz07uw8Ort2liRGFkIf9IjiajIyY/cjZS74MdNGwKURNV6ds6sMsvjJaOmk5T8c9pKUfQY
+Hhk/LcwYWgdcCWDW8FBHjs7GOhRCIRqtnVZ5VCUeTlN19dtMx9ITcFdfug7Pybtkql/+wcRuBr9
Wv6noYcJUD1bQdtNmx0/Pyua7wbDwEo6JiKP5E5lKPf/0I2ayWO+QgwnPQnmKYfY8ZK0nRQ/cuW7
egyY34O0AXptJSmzzmIUwPSNvfN9JqvjONU/CRWRPw696wmjM4C8b5DuIq8QzHyBM0P+RmwGCfFc
iFuDT1swxojzp3LXaFi6MkDpNVhXc4K3/YsuHcKSJgi2AGwMdCfwq3XwfCs1DWsTQ2PMqpBjEnKJ
UHx+lQ5z9xkQq5Nvv8lPQ1h90fjRyTi7JfEg71LVWXupiGzj4Y5QLvkhm8tk0Vm/SLHjUZi6qAGe
Xj1/g6Fa5tUOHh2PC3z8/jArb8THtJsZ6pjY/RIbTY19JtLsbj5CfBXc74R6gIGHz7gwSSZVlpHl
vTJP+tSQGA+XaIIrimXlcnX7+arCkzlzvglkXPxILituvsheBAJl2tHs/g/EXCxuvXo3/RDTpAuM
5KPEz/z1bb+BCMGn1lfDho247+ytzWJuruGqWWS61brH7KgLY5bCOpCQhmeGvej3dWFgLg4ciCJ/
WxV2uBbefyJTdqnUt/Yi667uhC/i5P1fU2RX4ceS1u8nhZq8lpBrUcO5RQ0aMaaDNY8J3l3Z86g/
/Fie0+eIookdyyVMbu30JjIn7RIEKm0669PNmrUYSQ9OfBtZh53+C6PVGuMOwnuqp/4doZqHmwhY
si5rVDEA6hyLF52OpI+Mfghs1f+xpDaqTNqFfxhL2gXOhRtWUdKEr4Jx4NPaH8wstfZkhJg/UAKN
h5qwFuX2tGATLjL2PB45h6pYHErXWn/S8roMThYjN4mb1uJa6tmHkr7JmcPkacBdK6snKzW2jxdM
fXH5UM6NmGdwQsasjOUsi+BBrDl6VR8gVb7LBF5Vt+C08ftanDipU1rP2BMeGvJcMFZNg2EFE2jb
OUsDLw8Vhlw8eF4SQZ9m0p4vKA6FdjZLdJlQD+c9knyoZgj5oLO7k9LxBjFfICvH2Ivjns0iFE+Z
l8KJTHhx0ZuwJFNxV/n/+cR8L6CE005tIUztofisiKrNN7UM1n795ZBKmmah3B8NHqwAgNj0e7T5
awM2xJv94nEwK/zFy6SsEPYrHy3Z5NRDMgUh2yFH37ngRSrAgfJPViAXqjZ3FBMmEiNKD0VO9Tcu
NirgZ3ubHdiE+3SrNfFSpJajxZrZnzIdN2tbOlcrXxr4PLxoxzUS4yKdUJEcZjD30V9SOUdrvn34
t8uLppLvy+Y7Uf2nT+Yc8CfZGk4rClW0GQ61BkkR+2vBeYwEb14AfZoS1eO5otuaVFSuCNPz14eX
Dqvnf7iaLQjnAMeNibNFUow3YLMQCQBiQFSh3Eo4FoAbtZjoQrNkxslaKiVM4SQWoDTZZ+hzmNwQ
CESKmqGlizP1UIoY0KW2GP7rK0WUCmmFbABtquMtacJ8OpIuWthcRtt33a7sJJ3cYFcWnGxCORvn
k9vPYkX2xeVNlMEiYcyFPRGNIeCQ7BNsTc/BgC4GwalybtY6wAeOdYjj8D+8v4AC04xQGHcVJeFX
qHbZGwcP2Hrx4Sa9pVbuST/4I4dQOS8491LLE6fJaKzZwcMihEisyZmRqmq5UDD8bDNNtDZH3oeH
43G5cHGyzXdFBogAtu9krlvs6T7G93O6vlka+boNEZH3Pee/7dZ+t2uFbf2NguLVBiXiz20QwN0a
k2m7mTvGrx1ADk1gLo8jjACJvU9pz6L1Ogtuo/bMu6A5JwyPD+cJMAKPaXIzaW5iTaUBsrW1blSl
xshIRhehhNBbaDv+ly67yqU0F141WJH3nsvMDxHog9R4IwFB7xXOvqdOj8tLnPiq5qfr3z7P372P
CKUpa0cOXqrpSVaDAKK8jhCRau75r/Dkkr+rycVi1egrRXBtGlPtZtIngYT7yc92vKRdj09gOdh0
d3Yans7jhIZlUSEWBcgfEqIwYcnPB5j0oHt0hBERh6OzfF2+zfxUMDIXDb/p4Ck5+6Ub5OW1FQIP
Kt8ZzrVhN6gpO4WYqWmRsRE9bUSeVb2ObC7L2UKuwf1jpqnT2fZS/PULCqlwjKDglQRgcKD4/e0Y
z1PY6ggdQA3DWSEr2ZidYzmN6oGwZOy0w54MX8BPZwuTfIOViofCVRRb5LWUvjRFYJNJttryuAjr
BvcwpiMNnAoa/db2rptPbtqxaE5NHu107vGt3TNC6RB4VO9Ef6MnwLo1khO2Ua2nksP6+/dDlZxc
hwbounUMDkdseVutnvPeIx/+dzPHXyAZk3aL7VkCpu44BFLU1vIGsssy666RBKmsRUS6B0c9XZ3s
50SCvJJ/AST+hoRXuVsXmDDeWjzsL4ifQDwgiv6fD3UfpLqkF75TvQSH9pLHN9nWz0TQU/4+TWFZ
dbbjInbydJ34OAEiuMC0rB77MRSLA+wqsYEOaaORER5VBIxkfNTAwH25O4A3ZdQuLB0IYjn+xkdm
jCo5m14q2RmCiL1DW+0vsW73jqbd7kaOTWnjF9T7AUIYx0CnJkY6mYudzycMOe057uP9fwVLZIPZ
kOB44xYipQZvidvAmcmOK6CIZwVO+CHab9qpHYu5BTE+baDxFzMvYFPziQqkWKKvBSouNHNG4+cg
9mIgoTWon+aoc81NnOblJ+i0Lq829+bCNcgduxbMT+suL8PCGRD/4RWNxvBLvgD6Au1IU55obDHA
BdHbg8bDaIdwmO9xxN9FWTSLJ7FTtW+5usLQLAGZHSr7Xc1U6ECBuVgXX1chim9vIxvxdrIsDns0
R/Z5ueh98zibTnMP+Do/Ierxg+1Z3qdgGff1fUAkEZZdsPtBSFZ1ELeunmE0G657JmfOkbTt09iC
eUHcNOqs+x2kE1IqkSFTSo9hljTNM5UtglZ6CHgniDVebJpBSbwCFOf53vtQT6eHydI2OwTBE9rn
51IxVb60Z813yPOkzKmZvo3/ZpPppLGYjHrRmL8eCd+JzsjNpJKERTmg9mR1e8IZzPe+PchDXYmi
bYQCKFOk03qvL8PU6eH0wkaQ+ieEOAxKGfJg3pBre/5BU8XoQ0HWGcUCZ5KSS3+JPZLP5JFtsc0I
RZDeE7zCjQmYermayyn6s/mxh4PgqedAThFHJtIFgFs+r5JrT1NwQ2cHI503mVc6mBXa2LdGK3KO
xayXVTQ6H5YoM7YrLQGAqVADZ2k/rFCEwdWw7isEIGhbZcBzAJHF8KvA2WTFwsPyNcdEmlzKr4By
V/o3cNnLNAtS5uKkr0SsjAOUhWVkFkNaJpP4EebolbmATy5jRik80dbkwMC5DHNipNVLPnGe/U5v
qnkLQkGj2SaTx8Ws8ghFTGgtbFvCETgeGD8Te/9rBXMrQmfOiswwBAwbyayUn5VYft4/ECX+xjpY
1MSRvXwX7hObIV0bf+0y46XbY2kI7Tmlq8gGhglk3I5LNlcFsKhYgrkF8O/eM3e2pdp/vEo5TPzM
Ag/H/Z5LQb190YqcBk7Vm2N6jhdM0NwklzPmmdm/VxsFWEc7mOmubbYQ1rozwC8drXgOaed2dR8y
1OKg5wI2f5OLKXMJyeMs+3QtZxhx5ZKyeNviJaTpPFrTQd/IihFNOi0wr7jolFPtgLFryaus7f9N
8upNLM61Y9C28IzEtCRSKxn6pKFkqec/VAjmASwRPR9ARkr0KF2dwn61OhlMRw8r4r4CQ1a1YNYT
Kadw94+jMq1ZPj7yN8x5cs2CIC0vth0ORMkiS1z0oKHmcbyxkh+YxZtHM5Cakkern4F0XB8kCsxH
RptAluNKDEDvyX0vz70QfMWEXcTRs2wx36ObH1Q6J2h7BPCFljKfdgFqvY7PUKZ5sslVvByYX3/n
nR8Mm6zIdhv8Oq6yl+YZdzPlvyMr0KsS+XC4bNsdzr9UZuOIc6ZSb040QyFOiWokiT/77DNUpyoA
joie1t8TKBdDnlSfS7kU0w9nNh1H5SPQLeXhObjEkw0JMuHmev8+XNwzzTthY11XrpokX4ehRegv
VBQQMyL2N0cHkj1MsaQ9Fk9i0Fbm5fqy/o8pGioP2fWN6kTSDELoe2S4EkDb1c+p63sTkc2pDdGX
OWE7MRT/M9gc/iuqpCQlxEpHIpPH1vNl66znpjG1eAEdxoifT5HL/otyOTpz7YYRpIgPOJRLs3Wf
zIsyXpbENwnTK+PPaCGTHu0wpi3iwFB1D+d1BWWXebk98iVfpvKrHl8zrVNefFj9+VhNhYAuXHjv
KLfze29W+iz3OTfucj5+Y1CimZrWF58jGLsqECYIuazt1kRQNuPbCiRgMYhUHmPSoD6IP6Rdn5tZ
q2bsECE/GjwsWduLcSoOi8II/oGZBJ+P4obylYGsJaFpNe1Rx5HufvC/Q9vaT9sZgq+SVDS60lUF
uUpXlaHwpyassQZFJ6mOJTStifBJPQHvWWLxo8RFzQ59hmLKKZXUmfQi/ZgTiIoi5arIv+TmRnaz
IoeP6Pksq6z3bQHtU/ze0SSeo0TZq49BrbPAghoZzUROJfW8qZv3xTWH+t33fO3286XtfLf6hPFh
TXBVncAhKVk7fTjTtQrOIpJ23FUdkpYfz2JCE8wY510KxnOQY4NyGFQwfBJe14jKrIaoJE22XUe1
W+lV4RLbtUZbhgstzZyF2iwgI2QygGqk08Y1JP+L+sBrPZY4HZOtvVI6V+oCCTubW1n+UvIQ0jE2
9e2XyGVNhf6taeejN79b9Z82x/TwMiMH5ksj0CdFIIqGj1CkCHJQBFD8KoCLha/AeA/wm5TBlCEX
61OoQge1GK6PWiQW+SqxaoKoOGXJt7+HJ45XLAhBuswdRzoWsHlyfUExWmyj20SajV6mbk8GQLj+
ntOHm0e/0pyD9QaqzFAs++h5MYDVGTK2lZOpj3M0LEs8Op4U8BDU3Xy0KXwUYqHhRncxciaXy2lM
g83q5HM0KPtSX6MlQ5etxVUYsICYjHgkgJzsPOClRJkbF/VEVCMx81KchjCo6rr7q07b6tk+uQSr
1C0M+Joi9NpKPjN8PMG17wEIvN8F5sFLbZLbawyz+guDBIAERChOveTKf+x6dCTeGDwaaAF2MXQJ
TIQNaRRBaHjWpPJmuB6IWZZ/ohWv9mV2JCfgLXrmwhr8oHgUYmWXjHSr8oodpQUgn7tRt9QfEEZ6
YoleaxT9pp9B+CJLVtZfSG0buaNYnZlEtfFMN4lWCUkPxr4dn0yI7l/ea0XAfgtM3AWyievXtZAn
ZvjWn5mCpbHCxFArFyYI5XMb3XDBVzY6jXeau4c5zoH/2Jxmuh57u6uX/Joa+sOyd7ONB7Bh4YdK
Wzu2wdvY7/MWHpbYJ008XXNZ/T2UjHXeDrz166Jo+888TsQy92mOukdkOMPzF8eFSMRNF9UDGkDl
BGW0pZu2bkOMxmRnHhh2RIXCoK81JEeq/WTjt3/2/yEh/TJvKaPkawoX99POQNhmBaWMKBNMHyxL
CqlaSNoQRM0Y7476YC198nATPwusqie6W9SrqDGrm4X0aOJ3ZiCec/sQ1fbtHHyPBb0R3Rm3CdLj
bOOHK8sGtPPaS8d7ZrPfx5y4XRJMFUP00siRmIvdJsl5f3HZgOhZv5YHvL3TUpsuW1pSdlqO2R/a
jtEJviMrXZMPuL+S1X7TvptbK8wPEUNDRgEEZSlXpebx15tUt/dNth5z/dovcLslqE4SdlGUC1Rf
eRsfdyeQBXaUrMvF6iU6t6wUrXS11PfYLpYSb2SE481VML4B5DqPf4bHZbJYqT6xJlP06bSA39DG
QmDOpn/H2HyCwGvQF4b4qCxuJJfYg1su491Wwm1IFBz8CrFBCZRYJAOQL7+ldLNHXH/6nkyrmgHl
p0vTCUlFWALTk7YJa16hUZJoUlcnb0Fg9EWJUNdTPoVwYE/PtX0QmXocX1U7P2GQaR4TK8D4npr6
Y2j4JBlyMFPXYQXkeXDR8aj1n2H2R1Fg6UigQQu+8pBYyySbApfU8MXMTjzKN0vn9VW50WJbaqqX
rgSl00+mmIftol2qeHVVC8T2E5TguBjbtK0/HC4S8LfN15JrthXwMjcXPec+8Qo6r4flRAbSgPXV
K9h/4i6EEXHvGiCCra0KSHC8BxXKafy1B42LmdneJiFBRfCdVPy8XuXiD829m1ePw3sXL/QqLEVi
qjwEzCuLWK5UGWvfHCPf1fryYf/3Wha4UBSRoAvKjHeWhhPkjlX/ZrOfcSgf/xzw9Ye6Wuyj+F2t
kYR4OlL+HjYqoAQDGARm2sZoke/XMpMG3STyXoOndlsL35u0qxAO6LzXx1w/xUsuLWbnJM080N/C
Amhdu+uKmlnhNZmgvhyOcCSXen4v+BO5oHfBjVTnvvfrz0TlQ0njG2ku7na8Ld5OB654q5W5XzKq
rRPq61NFcoId7u2t1Fpi8HJxWMu1kxS6R+Xw/ak+J2HXZs1uY4f3WLiqzNCDpruxwZLD5xygxQku
jitIT/7zOc37rOFdLg+yE/fPX8sGzg0pLBLh8ywsg1NcU8DrjD/inUYOIC4NaAeOPoj++NDPyBEK
q7gBeTBllYEK1A7EP4fbXKQjivlS/ZiYPqLdn7mLwgi6wIvF+HWLsm36Rr+DyzcKI9/YLtaq7tU8
XA8skZ33S8sv4WgUoExqlbo0Fw6ZziW6PACw6lpGxxKs79zBV27QtAjmuP8NSovH/8ryp+8UpDM+
PiwUUlNqrAxi6dUtdYo1OpzcM3S5o3UCr7WQNJA1TD2Q2H5ORNMCNbP0tzeRU2npxGyqnKA7JylC
paD14iM3kLA9//EXVj3TTZV+mrzIjO3biElecGmiZgDNkEmFFexiSsxyZ3ZbqLLs7kVGtXqUmVlv
F5N7uR2kSFkcpftltoa3NwSnCBuwYvc20H+u3epZLZKouOE9ldS/IXOukb/R8Rzd4iXIMqq6RbJj
+rOcfqBZRkhrVbhvzT3Rsfgy9kdvMi8Bm9h01O/lBO7OnN6qpW/LZxAkCn33/xxbUKm4dlrqwrFp
a4DUGijBWMiH6JWm5LiG7QgY/Z8FOyOi6WchlYWSL5S5y9QvQML0IQOec6g2Vk2UZkKTUEitsSBs
TBeRDq9NUpBnAI01QuRTsB/eg8IXlBWpfA6pTFnLrHsRkizcatjq5bU5bBUU7py8PzWfmpOtEGr3
oZW4v/jNj0pN8FgaziEJqr1VoWaoWs0rmLsmKh2v4bwUfL+B34LiiPXNVuWFjM8dqlTmQcGYIyaD
HhTm8pyaMcbxrw9J5vq1ZJmRIPol2bXxDGLovwIBaxLKGQZWWzVKNe7LanPbljp0DeGAmKsD94Iy
BJHeR+P3Rz7/41WwA/KnqEDWWEOljtOBly4imFg5rKTjIy1yhclRQ9BeyA1saFm4WzZNnSYzDHf/
PdnTrhDK5Tz5x+lY46edvbcVcyOGKUL4uruGTF+v3MKbUvxGVLMNMTedgXAJg85nsFRGnMUnxlzJ
orVN+ObnbpE31CajgwwdP8L2YrBWpKkLDZ9Qmr6atk69mPjwwKsMqjJvypgouXTAZQRX2nSULSj8
snUno2H0a0ikFuUNi6+TWuX8jnOJ94XqTeN4P9QoQtmho5+LtUchCuhHhPRQuqYbcMzi5Ez1KLkL
5WHQDd/GdJS/8FGzfHmfaJl+dpaNLkaQmEnzNLVteLep41/k6G0xuLzzsAeAEZ9qHGCipPw2nx1w
wy+1/0i20hWlBpHqbZmjBytX8z42HqhsFmzkwn92iaWlYvlDpDmAb/lKmUmG7IvAQDru7zkWUtmZ
BOssJA+TwSCOzW8O6OjmcoUURbiyP1mveXw+Hf61u+g0+043sqp80958zzfRn3BfdhMe8R1J7u2H
thfy+M72bbEFw6t7ssnG0cW8UvMGNYOquq8acc4dUbLitJPGfguRDElbIhOorsZM6OtV7iOlrWjl
QpC0e+9PiaeL0ZHbS5wcerNgj9Y1FMTsYuJz7oQwcAY9kzi8TBl3BrB20Iap6oWo6mpdzsedXl+v
XvQBfzf9Y27n/pQ8SYYvCtvpKYhAzUJOfBwNH/VO+2wlgf39jetQtfK7TKT7CtC/SZC7Ln/SzKI7
jc5Ht6L7bmY9jf4+MzTC0bfhCX/hEW7gFr8qNZohkFUEKGJEHydHXb5UaNqgTfBi4aeUUlzg+unF
/Z0I3WT/9VQKG9tW2PEmvOZXmWb/6DfNL1OJy0E031Do9N5a4YQsLjpe1jG8YKdLGSOGTSBwxd+S
jeenMszD8Z2NoJs3moQ4HQ7EjY9nsp9NuV4kVw+Q4Rv5KC/aTQ7q1LzWcHNA4qGDp9GbADt5d+gL
XqUdZ8JsfKGpulDPVz7/O7bCC7bVAe3JmqEBIOZPFl/jv82v3AXLqVNhB/t43TMTkfjE1OvBaxYJ
VpWZi1JtF+muIRASWir5QfFTjCRhsDvQuMgz/J/qKQU3LP6RGv6qLIORAHVmy6Km/hmS/KRtuLHS
XXHvAmHhodn+OC9XRr9WRvLdcU6lCNyonq411UNI4EdK1TVeJZbCBUvoslfx92v5GOBkzcTzyHZL
sSQNuBAeuVWGgYKV9rcgLBmpEwJfR1LKptfSpvPufoSltfQQidZmnQZW0Uo0hdYdHuDiWwmUpPuP
iveUlb1yZxzxrTkyMJbL9fPgl6NqFvT5I7T0Gym6LaI+paPmDrvwNAU1qe+akGbKyF1Ap5pA80Kn
+b/foZ9n24uyDcPqCBSOYmMr+k/LekPyvJkeOJZYGIT24yaYTWXRWSKq4+OllYxrH4bXSrRIRgYo
RYzZx76dP9ke8sodRog7+m9NkWlyyb7oGRTnD35ewu7tRayN6A2VePQq7oosZDQQLbzHl+M9eF6S
Q04A6GNAZ+sCUb9tqADAz3dbiqgws7aC84uJ1vhRwlKrIiI7j/SK9Ewt0WOLC7jQgoVGAyCCYado
PB2XsIYpVJxB+Btd2+ps89o8jVf1R5xrXuSvMH3/KiIRTTM3XAhfaX9NgcDXVk3F2PxJs/uCt8PA
sRpjYm6FPDxaxF5OJeGQxB8kvUX3pFxT+3dlv55tHP1NnvRX6LLnJHwO3E3oQrkOFdcRNyulth9N
MD8s8Gcag0m38ZcK1UXLuD4drC4YMttiCOX/+CA5TRcYe5B5JpM0KKAH+0pgpijJxrT+HNaOk75u
BC+TLIACoYAEfyq6WAflHboAoTfoTzh203O4LkB1p9lpkYFlNcpcg/+aMexFEmomaeleI50jzJHx
MP8OrEl/dhzuMCLD4RISBdF/ypASVjj28FqlIqFoQrSdi19L8zo4qWE50r1Pr8jJDeRN1qTLsvw7
mAYfy+GTFnykRdGZPPXk03Ox4J4jIGHkkntjL7q2olSfOyemcxGcUoxuLOAfJwSuZdtMJsA4X837
mZ6cuc5tk8bnhmfeeYKnNJ9JOUoWiq81GiOvQUBdW2qIl4L8Mr3woB9SkIGzmpgGVedKToj70sfx
0XD9mOJSD1dE98yyCHXuOR3h9PGsp3mFuyrvOwiHGnsgFvOtp3K+xA06dtF53XIcNNunvUSoG88Q
jaxUjw3eRA+8zKpa8xDkKEOORGkg2x0syy8/XQQ3vmqTVtIbscJVPzHovUrjmaxnpRW9v/smioEp
7hXlaEkOFvCby+R7M/+aiBGZRYHECyqxC/9qNkxxqdoQLZ5C269+VnxVkm9P840NZIh5MN+PjG7i
xoXKJJsCl8I3yWhox/NWREM5jg+iicgrllN+LIgbBEdHzl5XKBCHSnz+bxXrTggHksAnFMM5JT0g
sOEZ/nkpv/h5ZZofCf6t8nd7YjOLGm9ZYeU4X9B8cXXK6FjDvAwshc+jECINOHoNmuQu2KUtLlHe
MXt3fjQdzChZwZyoOzWkNN1T8I4pMp2vUDE8i154VtZlLVMox68cIhpFwAue9AgSrcuVwuT3RM++
363k+brRMIcZLETn3RDwjMUvPg5IFYTCXjvRPoEazcWeeohtbGZiCavLBIk2JjbRdG01tXLZVzfA
sG5Upti5IlHSkiL1d9AZUMYnR9jBJ7BrbU3NhZ1tagNPQLLdbgbY1U9NoqXVjs0Vm9InddFoL9Kt
3+wb1PZeJOAWg31YNzppZoSUiggaPTrQsBTgr08E1YHCvENeo0M/RLUzceBj/iR3M1g83A/96Bw+
gaCSdTQ4/em0xKckvZy5bX42Ra5lI4NIfd0f+66j5EtLxh3+Kxv94z3okZfkjXSzLX5xBpyfklFI
FrqYDtpfSwQwaEJDaSPYRDyG1YY8hl+UfVZYNHxSHqZqLnBcgToSe/cQdkbk5Oio2Mk+UJg7evbk
pgMStZ0C7+olEX4DMTqW2qrppVGr6270LJEarr7yLBii5fNU7TQbUvCVyYsRuR0GF8ZKpxgjKkgu
eIKieal8lLeHBNgsfQQjrqv3sLwUXfBBDFr7FofW0Ka9HF+vJwu/ERHVsMR3SeffEX6HOmiQIXMV
KrAQwaBL5tIxYGdlcQcwdBOVRTD52/RD2Xk/JwrB5VZFwT7t/etTJV+0vSz5Sf+GO/dRBuoN1ikF
rR5uwb0UJBVEwBoRjqcnS5SJ4sBJQSBQif6xjEeU/4RpClCvPIbv1zVcBu/onqnv1V5hXA5Ijgm+
CYt/n5xpUnYCYKdNQA9oWd0VqsGRSiZqQuFU1Qvx4l0JYaID+EBjOlkQ3ghRnMhUlMUwda+mbptF
l+oeOtaKies/bLZZT5PTCaMyEpfTiKQNwrydeXzKu/Z17SXMfplDXQh/DZA6ux1XJ6/084LQMnoD
+ow2jnPcHbwSZZxe6GwG5l/4NOyWkqFkBKRoXlBU+fYDuNOGVubQZ2BQpbUgXuz4rviEaC7dGiq3
2olkPx6Ufmo67o2sxlUF6GEXFo3QBz26fQHUhLxfP44FE1wWPnEiIlYfWz2mWl2u20vTmSG08WFr
F5a+agBJYO1jhdlvT4ZOIwtxcogNyuvF/pzvtp9CMK4dS+8p6Bd/VCXyKhlMm2p2sk+G95BY0qX5
/zRxK+44Nc66ecWYbxVfdXTPPjwD4pSMrP0nmJQEi56TUEucI9CoN1ptwo+UicaUT7bNpQPtIElx
uxh8iQhCPFBueo7L+nIRDbt5MgkVltSyKlJLTetm5IV3V7f5egCmp9BbKXA7J/hTMIXldf2rLmix
1F8I5Xino1s11Kl+y2zpCUEg0gPCvnVN/cSRV8cLjT31/YjqGqMNvEMuu3LNV59n1eCuNu/N1rWY
Sy+89lI/hGzXFF2JFKkd+NyocmViRSgVkDeAn++TLXrHySFHU1Mg9wY1Tjwo+V5GWY6w9DylzOcI
kUZ8jUbbACyvPuhqr1JK1ypqPcqRv8ABRSJ/mBZoEodjlazLf2bYSdMBkpKAOqqYtQiu2GvRmRW9
VHDkQrlB/Zzb53RlS2Q+xpvUtcRCU+UDpF3BrRP8P3YaUWIjzPuMTqBcqZa5hV2BZEZppe2RqLsQ
K6/dj4XBNn8Re54PAkluubaK/5wev3obce+StexA8Q844kL+QjeIw9E/A2UqYdqm7WCNNhDu1phH
/62EJsEGiGIYbHleHnPfLiUgCcFGl2bSTaIGMf7OPmV2rxhApu215QeU4ddhRcKKh5bgjkUv64g5
9UUtIQKKfKkpzeshswdR7P6M7YYQZzSwZZsLj73X5IRW8bS0jduDxslO32HU5B64TZrhEKz0LJ9O
0yXNn6SGElI5ePIJ6J6LGtZ8aNHmNXfEna+PadckZdlc5oiPuu5yb+qjFi6nKDBnAqeswzzQpeE+
Mc4CkSMC64R/dBe+pC548TToqt1hRpq/JNue8rv0etmST7drNEmCVG04cwgK2LiYBxjenYqh+W+T
gUosOEKf89VM+c3txnrcwlA+Yk/SMFthikteWmdXtmX3erDcElAmBqYFNcnNh1ARAGwFFczref/m
M84k2vTsz1gC/LB8bBamJE3/3YcOr1itzrJZc/CDb36lmjqLMrb1iXriyC+xOUZp3e4VyQc3X52I
nMCOD/NG5ZxHMApM0G+Hjyiv61NEvLDf0XpcUlmICUzAhCBkp0C7YoXXj3ad4Ca1spXVHCG2fnLn
zf+ytd/+h8YJN/bwBzuYo8gzaRZxyAaClLtzBwl8LyLXmWgXzyMwrXhdYjoHd8naOCZ87iHSGsZ+
YM5rZEK3QBezt3mkZcMaCmSMBIQqgWqxm0tmbgdcm+0z7X3nhKIojCRrHUVJFcPatW2/lLyGadD0
By4CuYVCe7r4/+gZJdSnfhabbuR+SDRU1QcJ2BgvMeNrdKWG26RzjwLY/7O5j3M+18sYEzyZ80kp
UhcOAIMk+fn7WOQ1KgxtWygOdA/CK7BVR8/s2vx/tbwSJwvG1mU7/6kJBArvz8oKVMR7OUWtnS4V
RxsoF4IyoHcZJlJsZ2qVrEejfkTkwEHhi8qr5iQJqS9RQQWmXStrc/NgQVOuHJHim2L9uKiv4LdX
xpsFTuwlOdXQjymRX3P8Lvd8IfwFKlTJ1lI1bDM8yZ0YtKpUtpEWoHYSkF2HK0HNNJwXwPVfqJrd
eCVUGi6bZsMoz8csrfa4qavVAI0m01Lb+Ji8i9bxf92r902592dU3KRBMA0jeVc4sXlO70mTbLgj
xIAL/fWm43PvC/9kr/EIfpIpFg4ul7eBvNya7YTvuBVQX7pCcpg8fymkPpmxsJdF6g3DP2IIFjy9
33Pzdods4HfbrUjV1d9PiiY3DW7gd1wl8tNgy/S/l+iUw/8LBELxQDDpZvPpyhirNXOM+ikS4c05
d0B9j9UN9U+36zCPWDyY887T4wkXDLBwL7EP6/KiVyxwT1IwcqP+ByxCusWjNHc8dIzZg3u8IehQ
w5czHigwqEcbzZKGt5S47MqLPnraXspxRm9CLYzFQwbVvY4G4PH5EjdvAaTQAKnji95cdDkndbcf
WVkWMyx7SI2Es4hk1mqXZllJqARZnSyRs0lO/iqZra1ZYxsShXJpdTkbDnTDWLQUIqHvYQ1kwhvJ
RVeW2kN3FDgtIRvcPY1PG3N6EQ2laNcoBu/gifR/65t07cU=
`protect end_protected


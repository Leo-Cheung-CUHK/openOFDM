

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
INaBf8vh5mCmDzf2yp77pxZAxQdyEQiT/vG2dEgvrFjseUnGc6ldwH4JvdnpZSpdf/ihioPyMNjl
u6ooyzv5TA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
S5XIZZtuFR/MZffuhwdnvE3H9oRWM4uXoaGZTa/Dyk62O+Wa0v41pjmZELCiR7uodZPFQfykZ6K9
2ZDMu8dB3afQRMs5lnd/53M1b9ke+MNEeZ/wzjUcsJghubnEAwzdWeW/0tlqST1WD9B/KCxYqwH5
Gj6IZTTFHAXcaVhnCT8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CM6IcdzP0PbD6yMSqylmi4JE2qpmxiNeI+prjGwJiD8e3Xsynu3PbGKJAOpOxtR1hT/3mpBcx1Rz
Fkz0QBh4wtE8fiziv1i+xi8T6cqC8ClamjrpZ//sn6dh7NvwSYik14MlwVuei4DZoZJZF63aoPUn
RXkQ13wtK+MkYKBcPVSZMFZmaCU6jMMBYclXzvRG1JqqZoa7mWFTeFZePUTXG7Wo12QaZ8GUi0AV
UIshoN25yn5e2Xr3FyuEtm5AvsZb+iLsgLeHBtKBnsVaHQphicgqwgwv6MQQF6ZNBgU/aACfibDS
3+n/mMMm8k1cj2bW6VCi7a+c8LmCf81NlJuLww==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ehl0CusS7+JNGq6HfhyaBMy68nccIdIGqixoEztEZfkCpXuUYsdqw6G9MIJdWdu0Ck2acV7K6IVg
rzb8/bNaDDVWp48kupToegTkOdwDkCejEqppido4BkJ+iEkjPniz+aJHlOlOwmauETy2hCMuuC57
oWDprzGWlsqbCjqzKrXmPYm6fNdcOa2DiOYstQaMFNbPU2ccrbLJAiYMHNDqtPNqWxKBsD67kiGf
2eOneDOmdmy7YkNsL+cx8MJc3BVUsYBrpAEsGyFMkmX8a8nYz8R/wlFQFGQAd/t5XrfxFNI58mj1
AHXbcAMhGKVq9YdKeU/vSXY/NwMqp12xJ1nUaw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
h/qRAwiPuqY/Zg/QWqbaYm8xWTi9SshYuPzyL0UME9ZDDF+C2CyGAugh9HzMdD0kZmT94TKmBgLR
dKP28nlE8VCCU5rvbjKxfn/wNtNKHCvZ1hns8CF7+pGuelhxGvXNmYKFw5co8+4grYFaDXeoZZR6
S5sjvhqtSVD3+qq4vYWRjT2Y/yes7L9dRsLq2D3iZ4xjgVHuIbOQLT/EUKW+9iYudT9Uy6YTwB+5
mSb0QK3YfZdGwZyXB4S3mdF9vNQHdW/rnACq3yngF+lprNkh3ooQKdGqtxtz8KSQxNZOAFE+koOw
h00o7AKpvDAp3uNguLvnNJH3rugOhh95b8Jatw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TsA04vIYHDZne2CBj5bWCBFH4MtNoFDCn/3DNEi0BwutuUf+X+lD9kAO3kl352WHjQbF79Ssm+PT
fCYpODgWdxSVbzaHFpITxCQ4HcIJhUeW5PC5tw09Tand68D6eg84qRguH+llbb5jdGJkJeTCf+Mx
pupkkLiDvNyTYWe+nqw=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rx9hgQkvaJJTJJcTjGFW1DrrWiT+xanrcMvFn0Z3KRXlZvf+SE7IQgGCiP7ZDA6T5z1Zv5nzS4h5
cVi+CvwC9UMZRWmLDAjzASJ2nx1g9BjbYe2vHAUmyurIiR6LSigTeM/9TlMv+fFwJbqwuH6FJ3/z
Vl4tIMk4NrqkMn/riOG87SjhesepM6kcQOBgDGzLTG14z3qeZG8OPzxgApfyubmX4qdD1oTgGm2u
Q4mQfFxEye6Jqkn4Rzjhifs/ieNYomHlK7R2/72QJj5j0WyYBIhvO+09izz299Z54ZP2ZXaRMfDT
lU4lQNqQU14PX9Yk9p7sy2PnK4vTwwF0CFIgSQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 296320)
`protect data_block
8L2kCVSgZH1+0liw5Dxxep4kn+2UVndFyTkZ4bYa/WIS0EJAH+sk8qiDBKnAFS+9wWoxZ+HkZId3
tf09NFRuGeyhktnaUUFpydG+RSsesj0/2Ch3m01d53bZSN4fFV6S52TY7bp20b675l425S0JRgBW
BWfszYvJEDWA0OXP89zIXDdIO+zwUWB+8TZTvGBvYJOtc5F7lSSex6k4q1ObV6h9Cqk9XAzMBcPp
5FLQFqGDe8F8TOFIAX26o+8hwwkiyIPkiHRKBeWAK7ietTo4Xpl3iyBjc2dZdMZQ3LOqq7A2H4ay
pqClY0QMJq5QboN6Tx9Is/1dJEk112xQsTjr6DGyU3/rLFv9xFw2zCpp/fFKmYkdzesby0r60l0Q
hclsFiRq91NPu6MBcNqd57ZRVUNRKMvzXcmtn2wGmdBKnizWfFhFX85Po1LIIz7bx0sXWn0zMTPF
QHUJoEs2rJQue2vQVVI4bJdz7dV4PNmHx/+HLCUG07cucN4tWZp4j7MKmAMQLSNh8nyULQmlfAqE
ahhJEDOmns2YJ8cnnl4L+E2M7zd37jySsj6V7as8B3QgEihpfKkKy9py7xh3JpgzC6KA9Y9Co+US
FCT8ar29G4tC5YpUoLjv9EeEjMFhpCS2BhVXIWIb3VJN6wVb9h/lQ5aXTTVKpJXPt9woOj8rbP8f
O4Pjzs/ArWWbAGpIlidD1tkheqfnk0srYd68eMtkVIwUv0lOAd//Er+7eqwBrhK6A6kLBDkYgnOj
G1MKFgvuBp86QCA+ZdoJfZ9v4SdHgSKyPmtB2uqFteSkM7R3f4BhAAD6dKe4e3XANVVTlKThFebf
cLcY0V0cf1ZNxMwINeNeCKsGG/sLh/AiKoz3VTgR5f7ZB/LwCUVKpCPjX9RKNA4gps/sKw3vBkXp
660DgLQKG2DEFN2oWsMp+Dkgz1GhVHek15VcMQoUhFVymz+5RQLTHpsRbiJHGnGI/u/00RPcZg30
tai3/F3BYE3t8y4pMFZtnW12aRBk4pAV9nY98D2N0DX4EfQi8UK/NW7yUXBn44Aa89lwy3wL2utg
wPBG5fZXAH2/j9Qpy4GqEFzlvRw//99G4LlY4wB578vdjBeJE1wyPRrhTcYYFJ2p9+KZbODnHn/o
KrLkpVJ1KKGcghlpzlZrYNw2dHfpp/ALd1idq0S/M3myP5FQgyFjnHBYrYrmCqWlHE3ASeNZT9Z1
lxoK7uQrAq7U64PQEBThUlJ5ljsL+6+qhhpfhvn1ROfADT2E8rE2wqOOfBIB767dJu4F2IzSA32F
W8A46VJiqg68nPc7+A3pWz2j4evB9pTD2Pi7lvfId1ACIFPeymld7KTIjYftWp1BLAm+jJ+njLn2
0G21e1s9ASnLDYZt5lCMuXQsTeOnYVJGfYkiXLyWEaxkuibe24RyywmeH08zCPJYzae9YJ+w9Tgp
1ss3Rpp6ae+3n0T0/onAeDqXHEei2/plsb51VjdM/sLlm23HKvZGSigA0AhHq35ciNrtRrBOsCPj
kQV2Joq4rkBP8ydxkho8rUpbildZdOamv5xpdWxEYkdzqgHRvlN3Udq4lHMAgzSG5w5GnMl6nuS1
6FM7qUcPZ39MVM38SADHmIDyMINwM24hlzWvc7HOoIUx73sYpLwrACnhi525x76m9dJUX8Qg9wob
S1LeK4PA/6/TgMb9Vsor44Y+B5syradM/dU9erPPMLWg69sb6zidgvd3B9xagCmwWAVgTJX0aSLS
pGiuXz4sGABVpjk1+5b2rAkNK3gbyutuGuHonegY7ru0cVDpyKRCuYnWq+OZ4RcAITAhDXKp+I1G
bFDjzepVJFjuRlZ6b5xev6wqaV1/PO1C/hYgaMHVTjZTJGZQdbkxb8PqmOHt9jE766zL3EWimf1X
AXObiu96wlPFOvnIaTcen9TSoNi/7wRu3yYYE4g4bMe/+SaI7PATIio3jJURxxaCoc+a1Rc0sebG
xktU9BpqItcgObC2T5+bfu50AjY7rJVJ3y4I3LEAwuBJrst67uGxd04ugiY32OmA7Kt25ITmS9si
gAvhQyOHiIDip3UQjeG15Dum5X+Ir5kgeUO9+5mcHY2ZTxk/e0cpZ3fAqp+MVhrUIWlcf1uQBfrA
YdJvu68Q/ORNLY+YMCWLp/7EA0VndXLlYixKMcVHLIqPoYn+cLBsY/MAwOEK4luyJrOyHnY5MHMI
1q52FOG1yWL/Or/LEZsQfIDRtSV80cj20oWthooa6i5sw8s5tVtZaEaTJ3Rj3BQ21FRcQhuE6UJ0
OJDxNCvq29BfG3D5/TrgNVxDCuzHhT/VdGkF9YexoDgeWhgOeW71ERtQH/SYRvuOLrWsY225IKVl
oNJQkBjqf1kqSdcdR5+GJ97ilIxe9OKqeMQuQoiFlFfuaJb6VgjVMiy4WNVCb6N8dMah9Mv1ghU5
U5mIy1rSdphwtzFygjk7hD+NwXoPmHJJl+l6gGXC02+WoH8cFChungMs4suobABJJjbm/T+gTXVz
C7PeFArE5Shrj99AVXs+oxY7DoRS+9Pp4NT1wb0uDSXgU02JtqJJV0kkzImTqna5kQwRqu2Kx7oN
CdmIdW1U2Igjwpg1IAtAt7jJSNgv9MbFSO3ibkeqGpUAu2fub52VExTp+pZ8oNt5FTVd9Au0KAV/
n4vq4X89gzIpRCA9GavOFiaexy3JNQKZUJU+diWn7wIz1iS1ttmEDlyPhvYaNbiebZOr5Y7km28s
yrVV+ES1OWqZR5me+9CTQsC5xXR9qPvRRGFGzlr8TqTOkBCXfLZKM9aXp9ETxxv2xeol8aQVNBdY
/2W+D2G94U/PUe9IeQ7Zrh2bHyiiZ9U/dBoRuW+1+nW/NoMOwSfWTwsA/hB5QZcmFgMMD0KxCxar
XFpPscGIV93ReIBgTY1MoEQVc6j+T/06msIUJWHAo1AmvodSNccgi9JvutVe/wXhMmiw4PyuEdIm
KO8440gSmlFvmjhJ4Qs8pmq1iTpeEh9hROt24t2RW6iKvRRvtZxrG/P7XXQx8GVlqUqohmB8DP5I
JNvdOUUmw/0veaBTB6iSRFk3kP7cg5Ek7KmX8OsSQasODavRhlTArD3tooU5VVmP5T0MpRBY1Bkn
2Gzuqzjyx2E/ekCG7Zk7pAiGG7Z2uy5tCOdBrHM1euNvgZxWDRVw3PHfHP7GWuTi5rmuCe6Yh+x1
+LRSQYOYS2y7aFmk0PF6FRpHVcJEfX00QC/bG/rgzVPTZZqQDR2GbiSBRUufKWdfLcZI+w4R5ZkK
J6NxgGArIQA5mqZ6BTUf6zubuh7abBhrgXpNeDADZihFd9pRp+phWIryH2NdkQdzwKKs53ufMkqJ
m3pUp+3CEIQLOfwGXTgjmb9bhnSL0sE/lwVdJzJhL2hAMqkqCXkp0fEe6BwJ9ehFtbVc7Fnjggt6
TSv796aHGMdMKmGpwv8uTKibtscAtUv1PVWEUpC6n0PbSbMxmDPzMy46XSI4nBEV+DyshOIHzTXk
DpugWjdLoxZReEPu6e9K8cA82f+08f8iWyLwPb6WzfGQFoiz2r+p4EpoPjqxLvy7CDZwIqGRcJ2g
zcuH8zStpEwwS87XgTyxkJbreId39YIVm7x5bS/ZMl/amJy3oB5KP5rtz4v63pMN4IWjRI+voY6E
cUYVhvWgoAY5Fn3EROjNCewwyHaMRWQgS9F0afnqgEG56OaOkvVTKBqjlDIoZp3+4aOy59dzCSEE
GwQyQmAysjmDImDmkThETtsh6lcPfukZ0p7bYwEjjJHPJsMExJx26MXMx6qKi3/B2Hjy1KwZ43Yt
ractYq1kTIIkdiJBwMRRUh34L0iYpm+xGw7gpRq6sUnEWiHI65gzvkLbyw9R2+Y59oKFGicDoBVb
KHtKrFGA/Lz5uD7ih8g5gFMC4Y7zydeIRG2vlvQIUghHhv0KCNfnq8r7W+Me/4IWapMQu3d27guL
a+duV24rvfCbErVo/bK5UQzB+xRhwwxIJLOMJ5i8QF7TH2ohhLfOsp0fAtvy7QAXisxv40XLDx9W
1leZ/PzPaA2bMMinjDSMx8JDrePbB9wEMzp/twi/TCy2yBu3F6uwoKqXqotToPPvyVTfWOaiDky1
oH5gzjzX0ZDBQngTjU0//zW8wLh0VW8URsdUPoTnxeL2M834hhXJcrmshQiCpW2MKBsPllYRGHms
mzy21HIbLvukTmIwz8T9aT8Iqf6yGLLUaLvXBZ1tOjWWPxsK2sUBk3Qrp6qGC527f72aiGBDbWT6
ClhNYn8uzA0flF0fkb1SI2N0WuutqqFiTvRWH7nE0j3fPgrv2ALif3eww5D8+FHCEHi/3ZlhO8Ud
7wZJ8hD2RF34jEjDbPaWqy/wyWew1G2o2OJE/YfDJZpcunN4LRpgMVWyoR+Go4OMwd1GuMPfBOCM
BUHjPkLZ6JymOOnXLrKc1PB3uFkDrLSOFNuHIHqMaYEzLeEdDQW6zFmCYM4hkxkV8kr1XFdh7rO5
0y1J2EMZKMygKjc8BLGAUgH93gx+ylhrMnO8zXipvGmjkPptMuscwLZrew+gpK7m59mc5BhPz/Pt
Bz0uflcStOWT+Im6C6I7EAJn7sZiVW+nAJR3nEno50gGvz/6jSMbcp85bU1SEgSbbxGES/mGA/HO
8dOVe6FM+UY7NIYMhUI+v3jL3AWYQH+vy8Uu/RERRAXYpeRkRvuaGR8F+VZG4oVOr1NnQRAfWyLO
vadOobCk4h+HUea8Zw4uuTsR3NZCcXRaBZ9Spm5ySXNU9wNbBZxZVT0x12/QLfh1eRxaGXmiVaPW
/AdEukPHc8dIZR3FTbDK3StbzaZkh7UNGbYhmKqLDFq8L+6xM54VEpnssMj6W6zKKxqjr+gboxQw
xQcJRUTJFVdtGYWUdnTYUOiXjoP0rIs98HICQ284PX/8wBcrfLgidthmaVCrs1drYFkFoZOA7r81
rSO9JOyVqb8AZbrjkU4iF0zAkrIOrhbDUaVA1m8b/0AcEt10ruAwLT9qfsOV/QDxm0Ds5anm4NKL
DEqS5x2CvatCqsqGx3hLXHk28qI6mPoeeNAJwO4blHFqhHXwkhtlZ8y1ZVU/+axo6DrxmSCDLn1x
RMNmVqLn8XgfXbS3G5L9N50mOI2FFSwgtohbePqQep/HN9Z9H5/OdLCyI+msEnMOowyfxRirBsEo
hLSVzFKqhHBGa8l2p/1xivK9Lcn4KcqVeLEGzWC4V67DxnFky0Ka6X8pMA/vSOd5LS+Ljq1uxtfD
2zO9h6HecVr7iK14DMuZ4cjErwS/kd1QpOcY5D3NYLUo4Rd3cxqOvn0gF/JOzuHHI7X+JzbRstme
t2mMZTDtG3y41aEARnRv/o0xZF/mf/04U/jTgL5wu6u+M+9du56dvQ1xNM51M6cncBGgOkGkHt0K
kxqyC/h++Vhrx7mToqFqvDyeIg0X7DXFH2ASCQD//kmwCh47pgIS+/1PwmKgW+YP8Y8+Ldb5odSA
GZVuQkNReELutxDZImDYyJ/rNqlugkKfK0Kpe4CV7SOMn5L59yRDzU4T4i+x20nX5iMHblfvO7py
2J/dp3mX0soq5MPwDiByOWPYhNSeZddsj8JT9Lm/YSAaqkFFEPwteZbWYvEwg5+iKPBAi8A6Guge
h/Y0FPPoAMtQW3HN/fS/YvaDGdDuvUqfXioNMgGiM4xFdokThuUhioa/xwHDxnN1NPtboYFVDGN8
NPHm7gCaXVrsA4XEw3dJG3XejVbnTI8Jy8Q+eyooDoTVXNV8lJPqOedXxVSNMgaUCMFkEd7GKZW7
EgP/o+gS7jFWL+OgKQG+JiHGMfOxuTduUFEI1EgQoiBde+JpfvdtOCel8yAaiwWx8Xk32TOQ01U2
WZNWtjUWZY+2ReH3Njg03jbKtehVdfzPMG5luQX3z+np3NpScxD5dI8q+eUuiidnqJjw/s8dK4MV
lsI0PbiJD5EngjkOAtbx55VP73d78tQsDxT9pF7Pd8aARw1elBKQufhuuwgu1sly5y2H0lsNCYgR
zoWCNIBw/ErvnLS90DZcamcLAypxhJw0oRvcEN3xS96mUH7ecdVGwIivrgh3PNBfy02RAjyUmV+B
RpKi/ZmAEphgKQTrTOs5S/qGuXLuKi6DcvSeLH97VXf4VoJt9mpLTqqJc0vI5SGuqwejJ/RIEIJ0
YoOGpXJ2rQ5qb4177xFp5r9LxYG+qhySTnMDf515aplBB3caHB6dIkG0hKjRdUrkwd8cjQTcn3iA
FrTeCsO+O9NL2Yleswopouj9xHjVYyxFljsNGhksxPA3p2h/JTBOy9B1Xkb0QM8tTJMCjKWDjMTo
WtzHdAJyQ4GtXAUutKnO7dl3iVNBWWVE9cSiQIJbeNO9DdqxChGY9aV8w3pAauvisL3hIjZ8SsCy
Nv3jR41tDuJPqgPpJ1Lew7BtTJFhKLBuos/GBttnhoaaU+4iWkO5NokgWpSiVS4uaXslpTsBNYTt
/hoDA9IGIAouLKcYAgt+U4b2l4SnoNU1FEviGO4/hvT7ceHuIKrq4krdH9w3fKJgIF3l4Oa9jMxj
cHPUDRJOL/TiK2432ofpZbTSZjpEuuSaWeojeh85vPE4f3NHCv04clgDrG/6pN2P2da+NlnB695V
D6Fj8L0C3Pn+6aelv7LImfJVhstVj7EShJ3V3K+/hFb8oHJzSVQ+0CqH67x2CCzEYRyJzE85V8wA
m9cpsg9kDUwavYHh/wKOtLeC2ACo6qzSxFlupE+/Y45g/JKa4x6DPfbgp55PvQKRAkgoEBXK74eq
Cu4zcfPIo+ibdiiskBUyT1upU6db1os4n+Ot/st/LZUUhjTIaLJ0wFNy7S5NkuTZ6Hld+BzJUfSI
m4g36cpplLbrnaCsF6aDviAcjSiK9I870G6jjFcSJkVbAMKiv8WpHOTD5PKNcS207wEIcX+F6AlD
fcniK/i1KV7fRzq7Wc49lpLjFSYueD8dZSCxUm2kgGwr3485XPIelFqc3ILxO6QWameK4KIUhXKP
TlDkECjUqrvD/hvV1Wwt9ZTv0VaAD9i961MqjHEAoed69EyVzo6JxwhHH9wK45yVHWiVNPlvp1Cs
xDVqcbZq0e9gKpDhwlee38bXNa4A+sp0lXgCb4xnV4x5EpO3SwCjMVTOmj0KAFvMvSxxqMbkyy+m
i0Ytm4T56n8wqe5RtXDd91hskNSfdNxdGwqW88M6ioSgptH4JTOGXQjxAgxeSzTR91bZyKbLgf0Q
9WpZfaWNMpjzpFVl9xWMZ9qluiDhPnSM6xnF5LGAFKktFRDhI2M7EfT2bb0Ye0uwNrFpOl6L9E1b
6Pw+cD5/xso6lgAo6TMdPSfWw5++mz0OG0xlL1HtP0Z8YPDgETBXjtMmDraBvhHvz3vU+7L7P0Pi
n8V+/PLhgkdT8kRm+oIRIP2aDbfIU3Vy8mfilceUE013EYYsEuR2VYMcUQGCiJuIkDzq+BAjLxJK
Dyi3H9yIDhxXmY+7GO1llqLGUakC+/EDt1eW9M/QfixdbOL8XUVHmJrghdkwQYgZ3reqnvf4cr1k
xcssSdXojmGBot+KiCrT7y9DiAInJrylActj++CwCO6PSZ24L8JMYp9IjkrwLHNIZGUMSBKmV8tm
wmRKAURHRGOQTEyJUW5Hb2qss77xq/jssxTVH69g5sYBVKwvaNuC3EwOBWcy/gRcwR+0iaMFqLFp
OzsbwEfVshXOeOoT72i2l/eWxuJy2hEcB/LVX69UYTz76YFCNZlByCtrAWxJY/8INIOfnfgfD4fw
9qgRf6nWJ2pN0/qPlvhd0YnI7HoGIAwZmQTLDplysZG/GKBQ/fnYTTqXDMCLj5ZtCJuk4Yj2FEaD
HMDE3XnOFrCMCbmNQc3TFWZcIcmnuzHTV1imNnJO9QUetNlvdmNrC8pG7mhi2HyhEQtRbCWlWwto
JlF9Q3h8adl2vFU0RfHcjoJfqLd1Qavl6WSj33TGfzveK2gWwMJOCjgw4yCi2xuTmvfqPWZNpMQ1
lEwadWBxkZXmU53w3viN1c4sTI1GdjqGQ7E85QCfDKS3/bF1SByvOkAtyI/PH6gNRt0ONpkGKR2T
Kzq//kUOtMNwc9V0sSxjoeGp0n++Fn6FCjayM7QdF/kG+H83q4dUXId88ANl1DI8LQs9pbvg5xdI
aYNHEp34joMVfngujMzj53X+fkkuoJ2aS/BBKhcZHP8aWyv/qVfz9q76O43XNzIhU8kwPGDP80/Y
0wclVrbHpKahyHQVhKUGPWWVdOl1LctgI0qQ+sEuEDR2NLm01a1QvmHuupoytiuOgX1+d9o/B4oa
F44jKDwSy+OeqcM7TSDLQMmpx4ZMVRVmTzUbcfQVer0a7Fjjc5k5odaSpeT6tk21p0TpbJxwPAIE
zwYYICkd0at/ATKbLNjeVNAUpBNyzO8k0PKqyUXRpDa97MzA4MBiDp/4mIYVzpetJFMvvD1zqnDQ
neETDUvwjDizXpnPPPgsLofrE6cV60fGWMqkjq7wPccuMomMZw+DvuNZ0310GqDpZvQzlpR7XJlb
KvuXUXqr4ZvTqYnHjeKcdWH2L9I23XGckT6ezA24wO4BKmvbEduU1cT3VV6Cg0Vo+TT41EhH/uyD
3N9oKPC9aiFLFUeP/zwPrMmIoYByzD2qRpw/R1tCbDr/iLSh6fOOSXouSQCy3AibmOi+W97d0fUm
RHB58/b2mAaMi6VOWgZ81EkWJ4KgdcSGnMWJpJ5TmaS0MxnQYGIqnbHT/yw72iFqMbIsFKDkTxyj
JmlqnKCRjOqsQ/8UVaEyespKpE4MPyM9sWqflrHdXdHQMLEKwO3J0OTUt4Nc5F0qNj3AftRW5uIm
znwAYufloyInClhqO67rexKL4Ru72Y4+lINl4zckV5WiYd6fQQTGpgqul8MXLhbdcaziHE5Xf+9X
oNzAKgpzgXyAZG/VTkjkBCYfWNqgr1yKo9+rzNKWiM0pYjtbbggFMoNlDj7nsB2FzNV0Kovgw71n
EoA6dEPzKOLjprsV5qMI4fgk1BpkPulIeQr9w+o8/++Zm2yl42F4S9XobgjLamqr9aU3y123epoG
AohYyAKhSeemFfkL0QfUrc0jEeY/LjjQLIzze2h96HNnR582dT/92+coylNK0jeIkhXvudKe8YKL
9VGh6YkkQH2/yhfXW1+spF9nat5bSBxLzGiFSsoN2vjgvyAbvyZUcexqk9mtxtK3UMxcY88fMvx/
pZyaG8emO04N45GG3X5l3R//spbn1Khi6J/J0EovjsXeKABNIyHNOoVaj2kMASgSNf4KOFnBbwwT
5tXOZdYa0FKbDB5i2lGq8IajA4kGtSosIxRRv5Amoyq1T1nZvHMfaBGgP1Yc1dUPAVeHMJ3SJ6iW
amteRlmlnYpVnY0ulfLmttNZOLL6wVQ4SBQzrA8qH7w3n3Oo395/yDEaxvW4ov7UigF35GTmKW8u
UwXMhdSCIonLRXjk340GfO0chZMJt9ry7ZpQkWpLmegpbONaq8na8+L8t+84JpVpBYCTBUHm5Is5
RYxGYcpri61Sn5LdVlXmbu8Ku7F9uLZloNXh16+APXFI1UhljspW+df80EKGxKUmFldt9wzaFYpk
UO/TiJ5uSKBZQxAfiGQingo39r7TT5nwlzfOoHQrKYZl379gcPpq+6TI9pOutC3RP/5DwF9+275u
KXd2Cn9O4fqmVVtrkn7SqHbC8oSkM1vHSkDTM9WwMwcKZSfJP19ct65MqzVUwpg4FXM3qejRHxWW
EPN8GbiosU3mO/jXUusuJSzarGf6Myf4S9O2ClRBGc+V7Lk1jO67ZL5zqXWy/qztS7eAg2IvFRgT
zT8TRs/sN1miLvNEGqap9QT5Onoscuvs2gwJxj3kHokmZqTp0DbTe14HRCtFxiI1oC0Ow4KrIMGG
QU/WgyyhHs57hmxJF2XI2Y5zR3jd4nPFf3YeOhcP2tvx9DQF0Xeqcmkx9mIVDSleNO7wyatnRBQJ
eT4AECQ1Ka0BDaegLm+Om3esWQKnOdZ1tUMGKZWYLcaP7EOUxkEkf48EoW4BdpgO4/YA52Q0PcDy
S4FXIb1LmTQYZ0Ppli8UUnC69bst8skLeOrwumcw+ET2Ujq3ClqFzs/qnOqe3kVz40mXH2jRYtMu
5Gf+pfPhsRSBMzgZ4MDXkkc5mz/XeGeEO6TnqWAd/+l1AK6XAIe8aAUHno4X29KyayX1WRmGJicp
Srqy7yMRSBlAvZZ2VaTb9jdhPugu/L9+6cw/xm7rbUy+kLc6dzWgpsGBEO8v2Wf+lLTnCBJLmbGm
erh9H0ySCUfKwdZsTM71XSryVRYzgUB2/htoj7x6Vz3br0zn0bB41XBv1E/CVaGQ40Xt6d+ugt6X
L2rRpnybGaFz22mm2HNTEAndF6mP86hbVfqyBF6+REfQEFT0ExA0hk+b5LtVwRGDunFVDig6VA8A
IGGCxjmu5c2ul1xfA+WeCD/vKXs6b5KqyzW5QdFI7/BR+B3WKYpIk8I5Fnm6Eg/9BwoxiZLDwQTP
CDHtp//svWeTy7c3Di7CAFJho3cqqZT3Oon+HwGwC8mUE02KPmmxaF6U39MbCmw0XU7gBkLT/bhx
JH0MHw7uFANw/uH8ce4YGnAS4fDk6X/Jk+c/IKRYXH/FHgPIMn4n9OAxttezpAXf3o7/mzeCGV4O
G0ouIZ0yBFBdfHbgnH9YlX0Q2CI9gcUyH3l6peBIDyXBlgWzedjPYl29bUQo0WxIN12nhk8LVbpb
uhd1s7k+elru7gya2ThwR2XTxUWZsUbhSpPSXrWn3JHlwcPyRnh1eyDVIJM2rn7iPg4FydDlTxdg
Trpyffuqr+BzB4ce9INsSsZR61cy7tYU0HDwDv8H5TfLjBc6BLFIsMvCwPeCqsi5CryrKbl6QViY
vFFtg2W1AX5lzFXgF9Pe5OlnMkge5OGmBiBP7oP7XTiTCYzmWpGOsHKbRFngxrrGVE3je3AMxUG9
FclK/6JQw/tT2R9JXgyDHr4PIbogSz9cSRedQRhUVoJgvV3d2nXjjy8wtENxal9eFVUTZLUDK+L1
KYb7QbyDIorCjIqV2cEBfySZKjczjaUMdjNoiLJmCN3csNDp0KtpYvTHLOMGS4ypm5VeK8DxauIv
Xul8uPFqp0lC1IuOh1QU2jhy0DqXsdH0tdL8yvVNb1KZrt1xtgLVeM8EmSNwnKLKLw9LxmY5d19H
iHMxkml+SfPGnXKx5VNyEQryuKIZhzRSfN6m4rjWz8DBmLj7PQ9YKMXu1rjhyBMoGBTMCOs93rE1
3j08DET/Bj08ZNvzmkoOC0qxgTh7muMK2WG2QAeytDKYZ+tQDnrT9ssURZa0LJANCYFm9er6ZHyd
Gw9u+ILzV0wdGTxMeAQX3Fo8r9RO9EmNRDEdi7eR7wgWkq7kRjWe3wjpomtvCZOSWjdhWXd29k1C
cTDVAcPQdVby3uTEN1cUi196aoAgXNcXId4s7HJfEEkotfBeoVPJjLSSRoIcL2gMMvlPB0IUk6RN
kqofWX0pbGn8IlWlQdaFiHeX+Ko4K2o8uIA2+uFDohj3AshcGgbY7MDjbSVee6ZaMtUjkFN2idkY
9/gEdQMtLSQY0NoIzjsX3ACzIe5H3jvfw7D/nFpKCHZtr/fvwiAOejYubSWGQQ8SUQdnrgnrUYOM
sZ4X/nLLsmU+9kCIl8fEb0XNpIjUlUQuQ14dMO3STXQlseuhGB9GHQSxiTY/qCegEcisRbPew5DC
1joY37MylKAf8YMmOmRALu848UYfTNkAbANkMQOP71zCX08QzCSzCBNNr6DK7CUrUFVavm1RBHta
Ianf1YjxNDAK2IAKDJ7XY74CmDd2JtgcHz3NFhOUUV43DtAI8+IDH7CDQUJC03kz+fswW81Jl0wH
Sa4vtuXjXb3L6jyquRuS9wi0ANgv1YNwn7W4I6gt5vBLtAz+jYjpVuw05g6WyAKQsAtr+er8bT6T
Z+17umTWfoV1kCtfkWiWQ3Qtt4+IhgGdtXpHBIiT7swCV8zRRnZa9AHWkIGn08zPyfG1JsQdab6T
cFZFZMbDnjC2FExiP+qo5FIKV2oXAmHdP4f+Xq3P94eryWDGJ1IeO0eonkjUKlNGrrvnER8Ujs9A
bIhfY6uqN3OCIckq/zmUbrqemBDPxVaLZwP3AAYGil3wdeWpr36E9WO7yulCICZ9GnusaebIKba1
+tDrfasAdsAnvQGaGrxxVTieIUsv35QUyI/E2JDN9L9rM+5aCei/37ZdLdIBFzbWLZyJY8OVmqPP
RrQIeIIBIbrGbaFoVI01dzab4GILJ8leWoKSJUaz6NFt5XJW7+f5rTGp/i2dfQ0wp7FnrNZHbiXQ
95uqxqfJOwgBmpEH6OUeqvNkPoZJX786MzAE+PQO7MZh9lR4G/rz5CWI4C2xydnQ0opNNYfsa6zZ
3QYqZygO7DvQTDDAo+WQvsRzRVEnQmPe/bdpaBPNBxoMIveBOm3v6pKBsZ2LKppxovDdLDSNRqkX
Qy0WjsC/SXfd6/t16vUwlAQgCNzxN/UsAnHngLa8AqdsdLXJg2iAfJzGJ+N4ZVkC+OE7aQPVOGQr
JjhCGLrab3XxL86CVSmHea9K00bk2uQ/qtwsVpGwDbAsRNZMoCbHvNb618Ac/J9qP37V9u2rr3bq
Iq1F5Df3si1WK1zvrnwqkJoAu+2Et1mngK+EKksmPWDDoWLEhbqp+zNgjIgbt6TKuWM0C/HaOOQn
gYkuUIfP6auBZ7ImHlSIObLQ23rX8kuPlqc+5D7BfcEFoSY4l+nvc5qRBR+5qMVOY5dEzattjmci
Obr3K5V2Bt7Ts2hqCVINxXOvsZIprWfXwxWfGSX2Le/TO/Os8EmIZkvI8eey/Aaslvg3KKCl+UB1
BobydSwE+MXZDYPGoyXa9SzelXw4A9ZbAbJLfUvCa1atNG0wMIkWExUszVuk0u1epe4B+cO82VYq
XM2Eu0jdpxLUHpx2sTgccIU/RbxtVAPBAFSo5Fb3EtK+x55nSwStRh0/V3IaT7WUcNFCbPVtckJl
U94FrVfAPMCJhSy8Pr8friGHrNyDNZShjZ26ETSZI4iS/9uzuA1e5kmPIG0OPfhb1w8xI/2A6xxw
qt+Y/pyqIGQlVv7qfN9Bk91l33bdkDWJZwi1nkKhkVMxKli91e2nmoS9nM6YQbpjPimu7aMRkNU0
FwQtkQysw+RU6citHJzaK1XodEvIJuIa4ZDqXzht5LgCxs/n1CVDG/31fM+Ovb7AoTD52DnFPNES
B0LHB5UcLQKdlM1P/xCdHemuWMBLLjLCLAl6aHrKEEwpLUjdX/bdwdlwP1bqydZAcjl3U7m8MGVF
pYHg4xjOvqotWq4fE0hLusszewgsYrYSyt0XopkBuVnpyfkwTQ6AwIKt5ap5Rp/w1uOOqvQ37KsV
bPo4aE6LbcW82JnzNS90aOFUysUxhMEBeHwAZnxMYZ6CYWE77+ZO2gD4iDjhKJO5E/Z5e6t7If2k
rJX2yIhffLooe/uU3SUtcSSnNfXYZJnK+dJIDX5pMD+j6gVX4z7e3psvzzhc6oC3z3WNqCMnZHpD
3wjlSDUhj1tZ6F354jRXhbuD9CAc4GwVJoXKA5cG4QIabqoPyYRVVCE0zOKpxG+iSCjRDZGnd2te
FI0n96H8j3QU4qNic/KRSabeoZXh3pgUOWl1AJO8mpzEqdCnS0CF0Gq/h6fq/JC39VuN4+iXWrgj
e3DdXT+IxaE9Zy/TdQA/FZ52SvRyzhDiG3YArZqshdcIATXMa0mVA7tU1rGlr/93cI9b8zqTK2f/
HCGicGVgu9VBVICWE8R4Nqtq9hP/f2JWeIQnjp56AXdBPyuUnnf5+ARM7oGok0h6JGgd8L0Kxr8j
FgPuIpos51eEB58fSX/Nd9CaZAdDxT//XhHeoAvn1Vs3UHxkbBLAhNue4A1OnIk/+XN4KTn/g5yB
Rh2djZSJePbq1y9CnbpsRu+hQYQUo4N8JbSPfyuIw9+6HGgkxrZogNTD7iXGFq1/kGVDP2YM9c+L
UMGkV3tXmz3ZfjFnngtDbCCEAfLR0xLvo01UoDQxLer96MLcodcEOqO8L2LTmJVCDrpsBSG9tLb+
INi8No5PT68+XsAYbwik4Bc+VrYnm65nyOtxbhHpy1e/oGXpuvcwVMddhzG/3Gyy9rsDzhE28zcy
tys/UEjlUM63S+FDwhAD0YtI0x3StGeQgkVTutPJMSrLzJ97jyUB2XSqNR1YdXU54YDYD2FSgJUU
So9lGUf6jEPiK87WFWtZS8DkVB3QKd7wPxtP0YB8cJeoRTxEoZ8Pzm+/ZslXrZZNS83QXisrLVf4
W1+Rsi/i6ZsQ22REGpZCLy5q+6p2jgsxo82f/R+ZS2SLiBSZAJBWoVyKWucnLWXR+urRP5kN2R+y
Y40+Nc/9QIx+J4eQQXZF3TQdpbcKIv8SjNGAfQmeqsIgBvcxMyvE+RZruUWw1jigtRJZkdsqsMSN
sHWVKz42ikWBLSFOOdQm30bUpabjDZNt+zorJKNod0pwtZt5hvBkxjH3ltf2h0+VVy4EdmEjvaL1
4NfOtoPw2nxZtXKqFmfjFlDkVBNHP5kkyx5+o+ULQx3CsJJXQwg3C7gqUWUyIGf74zgENjAuoCM4
WG8KAN860EPP6Sjs3V5WxpWQzxpJALhbFdWHurS2YU+Iw6SnlIMZqPCq+ogkbVtLDtScpZpYjk4F
VEdiMGCW7ENFoJWH3YYGJWd2XR3w5aEdga538PH22Zz+5JIGNkhG5QVJMcL/p1ljziy7pGizbFpD
gfN2nEPJilCn4k45kDWJrq278czHVAKhm7PPARcIyvJtgQrD2MPFs3HYF8sQTcuLWmIhOgvCAi9A
xnM94Mw82Oc8Knx4xWp4L72RnNNQi7vxiYVYBBWDsEGP73+HRq9RMzVBSWMOcW2neHBCP0cPCqL8
hxQ5HPEOG94ypi4OMzvECn+wk8sLQS9BNK3261+RJle+3gEZr2cebhfSDdKxQ1DY6zS1oPRnd7tt
xlX+e3ISY4vnN/XYOE3yu3MFajhYDo/aNm8kG4NIN0t3CiVWHHD2Gre3jCiZKbtPENFjH5G+eRPc
CIHy9Ri14oqGRsbHpedX7A6akdO0Q+/Zpd2t5k8kukrTQB0GWPDqc5Cr7CXMkbLqdMNUom1b3LSz
o4LhE4sb0tT73Wa0yy9THN2Mbb2vTiD1zg9sYprtYc/nuWmTE/uKBHvdL46DqRByPNynT8NeEcz8
fV4TbqzR/VjtoVzSBdLMiIJmoFES+FRjxCWbMPyEXNA9+iM6s0mwaiTmXkKq3ubhYNLrgAXZCmVy
+bl7YE3/WQSNzaFyXrR6cKL1k5AsY2j4jNpKZOp93vad7YqnxJo1/t+tUFw1tCl/tXpb1P465kAl
n7qRI/ieB/UEjuEomAIz9lxUVJBna1iZXviT2ImtpiUV+yEfh2SMwO24Xb78S69COYgCPSujUkQS
GXaOCv8xbRg6HuBrhGaRg7zV4x/5CKsvcqZbYtCiBIkPVxyqW0NDzV2Flu2bKjAxV1NXx9S7gn9d
IxWv+ckNO9CBetlfOBYEaxZNbRfWjRDvZCocmZSdufCSqUSLW/s21uH635fygMaQ5FOBMVVBXA64
7WLLORLL/0gorDUN4g6b7PcRGg/EMgCKaKG15bqLmqMts3fOLdzTER7vTRpDGzGrSGF09lrTpiVy
9LYIVuDhlVQai60eahRVEfqjbPmQtk71YVYla7KrRBxWVbEKxJ5gTqf6h5MeRF3G3y5VKLfyTBGd
UjNVH0n2Pq4Djmn9yrmQjsg/guROWNzApvI/Td1ggXRRSPrP7TSAFj3Pyv7J8e4lf1MJ+lCAStEK
+3j5q0Pns0xrKx8DJaRezux6nSLofcs0M+ZBle3GexRGbCt9/F/M1qeXxI1mW2q9H2YGdbjvtSva
Xa2Cf5aLTMVZimBY6h/HysaNZGfu+/MPSAZg7U/mmYX7hK92WtY7LABfS2OOlUWj5/sHunzGSC2n
VVkHGmfGOP1WmoDcNrzEPzF2MMLTtSNTEOyVd+Be+EMoVTGamO4LZCmh8gfXlPtQDf8fqQsXsoW2
PBtB40U1aYaND0VdNebnRyOIlxj8NmpBI3p4rCpljJ1vFfWADwgOzX9qTyKACHrbWYF/2c13YEKq
IS/t41zJHgXXp3BH/xZQWnyO1HlsZKvS2NYOg1CxVJUHbWGksNDQ197UTF3UW0ep3ubLKP8dBrqW
pMSUgJdUAGMqUiIDdFs3zRvpqvPsVKUolWcV2+Jzu2NHVQYI/7LmfH0RvviLM6oB+ZDeKB2VkdPz
e5a5IwTUjo9qH0fsFA0LlYkcAJRbhou+6+uA4EeOyK/3XoN92on69NGF4kLSbfPcXR9gp4En+P94
4eqWOPETtoreO69OdCntMgugbvRn79IJjH58g02faEOulzWjCqWatKmu/WdR5eBT7WAE8kBFHjKf
cDR7VfZWfL8YE3MYE+zi5p6x08VZsp3cNdu+4T/VX38pjaFVFRJPWXse9nNzwv/nISuGM+yQkY9r
jUYZuzXVy5bYNiyAZlRD60ioMG4c/idOGt30dBfBqR5aMnxhNI4YDFqYZJUkIexlfw52THaVsVKy
dtNcaFs7+wfxtE+p66ulkKbhZfvwQXFv9e51F8rGTxctsoxmeoE+xeiV6MrEtqZ0IBTp0rpMIXI/
Fu4FR6JuO+a513ls5BAUJv7+HAAhDZ5aFLdTQj43nowBkSc/Ad06AJOC3GWPYPkL5dcPnn5N3m5/
yVdYokG+oir2BUKVjBvtvOUuVaccWyDvAEmIeIldBzTq9QWHadXzrkMDSph/CVoLteh+o9BVfNfG
mRcTPqlBeP7NawC13f4XtFmBn1yJIugamqQPVrCHU/sDT2PB1m97csGdyJwYPmjxS94yS15uVl9R
pzy/drJdqcQCM1NWzvPtDN1eprXSDKMX+K3jfv6IKOP2RnwmhxXjGDrf0rznH7ePnOrwbchGX7zJ
Q+U3rSWH6BFepyHrzUOgksni5k3w652u1aaJZNiVk88zK3M0lilns1STVO2EvTOwcixw8Xl/a4xD
2caE2Z2/W9sEAbx2CfJ+CuWZ+QtFinjrR92qHT7rUE/Stth78fTjqvMADvudWHB6MhhgI6Mg0cnk
wxGzMr/shIOvurck8FcPFdh1gBI8crhQUnLQStnOHSmctEwR3QnpotX0rn4SIh+ZUzhKGbV20ka2
VnEqKgocR2hAmWIk9zNhl3CBA5kDeRtpE5aulD+F7193db42QvmvFUp5Kp+dojiyJsW7fmn+Ip/o
hRRtYEfHJz0E4BRnWnVA+VMw7+neYtyo2YIc5HJLEOP+aiJeKKGDlKE0ue6knGO+vwAv25Yaw7I2
ZTqKeUAhw+9cAX/Pc6dY7UUSWfE6sIeZ4xb8Wr+HEX4r0/VClQIjpNYX8FzkdY4+Z7eOLnRzmRp0
eGQcJDnLiD/9YrCPTUB7bptYFw7OSqnP12HLIIVtZXlvmQxvpQZyGfaD2zKPnLAwYJvkltLmHRGK
3ZERcuEQ7mTDOEBigxPdzem2ZTgsK27ITD4mvGdmuW/Y/ihw+CsdPM5pcjhdJkbLmw9AJsmSE7Fs
k2JtDG2yAsMJWBWIEZuyp1Pt+k2Y2o0Vf2hV37u/i8nGtYtE8MIIc/35RXNm5UyCJQPcAaJRiEWa
imdc0SQwFd5I3O4zhETZ39WusmLHxsB9605R4Qu/9zvv6M3BMJcJNuF5HOb5oVOnrgjUuWuiTkaA
jdYLqs96hse1bF+wXjJmPgd4PrpCWUFQQOsiCjOWReM7SP1GZvwgjvakFxBUyriEk6sDloRnEXKN
J5KegO5Cg5Ys7zdo7LW6vtIAp3GA/l5t4wAQbu/xBmgdi53+XW+JhdinJm4JhFb527IhgLP1lHwC
n9KjeDBYHbWRTo6cmwkWrPJ0N4na4k936aFSCyx6MNAsSuxBbp98VRUAV9B+p9z4qKrAECCjuqDO
3pucivaCBlDPer2281l6/fSsj3BeRxV+tgAwHKscA/w9ZdJQhlB1/nvWYDnCXvLMjjBRdmp+rDCA
wqYNYKZ4CSbk0dUGFztOc6NJlxbJyp11vyNA4CX4ZWj2cHEfDMYXNOyti9OQ7hLVF89Vi1mpwHsn
lpHXzAoG88Msg09PmxvOd6iujYjgzZTQqCFDJfyJCaH07+Mrn9RdMWnbgxCx4GoR8HwxqqgTTNr8
3ayGKAlu1bqMJ6iUNHGiMazjbdaK0hyuZO/Q/n92+ryx9ONgS3pDzkm7lpl+bi6887Eu8w1Gy4Ob
PQg1ix15aq9IDe6yNpNwk4/ITRsZC2c9BZzxdvoUpv0c/5mU5XfGtllNxFq85SVTpS21Q02joFGe
fGpR3JU2bQjDlxl6QYNXxyRfj9XV41qw8SYu/kB+ioi+Q4xn3NZ0IbEJnFZAyNk4DY7P+ZNTUEEf
zriz3R+Y18Q1TPtnGQGSdW/cOr29U/UGXZuvdOhC/zvjdR+/y6LGOjdgFT2q3ZeTnDWgbGaAOc/b
Yo1LSr2vgWJD5NIgt72UAsBwMTZOqtGNJqe3IrWYIXx4CYRi9nyqojkCZdNH7sYiZbTP8x3tg939
VruPH/onJmFDZPHgzNldxjNd5MVDPMtMosi+6JMbAnIP/3b6/AA7PSwU/jPrGQo0LI2W/o30Fv4U
DpASY3WVZrm6jf2RuRukQm/ZTypmL/GXjQutGBzjhK/xB1vKL3dYq6wvRDCqdojQLvZMffCBD/fg
1fpUyYfXpx++ZnggA5MlET89PeH6+pNdd61m3Gp9TSpH4hW60ULoEyFIkq4/Wgptd3qARPVU78ZD
t4UG8TUQlXUSETAYKyupi0e5h+aaeHyGuuMTtHjqdaLFubJhuIvIGZqlzRilZSQ7IwqxsmzFK+nm
RuBrd1hyz1QUN5m3LzIoKfD33d4d2iNsl57jOmf7LZ0Cq3sdGzAljc+CWAnF2rIwbw14ukqHQUsN
V/sICtPhcPElgy2gwtq8OCp2eR7Sq4UCy9aEg7ywzsZ2UY/58l4yp6piReAfLoTge2AeZPDb8cZ1
rw98sEoTnPkwbCQJK952pOJwg8j0ow3woYiyi47SvJnWz+rerTdthO8+F6vrooCESvIXUsMxKstq
QP5kIwcaOAzdkKdxLyOaFWF4oin1HE0iz1jZnYXXZHHKtHJW4ChfKHzmsfXVYY16PDSHysYbD9BH
jbIb9hCAaWzZEQprbipi0uSWUeosOhkeNqb/iRg4szk/Q7u17Vku+5RyAqPApBAXqeZzZTIz/0SF
Vu/LRAdPEX+dD+uWFsUe6dNE1LLIRG4TkzwLJ0q5vmmjS333wY0jE2NIWGt8yZxynAgPZku9sXdc
fCzfmCYzu734pqqn6vuk08NlKdZvP3GxGbaXFJ3tCtfuCMLcWd6zPxHPhvSw6ChUNs1aRsgfn9UH
9Cf6hVBgRieG78Z/fNs+kFqNjllubX780NRwBFlK0MlP2Exb/1HeGm2x0MJSEVm/zdt2192BO+1M
Sn9Hf8ILvHnCUnNrXAem7Z2H9jPQaFrMiVM9/FhqNrZjr8LVY0iRVgl175NKrsWTz48CsbMqtrMy
mYLxpMz34xNjJvp8O6+S2dnOU1uUaY7dVkk8UUUjHHC2YSMDhinmakPXcbvoI+9DHNdLDXHHdtr0
qOJkkJfOMHcFalQ2I3UEC/zeKkQQtu/FRte3Qgyh9u6ex64Grq7/rsaYc0KAJO+Tp/EtLWMc6L8N
/eytE1vDRpAmwswykW5Yl2FDaBpccXVPYFW8AgZHxGuKNSGW/bJIylR8NZKzgk1QyWZhGXCVxrQF
XZyOTbt0SPPr4LwsZh5Jp9VNeM9ln2bbQUPQGa8CCmBc91c/kdX9NHf+T5GK/2hz5G9UeBwsPqVD
GbrejyOdy1dBdGbIsqkQDJ8nDqNBZQUWSlqaAuaWBGjXwRHbR6LFIIRZvuOYlwLFw2fCYJMy45xx
7tl9mdHD0NzLxJgG4H0neaid7yAHhExFaNhOfoJns4nEAV/le0HFRWJ0cbKR6VT+ga2eI+oGOsTN
c8FTz6xwIdMjR+lczWTr1RIJxitBTJcAFkzIR0ZxYPLhg9hDGjc87MFOjGs1l58Zh3/zSDqNduad
8M7SEU7m1wJ5BbKpngc+tBsrA7q1W1gVwERLcT/ExmaFyt40shCkOhDnJNg0mDoP4mpn/iNrarL0
3TxZ0/FNRi3re8HT/CKHOy4tsXtnNkgj6fj2mxi09ZiIUBCmn8zXABdmpaz1SlbcL0iP5OXQT+V4
4ChY2qVjog9Yc5sKoc0p6ktW5UW+gcWEBRINMKxEIVqYxRSvV6ghitAo8h7gp1DLtzt0foJDvKVr
vPIU1kkcQBIF5q9rb6WIYaSFhpkWGkLvyJTWVLtWudfa+2CqOvi9TGccxvDQ+YMFV40IcI6ZC6Zy
mh7QeMhEsiqAfWGr2e4qH9BmNwOrqQ94Fvdbz8z9eiZd0GWM7zXir4977oWdxzWQJF7VxzGTJx4n
hOJ0wT4PAdix5z7+i+96WE4ZNjrsG9Ocprr1nTM29cfmoMBuz2nQj3qsCs89G3bpggphBmVtXRTU
GJ/X3UJofOAfIH43EBnSeOUtGDcu15Tkeq28SL9WPMy/5SER/tfyAmFjXLaZOERrmSlWx9R7QxWL
aRQqRtaLiirNY42GolvkWnhtrYdXK/uZ7zi1duSfMlpSTatkLAsXw52FZdA2u0iNuzP1zL6ueeeo
2NE5nvXwNYUfQV3FMwxP0oH21J27maBg1njsaOGXpP5U3Mw0Y8Sp54JvZSgcnsPZFY6QpkDSlr/q
/SOm8RJYFS5gDu4RvTA8DJb5SardyGMNrXkmKtXt0+BYYOtujuPXNhHXkAfHE/6qSZjJiTCSUfzq
2BeBh6Qqqle/dnmCoBFDOhsjj/TIpLkzeLLQPvVVnN9lYRkLKL0IB03Xko/+h621o+Aa9Ux5EWLI
1mMs9bDtqDO+17QUIoYvunmViy2bPLQ9AA8EQnWaq4VN9cbU2cffn+/Y36x9r3txi3QFNWZ1i/F6
tHvVTbtGdtxRxrdKlhuWl1B1dYVT4Btld9JZ2PIxRXh4ljHJ08cmuirlmM9G0RoEKcqhqFN6eJ9f
R5gxejYOcYRQy+MeOMeUkM5OPWWDia7lH3Ae7fGC08YSl5EL2IujKE9jUszS719pr6dXapNqnHt+
o9VZO1FluAGiw0JcJocOICDfVWSuDdLvNp/M0CeebOaIV7IGlyczG46CRi8M65rWTXqkEnUlEgcL
aESI1D4VTPYxWGd4y6iWC9VakpVLbFg4uHkO5MnWUesUahbqPYjcJPO6+5KLX4p6bjW7Q/LaDxb4
N8FfUK/gG3wcWwIjK48JV0BDXjSuqoi2Eo4U9fexGZG70h7lbWOf4K/EdYar0TCbf2VuuOEF6ZA3
z2tHgRzNGMWAY6B22xaHWC4qtOhXiNsOMpmMnVpP1rKFShY+EG9bJ6g/uLVw70sbycX+f0m8hv03
ftsZJMyYG+XgROWaRneSgIXUim8SHtte1lsgA+dceuCvLyjNa2sX0saFgl9CPY1RRiM6sK4U/zXI
88QMVcabVB9kP8Qqw3/5aj4ljsfqT4FewHHI9MJUQWhbHvt0tzoFx7ym/tmLluR6NoPxJefc5MFi
es9X1MCKif8KqKFzVFswUpHEjPdlj7rQNNa/jO6TIpZ18DcZMK8D12hMXLiVmWhkh1WGrDv8GXGe
g3ycVdqxmsyQoJLlNrIHTYnWAmGPRR5e+qClFPFtzUX85KzJjR8Cfi9yDnWxlO55OPs6A7Bxeg1d
VdLu+t2tVuO8BvzxLqwaLoLPSW2wlcR7crnkWWm+yk9OO5LzWJ6wZvWvJjGLH7VzOwr7AjtfvA3Q
ORDj5idl+e627cL4BhnplnbL5k8J1ZAoTH+H9/SBKdjiQrPDZHiIEkEymWQF1tddvHX6uSsv2ra1
WOHTOQbg7McqTY3XIQTd29JjwgNKiuDTp5M/xXDpz4/8CkuGpDWI+PKEyU6xXjHsHBJreX+ObYnY
MY6TQL4gEM79FT1mLwPopE8FxBKDi4kL/e/VP+MsO/3pEbV7C2uXACsQbJuzlIF79o2E6Y5b2T23
AUs8sf3/+bOrXlpk03DBKn8oqzwTt2yHTDEiw1LIG4epWp4tzv4AESgZxLHy1xbooa9hNXoMhNMu
vmG2+R3SUAeLETsGNrSbg8qgobnkvJszOFhFU1GuFuDmULvSsYM7CNcVoPbo4+xKPLa/iIOmdijF
+h+OijGF7JMmCDUgxSEtDFVARjglsIH8uO3mPPMnd53/akJD+bIT1ARLjnZKoWicAKWHia34qQP8
TQ1Dd+i7zpYVR22Sci35rUKcFHKKrDBkDJLAzFG58Sbhlccf6lcq0Q849295b2XUmuddtyhgoHwX
MTymDncSm7aETUHn3u0XPukUihaoNpftsONQR22qYOo+cC1sXMWfLH2UVcn2UdipzTCbjTsOtvU3
e+d3EIVZVmpQS+8h89v21DF1fqxadTqKIiHs7SnShzPChTdI81DX0kilIqv+lcm2ad94dYpY7wc6
SgrSy15JFDgiSbS5K/WnT0zfkQzx4k4hkY+75o+8aQu1x4K5FRFCpWrUhc9ylv8WgaOXZDsHR4LC
bBHeEIemebhDiPbxSoRTyMWn3tlaH8LEImEOMhKrXtzRdsNG1toaNq2XNonQ0x5rOhlZHrg3NpMO
EhYyHYp34MWlZx199LFtxqxkC9Ky9nriUWPHfz84nBK50hAg8Qtt2hOct5n8WEZHrzv15rOUCC10
hEUjnMY08JJIJDEnz5pi1u/AZOlZow0i3SvnBLDJyttMSli3xTA2XxSVi0CrA7c+y7WF/lg8J6xt
h3MOxl5AuwyaTNx4EKjbVRhKwpcChPTfxnzDjNhTC0fRTolOYBqVQpb+A1usvsyasOtMu32B9k+v
f3/60BjfCFZCn2C8zI05rYKsankjYH99oDHawU2aC8OR6M95ZcGYzU4OhH6TdujEAc4I/oQEVMSI
QV+8hYjV1wM5waE5VCJhLR5uf62rEtw8PEYumZBKEUs/gCYPDDrMkBJfr9bic2Wp5hjapfceSGbZ
nMikNAHx3XZzu88mVIQToNCb9L9Nw08T6+3e+te0ui6pDDIRihQnLoOkxLcsTZ+vimeB1Q3lwqir
z0XSlZx1JBGt5ORgPMHSSsr1/N6WZo+1lLhY2Pc4kQPiGeSgxZMjTvkVn1yTdRRC9GeONE7/h2HX
NI3oPgjOELtJXiGETkr4/3it4ceCTtOLPfRKN1HjuKBjcGtDRIGCz6JcDl55rKuAuepGZ+RMKqyA
J/mzB0DSSof/6HeytufeatH59AOBuGkhHu0U0evZpI1gM2r1LPVnE2qqT+L0jpx9QASS/vosHkoH
xjvhj1t3yM9hRMI7OSpHWMPlih/3mTUCQn1gFqxcO9SRfjxOIMtadExRpQgW+wtCFzCMQy5Y1n8h
eTQlZ0gKnBHupZJva8vDtON+3ABFRgonzNp8qi4d+czv0o277EqghNo+1yTrEQty2tkhz9HvsiJ0
Z+mLSoKk+QOzKHbI7zL6nGKekzzxRkCkzuCiIRdtg4oPgRfF1QGkeX7UaIk883httTqsxfsFWbV4
FaNYN3GArsrc2DQ9/esx1pLUJXBuM2JfK0y6zgQP2PkEkpphVCj50pDnjwxku0ZNjDtSn7TiKJIN
XiIiqQvFQVv0NDHNkUer/a9s+IRRRqMmRb7nE7XR1Qt2mhWyL30Q1YKlzY/5SU34oxcQ6sl1gUA5
hAPB5+VVLIh4MLwLXbevi+sMEeBDpBCnr7BNoDmlSfTAqLN9KiMQOk/sbzMXuIlsGSr3sQ/IGHjj
qAn9EYo0lbcVQVFxt+KCgZ4Wmti70yu5HMNMPKjSulUUueD0LMNuXQoWUJXONKUG1TFDp8YbpJaI
JTvVnyVdUmRY4o2/j96OqAi/OmeJQ18tBVO/GNVGmc5HGV0BnI3LLKt0zFN+yNjFQzmxKxD9X2DY
VE8QvNjZ8IPgWDSPZ9Z/G5k+ZqnNbyPUwzEPu55Y4EXpg5bFEkR1YFvi6j+sCbcGwQ0JuemQJpx0
lj5Bc6Dwj5QfTLdcpbTsFwNtlIsqZDzvGgxGa2BorgTbgeiL1h1jANCN2ps2+MP6ZbfqyjjoYVIl
XSs7767cx2xN8hxtyp00XPiTrlYHHk7rVyTuDL/aJRMFFN06Pz9zJJS9s7TUMWGogm6jbIa7Yrds
S2iJsmqL4aoDiof3RmLiw4O5aI8rD27CfRRQZ4ifT40BMTdVC08FVQwQl2YxLBQDZg7XijVJONZG
7diMbr+RWhmJKYxOCcEnEMBGIdg5dTUTkwBDBJjVF0rnXb6gu3tJMcTG0qO/HkHjYpwQcX8BbpGf
nGvQW6BnIB4O0ZUsy7qtoXXRoo29RLO38Q+xGDrsinZYmHPcyb1vdw2p+v2FaFKWTcphytQFw2NF
lhksfuoUBrw6sdnNiS8hjDODY4BdyW654fHXPJnWnQSAg4NYjoTADEvwlMxZ+zX++oSsMcyW666/
wIDTXfqBoPgjHlDylxw5WKfvHugy27py9gsnsk3v8x78Pg3q07BEqbfjVlzP+ZoC7Img+7lLAW4A
ymayD3dBtVhk6QcYDrV/2YYn0gRvmU7Mx2zLGabPPeas79jTZe1gbRQcgeUrboR2BTUEekocbmoo
RqxI63Y8M3NRb0RFDzn4T6SUDBsPrOKqygkYNgRiN8IaR2a5b1WMOc7BubQy0KTWhxtbZKPC/+F3
hFTfNik/PlcPwrHg8W8AWZ8A6zoVVOG0B7exjBcENIEGqgmLW3visIiWPi90PRrN+u5VizkZkw7v
0W0Kuj64Q/0rfMfl5N/DSlAEROFwo5P1I+qUXi8DwixW2QOR47bNdaim9CTxW9cMQPRYQOmtNiGI
nHwIWdGQ1uTsbabvcthXCbYSTRNC5/edsHAvYAA4K4m0AmqqCzHrFlNwt0hftnIy/JQZI6BwR/I4
d4iA8TkCLd1yEFvrEV3h8VA9e5JWgCxZWCzRZ/TqKqarrxfoqdwXuD/rgviKreXu8246Ig+Bpy/K
rG5ePZlf+Kgi3MhJsbJhjhb1ZkGi1H8l0O81uxts2MGhhuqXIJncbfPsmkKbDN+1kECYXDBGrgMM
YJHDE50pCJeb+pfEOMhZEcLmcWvUaoRJJK+d2Q6gQeahZ9F2rvE39mamdpEb8KV1GXcKK2CNxFyP
y4GOHSQdIVlVWHgEjiWd+g21QnMU97y/jNqUhKySup1k3IhVQTUuxAJ2NilJtip3gzEBBhQFdxKa
zKzYphCDA08upXKr66G6qtUCMO6XCG/kjg5EFVl6ZGJvJPv8Wd9mlwa9RHmNz7YZCjWnAh8yw1sZ
MG2xznlW2T8yYMXVdRW4GuhpzDErsF8fhkW+xrU2qUt8bdgnnfzYRWeHvoqM2ArVnYSNR3yXIPkd
L3svKPqE3oGyL0j0lhlejFj8Sz5tNp3kdsGsJGfTlKp7zEIvWO7nfx3M0TH1G1kXoyiiy3oAmdqk
EqsW0TqUSplsCTBbtP4Ijvbq+FBssGlrEVYlrMELLO2qWZ9fBtIKSDN/Q12o/1Q6VvYPCbnp2OCK
S+rtuHw7YQci86Tc4nbyhU8++ojOonUwmhP1Uc5z6Atq9s1x2cx84UEwLmlK2Kx7jcW04tNE7Lgo
T6D/tWp4/Il4MJ855+3G9D2V5iDXn6AJ47eqX71b5UDm1YMiYYWkDNgyIRtFO0OEjLgoeIMI3f6S
4IfrSXnl6XtV5lT3orehRVWAsPHN2fybY+GdTKqWh7mmnxGfa/kFjPmUUvViBdYjF2ulqRHmTbUl
QpKIFOsFBEP2I6zHgkJR9fSQARMkx7fGzIpAHEtKlyV+b/qPIf/B9yrZqO4FVYOOE0oUdHNh4dHG
lXiWZk2YRmbhYg4lAxPoK3T2TI59HAD9bESZSKPzLgjhxTSdTxiXsF8VnYMTkxi8JNJvIqfmz5cu
afteig335UsYOkFAnVgfPaoGKCE76Y2h+DU7QKEs+qKxo8n5wZAa60Gb7U4lWumscyQw2C2974nb
YkHPu6nocCncGdHhYV4fLq0ZiHWYg/bss6IbfGODb9ixmVaPq0HobXtN2roa2r1YJw4hHS+uUwjZ
rQBlRDr09iUxIkGrgvav8xAB6j1GgC+WJ6O6ab/nmotNyIdZ6mW9chqaoEpOXjYJf+5qtpE/VvjO
EUG3uLF3omG1cQVzCeC7MIVy38dsaRSaFYqHQWCBbZRxnCXebw2wUHYZzkmGQeRLk8cJR1cjDswV
VT2kfC9k5sJptfBV5Jzbz5kgrZ8iRyfrslJ92fq7IbUHlZk6TCm5qphDTDQsal0Hd76OBwpjF+dA
sZrgbswjIF8ti16DCSOv3MGX+eYRf77uBT4OzdRkjXoUL5HqoN7/iZE/KwDgSHsuQkp8wfYnO2Bh
fsTqVedV9X3nQWhYeFRQBoMxOWFerN5ZHfQn8DMihb+Vx9pLI/9w/Qzc/f7V8PJOtPcqpSO25sOi
uRBwaTlEZRsfsHvD0noHtq9mqUZxM1JI36EOQOS3Rv/Zr8UA2DrQtNMBDktWY/63aDtvcJFIgLt9
TTIcF4C6TVR6YhD1a7A6CzwJVNPsEtU9QnpSKZ7ayd4J63lYVqEPQaZ13B4KnJXHATd+xH5a8o6a
W0zYJzIdI3F/iBcCTmiKKTR3MS9OGep6bhw2ZrkegkVeli2piW0RZoOQtlrtwDRlr6s9Wp+7lUt1
nCOn8oC/nUjbcIFs685usQkdOREdU4sNE9/B1I21de55GbmRNkerVJHM4hCv+nFd3yuyvrojvKje
xZLr0eMTAyirtVP3JFA1cG3stRMHxqqZ3C3vTz9T4A5asv8enxjzZqvLam8IvhV6T96eKwBS+WHR
1ajObwSn4F16GPEVn983lek2RS29kEMbBakLJ5GE3uk5R/18AZogqvCxz0bNKY43yZbjM7k/lv6x
HhsrYTPxeaIPIh6EVlID0fSKYKBV8J7yhW245YW9XuZJLBo0FPdyhTDCp9da8MmUOrp6QotSNDnV
r1unfW4VksTVbwrVmy9F5EVdEaSclvf3yYw8D0QSeSIDDXbjfNLSF8qmR0/VrwSFRA3OBhG8UT7T
HbRmSTEn7sG+DZc6izB4ierCTUcOr0jI04mz1B7j2rW2jRLz7UdPSmkpSmatw9igcvBmWab/tbwD
qbZ85QgN6yX6Qpcn1UMnaxSipm7V6++vzMY2n9iTQ77u0dpbImc0UhGwyXRANYH9jEeXRJVfPCeU
8YYJrYc9VLWhYoQIcqZzVmcU18SeDK6Ug4YuTuyom+Rh3iUyTQ3YynSjvrLSc745tiNfP1JX6jfS
zfP1zwUTzAvn3jHk4Ux9bDCoFR2q7eKX8xRWfj8rjo9l+7NlnqTkcjnDV1NFqjBYfCEzHiTVG7md
s+9O6/k6Zg6tuSF1zkUwrDhnHwSu/8iqzwLQ1eCdQzc1Z3AooSnmmD5fFem8Ym6yjJOd51p3qClA
2hzfF/iFwuh72zOctxBrv6Mwyv+G9NxWgP0VgmQokfItJneZ95TSk/jir53XothE0T/4DtfqCSEr
WD1JRUSWbQz7y9obEg1edJy4T5bFiJQ9WgPxWn5fmvhzFKsV2OH2BTZIxz7tn59tkJgFCzFHvZQ0
D0n/bR2rQy89js9ROFLSlDTh9TJ4r1aVr9dktvAegnIPBuLTqLwQQJzApcokCcJfavhiD8gTGwg3
hArJoRBW4JRdkc6wW1ODmaJ9MKY29wYQSo1cL5V6c4BXWZ/HKqJOL1b+eH8ZWnmL4ex4lLiwpj6G
Kv6CA0LivDh8zkCJ/za2IT0UUr5iHPPWXcShLb0qhC1HM2oyz1vhKfQwdr05xAmt3TDrlncP5kb2
+/JVdiIJVp5O6nTVdAmlyfWCusJBLXeUXWRDmDD4uOLCkn4R9+ST5ZmOlkM+/uksRneMfikzoe3l
at2TJkNQ2e8Jylt3Kud6cyRf8Gi65uQ+3i/UDMRMryqjn+sOTZ/ow+CTxKop/qelS3oit5B3WbmZ
LGYCYml3RhgfqZzMrZXzBLhH3VXnYcj54uGcQrY9z9ey36N5JqR7MMgZ7MFj+dRxVqVfLBMZlqkN
eqtfdF+nhNQtHgxVAM8aJBemcY6DF65SB/PggwtE9UHPcFojIQzFbOtHvMECMB21zc9oorqWGU7R
+B85tvi2M6MEZ4NkfMJfnKDCn4eR/zQhj1iEn6nODu1Dl4hVgr78o9G76Qsv6mmxTwLdTXd7zhpL
pOToZRY76JgjY5XlfApKlRyOL5ZcQwEshgdEiFf/DTybj8rV+2idvrwcJa9NO+f8SSlNpDJqdXcj
9EJtvcgpHdpM9Sshyr2UNF4OACRFfVO37AilI5ETbfua86244JrenF64orJW53udZpO0WFDIgQq5
qum/Q5Al/ka3MjkhuzrHm8hqUaE0TY2w9KdBVQVR9kLKyIkRf5raUa+YThre3LviEfC4B+ONfXWj
jnzpHQv8RiawtjbvrDvRiQErlMuOCx3FS+qHi/Wd5mWyAoPlr89rMXfhR+5VqWKQqDVMmH/KVZ4c
+sS9u6SBp8BFB4NF+VZmNNhS5TcYklMsgolmJIbmdokLuamupgZXzFjjM9/yQJudg2gbXW8gatLc
+okZZBB+cQnQu/xLugWB82pEiXCcbt8ciKPAVijA4+BU1rjnX8kQsNY/S5I6KYPDCOxIsBXkJbtV
JR+gN3OYeqthlT/FZPABEsqYsrSXEvRLkpkjCgntJTOPprxcjQ3M4Ps+VdiGmXdCIhUJj3Rbf0FO
D9bux3kDcJVdbaWq696cP2aXuc9vgE5rcEuYtm+EYA1+Mabe0dpUzWQ71+zAGORV0jq/8XNMI2wE
H8jVw4EFrbao+joSeBbveVHFM0VzX+Vds0Bkx8nxiCt2zIwmrPwt4lV2upCPgnu9wHnDW6IztTu6
xECPebFm1BZmNALLY+wtJHIEXnC/5DfSperRjf8zwWJ7NzStYGGHz1EmrC9smD2wpxqkgHcGTbjL
cRQ3zJE0poA/AjXjUj/tg21HERtbuqLMpfaCS24A9Of/H9Dudk7JCzt5FNNZ3BZN1cVGQHBOmx5V
SP5LXXn3LXKKtJyrA3Yghe2apa5OsAV8qJj0zrlftMb7vvvX7hz4dEFxwtfQgqFtmMcnhV0i4dC5
63UXjuL6A1euLXzZKAFUpWGlr/N/5o349PjZ55vyPA+XI6PsDEApYOSd8tmJdKGi4X9vD/+2VN2P
QjJlCc022pEd7CrX0l4ResyxIMP0uBY0P2/AQ7TM9FiCVXslVejUQFVWzdwglW3lRjdg1HTat52h
oRFu/3vuwcnOzMQS6vxL3YRTjaRz5FG/iXvrEmZlJEjZwO7JpEurp0qQDiOSiwCNp3vHY3z3wweL
ZIRjpnLhkJ+QQBMODCjYDdj/qy8zDe7aGGKyBvV4jwnBbLfG8NzkdmUZ8EKA3VQNCJqmazT5K1Tw
eB6t9ufnSXdsy2ofTZojcKFWA9oyU4sXfbx3qR6hKHcuNgff2lskEtfDgvlAtTGTnYFrr8PIes/E
SAXtGtPM9lciGDIp7TjagbO2fzBwYofZIGySfnTljLRyew9BdEjmiHkrfAo0xQRodRfNIo1hb2Bw
yvfQc9/YiEGihDVODT2eErxcAq31NOL/m1DlD2R5+LBJI8Ip7gmluu17DUVWJgyddt4bRJOOnL7a
V9yC5D3G1ovV2656wAMlfSchh0XBVoOH0cFBSv/z1V9Khjp3oHYniDh5uynlSwBbiYAJXH9ltTdW
P2RANyNuekhTyeAGFUSSHfq0v1ovuRxZ3NFgpu9u4hhTWLx++PAo4G+EMczWdG5mLMrNRl24hS3x
8Kyp5r5uypvYsAwdfazxUxlBg9nPAF9Ox0PAU3zBPXoNYsvaUkYiS/x8U9fc/ZM4q3t8p+P4rBpI
Z+SgaLsOqH95dW/xEYFmZgHdzL39R3R0fksdA7fIR/Bl1mQU6aljaAYjvsOtp510QO5IaMcHqXGB
Rs3smsYL5Kb62sAc9Vt4jANbR8Z672kwhUy+qlI83dFI/132jZ4glh5XzBpkZbkYQ8BfLgb4KuMi
s3LX8vKm1OrLjSOtndJHU6J0MndEoiiO7CEfL6/07E6vhEu6McO50+M9WCNrumK6ZddEaDembaRT
gwIBYge+HR10W45DNMYK+6FwNNBVsA8dAlVGRIlGkQA+jGWm2hhd2igpkLhKiFuQlycw/BN+97QK
45M9nmiEM3e2fx9aBy9cl5afBCEF4F88DsZnGjkIIynbV8bYolMu2jNJBR87b5FxAvhGp1qR5pY7
uomnUB7tOp+HIWPbVNo4SygnUvTVp4lnCDUkeKjhGJMkTFppHHAUiDqlAPdniBh17MhOq0QGuaXC
HdVQdKKSJZlC0BHMrZURl41kKve4E8Mt38ZE21vTvrPygl/6PaDu4EqwU9rByjJl98FI9HmC1dfm
hoKC9owXFq7cTOIFcbkQImtZHyXSgdn7aVLooJSTHV2n3f7ALH+3Ua2pdNrBCGrFm/ohVa/9RSBu
73o454R8Q1lkUwpmWkuihE/Roc9QoYnz/7GQYydXRpDb1sjuZ339eGbKTFH1KQa1RTdDz1l8rzpW
GA9Lp3SNQBBapTQuJt8oHZ7Zu/dI+wR8NDdweRcXkhHpRdDELVcxcZn4zsVuqAAYnS4IwCrQ+efo
x/XyCABNmb8XZSGF0ULzoZZQHF5CXLKNxIyutccSDKjpunxjR/ZLhm3CVuPSoi1xvFAL+KaLHzzm
0arDkmLnu2oHYRx4d0ZoKmLgeTLZUJwGXhylwrke6vT0mCDrB8xQyAsySEHKzgAXfluiF9qcj3dw
StRoLbON6IDJGRURkl/AuchIbU5XQ7PADUagmlKdaQ8SgxlH8Awb05qVNb2UguSPsi/ppA5HI9UX
3tH0efGN4AoYjLRFiQ04RpNN/AVDn1zfUXdlzaaIoE4yInlH4BFaAIvuz/KZX+1H5gpOKMlFvXb+
WlmqI50fILkdy1iwUfNXmu8V34BsG6Z/G0wTUBf9pZ8REoQvbL+nEMLCWChuoyPIdo61PZdL4+b8
tATjj/ENU8dfZn8FSjuWYGvPMcgYFZHyKAfgtR/s0OZKGkaR93fx4aT2PrYWoeBN3FV3XCHJTs/U
d8dmZDnry1yEr5d7hc4ER2fyv8C0/v7iLkUI+eJI25mQzSQ/K0PDbzfX+rY6SgEN2MH1xBjcRw5K
7yFcUBLZXJHUXjeHK2ts4ePeV5Li5XAwhhQa+YrTEQLF29E1W3ALpwqzzDdAOR2dg+fzqVzDQvI6
7ydbly2A2vXiQKN0Fef+lFcH2AxrIUJnrJP/RrHUx2LNI97edvm4qkp7R5qzCbjdoDpQBeUaJGum
pWliF+1RExbXLukaT2nfBdXSTaT1Kv34eTORz6cA/iwmxhXXthZrCIfaePdF5p++neLpgC/339so
1hjugC7nPo6rGzDP+mKjSn3K6P8G5i29SAnmfhlApx520jzex11RFgZqZYN7pfzlfG9B2vRG08Dh
D6eMfFXCMtn6cYQQP0wJ9bXYb1FqKBH1Qyv1WtI28DSyKXBvh9ekhjff1TY3DU5cssCKpugwuM3G
Qfd4BafXUtMZiuzQi/lST/4N8bZH7w+L/L400toL+q5d7YsA5uzFseymz0HsJIZT0+LNV4t1mDYL
ULTrt6S7Pd9fL/0HatRlxh2vm+SAfk2iP5EgiXL9XcBoWsQOtuIs26gKS28gpIuxIirHJZi+wuzd
UyXRZyCYMwBoraNg/bx0I1hIs80mhNBIF+5khzuUZtL9Qu5ZSZ+cc6WhKY2jtHqMb3IFdjDWAnXn
bcHl4bVy16dTEin5OREhqP2XoXIFZuXP2QISdNuSI83PB9VTa7wWPEe863clw0sRElZU2KE90NNd
PSbQqy5/9qS4cHIYUYfNPav+GokuJeLZ/dDug76SlNmhDhNa8HHCV89eyHl8+mgJPsv9hQqtqIHR
Dsu02obAwoj670BpIhOCYIZpxYRNWKKxHK4yyYJW2bpozV3Rcd07o4K9fFoT0Jpy1KuK4y2xtjCB
jZhFPgN1TikBtJ3gNUreOvOPJEf6kWm4QQ6gifZBx4G2mFchqb+NynaTjv70ZEuJOvK0rcRq9k4q
BaOHrpTMu68Tl5RtejMYhyoI5UjrA2ibhs1rmz/LETFLK7oGEJbpcHIZapVEjpkDKhjz5jUZqFXE
qzza0rNdnyGNJ02xbP7Sn56oF30mUKDurAsxI9CL7VBqkl/TzpuwGAKD+e6bUtQ+27XPF4ZrHxmp
V0oLUxXUVoc9zn/61o2KWYe8DBgI/83NFGxUROGegTATORK55NpO0YE+YBT3CY+Wud2MVMv3j03i
GrEHLR9QHRX3J3Z04PS3MnUKb20NbWDCEWVwZKN01WaXBENkvvWAYENKgvQ7v31ihSBUOlF3vCm5
wj9WZ0evYW/SZklAzAjCUBMb9aDD0CBDYvwKB/BiB6w7hLUfoY/A/sXw/OLwO+lknIoyn1/uVRAU
7XVZnq+hF6LdPoz/BcHGSt1uIvoVabbGalNPIybLrrqdrkEZZEwbIaXvXz9JmDp8MaR4Dn/aFFic
jLyozwQ65JdccWucxiXlZ7rN/DYKyupW4x78JJSTXIKXkwfLbH6eXsdY4QXKmhfeVnp51L5uDdAH
wwi0SQ2wyMKBcwxIdec67HybOioSz0OViYgSpGLezAT80+q0QfPAiyTPuR7TmkgloUh5GqUauoz/
sjqDPYbzJerES5jK+IY8NGNXy/fsks+DDIlI37tmJ+46Pk/3ekHzZTSv6dI+bq+IQt/jFxxjUaEs
+y3OD3ZzuRiCuMpbSLxJmCBcQBC8boL4NLNP3u1g3o2WtJvhjjCD9nUzI7NwcZyr4xQz3lQGcyq4
ISfYdKrTJHqMCDAc1tRf3qHYnk98V9/PlZTJhVaaPv5f+pDaHO7JizhbspMZHhjRlzEPOOh90sFE
fjRpaWtne38s/gSPJcYLccWB1PYpePtIOjsvTy7vEkSYBN68aTdcKgVV5fSaTUQJK0V3CiT4vbrp
AGmIyv+eKPqEHsvdGChgaN1JnhBv2aMChgDpTCB0SjntXfp38Ta0veQkvz0Lp1cQYktl4VouIpUB
t0YydvvBBryQSHAk6b21fPkwrm+iyQc2aYzTbM2lKabwLoixTJkNZnYDDF1lyve+QXn4/wKVtS1p
eLwTgJZrB/LSf3eGHYs45fgTMm6FyzKvFqV8UpE7dQellaYbuAj7/lnXhmH5hOd/VBHJZgrH1P9R
iLRGKjNIPBq/tRGO3RzU3mRj5y+hiYjd6Hzn4R8DjgeVjLBAT+2gn3YKKSh2dtRN2NnqxHyMKivM
i0LN7DCblOtly8HdTQXxX2F4tyOM2Y7Nauy5qaA/4QwukFnTcU6FwcwszNz9O6tThlN3VtfjWXjx
pIelQvfWNrBNAOeupOQNyJFtvwKghyyqmzDHz5SSMNA85ryDquFpkmSlu8GF14MJd6Hs7PzFoR9r
Kv3KcVXWFFsSqZIrUDS/rG+TvOvM2coCV+WfRQUi2PcJmYTxwR5h9R4cO8bd0MP6SyEEOlwg40Qa
toW5olDmzqDMmGoG/cnKOZkk9LaCdOcqg/cRRtqk4/Al+maa9AoB0O3PEQp7RMs+Z9ybcYOEpPmc
R2AjwvPresjEaJ4UY59m0ac1xfuo2Qq5YtEVM3hA2URTKbZ4nFeqW1Wo2/Uzy9jWjtVYmYn2SRZP
HlzdY7dzd0kpxHat38TioOa9JccICNtsv1byRWm72dulF3rEDpUQNhFPuLQt/B9J25jtUCsT8hFU
Y6I8jrN72qdc0S+5nGKCjE4G7V7rIwRVw1WubJ6mTT9H3u2JZJeI7m46+KghgYv7LH4C2ZbHocL/
kgunEHSnS0OF/tHp8a8L4nUHMUV5b69JlouEo2Irgy58vmynQx1jWshn/A1PLK9HHk182zlVOgQk
cu1B7lxwq54zE34CD0nfJ2QNDSbGPyf9m5hWyewdCPxlFEGr8kst0VzsDCLIJlzClii/gdXAof4J
Hji1yh6NsqAnCU2j80GhhqpWDeR9O4/CzFHaEu1JZDKU/UvZB9G68cWkK26hv+Su/aUnvmLkyzBg
hiWDVF4MyBTJZamEclOKgoA+r7oOiR01oax2FkeSXTYRhh/escg5gIwCpRqXQCrgaD0mT2YDfFbJ
RgQnDevoaw7ZRvHzMr3/WCSzdP5nruk/ssbYKFnzbKe48ktEII7kOlqkhdtWmcgMJ75SuNCj9hqZ
+3lsiJFcfgzmKKHSWXsSeIDah/dph1UWX8zirabJx+j5ySHe2BLGIs2i5KtIJCCiQi+3J1MQwGSp
ZFljp+4BK2+DptNCNbLwAbLPTeKWo8+9fO4AvW39gcSkOBVcxK3n7ykmo7d+4H8wnRVhv0fh61eT
exJe86IXp2nCfa/Bk0Bx5l4axfxXJYUKvW0AluKY4gD9cAzoi5IVZygJ367K21LP8Cyuh4Fimsg6
8uOErZ5PtrchaK3X3qg8BcuKE2ENpjAKJxc2IfMNfe8IksJ68p3cmIzTyOf9I9PwuJBesb1gtf/1
EenQxTgpON3XYbxnsUQtVgyrGdHNnhGX8zHcuxsT7BX6o+jRQTevqjwj3hkqtAmDuBNOYsX+/Pte
0D15X74NZ2LtiRoJITYzRf3MZwir+88CvWL/mujUtFtsBpidw3lejv4DaTpZ6vnfBwjW9hXPvbkD
cTbdnIjVADuJMuXujFDw6M2JBcXo+cbak0DhcTH2Dl8IMAmmKNF+FbSGoyPWGK9OJ7yEzGuYjslV
8y5xPGLn4YOhyR3zRZ/0oRFQWYGh51fQ/RO5sQTrjC53SXDYUBz5Q1EcepwBQVF0A+bJBMFRlBRQ
4GQF3oAbGnL8HktbYMDqDYOIz4D2XS9oHTYveVrkqwB1SghR3zK0vekoQlkRq4JqW6XKXIvRskpf
vvED9YXSRRXA+yIwcmL7knI5ghoUKvlGmRisa+T0WAKOLgzX5ZCWonOT4E7mvo8MgoMDJD01OjGB
1zkgkg6zg1t85cOHFADY9pko+LNPmMEKSPMecUc+pIP+Ar/LVuLnIUNAjnRjQwHLyacx7sdzRGlW
dlrW417xLOV4/erEZ49Yp5yxn2XEf+B1CHwakcb4qzGBC8PaZ0C7lwKtX9nP25sMKERrI+f8/PPl
8wxO69tpo2uAdtbmuMRnC9C266PPAXsCFdxzpOe22WszbOJQkB7dpgyaRdh71kk2QEcaCD0tZ2Ic
Kz/iXqvG6cHIT7z/RJnled3p32uoHCnGqPlKyE8AIVNAAyhcSzgrWq67ObFCKPwgwo2MZfORk1L/
YH1YKD5PaaBdbodMxG7e4DSHGER4GsL1j6wyVcole3L4czaZ/zmaX4UWLAY3bpCqI4FmS2g2zb2l
TG5ar0lsE/th4vYBTVRgaGxCtIaMfJ/XpPIpapt/cg7RrlE6KMSbgAcebGrFfteOIyFm1FJQsKQT
A1haphXkRsuzXrK8orJeOnb/FoG8sak9pDzgPJ+FevfqH4bwNtJYPdblEyv1xRcgVknpN24G4Tts
35SwFd9xVtBr2psJPL6zMkB8gpwaDyyzW0dDPFR7GbrPJ3SHMTqHrDb/wEI13UUwhJQY2fTLbD7y
WRnNmibEz/42s3vChd8U9Q3KYC+nQqbtQq06tlrU0l13TVWryoHJBGwpwT3Y9LsA9DCaUEQ93I1T
xJYeU1leYEISq7CEJh7FrVGd0VAPqBn9gbB3blDcjk7LxwCoAJChO+bFj3TR4YcR7gDNt0lt+/nj
l6rAzVQFOS8imu5xGwr/ZjV2Gt0afG9O0RRqd/TTesny/Sm21WekBLacBJPkzjN4ZwhuKVUFrN8C
T1uICYx+jxqYE1x5xJcbVOW38FezJ03YuyHhp56m915zsRJv7QFycYgoM0J5CCBQ93CeNC3+omNV
v1sri37cFEDkMnyIfhk8tn5zM+jSnnnK1/dkqWGzZr5lXaaLYNxm5TwqT81HMua/rw/cf3+TzT5c
+5inK5Q7sDfzHFmKRDAalSPgO1qjJRAi36UOtyNNxhD7dPfWoViYlfzEnrQZ08WGX75f3en7zNfl
43L5jOWcay+B+Inr+6STeoyw3vYRtiRdZt4Aomq8ZCsWZ0ec2tl3o/P7qRszxj6P05YSAETVb12H
DLu5hwczirnNJrKZ3P55tgBKp9glPgMG1fLV++gqA7pnVr7JiH+bdeFebtM1HKj7zTAhs3ZW+tlH
5UNmu42Q82sE8mhWy27Tq2RFIwH/t82tzwW3Gvhv4zTDImCZCixaZ/6KnxR4D0m/LHcW/1uOjPpS
ETzKXHEfn46QQFJJ6QNB66j2ac+t9zrcro23dqV2ev55EWPRV/Pb4ToEe3Fngr9Fh+BH6RSg19sn
fIMsirYEUJMhrpqBgRT8bT7Cqntk7VWwcZZ+j7IA5mZBdzxs8gNy6El7vRM+v6PWNaCKecdVS2EM
tjF0pydB8pqKVw9HzCGEa2NJpWHPFMYtStSbxpoxpPJoweD9lZTgXwYabwOH2oJJh/3s4sxdoaC0
+ND02xEG7RINlSU6cFlhZUc+TbeEKF1cnVMyoi3yeMRxdb3kwSN79th/CpJmaka0hjSCDCbcaW38
0FTwqxfoOVJG+N7uhjux7qqs7klbynD2GY+Iylaf+WwyvFT2ge/BJaz01FUJrfMsHLZzI0Q8DJ/4
3IEw46Ow3+h4CnShdxp26HNyh2gBdbVThOj8p1vb7ZwvHm8JMoFIqh34sUcud6uXtJ/jHWwTcu5W
o4nunfTXh1dt21y9D/Eku0nE+oNyCTdxKsCWhMPsvGOAvnrWdE8/fjJJLG7K3bbjPqM+CYVyivq2
pI2HwH4ZSyA+FZqVgx1NNjDtQ3XL9UhyXRqtb9cf/yagMCL9NxcONrjFEnQZ0OOfLcgTuF01xX5o
RMg9NcU88ScN3jPeE8WOx3HwbFehJzp0sBv4E8J3RSDXFUP+1zar2S0LsoX37vjohf4whglCnfwe
bbdfWBL51TnPimK8wfP3mYEo+Byn7Daj14Sk32sAEDHHocuH3gfiPB+IM0gI3vPSAGuG70YBXRkb
rG2t4LNhXDEJUz+l+KAn/2IT3V8EiamEewVdvox5RoXUSw7ZOB1dGjfi9fgGpeiSSob/ujtq9J71
B+GzJQwpkAb/+CnXIqK0WvTaeCMl0GNbPanz9QkPqQZoKf0UAAoSYJhFn4Cbdtix9/HIH0AGC6nx
GiWCdWO2sA0wpaRYpBObUUEGEWoF0dSvIrigRHel3lu/4kYwCQosm83XFOxblB6xLBsf8aKUj7PP
Tg8bWSE9OIZBoPKCw3edxq6s3nPsvDlga816iilUk7W9ia8vQmhQTVQR4PqcAcibNktog2woWhIV
n9GHh77kDU1IXaDnMCEOl6rfDaCSL2eH8xt/GgZjE/x/VroQyWz98nAdTrhC/HgK04/POnA1B0bZ
S/YWT3fwdZqoHIUJPOB/Y706RbDPZi+/VICemTF3iNfX1+r9b+g2gqFxwmJ/XTgrA8eljOEg1SY6
KSgZtQhdkOWuO3m51KLXwijR/QARIuUCtAFzB09bUySI4J0g7h1EPr3JF6QDq0dO0yDka0Dozhyc
nHJEmxd4lzFy8OJ0j9mDN2Ly5H7gSwXhUISUOW6Ke8JDH1FJnrpfl5S6UMOd8tVgXkasEW/7UPns
IeQQx7/ahHjNUWGpRPGvmVxKGWjqV+efqGWQMzPOKvhj9z5b4hlwoJySGTgn0x0Vr34H0SVTr+YN
oEU1B7rfyiLB4O0H6VLWDeS0NiqnFsuv9sFWx8FzS0XaiVNPCcYUIf/ukYIdtL8Fq++flL7nJtAh
0DkfBPFjGE7M/ziUbwipH09R3XY+ZvPLfvaVEJhPIKnvaM6jxypeObT3+QNAdUkmpD6liGcDJFm7
t2IoC1dS4XG3n5MoDJWCthp6DDN7nZZsbxgy1wC6Kn0BNcLmcMSQVDl0kMGw4Qu1w9wXGtUStmY9
kWzKUDQst6Xd3cFN4GlznxjoDtNH3gb6aT2FNaNnEQRHOGaiE+264OAKpge1abx9DJtriiJtNCey
/Vrj1Kt+kF6w7dLfOxvO368U3KOYxicU5dH67hYcOQGTscDBG27xFLD4OeL5j2x2D1v9oKmNQAmF
QBjr0d7OVsi7NyoVfZabiyTalkUZmhO8fa6vjOTE9kLUU72EON3hfZENhba5yNtNU0o7TB141Ijt
97R7AalEgsxD0hFfWzTfpzdyv1E6KvrQPbw8vPJH2MPtWC01lP4R2FlGOabz55Psa3T8svFn+qb5
+bfUdSSsjtcJjgPvNCYrdDjcONat2gbK5294Ku8Q2ugm/mYvgFffBGz0pXOJsY91cNIJLCbe5hMF
APP/DOSqOOpjxVGYFAxIGtbbgoas4c+4q4Sf0aY1FSwf9FQFiwTJdtusF7wuej0oQdWO9YFwML34
kPrKFDBW8ov28IN0N1inISgLAxC/7PGoQhCyUMP/pSEyI1WHRVcoqJz6WciX+LCCIsEDpPnoExi7
fLGmIEEEFfcoID1VAK68ZKnNS60GCNg8A+ggTGd/ne8Q8K+lo8B+5Evcg3VIF31WzkRP7b9ex4MN
3tKfG1N1m9bLgmcCLFtc4kzEl5QUTseuwuMAW1DqGImck7vSaY23v50XZf7NlgMDSL8yQex/AzJV
LwOcGgKFFIYQJGaLdjIMYxR/JsanDdhei3Z+nlPop2JUemhtXgde8cFBHJnsHmPOP3mbzwO8ch0S
yXyBKRyeCi35PZn1al1qvmW9BGlO4Je2kwYqbp62wqUqQ4oYHlhEHQk28ClSxmU5Q1R5UMe6+sl2
XdJbtjISvIAmPzlNbVdht2L0da2GP+4hBMWsPgZw3BQZL9K8fLJF2wdAVY7HbJvUrgfSDRouDCMv
yS6/4KRmNeEFenC0+iJ/4ok6Kn748zzg7Mxff/b7eb4qqaZwZeoOGSclSKVBG5vIGpcvcvAL4JFE
UpVLOUN9XFSjUwgc0bNBiSwYyqrjbahOnrh2KtpTZsKpvhC5/BkKX8pnGKr7599eTKV699wM5V2l
2ipwggdLd03UyvOpTba8y6vGNF5377NVO8OJtPiCcO3Jf4yJMlRs+mLB6DuhXE8eIG22MwSipZIe
HRIHwmP2tlT67gL3nEym8MLRHnPzpwxOBJMxT+7v3cZ8BoezCmJb9efuwbV0DXTG9cvbu5oZkqKy
jPysnfaUO+7gYPwwQpXUyNCYaeelsuJ6q5TilIXqNH5J7qcfqSSn9f2D9ldbUuV0OPmB5cYSrDyU
qIAu1NXXLMqJ5tA2ZzAD9uhOKCx4wH1HFMY6xGlrsS+/gF5iPjU/TjgmvbUXJJ3Ba5q7pqDhTbOa
Q//BnEeFUcwN5LWp1/ZZTXEWmLtvgjN6o+A+Vci5PE+hOlYBVTVY8bstsZWVzauE0hPk0Akr9W9x
EvJ7kmc6YR4mz8Hjv1CY1C1PpdEGTyIDN9qZWJHWJvQOsgi5RGk1ilRke8Ct481f2ar9spGQIZR7
CyfKm6zRoiqeVKRQPC4GbTsqTh0px1/CHccOWKDptxSf2WV9na6l7Oe2+FNlo3DPx+4B6JGEkiYU
mP8Milam71UywVbDIarhS2x14s1J8mW8VDWRm+Mn3bapNQ3lPpDUZkS8Sb4sMidKal2l+xluFvxS
z6gNzsi1iKmlfl/O4zYbrbBMexJ5sq/WTMjJ6LeDZ3yHNVCmxgukOQeTL/NTL+guFelHt9QEw4Gf
FRrA/zna+bcciKfSRfaAkXR7QPGvkshC+nkUSlsuCtvlGlrypmib+eqW0EBoNV5RYxlV10i1uXen
9aZNBgEj1Qec9kYzs01dME7r1nD3mO01pPpONy0sOFBpUMsd33lK0p0+d2HxoLhPbvi71cdIcQme
Zh1S2ze6qPk1CSj3puYy7CkXWX+NwRMUqLUSPgwo9kLA+NJwBtaH/bVEus+xqT0Iv0F2JyKz7Zy0
F+imeGwTkZQMVWz5gt4UTSOwclPmjqFNtsPJ2madOAJSQ8HlfuYNX20HoCtheBeC7eH92tSHYEzB
kCqQvJG+v8w+D3zqtvwK2QvTwXxRCrf0C2UVw9e7nqffb2uosaSF25ZdQ/KOOxCmrtfyrcg7ynfF
CM+nmUu7uNP/oqaWGwwl2AloM9hxEmfVwOr9/N9UWxPNg4JTprf8RltTBCgjL38ZY96GzHGVPYj6
nyUOZBOxmQNUqwXzM/1CdZ9Cr+O92M24A2/QO4GjICjXV91GTsB/dF8sB4WC3yUi85jTLxSWRi33
rQRxFFkGFndFCIDcpDX2wt5oPjukt7tZZTodDSKLheCfZHsymNdKNYnAILgZX1K1sfqsSCQ3rsay
1SE4Aao16bZbCbuGyBCdGLsSLJesNPqRDgY7ZdKAjqDh5n/JS3s+fpacIW5AnKizByp+nqQLVfw9
IyiNjvTywUxEefKI35KRcQ3bEfw3gwNQdfOztq5mA2LWW8obJ3FXA8HfI64DUHcXX/prOe9d0zS+
jyKE9v/kEToELM3TrO5g9NkkYoz1TmtLCf3i63x942lkxftorjLtLZB6cixot30rUsCXR3XvYuUL
yH/UZGnKPYE6KJkEmkRkWtvqkh7NP1DZ9zVNuCUaCzRM2arny1H9nD1bt97FI81U+rcd3X5nnW38
P7e9GxIVKdaD+sbK2iuFzXAWT5cO4bgAG6AETnNgp3ug7dYri2bxcX2+8Va3ozG2JDBtWbAYq6az
JxlyMLwJ6cp3ie/g8ly/OfGmazfSZJ7nv4unjfm6EEVKjQ7cEfID+MgaaJ7jcNhodA3FLmTg7F+Q
KMEw537exxFyaY35iG7SfU99EDwxsbUd5bR4VQkAq5mSGXBpmzPMm+ECUeAcOp9/zNbDgLRj6n5u
CSEIV64QuyuNTtXGtJ2MjJ1v0aJ4AXYR55YO4ThNqqoAqDN0KwIRxwBJMR40OBf02SoHv0ZFkwb5
crcaVadKyPFEdJJ7gsFan6jdwog3+qFjzQH14z9ISnwTdY5+2BSm6OdPT5ZJWXosXLK2rh7iABOA
oYElkFbn51ab42r5TlAsrUShItU4znb8lDfF218BEorU82Jt1jvfSHCwbL06f5PjC3yznDoXe5Nl
cA1K4dqM16lyFcwnvk7/n+vdmF8pfmytovLPCSfqZewEVxoopby9+ZUiULltuHwMaDiwK6X2+i+e
7sl/kjv68sB8LRSct+vBBJwQasuiu7fidVACFiBRxy+9tfP/GmGYI/dDonPasKs0tzeSx3MmWYHn
BgMptdMMtz8hsU1VOG6tLWDkGzzsDIUIc9TylJLtnyYTNNhp96UIGidLQb/d9P+CEVCiB/RM59X/
aBn/pPPDJ/8I0XGqf6ecr5nDHstIpDlBBDLPT1PVBP9SZo6D1BhvLnIlOlTvUK/kI+xHMWcXf7f7
le1lj2ftQnrZr07uZa+v8korAJlG1fDAHOD4Q75xyrNQ3vPXdI9g7BxdlGU8TNBaW8npC+5pLcD1
tFT29J+Iqzv2x219/8WASDBx5GfZ1Xx6rec5+NOfC6eeO6eCybYK+mPa6sd9jcOODKjsiD08159s
oavrKoypHRMC5P9ZeoDDA5ak8XiikT9bIsi2Ok8/HXnZlO1OlBwCAYyhSPtuB/lVqzWx3tvkjSYX
xF4dqMu1RGYWsjnvHuLPUyekVWj5L02WVfpAqbsmBM4qcV5aaJKSkp2phZfYffHYVoT2ynGafSSJ
F3umwuDPi0uQ6PWbqm4xEX+lqYdfYLkQjdY2mcvkbiY0UN20BUHzubBLmTikVXoFwYPgMFC7wppV
tKhiY9uncXoXzoBVkl77a0wvDTBYkoU/jAtOEprbaYK2xHAA1+j4E75XAms9upSZ8Vn9b8sE7KVD
3W60iB8ZVLKIGFgi0KvVDpdqYrl5kZLyiWTz8PYN7xfUOrK5Z3iOnPYyG/cTIHfU9CakGCL0/A1c
R/hJVhD+xBi0DFkEx5ioWmJfT5aV5cuYDj/5OLy+enYloMUS5NtuE8PoWY20H5KLGw3qz/xy0xKH
E7+zyZUIK7+jnZRKDQLfMjLkcNtkGkrI3f9xgLFw+KOZCVxa6QzcmZoLBF1Iyrm16/9UFhDs9c+x
wUlP0/nXq7ivDFBXWUqF+ZK6h5WNPLOycwBtXlT+kyrzxkuJku4C+YSvOgM8j16vXvEa8loinOqU
cTwcwd/8h2LAFFczlAjLCScD+OTKBvMwrcMZnQKdbUF4IrXQVljgCdG9A0ph0iZwj8icdfpikT2a
hdDC8yBfQYnZGhgYS2Mq6fYQ34h8ULqhKVIB4IYS7r3UaKrqo4Sx9/aM+GDFZ3DKT59WSdd18wm/
L6PerdItvk1/44obusberv5911FOP4MKutd8yzIG6gWn+oRtOcEuB9uhya00FWiHg6o3llrjEgiZ
3EY1JuDs5StQyfvus48aGQwrAJ0ReEpPEH22VFYkh0jGitnaSPT/zDCwe5RKa4OTgsaiLS8dCC4Q
Wv8xYg0CT8cYliW/WJpLYmo5DnIXZ4juKCXMfYZP/IeBgsowG9/fuUr3CqKEerQ3Cumwl+zZUGsI
Xj9GPQ0Iaatqu7/Odqf2aAPfubJ5WUKImyNulZUT1yxJtLDOmtZ+xuPw4T1Rfm+pwpmXoo6v1jCW
Vp5JKNKjrVI9MAnW9zhObNLYOi0vcJgQIBa1ELJaDgTV6O6L2N3swpvxBCC517tD/vWGCw0oKEIh
+BGyiB3roLLBwASoKq3tnIMAUIB0TaRkxd/pB9bRUl+qzjQ98D5X0SobXM7OzIp43L7KDhgztWta
4KvTCHmKCahAKcrCbLZdd9t/Ue931X/9xS05nSdvdAG72/g6LPJTXmobprQQkTrL4LFuDfEZFZo8
DW39sW/iQQAVANNuNQRyus4JTTkzi3Lr3gJwb79Dao0Q9bBeCDKvknwM1okA+GWbsdFINTxWGO4Q
hUOQm2zmR86OaQytg4iKnHXD2acbpWmF1H5mUdPiLTDIoCUTTyrsHy6nl4peMIXTdKT+D3/vNmzh
YA5Mt6tVslLCLg74vJeAAvfJ52t4S0179UMVex9C4GcaVJIMARHZLaS7+XXUDS/wIaaOqco4ERfA
xjz+zCKudGGZRuJQQho0wcLaDFg5l9f6QEARDgGnfRMYMjkz4BugOdulregcivUV91PYe4iHkt0F
5fV04vzGIKh0SHF3PF9poALIlXW4QRQExeg8RNq3bh0iRhY2PJvi2NFWHzjfe+Avq6+opq/VFj/6
aTIkem7PPwS75yt///aLHVFmrfQj8tB+RwQ7veKc+WgWaTbPJ6Mgz0oYDSizN+gzU18G/9gJrfGP
mCEj1jjLAadDQJjIjXjBgBgjHF5Lqd1hHu3TPiQTibecY1oRVl/Xn2jOBvS1FrV3KVjeMPHHV9V9
sXbIx7aD7FcQ496UuhMnbrLE4XF1rkuf2VDLMhMbvSA465zBCC48CfNgUhLKXuYmPGGImjRq+nKj
/ekGP/s0f+7AzdLAtIGOB5jmRCdsrReT+B8zDe7slCXxy5QGeoen4StOCQqtTGFgtM+Gaha+K0Ld
i91l+Nn6iyQhCUGj1ZIQMIWerg1TT5EKyEOhOWQT1C2+xs2nixwnV0mXlTtMP62vJj1KDhsREIPs
qC+AN+bu5dTuYQiE6FiA5re6+VxNOirDTA34an3ExCmERQ3m5wjsrn33NLj5Zijv+rxfRURbXn76
lE4UPdkSpcYDMqEid/nFBnSFotoinl0Uh3wZr8F4+qwfRqZIcZ9p0BR2bDOlrHXnTTncJo/AUPnz
bMgbyQPBuaR7A4Ho/mmTOfnVu/lrC06moyJBCZtW3q3B1DrcEUqLjLDzzmLqPDj+BkxOcico79FG
hR686MABQvvz26QSmKQQWHpa1eeDPcOE2peACuNkf6ZbfoAkSKnqkBwrRUZox+ZoFXhZs1q6rdlJ
McJW+Dbj6zF8YGusaH0slrmUpD+cvUvgrM7A2DxqNXqLhhUWWhqmNmas2CtNqxSEAxsipPTqqy4x
hAMRFLoHqm3Uzw30t9ae3g2VGkbjx/XHWGGrkZfpa0Pkign4yUcy6hf+z8Ral5eswSIWIusoVbxu
XKxw8uG/MqEqKQ77OwW6w2pKDQgo1qcqBZLom80pYRYrWxqau7N8jSqnaCpiatDgOZBOs5Y1HBfY
U9Ny2FYbOUo9QrkViVSu5H7ECCDY2/vrCB721tm0HRFxHvxBlxqZirJop/7+tBXQo0H2vXnUlrEw
Tdy4PM/7pOmU1smF4uEZParS2+0Y7M7dmzGDH8yT3CW4NLcr8nu2MymqswHYkcfgRtziDPLi7+Mx
Qgm1ef71XUFH4fglXKUqbNaiCnycwiiNfaTB6dOX4MD8I6zBXu8vn4LsUDm/sT6BzCO2pPiNQpPC
hgjcknPCzzFIhv86kHFe0+cFQGNedh4/gjyA1N1iVdzCVJWCPslAv3xeKKvmvrNXHPaINAfCC6xR
XgggYPqX8jEG8GbFT3DBya8J3lLamNIoggbNXckprTCLa6VMCgWucghdKZkB+GaPUpXYWXFPzQXw
NH1OUSzEU6EWrlvp3EPWWi2d+9QBprO2d2RXeIr9BxSKfDR57mzBrn+tQT8yzaY7Y/RJrkDNNzwB
gPQaQwq8j0hfRjbXi32pvtB96CiwT+59s79cYfB7P9Pw1FywU9huWj0yGkHiz9/oIzsEtIpJT4f6
7dDXmg1+tJPWz2niUG7v72OnBk1P5Kvlj3CuFeeB9w/GxEjSZZqPp8j0yNNg/Rzvu9d0NqqDopoH
yl4zFtZAqJjXQYySm10OFHEVDtDnsCWuEhCk6UmCju5Q0R87CGlgzuzEu4US+ucY0lMtV9yb8r5V
tLxjOtR80WL3w0u9GTrNOVbqTttYgFOuxGJtBP7aC16RuVi5ePsrClpSvIpMdZgG8BzPCILFmEjR
yM18OCYaGjpzTr47hwrkZO45po0qvGKBc+USU2xuEHKnWFuqKOc5pkkdfuCW7bc8GLk2EgsrZrMk
MVR/JNXlgJObR5hHknQWV3IZY1yCfs5adF3pKb23olw1XM42sVNOmWTTWSQux4pL8MQhC0NY/ZD1
DPlvd9EE40X31n2drn68/3Kz8j1JkD4t6uASkOi6albVAEYxX39x5KEz63ExbeEnXS5Ue25hsWHw
N5bcWyjgwhuaB6Liu9/2P/zyVMS9bqmPzF3RR4dp8pn1lsHjzKc1tr10DZN8QOeaX8hTjgBMNoN5
K8IuSFEPvEoaDSTXLUPCXr8rRcxoDUF51rKqQ31JNOjxAS2sctIkPCnYxBzqcX0LU4dzY+Y6PtT5
zr3I+aj98G+DrucOIsfRwZYZFtYQX/DwQKvIFUs/OgC5/a28L1yQkLG59hxb2uOvjS5ijoVrVhQI
hGzkDoUuyjS8tSs7gG0tVhJsZKRqsMjLlt5vMVbPquc5UrstTdS6gwSog9sOTXSrtAUn7A5O7xL9
uVYa/aweElSXqKaawyq50vy9oY9WAhpazfX5vIX7xa6yofKEqtuFVii+ptfz39ezcKQnUfO9NwxG
kmyFiMZI3EA5F7qg+uHfbTxq5/6p0pyNmwqnQ89wDsoWuu8MDLF86RBnlRu3HuBVWWkPI9l9mHFp
GsRQwjRFcI66BHUPCg//RTFBntuQUypVHyoPXLlOxblLl8CU2lbAv8qUr2oaj/xQcGaK6cKHZ8Gc
P+92znewKU+pGo9MJKf9qJOE0DKleC/+L7ZBMrrnicHAN1Vbj1U43mj6euGithZQHrxF9lUOWxNp
qCYWZQGJ9Ghx2Jmpw75zp2FiydcZxrtjO3Pc389W6MWlOIv3mv+MxdmVzQ8RMgXSI/D2KKKWJoGo
Xzj/pt87z6x19GHqkEYtnTRqhciQ+11DyBF+8/G/QjIEy9+ysMD5/EIFiDpt9smWHpBHjnqyoCNw
fT4fxZCwiSntAvACmqDGeB3OM7HPMFb4LikSpzdGFzgb4Ut3AeNw7KAdkCfGJ7x3zQK2EElvsOpZ
wlxiVKF/fIi6lyBE1+WwDg1xHwl6P7kAuMwV1ON1DC+YhPxinpG3MPf2BM3Rmc/TAKsOYkH7RBeu
HdxgXexbOEIMJQUkHWnq48FnpDDlyUkP64e/TrD4GpOKsH+FQKPomnavEY2xMNEh4AETfTTs70TX
vsvHUudHR5onIGfAGLnU2vhlf5pVUqBs2wd567Tyo7cXeAYJFPB6SfQ8m0r8NKhofjEJkza3ewpk
Xq98Sz5lYYTwTZREQaxpnwP3cbRu+NIn4ykOxmqEODuEqoHeHPCOyvW1ODyalL3qwOLsnIV2ll2O
fnUVQUg9yQWA3xPR0EfrjaRDDX4HJa1Eye43UhozbdyaQ/aYx7M6yh5pc5nmyTKxiHAgbqKdlViW
iTSCB1eLfPXB1U8HvabKe+EClJ+DLcb61kuIr1EZR8j3nAkBXClIr4KHtCydGY5lOGNXisU1KeRy
lFkJsEbduKA5hdiFm7P9hJXvhbJf2JDnqeHa5h3d9IYsPyrUZrnQiydXBy5e9SE6/gdkymddgh1h
QnNRLMAjVrZNWtft+h9IPfH93L11upShKLu73e0K0LcWh1cxxVGfwGEihXP7o0wF844gWWAp4llq
cqM3miWs2dk96aa2t19snXHDvIwnPOlVJwC4PgnUrjx8VJvSO6vvDh6uhyGQxBbCqTlL24j6K2QW
KCzjnl2OzKlkkG3pzuyQol7DncGbnxnggDScUwDaZOXZmqTSxMey+B5BB2xR09wSPM6X/lMNA51Z
iEgmfZcUkGxlGyyyyA0NBW0DtWPLpavOtQ141rb2pPhErIr1pSmsjQlz/QNUGdlD7NyPeMDti8A/
QG7Od/XBQupg92Ix/rk57mZgO/ooJHbG0arLG9XW3CcxJbM/HxJxeCuOKoCmSOJKDY0efc/FOw7I
7n5r6oGEi6b0KTEvOA6EjUi1JBZa/bvvV5qP7+xO6XIVACwIUKJr7ojEMvATWYU2B/mppJbIsq6o
1g0+f800mBXfF8STWWh+svEZuqeAlu4eK1oUkTX0do4BvzYPkT6DqIkFdEdt/D6qRvlTRCHSVJ/e
YjPw+ASM5aWSUJB6goGd58LQo8E/yvl1jQPmJU9kZ7ZtV2BzAzl9pDQeuDM9HK2zrd7ATEr2cMqZ
AiitF4yY0tU+NLRuX++aI2PAMIEt3z3oUa9vhkFaZosirOIG+uayNCEOgzmf460PwtiaZTQl5bME
VD1ncjMpC1zkcJ3SxcUCMQmWw/SA5Zcvmnt/O1GwyirYdPdtZmc1Y7qx9S19HRiXvctcBlMX7OTZ
ZojAh1OPGhLX71AiZF+gD9gwpduJIBPGddFChfbD/X23oMo7Im7BDa6cPShY64v8P9nb8UnN4X0B
kKi3/eZG3XWUJxB516PcYpMBcSPhnbE0rnU7jcHgjsSrzkRPZa9J7s50l93Pt6wUsA6Eq35udaOI
xXhPGkloqrRUdT4KCT75vdalsDPpPfe9WxfmTQn34I83zAkUIdXj2TPrGcHMbWIhkDxW25IhUmdn
QhsHFFEfXVdgU0nlanWMxFt6ULG+FpVDyJWF2nlLkVNPxLlb3ugAyOIC1u8lxwpEMc0fa5uuiTPG
yIM+/5iujBd3U0bSZMJt3CRZAU0oYytRl1ux5PIMMhp/aX0rwQgEjG853stDBPMaUS/Un6U6FWC1
7Fd2QJHVlkFvMakUfh/5VceKoEYjauMPR/oaIlCuZzDDrgwCn3rPHyb+QphbYamYdbocKY1csxxh
DwC/NDzldxPQyqvi3UB3VcShoByGteZjMZe8gYQgrHDrgUFnpskFuvu4cbWoplcaNQsBUp58M0L5
qtiJvxheA+MXbS8jvx2yHfkfW+UnDzLWNTX+qXaLPl6V2x/eKqs0fWsk4/pz2wCGjeLtli6hvcUg
Tp8DOOy1rHe9agUwtfVaeDUGdpFg8v30mjpHD6GmWQ/asUynxjXwbmLrGD8TWX9GK1yeeg3gGCZb
VfHvqaD1r7Cl5wFh1vuN0D+uvsK54fFDekcuWnLeqSyXP9He5rp8bP9eKV/YdTsOPAtHeBdmuk3V
iaaYHfqBj8ioE7rpw++RVGRNcB1YpKHAlgdZmkHTuZGMNDuTCOQ0P14CkNL1EbM6CmHCBHN1mTJw
8uBahwMypj8hxXvkOjzrH1OjHdrmbYyCotoaO40FGj5BHyYUq6QW45aljUXE6zTrgTRYW2SO1TZk
NU3lPiupU4zHzNrws1Ka9DUMYQHQD9Vco66FPKLdMDWprPyUwpgnFIVVMDcQxGH9SIs3fvlHICyF
l/BtZzL2DW49sSQN9K5gNbC6Y0CinEsE8NnB0TiUYHIn3wYpy89oyb+M6CrWEsmSrbY5Za8IzxIR
cacjOcAWsPM0ip6OOvD/jDAW/iTFHTU8Gq4re7QeX/kUQI5Z6nrvcMpz+24qPdLbHzjNjbtORjtq
evKGJOYfJnpNMh/tX6SD993d5RgnqqMpxMp4Oua8xMTK7zCg9uq3xpESeQ+YnR8wpj44eawkK84c
en7O1wI0hpQH2RdpCX/tYTlFMaHHnDdFjpGylgIYOwcr/x/PC96k361MTU+65VRPcXASNyc/ms3f
fMjDobyhMDVKKSrcQfjD1xIl9M7xkIHn9pGYg6bdfisI/4U185CUPaZuSnx7ZzQ9O9LwSxMv7IWA
m9GzywP4whSph5gtdusZPuNvA1vYsRNXS/YH78D06xfObi7x5hd8fBgrPeBPyL64iJ4LoWQB2aSd
DLcu+FKfgfb4JdUyRe0lDaY1yu7fE6RAOpE414dVJXK/zl9fEehFEmZmUtZePYnITvdlLfX5bqKV
jOF/JQs4676HDfl0diYuk0MnG4nsBOaIZ9iMId3NubLRfyiBpnLysA63qG0BrDtVsj6xqCji+lFW
eLOkFpFHq7zJIgAvW80YM+IqqAmVlZ0JWykdPYaxjpNloZeOMLTwN+FmxrL2ngLGg80CAvf1taid
7iEfz3YhBYQ/u9boABvklvtXEJ/B4VZ4cVa52v1pyQerNR0NHQXwyhApioLq+5p4KLmumeFm9hYw
GCiOcGeSvofGU85Rr0suVMfEIDHiam2DETbCjBbZzHn7fWx1IXy/sDQBUPMjIbmmWXJ7LE+tp+Xm
5nn+4phr9GGZZl7d96K2VRakDDCQX4JiCCdJ3JMkG01VD/VJWKEwjxTaLCYZbYx76HSAMYdp6WLl
v6DgPqdbNFCIVSWSfU7sKo2KaEvR+B3mSFcMK4y63BjAoeV+guohA74q0BJDxG05utxwupm3jQ+9
hkk674SC2PW9DlliyeRvGoI7YwUDHrzcUx3BhpEepkkxuIlhaOcT6mv2VLvhdVWq1Kn13AVWtA2g
GSu7kdCVuT5HzxJ7RN7omzsGr/9YUx8TGomjalddK1MK5QMqIPwSwpH8RgyfS6GHoG7Boxnv7Wbs
shdOKr2j1d3OXjHaOKq4qfH53XpHKMAbfaSf5bFCZuRXAjGSyQebZFvYOz5NRXIeCw24zRiRk69o
b4OALd4lBLrW9vfi9DrW2qfuXSc3TeuJRekzbRDjc2JJafyU20pBIqKd9hUXLcwAJyL+0Zimw3Ez
aOCrsnoMVyKQ+Mo8ImqGJclxu1Hsdj67q+phO5aGTY+ChmtNYlB2nUdv9FfXK6ac2aYtMEOsZmsH
GvKGq0n5E5gphB6kZvd60r544xSou1v2neRdzVAsRHMRpRyhk1EtfwmvWZvlreXGDhW86hJo4eNq
kcVqnE2qaCsrN3LYiFQtaLkqnjtIPjrRFPRMVDgFXlUI2vvzoWd3TBBWGfaQPXlISX8AUggrqSOp
NegI9NiQQvbap+Nc7xQI4pQtcjL29M66cNQ6cWXpKSQauu4VBAyz1WmCGz3NTJChm7fkK0aoz2YW
bMUTFmzciTzxJb9w7S3os3SHPbTbvy29NsMOgfXGg41R1xGHj6gECyWs7JT7Pz8Ys57Hhn7mwSfZ
iauxPjP/QPz+1N7YAmmuKTOWLyPSio5rO4i6nVJCRvRyhZORBAKsKjEK0C+v14ZmvrqiExSPyuIQ
oWpBC3LYAKdlwmcMA7PdHM4bWpcOJ5PK4WSeG7kOVxRqVy/vm358YeSmm/ciFze23rzOzAfDuVYP
IWIYzo2RSnwpZ+rwVOSBRqVaD+RKSmLl5ntg0HL/cZlet09gJYdsrsg3rHffw8LQUK4LlMGkXoKJ
Jx9hfFWMpE06dBSZfCu9WHEsQxq3NeXmEHyTMirbaK4N5THnPzEcIFC9xtSqrwYLeErABmXubZSI
RzY9IGJqj/3Q/pYYePoR7IPCzCbfxj9FsAAhQSUGTTE+XWPTqzb+42/tlQTwnSHhzvd1hqg8q05l
i3Z4DSPGNWWdWmqGH8NrvM/WtwzJeA0ZskD+EOxTMunCsKC8iS9U6xHylNZuzVknRFm+W011xnAE
1tVi8z5kMVExfjA2pk3D8n6qa0h29MvhGLEoym2Jmjf6UPyg8VrvB/C1rCMWgLBPqUp+DUy/PDgz
v43AsX+R132+Y4xSG+DP815qSPB+euExjzsZydUgnKkf00MRjUrQvHh7uRjzNxqzyxVywrD7pWqV
44RQMDvVpVw+eWHszZ/deLuUr1SE/ZDgMtzDTTkW3Hg3BWe9UgyucWTw8p5NxBLGXwSkj0OyyPMX
wQXOha1eJiavYzDD0qJok3EpJWPA0V13XPh68T1Rode3QZBk6L5uh0FyfZLKD99f4jH9qsaCl5T/
eGEU2Z/z8JTf/KNbOt9+OQwiAnYaNKUlSI6t93ATgNjYEjDF/5F1YCPblLfZDZ/bJSHEmkCorM4B
V0hjIIdSyILMd54BvxUHpp0h1UasHtlp5uOxFhhf3wmuwR1WUcUvpJqmmcduFbeN41oYRoqeLp1q
niBGrBJmiEYluLnQEp9GUVpSu6TsICybgqbFNiz95ydSlmct3K9Qu8mePtcOOxDc1dbP5K5jinDt
vFefMgaFdIhn1IB2poxhQVkaQL5STSSRnP5gvUORsBS785uLNzDGtbilOYgLwn98S6rSP1WjzRu5
QBAhdJZKPLTl7MMLJ8nSSgXjLgud+2pDEW5LHN89qzqhmb4GqmHG+3+/qmJSk811RZvVwo104LWh
JQew4Jm+bLp4V2cT9zbj/CfXftOybUHVP4cfm8g42okcjZjDK7VlvzuIEQkAkwkn8ogcQG69XzWv
vWEPKSiOPYbc7uZN1vFom16EigaYVEKac23r8eKc0Uvkrv+r1+sShIO5+N1r7ID6PqnPaipu91vu
6ril0Mz3BnRbrkCZM1D682Led2qT7DrMkDjUXuybSMn4u9G6TExOEYWVThotb8M2ZUr3wMSyzfFH
VKO/rIjWLUAGVYI8gzw+ydWiPJMLzLmdF9BtSD1zz+ikk3q2VoMG2LZ1c+Qs1gjs9A3fVcr/D7L+
GS3tJP/WzJJt0s/1TAPCddrOc9zq3S+ytuuGf34uF33U8xbeo8PBCknGrIUCkNTUxF8JNlm1DMyE
eadR7K1XmuZU2kHY/+7AFUN0GFihplc5nvFRJsFTmdtXHXluFLjZlQQUcbd2DaXEkAplV71O45jH
8gOjQ5fpA4eWc+7izMtfY3SyoC6LufNIJyP1GiYfkQlou4zqySdu4Di1PoJwgyOtoWlSFWEGUZ0m
e8bR42teQBXxablNgIwqJ7W0lZxr1pE/oENnG3dQuurjLixP5c5un3MjZ575P/TR2ZK4jVd3rFeV
OaC44oZyxoQcFqm7pQNTQyNzRPRZq3/AAmGIKxe+oC3Nl3T4f5/sufqbe1sq04Vj2HanhNIl4Gs3
1hp5V4MjIzIJKtvW1YVyJxwy9cTFnpjM2qtoHDFnVdHSl3/BB2VYchboQRoEpuEhGhkEucs59vK2
zO/XBFilyZ3a+1NErn07eZsOyPhehgMoz0tzmdTojTDXSRpVSMKhT64OqShPiqNJ6NgDBDTjsTCt
5mp27rW3ann0WWKOeCMtJD+GRnBECzvO5LBtMrhLMebzFXjENkWGLGDA/iCGDYYNdfYBoDG39LvI
x9MR/+z3CcBAggXrbBaq+/l+v+sd7DIJagc01eUl6VSxfArtdTJ3cNGcNmU68rxXyP0JTxUcJhTj
u85emAI53That5cOOdn8aUEMdrqllhr5LP7692M3pWQlunVSeH4jLfHqCz1uaqL2dAasmXavDP7g
LjsPMtBZ7Fbz81v/pWsF08e54C4maYVbNwRFxmWyBW/ECf6hhLt8YtdAAAYJ6p3Fu7SDw0zaxftd
f0sJPdF12ECWYyVSc7Y8XqvUHD4Gie2FxFNe3E+pr8SxBASbEqNX231kPL86IICOQB8cXdhF1elF
DBVxJ1brfnt2b63xBplXAK+XbRunLaifMJeqNga2aQR2BgSuDPLe79sHoVJd+uKtATRnxSu1/ouz
8J+sD8/YZkLbQxjvu5RNtLUHQco+YKeMOnqxIjcltPUiWnA2jR15kieZVgCU4ZkhfN+FezpRljnJ
KJz+ZS7XwI67FqRbIuFKsGbg0i+D9ae3LGTFEAfV0+8mJCzSkgP4UN8X0p8wjB3xiGdpipTo3fw3
lBBXWvLC51LU5NfVudZg48CLVYvbA3LllqKApy68EgaM0cMXGNuvT7aZ2SXVcdVbAoym/RO+SzFL
YTxHMSPMR7rpciQVgZZqbQ/Ku2oF/JDmIpk/18VHQq/G23ssIUWUPpyFizImq/jLNopLfV9mlHBJ
u3o3bD/ISZLDvG2GD4XPTm4MosDl4bHP7L5EpDd0ASNbn/BSSOTjscyWPxbayUZ6NPL5VazzQyVE
ygzwYFYNpfYgmicYdAJnky8+jcVKP+NM9GZUKqimFpn9eF6QT/6yc9e4Lsf5EsKYcuhZQQesjn1U
4prD1asxjuUDm74dkd/HoxCqdzd3MuBo/5V5YcqrBUk6Kq1X2UPbFG4ZBAz+48dy1+cZo74RyGdo
HR7tfZXkuGGNwMtzqVqxzmgITGAvel5Ypu8XnkiLbbOvkiAb9xy3wWS3X3vaUUuGGh9L8uUzqaDV
nA5jCQpTqf7JWXpQ3on3ilisAJ8/HyQfsSDG6ur2PAVUJ+YE3yrOhRoejrPnS8rgLa6CDlIi0kFu
efVGwzeOz3W556GRo1btmRmoypq47gUC+a3qzWKOkI6TFcG2gMxTi5LDYt6pwMwqlNJLn6r/yOc/
A6owe9+tf8igMfD9u+Y+TgljYYeDje0ll0vGHZAcHGYEbD/7WOKDA84iLwNKNS+0rWItYCRKDqPJ
0v7JkB9aWu4gcRiP5jOqpeieESvzybSn7Pa4jloKYoOUyBII2mQGbbbNjVUqhHslAMcm4Aw2696x
esQRfRI37VtmVBF9JFPS7QU5ICkQzDXM0FmSSgBYi6SC3h3i45Y7qLNYgL0c39XN+wE0NPVBnYZM
vZ//62s9+AD9/22JeiHIHILX1vbk7FrmuuS6zzC8ZPxp+afg5rRv4z6WoZpQ0JfgazsO3+e4g8n2
js1DGQmPX7Eg/kwgIUDA8eaOZIJwCwRnQ0iOWa/HnlUc0YOZhjDlRxBy8Tk2h2q8mJOfleXM0Sf4
iI2IbAcaYwHxBR+J1kheVNnSpynPvDr1DWNCB2p/hiwr/NwGxbh5G5EWbM6aalhjsvKQ6L6CKLZD
IMBQJeNGfIyq7NJU5ZBdwELMefmAhYUHqWBOkYkjFb5GEzwr22PpEuWMS+Y56MXAECywLYl6pC6j
+EFV9GbJ51Ldmz7JA+4eJL/PX6CdH2soIqD3LcQZhdhaTGrceUAYOPiFziGj4a4iUDvEqlPYefhB
DBeZK8K7UBIisjG50UqMjCHbig69y2BRJX5JVPAAqbyoV9/nnnxHsgd3AXjkKtIAIgnCLsgviJ0B
qrqq+n7RayzqYBKDAGz8Pv0RdVimcmVB5vj6DSeBWZXxrAx0fB8U3YGe+gh3Ql7ywvHSj5jrDzvQ
OcZH6FR+Wb2UbcXpa/P8atNqRNIkygQirtCFRlxXGQFb3HIWMJudBezOH47XoO2gQ99sYkvR3fBp
m7RaElj99nrqudkO7gUWUgY3EMqMxTUw1K7lwbLnzwBBfE93oLHJs5MzE6Lr044Y/Bfn51FJBxEj
atTYzuekHjG0ATFE8AkYWCrziQcGmSutt8nZz/RGuvotP8JYDLrJFRrzaR64EJ6L1G3OxQh8tOUS
2IQnNADEJW4Cav56VIMNlHFo3zmyfO+zOK/y6W9fYli+SsHhXZRklADf2Vm5dubrD5ir89p1M5iH
hbNdqsml1zupnhBCvDYT6xmJrNFtPHtYp6gLtR4VZu0Nix+Pmr3dfUKMeX40/InPIEmxxV7hTDbs
jcmDp9XwhAPBWICdaXGxOAIynI5KDNzbAfdDCiM1JIgzOpGpwrQldsCSGcyHWg1dsyQrx7RvGymf
YRCPqoL88kc0wDW2cXjhY13wpNA+EduKPLZViYOLjZ6JGus14HMdmKTEbceDYyEhJK959luVUwf/
K2tf+np/+uf8tLP8s6IcQt7WTESzUz1vaATVQGtU+f1EQAUXpJg2l3fTBMGwkR89vSnBjEonW325
GsVvYmyg8Ga+BThTyby+5qpg3JUAXy9zI8jJIMSu3NgXWcDC6nCsd/w9ZlN2s8ZZKwoRc0R01r0X
XQO1Gk9DjsWxYlbUPb8rGSW4MZEHNFlVhWhHyQSY5TXLu+DCDmnoKSKrvVvODI1OATVt38l4CL+K
jKTqo8v7YqJMfeWOJ8aBnbkyXBfztURArqE0N4bhmE5fDHNPPBUs18tVaJKNwsGpZl44/fGorUwY
XoAbrQy14MYC2Pjpo6d1ufsl02Z/ggb47pWNqoAm86WWBbWLHA2SQNSz5D6Evh8QMz2rhXnIFWLd
BjSPH6b/u87mOb/RoSG7WTyrjPFOhL6zLZjdLIoitQ3pD4vmLWU1PdjsoYgOTMZuM/o0I3jCguzl
H3Z/ieqhK2N08xrcHCCnRHQ8/h5hM75+Ue9LooA96YI6sds0cR1EC5BClJ9VRWpV74bewnDIqpW3
RtUSd1jZGg4x7qDRXcnvj2LpBI81dU7rBr+SCQhB1AOnoO9/ZZlKM8dAfxOuMwOqVmKd28AZPPPw
08fsaiHeDwdTWRv067re8KBVPjRGCJGwvcH4p1MmRB5vCU3DPx/bnfg26M87vXsYF7OB+/pm110F
1+4IjdMZhD8b19LhjuXMKOt42DuN0QTZn+Y1wWg/tHU8oPd/KF1lyfUfW/PP6JfM+5H6orWGOWpj
8768IiCYc6j2QBMCVDJlkcmFevHE4Lvu+PQshsbzatDDi6G3c7HSlUAipib/d+JFflbSCmV9GFSp
veuu4Jx2MsTkmVfOrxZeVSa9VkPd3dErO2FL+8LxuOBoKVvO42NBGutbmx6mue8LLVwhYOMo9LFa
jObYX8JoRMPJ70gw7ldguOpQqRU4nLm1FtH2evsSt4XWsotYhjYKE4GEG/e6grFkmbsOcV2Go0rj
ccYTf2fRPyhIs8DkvsykxJppnjPEGSwXRlaP9y4usTGzBcC7DJYtf58UvkFUCOwrroRQ/ybj2hW/
LzCkiqkBgiCtnAi9NYpYixe4LJ1DrhZyHgSQYKSKT2T1c5woq5HWIh5S2+8HJV1V/gKEL04Gvkyn
xeg+Vb/yrmgkk/lHQ5Us9LXDTYpPeUPfbwoVboKIM4wLU/dkJasV8st4E1B964Nblv2puJUipFpT
oxXGqSnoFzkIg3JNdGfBtMsyGAP6+ab4H7VYrO1jcloyW1LA8vjZo41WvSG0W7KN1q8MxYj1PYoB
TIIBNOtD2DaungW/QyEbx5OzaZVhRWnFNPvNy/xiHikHjwXLXz2q+NNeYUgM1pHzDzfMBKSFP1np
dyVy5Rcbkv2YL0B5QaG9MmXoEiOHhoSVjFr3ViAn/9Y0EGNVlbjbNbkqY8b7HRjXfLPViu/cCDS/
bBThu2LAKEjIaWLxSTGlhWccGolJlYIiqK81AxVvzOn/q2tB+UtZhn6Krru41+JB/9MRfBwleIPI
hnIj4O7bNWFv911JTZPHdtjSbxybuIwCYDoWHdHuBXfsXXZSnCEwiKkwcLw9G1Xz3KUv/8reS1LV
frv0grle7SPqerOcEYV6w4S2nYwZEr4IUkPKpKShPwpmcDpI4I7mtvfmoZnviHdtvFNLoikF2fsN
BYRfK59gxkUbDDEsFl13w7pCZbYV3nmrAZBE3cCvkIthDdC8/Spcddwn4mmErENgCzF5k/YAL6Ec
MOm8lSvJLh4lX4Y2L6R40tR+n/eNaD2UUxRLRN2nKaezt5BcRHci7yBnyLNbXYnCAHSBW6xHQTKH
fI+Qkbaw3TNQAANCPicT9Yq0n+k0hR5crNm4bRMmv+n+gnZzuHaw7Y2w3uhT+zBLoJa+wgD1bGzf
aMSFj+01rBHAI649kXKSTU5h+5ik71Q+atHWPAFLGtxDpjwybdi1FaWzHiUVT28vk2z6//2KuKIy
sZs93tnSSf7d/xYL1cZMaiefhNJfZv5qyUKHthAzq6hBJsxiyK9eoZ8u3tDuusg41P8Nf+t92vbe
PFegrkn5F2vAny+jN5RRJVo/+GWoHnepDxt/y4F7MiDTWt8PgWg1nfh1LYzYWvI22TxB1BpYHo/E
xrBjiolRqMwTGqm7rklw+W+yVyJ/R2E2pKeBDrl2hXeS026qvksuIuI8h7y4EBoFYyfD2wJKiHRl
FJ48OPA1hcLhnC8pi6lBiqKR2m8I//Frr87XAH95CFnFkrVPcUsyc8wVfE9T7gTj7znRghogCyXz
j7fjwPS3PnmpABehUV8Lqr5XBzyL97Bj0tIJUD8a+P+h7io90WiMvUeMcFwhCEIJ6LiFkihaOFqt
49SQLWC1/GX3/mQmn1FZ9I/gXzMLvk5EPTJFGs8JQr9iPGDRYSApce1VuDo4QLTEBgkiUJM54WXZ
WYR1yktcc3+OSTHsQGeffcxs/0M6sGbI3pV7nLLK6ziDD1l97ul/ccwJo0YL6iCkG8kDg3aRn4Wq
AWO3d8lBWkkei1JB9PTuZ8ynkqu+eoG3Ybsv22BrR+bknxHOcLxqE97D1ardD+48nsIdYEC5m12+
1QCo24cbr4ngcmQhZAagaAlK2xsKZOWFP/hmSHC7azF6LK/yBBvvP+uj+jFi5+S/zwg5m8u1bSov
MhcsZKQrHomrFLuqHEQ7lvYk6/L0nWyyzdPAt3QRL672Ufjbkax4Jpj6A4TZqXLlHU58QHACyOPU
cu+0wWkD5ASLVie+0xJG3CmStRMigWanC6XvNBOIymOUHFIf+O5Hl205heS1CXSaO6zUBBPYbFJr
E4fC72IJBfR0/kRVHtSbvKjDZScsaTA/tvMpjAbcCCXC/u7vpbokR0sYyqdCEJmoHA8v18KkT22W
pVbfxtWNWVAqdWqvpBzz4pUmcqk8n2wd4Fy56RyoSg2vyCCESs1xfFbcdrUpEYUpMLTQpg7q6A0X
48V/4ZY8R2d1bLiAIzZxl367v3K+NH1G/IAvkOAnrM+ytxM7+OQeN4B6lwZbKDpMoYW1BDDgJ2Jo
tXy5xrLYvltbA8q/6wpcD68+d/D+SlodU4/1ztxcv0LdwfV6vtDjuvXoq+IsmoHqcKPMHJWaofNg
JAfmxve48GEhPfYOSjEQeNJOo3/ynb+m+gnKDDDDbwdKnsyZAAgSEKrPtvdEmUDpLp/JGiBhu3YX
nnLLJquELHb+yOuoCWZ0YBMmWQvwQgbCuAcHunO3KVty203VKu9Kd+DbfOB8rGY9SsLQHpOM5ylU
EgruSDSjuSeklxUN4uBR2oD8uCev9oFv39a9y0Z0Vl7w2fT5B6uH2kJnJ9mg2r/nPfRpuFWvQdba
XCBzqzFIaoyaUe2JDdWU1Ug1EA1fJaDtZc9gO2fvoMeBKLWtMTJaNAAnWsY9FE4m43fg7ozWTIu1
fgH20FW1Uux89ezC7mmkxLfacMGoh+nAN1+cEcrbJzuFTuchYevSQyDHK7dMEaCFmWD156iJTHvf
YGNxScfEdRoPa65KfVlZzDuOyBHJOyfGXCTOm/bLfqqOiQp3AjRKc+bDf+pjyIy73EGTjZLl8HWB
5rLNVks1+7rsrqZ6Ed12YJim0nykQy8Q/lhzWw5igbQriWDD5Ic/8KU9d/0WK3XVDVkJy5otnv3D
7hlb5sT+ftADZ3L3tsnI0pj43HBZ5nKPoc21a4agjfpTqNCble8lG+YRBDZXsbu5xGNisFSuB4Uy
NLtqPf8Fj/G27XzJifnxY/UbrMm4EU6U1Pa7xOmhRc1DuUBylFyxeHn6rnTu0VHm/wujwoLjnAIC
ojGVHG5XJ7N6CvxlSTkfmO/t+2OJvmeCBtZS8/xOiJXjKYWTYqK5iIXsQubAYBy9RMyiBjxcSIF6
N+jFQu4h3mX5LSgC6SxO1f1BFNTsZdmSmSQqhSdmDWXHZJSSQqr1U4X8xI45x5YwfXdneiPTieXO
CV5sVUWN75KGh80mrRlwI7jo+j44zhtWxf5CDELgIWYElSIN/QJylAMQa3x6z2PRrzMDmqedm2/F
BMsrSCXyiIrOpU+0Q7L9lO2PPNkPH94jWCeaCWi/4MrTuOjj2SytiBK1mhKRFaaYAiq+MlxdcaEY
30nQd31e+s3N/evrwJGu5NJW3Lpv9Mv1VUkueTOCNWgUPQ03WO9h2Azk3vJ1x7+ivp0pJUM04lGq
6xYxSbe2DVoxly8Idl+o7D8AAOlE12cbusWWB53sQpHj4SNVju3+WbKbH4+jIq8+OVCdQfxI3VY2
jhuV+9+J7mgBPV0CvK9OU39hPNoEd7BVxl8DzSRHRGHx9Z+trWFFRuWVtQdOCSxMEUYGsCzs304P
owdw6XfQ/2Cs1sEbc9mJYoqZPoBAqudO/IaDQFNg8MSPo3ZsXdC/Qpdaq3Bir8wv0vazOZ2T34aS
uBhurRdKejFiYGsJHyHUFrOZbLkSUbxRv0QZo3/5DMtceBkwpULL+pjzD9xvUulmqAVAtaH/f6a6
YkNlJmKI+yvbbSl6675+cMA6jkUVOaiTyI+MkajAzsA8Jvekiu7eQqthjfFbcgrOc/Jox1BlfhJD
rcBWqCGpDZ+8MgwUa9WyJd3iggzMsv3on2r7INdbL2//aNu9Ujh0CVsjKJBqD8NrNgBB1dzkDfV1
EO/efdxlPIdqYlvf8qXn+ReyE3g5+YmM7ZPstlADI9WyFbYp/lqNKrgGh0eRxDLHbMjE+ZD3MZel
qQ3dtdQvtq7Ce3OOb5HDDDO5HbDAHnQKqGHaM4h9/HBWB4n05Zk+h5NhA/V9YJbpiqkfROTiN/qA
AHR9Vx31Ebxr9zYMBjTuJutZg91Qx7UM0MI8F6aJ+zk82jSqRpsMXeZmBACLJ3WInNLt72PBrcY0
qYNQDmCu4OBhqsiCHhUHSge5sR+SHeq1q0sco6tlyYejw4d1vEMOIKmUNo9PgjUf4Ze7rnzRZ3c7
m5/88NLooK+RPLzyGIp9INZUeXPfCiC74terzgBPl1dGNYO4S1Sb6Z/LKSzM/NvMDRHuOb3mFKzR
bv7GluVjYNYnRTpQagWEYQ9vimpQoA45mRFNWzR4Dl3I583YoLXNvmDj1OW6H9LTot9gVhg0qgIX
Wqqrl48dgTLx3d2ibCqHbEZNebgNimizXkYBdUsKjwGwGdwjzxuV+kyN7ut2DWroP6TOaTfZjFK3
qiqvayedazlzshgk4f+5f66HNXa4Be6LNErDZ8djOV5UGcMKcbEpDSCsMD1fzbb5aq7l1Y/HsmXk
3bdl8y/nkIpCB9NQW5oTLNUgxAIwvKf7IwZJKcgA/0RW8OFWHkqZWo9w1UvAfm4VIqi/sUspgyE9
yn3A4MOr8SvcLFZurx7tYyc+/ipc5bFe/avAIVi5IEIJj7FWCBVqKtvzRvMGw3jS8H9w2VTM5bRY
S03XrtngWE0/SeG2Rh+eHQ8ivFeqQEJL6T641+mhU+euS3pE7eW17x7540aE9zvRu+Hc+PvsJpOd
gRWwkLQiBTkZrDFFttGnkPXL4q3EakIYxrIzQ3Ws7WKLmxiLyomj7O72IFV3FQ1GEtJlKYklKfk+
36yAQ6AQnCW+pMXhxRz1XN+wL7xoacNQZwVQrHMhSTcOzCKK2zmjGZoiqz7OtZZXZHJeQ5eTCbQq
H/yXd/dD778lg59gtfNKqpIMbNVUpcYyu4baUQaS6d3h65dPbrL4pXYhHxidgJJKCVhT3SNbsUZ8
7X02d7tY4T9d3ATO6chWm1DwMNrWCUy8GA9wnj+0Zgdngtgra2hgTHkyhJ64W1Jf/6LImjanKg1q
ye5u0amnZ/JGMbHWQVw5VN1v6A0AHrIX+hsgpYdvTB5IBiasrxQYSNc3v43o5017v0tblBi3/wWO
aN8jIiDpMNA3UoqWcVPJU+g0fiPweo5g64y+MJSRNtRmCMpONfq5YKD8p5kKpM4jYxqwQdkXk+5M
ISqqef7zyGnczW6cY0lZHq35/ejgkRzUzB3tumiFcErDw7cNUcXBWY/zFiMAt/gFTucfEVtdXkGW
4H0tQHYs8tFXtxRGfzPQZllLAQoUwp21H9lsyCSMh/2ilPWHDBlwAugWX5S33fyiMCqcylUSces8
tlKeLzJQ9f7gAZZOoWbdIcb6/2SgE/D4iUNwyDAdqFDMPYK8yAMKSYRXi7rTKaBFlOSK/FiksAiB
u38c4JahhNMfn+WNFQij6b0+QJzz35CSr1vMZuedz89+1hQjUsSscKyv8/cog3GHDdrYk300hZ/Q
lz9b2Ijs4SSjJ1XtIud8f9i0Rn19F485PCzMLzWBRj6ZkvUESIdv84h5zBh3XGeBL3oUjpVpobs2
hCKjE91pL4Jj8jx3xIqnhdaxZNWj37yUeqOCYv87ZhLStHYHuzK0sVJOLyu2OmwYJWBHks5Sknrv
CNqZy+iROQTgnJrdV82HDcfH+Uv8boELYAT51HcAHSMLcIS4E4T2ftf2yBqX2Kgo77U249fg+ZsQ
lpSKdMG7nUWrF/NytMgug1sGr2u0VT8FgPFol1wJl7wNPyhVxyUu7Gpxkss7hVtbCrZhmQXNejKx
/b6RPaASeaXTBDwuNG9oqnK9waYsEVaToqNtJl1jSBOmu5Y69Rt++Gbvl/d1mMESq+iXi+nKyJTK
gvG+LKF240GK/1isPJfUWbO47pK0cO1kHADfif0P6SPSu/NCCj927urIG+p/VglfSPFPpsn6ZSnb
MrW9WSO989jbbOjjQ63mf8vHIR7HsGO5WgI9EX5L4v2G3AhKF6peNWkUt5fbvzh9B2PtJL8RhVb1
sj8fgmraaPwdWHXIAeZ3O94SOWNi1m2DbDa8RJ94dvOS/mK2NT9ZyLZENG4mOPsRuXw+u6mPL0P1
JaRul16UvDMtLoG/dmARi5ECiShr4ezjpc/FSUMlatxEUiAEnDktE9Lm/x8TYCa6YOMh7KuUjvx+
0YBeI5dIS1AYHDMeEPCw8s+KdyQ4iKHoQHb23PuzSvYmwyTUmqlxPF4lNwR4m7rb+/Bawifv4jIH
n0FMPWV+O3nvrN54jBr9KRZfFypTvIxmXpy52pTtu2Jb6BovE6RjngYYxNTLRRzfmluYWFlLMLtg
IMLNWZOE/NpwOD9JVcBixLIg7enGBFcH+EYkdPppxP7KfyGU1sgU1qOJfwbqIafCqNv20Vr3HFev
OBMz/k2pLRy06wdbJ2vLgehyYZ67o6aZts8iGD1jkE8rjWGcwnOXkh+Bw7G2oEulvNluP12YWIzY
TcViFq5G3k7h+wPHVHdXHEnlrZmVSbdzC61GE+DU05R4O3HYsAkb96Pr3aPFaOqKB/s/tgWzTD0V
yfuwHC1eHa8rJGFlBx2NKojcq8vCswkxPYeAJt1w9XN9mRruM6QxL9vTYdxqtfsg+1/BIh6b1QGj
4z0rXYt6YqrL9yjePW2PataXK9+f5X8efId+aJr7t0XF4QjtW+6JplfUpvRlgG1GG31isSNdus0u
+RI2ILnKVSpQZFNIvc3Dcoe7t7DVsrC3ufxE/pM13kygFOlgIQA2m6LVcOX9vBPy08ah/5vUJXpY
5TDHnncoU5ip6ci6fCC3NQgLRBvAsk0ED3wUyJFTiMQ97Z9bP9BpxV0cPJuO3k3dWd5v2Nf5M6Qq
cNMS7B2RFEPKcKetXokaXCVrlLWoBjFkGZgwIs6mnno78izR8CclwK393J65zU/OfhSH6Dt00J3v
F/pV822teyonvZ03CcySntNvx7AESWBA/MSprVJW9OCorqYnLbPLc7enc8T1WaM5VckSC9NH7Zh9
PJz9rCaq9QoRJp6UIZUmFbEmbJnlS/j2OhF5FhHi5/OyBkiWR30NTBdFJzByP+1a1+4qElc4UNqx
VqNPOVbazJs06+Cv8wHSAgSwYS8px69yH2k63uiA7ad7trLt1eGpjZ0QhnI1g/+cjhoBhiaYMCkM
yQNvReO7EY0+ITlYJ+1E76t99hQdfBblUOiPNJjSTXqnw+gOKRrYyCn/zGHHtRQWuFG312D7dcbz
/zyGx5rbi/Vo6I6Tc/bMSgQkr3xgm/tScGczW/ock0cAmMelzOkaXas4VaJ8KEBdUs0mTRsY+rEI
4ixf/u11I8n8By8cGVN9mBDhlEis/kgw6j5hogPDFFGBdMJAdGtLqjD6cbwT/IOM+sjM5irwplk/
a1LQeQwRcl5AxBtKIvBHeSOzj9bvaTF5KUdkA+7g6LvXaLYptKrvzfqgn9PRzEJF3sNSLxEqDauZ
oiDHEWayEDFCnVVPtKrT2YnwYW30OH4Of087lTOKEGyBZOfb3ef2gao8yHaaaqWl8YWrNNx1i1vY
Ikanh5Mqz1AHyPPVuyfkXNj3D6IaD1ipivpM1l+TI0HDvPTbt3N+kBO1x/VvZ3H7/xfJVYLNBDIQ
lP2RCoybEJwAkGbPScOuJg12yn4zolhdwzBovAx3ZhKXqM/lcD7E5EV70s+LIU7vr8ZMZjQaDLBS
WXnKK5ReY/R4QSHaUqa6xDv+sOO6f+5QIOY07dHuXC04AYrwky8heFFXqGkc5dWjgXcUZ9Ja93t2
LV5N0Z3cCtlfMgYcFoolTs5YENuk9p/VM7DkfKDxodXVYOPk2W2qOhaW5n4kAPHLIT5SIaSXRBm1
zVyn3V0KpbNPch9em3zfiO3TzPJRIZLkoM0AP6RxLqPskctmnh00XKFR7CRf/T7NKiZxiwLSV7dT
XoTNzNSrZPcj9zyyrz0hXJtzWe0nPVLVggoNHAmg2Co64nLOlIkUJBhiAwJCxc4OiMKj//SPvF+3
Nt2pKH92jw+Cu7NUDEWmrqvEbdPv10H+HWH2arPWnzwVipZbMGhTU+6Dkx/vkcdf+fLDIhwMijtG
OsGnfrWNGRR7itE4BXBwFznKyxztVYveThqBEeLv/hf+Gqewn1plGzHHmV2WH8MX08TP8Nqc6eyb
mEjREO/jH8yaVjYhI4jkMEUogPH3q++PmDqJwtUvZI3A9sDcr3UdOgoJtAj878hUdvYscXRzK/V7
Rr9Ms6d9CdKu4GCNX9XI/OssvY0Fv5YnsC4/kGshOX8A0FsHkG9koXxjOkhlJnasn8g/6eSAuces
nwWRQNYzPt/a/OloRH16QkuHig72ESoaYZz0rkjgnp1GFToqoeHkrkutEh+ouWG28t2rDzMi/36F
uudo9lLvyfeNETr4kgIKo6x46XhLWmChdrLdI5ubJLD16dJeHHtJH3JKvnPWivBsnglYKZI7fTe4
5KW9zbCVgCCmNa8RoUwDGkvtH4yxKiF0pKDKY0s8CrI11z4DBxM7vXakjX9J/zcwegfjNN1/5dTw
ENwoRukQUJDVMrpuoYNjznZV8WtKS0PdAVRvkVniYtnPVnuKu/v5B7qBukvgvwuKq+ENr3zV0miG
lNsK3MoWIpE8ZpWhPLE+rnH/tjh0M7EUXen7RfzLQKDFObV3isdV9B+T1/xmEVK57qPd6SBhsfWi
UVocRSEmfT0q1w10RoqeI4wGFJpX3TtF1qmXkl7H4Wfjb4mKBWK+SFGFp9VdZ6Bovy/UfFPHZ5rZ
/eUi5XA2ZVFlBPhQ+dO+G8Rr1LAKl0dN5UgzgP4xaVj4CSBMNYvFH58AsB9688AlDT5O1uVcjToa
xGT2/RC/bLegB+fYww7yKtwe3SF5goaSuEYt4UeCIJsLRZRHI6orcSBVQqDq7HCoKFeU3DxY1Clu
GiZsE4+WRgdeFGgeGPwsRM+I8/1ZWVu1mG9RxILNodR7edsebQVayxwusJJkSvQ4SiYGItTYqD/n
tlc7DOUYGF9h/Q4agwMSiS/OkF7AkImQSe3hWjKKGeNiEUXQzPKV7vpSoXrMiasikqtCzoBNvcEs
yCas2NmZACrJzDW6sRtCTYOfHQKMHVczUkkjAampKxdTtifvQ4Nd1NEzUPa10HEoryswvnrYIgPc
1iMGvpEyV5zH2F5JkMSXdv0/HSrC8MjTN55zhb9USNU6KQtMoskguFVOZjWvFp+S7nM8oPHsRZsv
//z4h39R7Kn54CRSjWyWRHB+fVXQEY/eIfN+34gUbVVe+xiJTiyPGDOkwXsfJy9dRUhSUYlpDHlG
OJgnDyrqdHAiKz75/+6mNtL4AkVgDtSXqOSfJO983qnPB3uOkD0vyRIAr0xvADWojaUbbL7wR1Ua
2/tE4NTcUeh7mAXWlX2aNE3Mp95RpNvI1RSTh2hEPA0etyc2oSsiw2AAypEtrhAXY6I+D/cCkkdr
CUnA2CmqileDgBe1KMy6EHgNNz2jrdDtc1m6+JSDoXGVdCpSoaG08xSpMB3PYqxZD7NmxMO4zhvV
YFVVyKaVpduGPCIZCVU3dxe9NCNu513nYnpb9ErqsVmsNLfRvOlV8n6cbDLpYzwS05rd53BTotF1
QW/X25WpOw5M243Zs1OXh+9W0S+cJcHHyfui+X4aJShi8J+YMu7EARRa4toYYwpeXb1k0Czv172M
QxmdsboV4NrJxhbmRqek+BXQlVthshPcyGBEINGTC1rfcXuPRymPdd3W3DchVEI7GOrquNiFukdN
1NVgzbT4Mg5BOeJqZZxdKZBUoUkb2fLZgFC6MyPdangxkQKZfRhvgm+on9hTOjxs/kNHSozEEIWD
MUTHNP1yH1iAWH27CWgERd8Xg4WA9JcFFZcvKbi//dLzGNBNnXSxyjRf0/BOba+0kjpAa8xCcdpT
oUb1R+kpl+MbTQ7+drOANhSIghvF3mFpmglPTW+GKID/C/AlAusXxObt80kKa404UCPUElnp0PYi
BqPlCxQ/pIzCNTUmdbONi/Lt7NoPY3MJy7/2kawqo7MR/oksN2Yw/DCNdncLHRCHJht4/iwlDC/x
wM0sCm9vljtpzYUTWhycmWtYv/4llvJNhjE51gk9JmbQ8sb5ubq87yhk0y2uX3mLiexUsbGgUxo9
uJieIiQh5LFFV+7u8Wkbt93HJ9fEeRajmHuW8lCrk6M/QYrLn20On+3K8pF+ibj4uHIyQ0UpjYgt
2zzbD6/3/oFiD88yb0SlSs6A5FucYiAzR5IvIE17ejrDegtP2+NmGm171B8/EVwMvA/cXWWi6vLw
lmw1hpC3bukYxX9NK0FiiJtlji83HYdU9tCGsRa2GIunR0UtKpLejqu3xP64cYGjG1ogKUiKzUPi
214AKtSgYx1sBrtxd5OGNnM3pbSxs6wyFs8uoHNn2KRBfsFyhxO+gvwDo7OV8DluDH6zV5R9UosF
ICoZBC99l7tZNmmoMquj+aOwsrRDXtnnMbTV1SMmMRmvUJLPFBJPMwzaLhVusadVLAjkhJ6z8Hhu
FmLsFmDvJJCI638gX5x6lx0fB0mDgl5WnUPd59TY1FvLm3AAgCZTDTewsGe5C6zavlMbHgX1lxJB
9ZP3hpGxzOGF1xJmW0jUaiQI+MHcGwBJd+QsuaRfZYahl4hWKOxATT72bx7YyXUv8a6UL9eqsuKZ
vHDVrVUUirWeuWsItwKLDt2qIfVczi/4MldqRIP2dg15+pT9J85/BYJkTFJqfa0Iw4IJB090dTEl
4MGq2p50QKsSU+7DoYV1DTwTb8VEHaeVYgrMwIdoOuvuE+74sYRI/CeSE9VksgaZjY+97VUA0KTS
3Chk6VRxN0cuBAGATMoLd/zejf5LDyWuRkMkteGQ7wS8r1MdM+ba3rvZpy/vuzi9qy0W8k1gmCYe
W2pxiIHz9YsaF3zWyCvwAvh8QR+IepzbAtKo1694RN9gnpzil6FApznvSeSAz5L37MKt4HRl5hI3
FDmoPTEGIVUnUh5Pq59pDAKAVjLyiayqsIg3fVt2G2KITKUupl0tPmM90wmHnhhpVeqZC59+FiXt
V3c8iqFuHF7S90t7lwcZwXuyWAS0jVLwz97RJ1GU1sizIF7aBzIe2UPGrFtHFOdAjYsmfYzK+PvB
m81yzhsIH2QA5Ce4pHFXFQ1BqO4KovsiFdX+JX/WR7/ROjbEC72sQ1Pgvun+wpv06uo5Tck1sNN+
4arqTsKxgKSbcqApmvD3xkpZPeF9Ko4u+EbiUVG+NnnAJboXEFPTvHqiFT+LwQoIgqaU0rpn5P/U
NBukO8IYbNo5nnzkQo6+FfFfEGl49XszwxLRTdh/l+9GLIxUI19+Yxg4+xnb0PJwj4DHc1I3TX1B
0spq40M+CO4+VTug/PBwb87Ti38YifgzoaN0dLsfJ50zUgdTwZqwPxfnWDuKsy3HYFKnyZrrWiov
NkOkHAX3pFXvOE9oAZXHJG7H3puzj2kDL3Zt/5rQCImK5GkXi2vrhZPVDw/X0EKTBJQ6emUKvDR0
bZWl7CWLwBa0dIHIEKtH1mP10TdDSJ5v/kLcaKXgR+Cyl9FRXbhU8q2XHDRNmkkG2e0YL90FYloI
mKidasAG2RK0+ZKVjHJrHM+vIEbFUhGT3OIedKwT3+2Gj2ESkVcf7Cj78wxRcgw0ow5yzTyHMP6s
znEgVAK/4zym4ebgCD9wLvJ2y6QvorqXzmIN89xcthdq2NpU325KGOdR+tkpMQmIlbcQ7H9qLWsx
VWVvbXRraf3uy9XefDT6SVBIpyzQbj3pIwMCG8neA6bPPcPncJpvidduMDwoInrCM/GmMBTkig6V
OvKxp+/S3MKJ/V7E3Sy3eXhHN2Iok8cC133ThaVtvrhWprViqaUYvwl72GVADVqopniYqy/g0nIQ
KIVjdj4QFgKOqCYBCBJIa9x7+G1DS3+A1rwhap66Jtp0B1EAOLTC6rm7rH04MmBhHLOUFmPU4raT
c15H31xsB8jgiaXsGigvmIjMDVJdRHz36dxHEtyTL2aV/yRkYpgtztNPsppEFyqLHAhV0r/h1sJR
oSTj25KoLTYXBfJaMiSXb74PPafly7yoDMkG+0rKBY8Nqqyb8DWWpa0t4ojc667keS85j7iT4wXU
ec+1LtEHqga8G0Y1sa5RO2aXq6qfDiSP2Ua/yzdlugGrfEwlDyHNRZazwowmfUOdov2ed+xF9FWc
nLI0ZzhCEhr6Hy+5DDL2Z51O/iEqIgCPms0vaVtkQK2INnZn1+eZ54vNUJFh+GNZReSvO2zMUXOP
U/Vz+2a3/qhiDVGx/UN12Osr23GVteF1WHUPZpIQ7HBxyAqT2tqx5unwfMKpbPShTnNFsaL3sqat
gFV+V2pfU4buaHllCC+eIvPYMbZU2NgMJuAi8PoLGuNJdbaAm4weKWJi0jESVXR9fT2m0PfLrGWL
kpthu1EkiKTXJgMpukcXWuduhTFskSj77AG7k7FeFehGufKoxrhUT0FCqpPOxGnVrsjf4pyWsT26
vGv/tdX9bQ5hfJkjnu1P/qy2nZkgxL6tAIR53E/xj1BUpsU6Osc6cdJE4pgf6oEQBXWkrLh6AyIJ
VJ2HIi4sXy61R1zC0JUjbwn3G9jCcdn+7B/HR3klFDR6X7DSGUxvCu2UGKO+A9KFoBxlXIlqGyKH
Gbt/OgHl59QLTcoJrBXBUgcOV3ZctAMBQ/PesIBiUxIP3wemtSO4SuRGmSbfFcMzl/3kLZ9DUtet
rnVt1td8DgUGcIMrpyWy/X9SDbQ8CUqG1YW7PpLuY0XpHpAbp19DWZVxvW+snINrgAqQWjqlXPIn
1xIi/3TwisMhYtPOd27+BB0YbO1DKUP8x4V87kJzFjgCzrmG+j7bycZAynh/hsU/NfHuUHiJ6M6F
60bS2ePLk09fEFEfKYh0HMA53dEy6X+rhbCE3PKVRqrnRUFy1dojs/gpT7KH+UEMWRu6CA1efxNs
UMwutaFRw+UehJP+Da9YxLEdoqUonBHfKzsuRBnrpCLGR9K1Qio0TnOmNESCo2llULs5b/1VyUHp
raCUMkRBcHhTBotaY4KZ6jrGzyAicfsZbq0AVMZ8+8OCDkMO6ukGUmMPlLA0Pv2LUwTB8hcBTGHJ
pW8oCPa2Kz+XneLOAwfiX1K0ibxmLemKGz/s1oci8twCN0Cj3accPLaQSbybYL+a22G9e/c/Xs6y
fxpqjttXAlQsuGGAW4rAQCcX5LP7Z5IXsO6sHY79kRPAtGypBSphlhxCR5QqXnQ0OqxTam+BSsgj
NCq9BDDRQjNWHKXL4dgySMJDc9yorOVf7U8mTLsAws/j2O7LvVBLS3JOBJJFmKRbmuIxB1DlXaOV
/1a1uSHgunCYBUjtZPQOZNYy14V4dEG1VLKvXoyIGxknPXmdbbMfabDI0gOKgQVmQCIPLsjb6GBH
SWSt/vN9nmwslZJ9nvLSlYfX3kZfMHj+Qw+1fEsAcbze3aXkAy76WV3pYajt3hWUgibbwX7iequX
J1vXKeKonpPKjbjIIS/XmG66D3dreToi/0ujPDoEVXYJ2dCgt/fa9mKvBddCkaga569SoUazuJtZ
l35C3l9ciN9/BSg8rigQraTOfANRL3MS6wODIDtlXiLvODsIdc30Irk+CXuxKaoD5l1iiFarXWkt
u9VOweUndwzcTpCkziuuYEugo7lw39XZzrbQ1C2c+gzcGJT5gDfDRtJeuNfNKQC7IiG9tkylfci7
+PzcORJvL7prpfFKllpPrfcin7q/7pnBwRJQ+PfuS0r2NlMYYa1v+1QFxUlOGcamAkPtWt8LVoeS
D1b1o0CIh1KVkJEkGR8LEdfIhq64LwV6MKTP2GnXMhN5lBcmXgnPe+WlQ4lwvkNWZQUDurW+R+Lw
SlexblnbScfordlXqt9pAba2vkOujPk07gnXPx3B8j4WxETmkhkJA+f2aVLzRG37D7bl8LimCaO6
Y7oFNxaK3RP7RlgvXtlUr+ChAqhoiWiYLI4dYYkrnQKQXfBRSO77IuCzS9skf98LtQnUGgMS4B81
+SNyGvGNd0UBLJsOeO4DX8eqxUrDDiEQFKrWRh+Ao8Yo73yGigipz4xlONAscrcqr3MFd75Tz/xy
XXspjVvR3RF0uwgupLyCFUP81LuaOaPdryB6lxheFy7E2F21xSr2Q0khroZmkoZ1JLDVOIRPvo39
Tjs/HSePxqy827e4oB8lc2M+wK3sWQEAZqQ4IeU1gvz2Dl4oMothV1q94XamwujcoomzZPXcj12H
1Rwl6nP3YRsQA2oB8qYDqecrrqM9PdUnRGi+d8uMeqO+IvKVObk68jXNVvyfP3+BBTsf7HbqQCUX
eASChS5MQsxFU39423ClGVEM546bZ4/xfK2G9ubd91ijcrlhVicczEFnKnNV376zpOPQXfnCFdYI
gHRcoeTj/GMHYTHXTxsU8FSgmMB2rsEdu0wuKfvBevoN5R5e9JSJWS7S+sDl/DFmfjEwcDIHiRXJ
5EP4I6VzIDOP/MLYiMhVES9BJu4DQFRFqINX69s0v2V8aN5aE9gLyG1T++5P2kg+6zGz0fDF+pfr
bBjH1gVLoNweIKbWbZb72WQjpkP4wjmQl6vuJowtE6H+PBkjKqiiqkcRkqmgc+gPah3UsGafAw6M
c6yEVC/mmAQP7gagSIBort177d+makocwIpJ5CRAOroC/5oQJA4GCXuUIQuIhA8EW+JUU8R2WaU3
p8EN6O2rUijiTSW1gvPB1tOgtER+hZpjHq0DCAkCOtMFP7WP40LTn9NmOud6ndm0r8wtwqdQSO1d
iHXfbSfZsTYiIh+fV9iZGkXq19jHP9PaLEaE9719caTGJ+YzCiQ+EQN0Bvy9cKxgQi54ZWc8GBVV
BYJG+ZqqffOwk1hnJAc2st21L1kz7BAjARIRKbmOqhmsiAAlfmKac6EwRpPnsy5ny2N+UjSwAPi8
hPHZ9oN91EJwGvv/JS7eC7n4v1nYdl/hll3olPXwskmKRjq/gMJ/l1s4JfZtIO33z4M+EyDw9fnk
c95bko6TFTw9qfW+TsmB6g52g2vp3ZCctnse53WCJxu1gkI3OtF34AvpRtakfMlg4C8CbjS5D+SH
k4S+juzGVKULmj9mJnKTjjHd2GR6mVrg1hGG2wwqvdeB8Sub/O3LEDFi8OL0I1kGo6I9rAqNRNZ0
oIJyOTati5h/TQw96p7iKFD+2Z4Nm874NRPIfbCXqE7F5F4WnQxfHz49V384HhhEJD6N2VuCN0Tu
TD5pRQgHXyFtqjqYSAPSV99rrBxqqjT451W5/Qwyw8c2DuH6CYtocUJ6Rwabd9AhQryBnQaZ2n5O
7NVAoshGFrtIo7SxxfSXF+nEna1zl4IDDm2lRLzP9TNfOdKPsqyi/gqmY7NLghODo/mkFO5cTZMd
BHGOa3h2j90yUqSpYTAwRK4ZpR2WEYTg/AodpbEtRAW9+qV/A/l64Y5hZOXcJPNArHbaw44ujJy3
PWWuisimErSTb3nDGMwWW+jFAC2+6li7N+59SDQtrYmWcT5JmK7Rqbe0kPsPbQ/I0pG8Cllear5O
VruA1riC+Ce7YUG3qsWXRXDaPg2p9HqviK8AlIsIg2CHqGCQ8R/jWC2Q79nCF16jiABLQzvmWwFy
7te7UCXcceTgGppsJHaX8tfQeFT1PYKMXbPm08TqgRDdvHtxOUoYbVN4CESpxzfsuI5PTXG6PEFz
vZhsF0pkKcsp6AQIrV1X2P1ILEGcKlR5q/x+3tX1JTQmPA6R/17vUmIYuDG5jHjat+qcfj80kSpp
RHwNT8eXgQcn9DspzdzH1rs7p9KYAoARkVFvXKQNPhKvvL2ME3i0EOSmev7RzQqlGKwE80Dg4gkO
HmxZLVEj7jWXXcLXaDViLdmUfc/chqItyQNrR2Q0Is7/jcL5SsWJYsy0B77lTzadOXGM2nYVdgJB
/Bwh4q4GvQN9XBT58h6Ab3+thk1FEugU/GkEjlKvvqy3I0drco/xvMoXWamqyGevbdsS8ivOtq6m
KyFh9VW+DStclfic5Ta3GkIZUx4mfwJjST+5rR/GxPEF3DnUjmn6TRd+b5WAXf2qiTzXuJhJRIDD
Q3CvjNWqhZAfi1SlKhumFdjyokgBiy5e7RWiPuXib6VBTDtT2pS4OcpS679jHM0DclHskj+jR0kL
SnYJCqb34rUDY2xJekoHMNaw8m2B7iWlntcVAJ6s8IO9JOKiV3jizE5T1kGOZNBn2aUZJoSbRMT1
ItcAHqacOw2A4cdE9OeKgB7+Jok55F6TluId2DEbCZynZLsirfWZELFoI7hbdLtCcaJ0+1GDE8fg
Ws+a7reIk7oP9qeuJbkawic2ccxvAOMF3wqdk+NmuQkX4U+5gzvLNrRpbMyJsCRzLb84a3quhflI
g6MKrUcDx/GsEpeUSqdH89uOyHLGp47aL8lKUBiIhoQKYe63e48IDDCwTMm1Hf19Mba3Cc3NfIRb
pHGXXjNFxlQ1TYNQrUBgZTgn7IuzufHDdctDcrwH59bI2Yo45jf1bZUChyjHLpCSEl9fweCSiuZc
KMdX1pAWOiJbLwF66Ub2T4FiwWlMm0F7b8A215qJhRBV6bfsPZXSK1jv9C5Fy29eBo9zFsbrM9CM
6uuveRTT/7fdRcZIxkSe37NFf7MSmKz8VNwCExgrxAv7+x9cZwaajk+GT7nkAygjSaQ/xxjuLTm3
7Z180kQiJ0iCWweDe+WPLFAazXW/zDme3Re4sFHR9RD3gw/yvy9x1hdQG5yx3Oh5RLTl/9ECtwP8
sZpYWN/9uzPTwdVr3zcKdea00QQhNqfhkcQaKuXFTYAhpPxDUfN7fZ8emek/NcCJyIz9NHBrj7Yw
gkqF2KkW8/0xoSiLAN/9+Ka94jpjhxL2j+1FwbkroItGRfyM4Rd0bIoAhafZVPtFGQUINfd8L/Lh
Pu3vBGD2ZhxV0eqk0Hv16qZcpujqss8B+xMowNkeOGGPB09S9y/VIdsVXsrhCWT/4Cl61g6j22wl
aLj/NJ5SN8VVbIAEbqel5fgNHuLFORjj6C7jOwSRC0ZMr/pVaUL2+Z5CVMYIzUByuJO4A5j67BTE
De/+vl+8ba42qs27M0CGJQLGVeG+TuaVe5orQLhfLyIYzIblNUVLB+ziFcWuBoNJCHPc25L3Dvrj
uOkItgqIAYq2eQ+H2dIeml4foSRs1eFQVezCb3pSYgalTJMfIs6D+CuDI17IT2Uu1rrMhuANjzt8
HYvDnI8+dHkxzEm+0eljKoC1aC/YBr/MU1yl2V9n+2/GyZkURxLWI0lXekdGOFfj3UfaTJLvgE4h
o9qQiysaEYNB7CWZNFQP0St7xxgGJGNsJ+u6EHDXpPardcMTTFUNU8e3Ene2EUiRnaXZoKW8MIIp
fQmzKkQDG2hgLHNPzE4OX/1Fbklfn/hLtY+iCsdk8tS9y53/hi9T51sjOEyQTfLGeuiZBNqN1S/E
CG77bb//atMQlkRLSz2y9XmvvR/jzEjjPgqB5pHifqrO+UZ1CqgC4Bfx0r0drKPiA/hYBzKp+9uc
hYlDczaHRjqzrJD8ab8SUohh2zgj3SlBa7I58njEc+P9cw4eGt9HwFMcJddWDmH7Qwy8hgIjNp/W
LDAStJ4q0VJiRxFRxxW3+076l4Dz+3n3JRvMzPBop0DBm/WX+SGR2wGFm8qpkHTap+ddBKqzhlX1
tQX6KTON6G9KhQxoA2FgisLPk02qftRFEtLDyvguJcPNrxxBD9qowpiNnRveiwUK/ikiBwKnUrcp
jgDOaehe+DR3egtvOuCuCm53sz50hImc2w1QwFc4eWw0XUSuTYiVy6+Hu24GW92XaiFuQJKENzQ0
USb4PTC1hcpi1XH0eORnIrPy1RvhO+I05+MjvhA1j3sVjw9xwjuUcRSXDa2XaSbCMIMfhb/KRYg5
YuzsLpYgz24FO/ktNj0DP2tHimX5ipuYXhIXxPM/os1sAQkVX9Kxt3pONg4outI5+f7jXnsWH9lB
kgvDs5qr328hi/7umOTUvwpy7gJTavegn0y2sSiC4e+r7GxUZ1SpfSWTaAhCysKBmcbQnjcAX1Tl
dEpnoWrOjC3ts1pxUClRWt8DAPVlNquXn38IJqlDe7v2ZzYv6ow4eIlwyLjxwCOWMFndYKznLIQ5
sfY5GU6ReGBFak4wD7nWcAyRSfMuMmV7SL1zQRAOrMP/ksnNXuOjr8Zw3oitHlrRt93iAPBkRhXT
FOAOAOixHeWnNixG/VwpMh6UzgVlTq/C//VstQsTaejqhzG+4Sg495AXJyC64FPVHa4TKziYMHjI
xZXvTISIFORrAFZ49CBNbUp50VeSZPcbSpJn3JFtZcB7HDHQNNf0NIHJ8f/TnbpC8Nr95HGIFzGU
pk0yVraIkIYUJc3eG+Mo2bQEnWtvyiyb7LVOcidex28nVo3DYDNWuGC2+udkMfPO0+skfLzSJEGo
UFACsI2yytLTpNipM6cqcsCYKVGPT0sJ1F8oX9V2xm5SaCbLLnMzgm9KLSvFGoic318DBPn+QQg1
+mUO9stT45zxn0LlBqXsG+eCyXw1OtLsCwLwQHmC4EvjRAUvVb5GwAAdj876vZSmfFnBV6yJqgPw
JxQitczT9PpO2t9NZyeSJm3yy4zpZp48MrHowwYLQl0uRE02yBoBLeiJWZntc1clXqfd8LqPyP+z
aZe5fOlvx1sbOMktZIvHipMgSsIvwbH5dbNjWew4eh1nyLFgPZM9NhisjdasSVxioY7ga6htZEA3
HMArb0qbyytQmXqAnHC3tHMqDZ9atlUlDL+1T9vB5ie6F9wdIq1CT5o5gQXWWZ+Q3atEFnttIqdz
Dhcy7dZou/fQk8cwLeQwdoASrBNv9cMJPmTj6ngLhxyHropjCMguD9VeOU7Umn02hAxgxDPByrUy
pI8ghno5y52XzAI89dDmPbZ8incJXSivQxT5fzk4AHF+e/8UVvyRcQa84u5VLZqNhq13f+ivc2DZ
cxNqucYXrPFS7uZ6ayqr1GivOhZU1FysAtZdvaQs+RnTNk3BO7nfjv0IeynD9EwTDOf/TUGV7Bjf
xmrCiKInQH62bzHnDj+PiYdPD+WjlELw8k7jFMLc9l8I1xItuao3dZJjpAs2vsGglrRgsqRWxiD2
NCraokeYOXZ3iVGaDYdEFhaDiiOHaAtOA0RleqQs7CnDDJDIEIv0Ww94tF3jMRlpacgwGMX9PLu/
7+tQzrs/R4GS+00b1bomSRpZopYM0xV5HwAdPg0pHtOR8gjc0uxrWxrOhoneK0vOEp7HB68xNfkR
uSCJIctimTtRRvKvNFve2Gu0t0kZrS5HAPapOqwUwTI7soUDQrWucTgR913OCc5HXUWAxrlQ5dV+
8hugwtc9ZYXlFkJejVD7/go7KWt+jPOVpLJ+MunICSdlARMhQt1uKQeGQQWyF+jqxDO/g9GN2MoW
ZIRFD11IqyTbAvfz4M3bNObdafF6LLA18PzMgJJujduBGIseT5bW12dP0S0gMTIqJd9e/ohfyxkG
MTIlI4Dgjb956ZuDSGznKG3FIxsldnqh41f6MNyVIlv5hTe5oYu4IfxKR0Msvs+HEi34n93EYstH
imPXt5q0Yne3a1KmjuIzs2DGkC/1InmErj8Iyen+V/nQbG7+7W9hJ0N0bh+8iyjVG/0KLWaw03x3
+i8wEWFuHyDEpYb2h4qjtS04DVuUMmesvJJcbuGfLzMYqAagFk6wtIQq6R6nX2XvZ+wVluRNuZvy
WxsbcFKZ9ZLQFYrWZ3WhxPeGrFSVIZgOD637j8JvrmPPmhsayDIDPkG2Oabg5PX1LWsH/MWyEBbR
kpcU/e+KmUCwpqNKwANx6g5dzzAmh4dyiaXkeA7BNeVPZ3fHL7YN2n78HGJLbsCBGGvnkdJkCSOb
A2VDWBvbx4sR+DqmkC24AIEGjIvEtsLuTudy3GkbPlVtGoE5roLwfzIMv+5naNqhDrwNGvGgB5jW
b5GJOQ/+h1Ddb24jzfamBcmZwk7RwwGACiiZdmyXZ369Q4pNOCjYY1k8GTrbNy18ocgIqRpbOfap
AMJhLVdekL2bKoUNtWSp7Y5v10R4ra3v5n8Psi0mV2IKT4vrv/9Oe5L2oqsRdOevNDyT/AgL+jUQ
Y3qOlTATo0jvu8kXqdakc0iScaYqjcjLxnuf8NJMANTeSZAvOmWl3nRM2l+IatHBJUfRY/YijB47
qRZ6cFt2PyqyCGzs0Y/dxb7ZpRw42H4OH25tGGet2bY/kUR4uEmevWivAlfFFR0gZnVmNB2c7ch8
CgPm+GY4xxMiLct/xh8btD+bGIv7Nfg9ITRDK4bQY7xZAPaA5BDsaaFx2opjLiE8AvCmjwY0X6sm
4k7poJ8gsDLdDhGNopZudEODdjPfVierHcMmXJyNh7W4vZP7SjdjpmuDaqiYzA60GSdV7PXTpoB0
PFfOOlhkuDXn5CCz7huAF5jiueubcaBYL61S6oRAR9ssPav039HGeeBx8zlyeWC9DwiyWIqR3IEX
XTZeWW6JBS3t/XfPjJAxOxle5nSJBnXsgBo2m6xz1r6uI2yksK39f1Ts6p7x0HBD3cgUoCFwxBQF
3te2T9Z2H8L8o0NAMGdQwNG60wiDTJm73su4qm6ROtLzdgpV7wB0lEmn9lSXHzn8YMIby9l+gbe9
2Gio+IvFJj1KyYtVYKRBQ8IlHRq+IHcygwO567amKVTP5s/NY4msD5lDPQS6lVGq37Gyt5W4r0kx
HRqqS83RSxsRgLmbwELUz6s1o2Ad+Xo4Ik3/gI3DWPfvhayK9BJ4DB7sIar1e3BZ7OF4kFJQvbdS
KxvEiMtojLuoueUfutKqkA7jJ0+M19Y+rqDBliGcjMe1vWRJVZikfDfsEJfajPyho9IQGOCf8FOE
G+OyxQu1K5L85HnPBwBDCdLk8uCyz6WP0zrs672QoCLww1VIm4t9ysdNeRF7WfahfeoIizOx0vI+
bh1HSIyLWQnGmLLXDqeziz6JaLJSCL4m17m9jCGQB5CVpgI+V1KCBkN8CA3n7Q9G7Eh58W/Lzhhz
+x7SBTl9ToPiFWmRHpbsbemng3BkwEWJtnIBRCGzZyEOdNUE/Vugtax8UACBMA+0H/A8g+tM1Smw
LNHL7HciYkDUd2IzWnb58nmqXDnVgDxZKjLvAtHExl3r8/li0HxD+selva9taKugYOHysX6ck41A
oOwY9QHpuwD2133ag9VRjIr7Opo3yNuimm6M5KbVM7c/YWxY5FH9V8w2RpdgHGncNIi4Z5RoCwGN
wz+fypcQjuffOsVT29kgZ+7hWt64X1QBBEQcyR880l5jz9B5/425GbTiQcgFmuUykdRYNlLPq21f
+fEyT3ftJYsJqHjfgBS1t57YcMR7NP2D6D3N2wz+e9RXvR8ntlMzi6M04MmG9kvle+viImaOP3OZ
fctTv3Bghdq1pwdJ91rLzbLZI2Atcw+nQDNMxJQagSqHBzG04Vh1Syp0kaA67KzCG2rsy9TdKdDy
tBsE0xSJKuLF7JgzIdAWGKjR2waE2t/9+ABGFybdB6DwfbzwQVCJDQT+/yZxKVr6Bi7KLaGPsfxE
bCHSWet5RgB9NH0x1xnKESftppD+L1yPRztiKjqEBaGE5bSL8rKDCzElxEeopuy1ZfrqtUYBcvu0
JUVFoOJbIsqdHW5QrdPaxmXWZubOVxAKxtCWHl/ln3R96Utx3XXeJrG0QZRLGc6pn4d3n22IZ57h
rgzBUwXp7uFe7/Tnwjzqc6TQCj/VmNfsIrJmoKWzEwvBdSIzGfCz0nfx/3LNjm+F4alhnm6WbT7/
7R6v6ab3l98E5XutYR/WcpJSMx1jKqRWVI/Q7te5Ov6d3mDR/LJBptGkHvRnx+HQSGEu8gF5CwTj
AlBUNMoAq5xNXTWu9M/aS03lSVEJRYzecG+0CUYG+JjZmAmP0zAVL+6Wu37lXW3zMZ5wQVylrSKm
MxkS0EEtsLhtWeFsDme67wBD+te0ZyH5hB7u1VtK/70EjG+BCkgGjxWIGLw0XhdK9WRXarwURkNw
Pkar4rkAsOA6mP4+KO2xAsfHph50OYtUB0DF5NOAelnMRZSoKxi4Dz75hazTy+Y/tmk7j+m4zIoc
x+QSCZm9J1OhAvOQSOAfQ8WWBdcXWpQF0yvD3RHIAsoeuWDD67YHNagbKutC31ADzhErk/wXy+EF
BId6tISkmnzZOGx7XYiz4/h+0MRNsqm1M9wrDP0iPU31jfX1r7k/jLSHCXocib1cGtU1G6DaUya5
GqN/KCXNOTeIu5o0lT1kz/HtOLd2AU0BKsvNOTyQNkZhJT1/nlnG50t99idFdm1aaGMHxUY+21So
oNzQ/nrel47IONWbsdLiJdJ632DXXg3aqeU28c9kneU9WXTgyeslA+xfo+JaNseEtXY+S3vmRw16
92dh4hGEgaTv6D3urlBrxqRbI4eV42rWlDgbXAxphPpmn7/kBDo2Lopc3gmCPlRATaR/JWSwWKhz
W92qY/VvJLYbzzTFQc2H4AV7UwKCixD0A4Mr7z1YRJjGc6id35wAQvjDdUqn8biSeu9tgNLanvAZ
yrFZp9SEUOq/Z/MUDwSUviZA8wfr+Ekjs3YihbSP/LNk1g4AdHN4ZNitMNclCqzFEPvHb9jh7hFW
4XPu/C+CAMcnKoqf1b1AWwQl2x2Wo0acFCE911BgME1tR7in+GdyoAkOq7wJwyynwR1+sFcTHFFl
BjClvH0f+mX8w2QLQv/zIgk6/DbmNiSdKk49dVZF9zsp9VIq8B9i8jlhO12i6HECGcPItXJ6G3r5
X8mkrK8WwQYv7DpwLlcoKAiBxwZMdLx3pDDu5IZq6woMIxX40MEyJU6g15T0e2BK6c313RGXfon3
n09Hr4NSP/vsPdrMRVpF56Mg1LmYmFCnnbh5up8ORisc8XWpI6dI+08dawUiI+/CqogxwLwuAqU4
gVHi/iaf+qt+Zz7TJnn7kYR22JYgo4tYvcui0hZaCoitTXBFQZ3LbPNaw+hBIY1F2QWECTnw3xok
SBykcXXBs0Z2DbuOCWxmBfuSqQ3gxK0pdpabHlQCtrpeMEdL+CThptWsj1zElHBUcugbguTMpg85
Eapf81I/bDZqhF8XaHJQepAMkC/vgnUcdbT9bM2DTBnQBpiaxLNPUgrkoLl5l+dvHk1TLXvnc2gj
YGYJfqwXiDEDKA0L5E4gdCdQeb0RkS5IVNRWdTT0XIEiDjnDGQUFldeVrPuRaBC/K9ek9lVunbTy
tb0LlGhqUBNMomLFqWKmictr/0S8d1jToAN7TZIkKiS108nzbK0cvTcwdCo9ETXeyJSj4sPifMOi
j7jmfNMHZeL8wvUUNK7lzuIYRG4fW0y4qL8Ag/e0nQE30IJAAKJPnobv5CW5GWbjJ6XWMJGdqp6c
D1zL/mJklkB97p7dZJY/2xbrwa+sGOfkhIEldMW0D0SW2uWFtdGFWFLSphCivej9r5lkRE1mK0eK
DC5cjsHsWcnzMifkCIyyGEn7uvjULROcHX2aw4c5D77qogjMfSV1w5h0YQH2xw+l7YTQNebZDF+c
0uqTcmOxM5vNYcRAQ6k9MZziH9zJmj/bnOvizv1aY5uBJsKo2lTgeMr/lTgmVCC8m62htqw5mslu
pC0TqwmkJoSL1MrQRtvBN2NYAnOt91FfLDCHP34DTzyDfcJfHVZjPlWHT33tCEFbAuD0lYxf7jRy
6/os9BUnzQmCh3yiGLx3il3To3lqcC/zdEeisH/CkEB8SQWT4VSxksmrmsgqjToIhs/E+J6bRsvM
i0iz9xwbt5uoWcAUeTCU8kKIJqTAiLRsRdmIRztw0ILGzp8OfUybbUfAjlokf2SsDhxSsTXTzQL4
OrlHKXFdWxnGGowaEaUU8Kc9Jpeh2htXWMLK05nRy/1zoGbF3QbzQGpl87E0T5lnVb6kNdIV1UDu
N/wORPcIfEe/yPbrXg+eT7eDRikw609AR0kDK4CGMKNYhkFiwvI8V3zHf6yXjAiFlHMuch/01vUA
7NWmYa6b8uuAtCpIBGbIlpFRsMUJ2cvfBmqHQEOIqFL5OQaKJCuy2/i2nIWvsx6kg+IIWPz0n7bK
T2mE8dlpnnWhTVcJ2SVeAUtTlcRvpGCtbg9Bs20DdXtPu+Cjy7k0ACE0uUOJ1LePK8OXhnoFyonQ
h19zNZQaW+JnoDA3WYlHLLwvNjLEsHFF0ZJPcdRYbrL/fY5EvMe1v+8w0jRrzTQsNT5oij1iM2Uz
5vSpCLLf2sEkncyVKHZBbFGVBmtak1QWYmFZW6g433AM9YxwAlPA7v1g60RjZEgqxck1n1VVIH62
RGq9RETFGktvOsog/F+VVtyBB+7Fh5J7fh9VN+hb28iPyOLGnitcCqVxMePK7/VkuXZfwjv7JBBz
P5iSJBfpDTBGGSFR3H5m39g1519890iLDlUcZZXV3ObqKrnisCOv2l3iMsoPzbmk5bqocdG51kog
GPVy675B2HuAXxuFnB7oQPxVBt7OCyjbaSuhYIzXesEF1AOGctwIUtLBjJDxluwqa5k1MzxJ8Nqq
9qd5jsEExOMKGrspM6PbLwzzwR+sUeidxY2kTWZDMiCDt54mpR+E3VqJzWhF4f4mGE8LigpS7wiS
EMJ4IyBYdHeht3MjBzb5ynI7b1T5tD7Lfc3dttLeVjUMOTOCbxlC80qZzsCVeI6YkBznMPy7xb/n
0wA+3QNDqinnrFMH9p4RXLkAeg4YqfziH/UDMj2cWN5E9kRgWh5FA9FIXoImIfmPT4z+/RvYDOMW
W09IB99up+zmK6JWXItBKSmun1ePnJ9S3C4PZ6sgVNQZZVG6idKitUfHYIdL69pAbuDoIBw8nzFT
URJvZ4rSg4wig5qh6h6X0eIaGNrZPodeuj9hwrFCSHVxitzOTAga/cvXO0YwYYTNI9EgoG8cHV/V
SPEnWzpVH5kk2afxiMFZHVWyMsrsVPrX1BWwZxZa//AGbgNduvDVC3WQSQJtKnSUvcUv7xElGENz
gi1UB2NvfaIk61kcZ335yZpKgtTAfSa493aAUGF8+vNwgxQxIxht7TJ/xRgmFTgduUZD8e2+9Ite
08brT1IaY8KfFDwYj3See39huYuENERCMFmAGY+6k2uEmDeV/4jdkuw+GdHiQeVHY6JdafF9g9ti
4vev6i8vlXE0mYeJwuO1gWOQDb+9rMDlCG247KBcXRPOQ3/IvxQG/Y+fJIs1vPEtK3RAXadfyt3b
3IlTiE5Ib2/vdlwgpiaHvLjLKAubNTwpZwD8MjTymSb4AFt0o2R6vXinWsh0jmivh7tbQyFI9NM0
6W01ASSS450il6P+602obBq0oivsOT3AHKJAiE0uadgg5PDdoFT+aNd22BcK02n0XrQSE+VMCa7O
QmuOrrFR/enheXMt9mdkjCTMhU944DO83fqobeXpOREQuagIJpuva76qUd4S11ajC09EN8rwOSb9
QZCSrZek+wITYEU1h39G6wwqaLsnK6MkaYxJHz4zzZWnASifimusrco+WQ+8p38BMPIwEMb7AUpt
wFmHNawm9Ahr7Oqke5+9U6nhGvNx3T4mgwFRx3FZtvB30B5H4mwTff51teWE8QFIH6PYtfpl6OpR
gjxFhCYVR7J00jeifbcufGQ+QKct/my0C3A70ib7usAwKNCnnivEQR34UY3nDoTpPG68DKL3sJ+k
2JrgNW7mfKq8ToR4dlObD2pHC6CuTQGZYRGc9XLdLwfeVfjWItNkakR5W+ZWIILkjSO0XkoKEx0Y
eB/IAbKJGYrYYH0VGCH2W+ManWUL02s2LduocSynzFVZ4OZdP7WqIdLYGR/CM4CGa4InMzsCLb5v
MTSa6qRCQFbKC/giwcmy+WKkGfAbU8hUP3NepOMyxU8QTgKHVdwHHZya475P4qFkwUJsFitlBN+c
l+pVdrZ/4pTVE7kIQ1E/ZUI3Ly+IkO4CUgQl1fkCPGvviW/fqT8gPwXjJdFX3nuCW1bRnEyW8FGq
Wmarhf1UPLtQg1b3G7ZMhOyVwwMajha1NzyKCcvidMUk3Y0HgIWZXHbELQjUukBsvtG5ojcoZ6B4
1eQ1b/FD5k8NdYrXQQMSgg6ZPpmrTmisKIbJjtBlcvDk3ME06FkN6HJgUgqe3bl9WYbc2ipV9AmH
kP76XT3zK8JZovW00YrIsLT5v1HAXY0flTl8rW1KywNlym4+H5RlXtocHVTyB8ydLh8WMdgsIapI
gcWuXgUfJVcEPRv/QS/ca1vzsIkEPLSBjPuCCGcqMLk4QZEaZdZYVV1/1n1hg5mV+CdUIaMwuGa+
mhzbkjIUZyCtWKkcB7lmf6DXX1Iy9/ZBtILRfDdq9g7zwT0hF4aGdKLoJxlf6QFXUNKRYkGGod26
/FAth9p7HRETPBUeYTHMS2RULt90tSZClK12MSjnfP7PKpOKXFYWv+KE8R8jPdVBYtTb495WzEaf
F01Mi9dsr4Y/rYzR9gcHDmntTwq5YDOH01fpmfQktLO4uQ0J5KCVS7mOzn2bRdeTwGkL0RfbEjat
gP6AWm3SxgKi9oocIXWrCM0N3ym8+akYgtB6DuliwohXLvJqL7C21GaJsSMIL1QzcwVcyDyky1uo
aYHfLqqwqoGiCd/i/qrOStiHORFgL9F1KLglRLxnpmg2z5hQdD5a7I5ByyBmZSIohXaBvOmWUr36
ZwiTukFTIRiI8fyPXaFSYiHf7sUUaE+fZ/MMloNUu8uaoxA0u3LUx31J3LyXxNoDEaKgsKwXe15L
z0RjLRZpNlEAmYC5ibVxLSyEvQ7+E88TwZrvvvkt4OPegv0XXRdJymhZ4/Y6R8E0iBfYeZQBba9O
r0qyqCWZqzPnk9La/WBuvsibs3NLPtJPxkEnuxrt/9Fzv37YSX6Nexdxnzg/FDTzLj8ogASIjc+y
Xt9FgbUohX2TbcgQ/A6qjL1BSc62r0B7gljhjM3OKZg9iAaqWW3Oe0n0M53WZZgYBV6yCKW985MC
/wvG67l/Qo8k00EDf4xM2R5UZiCjJKibZXteP+MfjGX/HADtEfgcmEqnoEaPxpevsBA6DWSKnDYe
ei/5YMoYRrsNpYiT4kLoYWnaMBeGQheJz0UXYR6neXEcaw2mstKG9SkvCkKlTkQqXTOny4j/qPae
baCt6iwAWf4GmLDPsc4IG46PO1hnzV2Q2Ae00WOXN2DhdMn0EJeBZM0yAwqtp8Unjm6RvbeGdPB+
IJbHUAZkvIgRyBY5oT3zaVoOCrkbjw2V7Yp9CtepOavoW5oUqxHZ+crtVw2gDxC7g8GjHLrtHLRY
1AGNK8nhpLA6KniCB7e9pLsv9IX65z6dAfQQemQUaOTRRE5vDibsB5tv8UBkBXlAP80W/wEmPRde
j9xPbG/QKMLy1xri8IK0UgAM12kw/OBgNgartBy3lZIyq0xQ6wH6x0yNMRvXsxWRV0SgoiqaKD+y
SXX/vwiCkB/zd2pS/FjozvpBLclOVl+pvzTbefQRiMCFlc1To9cHWew4Ihv97pT7YfpT1vcRXNyq
sp0N0jpbAIRUI08qmlOp2UhK07pTTTNTPln3q+riinbSCRcisPpfXVjbSyuVXU9n5mEPM6EkA+G0
3czEPJzkyaRFvBvrM4WZ1kJA5S630qnan1+0XBQNdcsKuItd3s45fve9ejgdW9p47TO5F+I1xNcv
HqiY+5SrltjWnbIOjkpp4U9PCjUi5XxnKYcevIFzViBwdR5Nf7MfHfwmV3J3nxO7l4uU3N+b27Ao
hRj33Os628zb9UnM7gdQfIpLdhfSRWg0pcnnUgs4hfQZ0W301ZDaecC5uoJ9cfjnrOGRqGAGFvsW
53sEYuZKHtu5lKAEXC/5lqpwSkl/GCx8Ftj7veHkc97Kx6J6lLkkl9EQ3rj2dcq4CVhLmnv972Hh
9mcQHjAEH8P6Hpu/yq1ip3dDayCrqa0X3EtyrluJuwHYkqvOhF6nRW+JVUd+18kCLGoky+CjBow6
kAGJnLxy9PTrL/Ex5Z+LBy4FNi7fEktfZuNRdchhRjLDqVbPwKlLPqzDOh/P/oE5jVggasfRfoj9
KdaZAbOVTr009IbzIPIsdzGLcPUQVPPW53P8+PWw/WvdcGid/HssLUAB5Hix517Eq5566lbk5Imb
m7/5O8nAbId5yM+JDj6levAx3Qk3XeYgDo5NQ1YMVidGL0ptzGKNW9LXB4HrTjo+JY7wA5yFcaPd
kowwUJrtpWuuyBoT5glleT5CGHWVg63uIMiO4O7FGUn69fkEwcdhbyDFb27GOg3sWlFWqjlCt4PJ
uEZX38AcLkpykZGaokcyiWGB05KgnfA7D6ImOHoSwuRINIAuQnesDSZzgs4/sDClR7gpLoc2ueUc
A1p8LNuKAULtsjFZ7h5ZW6wz3WQGWDG4d+uvWGqzL9ONnUd8yAh9B8KvZd1cjWukyyABPBwO185G
vMVhMPpY5S4Pdus+/S5PdELm5fzOvI+aqcCHqnDOAZIxNufW0R0IeuPt3/hJXZsLZVNFXnLDLftI
gDfSQ2ek47uvEHwzxiwKcHo1dfH0/zVu9imHiNxDGwHqmAlYJzdo3cxs/sBo/+oX9zTTMTzixL8S
Eu8g7vdRpfhB40Sn6B2qqU7Gj/xKqwExlnzo4S7mlHIXgqrizsokD0adTrwTbQndpUjhgJjWIjBE
nkRnKlPw4ZY8ei7nNkEWdSQ0GAsfoddKwXwJ0CzFVE/9lNOuZE6BECDToc0dcHTWPxxY8dHhokXH
iyT2tIH1hc2PuRHtoW+PYI/cv2t6NVQSJFIaRCEred/6Bb8FK+ertrIoY9bh/+2o2VkMBi6jgDNy
wKpnZAfxzpVTnSoluA+3PPPjNiQRFOmyDjmAVEp4fUSVYuX2x8eVP87QXnphadMYzAHh40047L5y
Onl/EfePDg9fzR0r/sXIGdZHu9CCFRnXff8AAdMJUfnaXl5VLmFyKaiXrnfTQUWZwiyjJP1E0Tu4
inipT5OENKq5fK3YKTnhk5XWLg9RyyANozyaAIqnQy8L8X3u++4/wSmiwm4GmUUbqTEpv6tMiSie
/mmiNSddqhYNXXduCKEX15yk94SUIyzK/WvGkfRmKg0LRJ/Oc1BAYUwJnm3reeISzvEtpN+darIC
VaRkp1zVkLB9KTZ7KpF/EPAn5RnE1Co6CEltcqPdWxVZVifuVIZJxkixOa3xjUEVu/udw3M/vVFP
dfmleQ1r4c7bVk1vkFrTouNyZoPwaTIcg+8wDVDqU13TB6/8TbeYjt19EeJR6/6LjuWEfUmXU4Mu
bUsNemAfR5TCp1IWHR91k+SUHTMZKhpE4eugsky0TUHChiMmBWgsNjos8LTxL+RXAtBIeruVvQA0
RZ0KIn9fmmNO0xaQBXf+T8r+ZOCPtVKhfyjqgEIjOISChOlbLVSh2jAZwqC2qYFyM63PUP0eZacw
lu4Igyv643J2tqHJHyNbtPSfPNvbu6u43a2Qohc9nTktoJAGwX2kXNzRdVo7/mrJNtbMRdYpZuPJ
FRTJGZjiNC+JRA3kjr9YIObvDb2zz8Qr9wSrhP46jWx3K9SejAkndNETU6Ax9oWugGatjjI9VYGV
Ielld2EEJtV0nwjI0aWlfqE32YDQqAr++TYeJY6lvKZ6ohtVNKyQylabtbozw2Pe3hkgxrF2ER0i
Ustqas6hFl8kRpVyQx4Kh68rLrCtNXTmZbYASVna9+kCDz8m7oQY89gk27C1IeN4Av1Pb2oi9KAH
zQ/Y8hRlousMAeQnO3B+DxppFV/rOBP+XdNbum6wda+4QPuSXWa2F4xT6LAK3KF7agctqaWzgJlF
lwEQtFxw9lMzbN3NFV9AspvtRAJYKrGUPDPUQvUAxACHYxGDAsFykrD3+BwYJ4k6Gu0TRm5+2112
r5y+B4eW6k5VzRPA+lUUGvQTd/hiiUxdvIDZMPgdyqoykO6FROXtaEatmLTTgtb97P0N25djZT9c
eYpFgWkihL/RCi7Fsdwv0fGqowGn/kX2Zn6b4MDVYWCRiYGgERDUbLyjS+hZ33q1CKrZVf/eo/Sz
Q4GtZ4YEfB9IocpKB1C1CnD12YuX+5OTCh8ISCx+D0Slbp2wvufFw0Js3qOvKqHvXefoKnO4FD0O
tYKAO+g4o/OPfYJWuNYzP8jYq2JaXCDjCB+Ne+SXUz0M1TSyHmMr2jOCpKZusUR57tkCW1wi+rgc
72thstpBG1qsyUoR2f/aLdsLezmv8qGfcc4rJmytnV5Tfw6MoXlDhPOFWzT1N2+NJz6iDUD2sWEH
ApbA2u/0CxgxLIDkehUdQf4XlZaWavxhFTfbVIYPLh+wwajkGmHpFvJIPxha+jUlkDhOMghtyowy
6aq8EjuSsXQiPygoGkbS/gu7R1RYg6yZDSz+yZdgzKD5UySXqUtErRmbYnZ6U9uJuk2tCBjjEalv
srsyMxTD2/PBuICB6oa4DPtwOdzL3q0ZkqWnsPwyvH0nEjFKQJwWioI/C7ajNEw8AGHVgk/lNFmM
GC8AFGQm8dTgi1jD7BQZwx73POrBNgAe3S7GA5ZRIlc0Iv3sob8+WyGbaOTNOBjLPfrg5hRlPJVa
dbUXp/TLnv44D7wmNjzMCpSWIiNw6OkPTqJok0gDbYLyDRP4FQ08wtTZ869gAOKFLn3YJyfmQuxd
UeKMKs/uAPGAluYuFCbV8QHV8ywUXpOv+P/40nkhh9tSdaNsISJCFG4WtYISkN19W6rklYM8B6xG
BrfdOgzL127dQjxsSRSkHQ03r5ScEH3FFVKs1l0e+XJZjfjk/5oUs6QHvpAUPmHSjHp25SQ1Ssb/
qj4gZvziusqs4fMW7BkperQO7IXUg8QW8plehzfn8OrDYT6JUv12+u9GABxGmF1rwR8gUHg1+fUD
osDy83gaCsSfBDp7DSRS6FxQGLS3GC4Q5w+HTzqD/fEZkq/JlsaG9NT2B1Dcwdhxp8kv7NoAYPiK
HuHzeBamSe5pF5KnE4GNZSRkntSkuZGabwqNUQZiXbfaJ4xf/CdpMTAZki7MSBbKq19WnlR94tjR
ZtDqJn084VISUTlGmEojSQPf3DlacioEGdyk+P3KjhBfsBusQ124cfl/rQ2eTtIYV6GqRZmcoNq0
IVxizBiDlz++CGZgyfMPXvVl+5T6Jbx+J4ViO9OWmNfVxkZn3Az2NNxuJShJ4M7NQ6LWk/qrfALw
tAtVmVt0LIUc/bxb0nFFOivvkHQalcFPgqHjhPIG2hxVbIFjKPAr+IbEXD018kZ/mtT15KSIyif7
0xrtQfV9Zj52yyUxqHcmeI3b0UvwOx6Tq2u5YKGefa+AXFNxAFg1seo0y7M3Q2sh6UoBW0A5ll3t
IDXmG/xQU9bpauhtowKCxsVnG6CBcTocQl3J5ZmEspD0hu0ytE8CGMGMSnPrjB9dVNDMEjxWVUhp
VHfqxjZGzgj+kvy4zT2PYTs3D/4LgF++yhMhpYhFIkqcu/4G2vzCwAlAH9H0yt40Vd3x1Zmw37Ot
wohN2UQEwKB2QM7RKirKU8gkpa86gBbmAufHPDsYlf6gL0n4tEMSw6RCgAaBHnBnZDviFhqN/hq6
IaNlI9rqfUYkbJcfsrZbUmVSkr9T1hnsoe5HWHK4o/THoFbdPj5kFgGesG9wcyyl5z45aX5qnjTf
5R3lh9C0Dr7vM/ikbtdwWEUznMMKdbOVZVz1SWwAvb9DU6QX1wzVNDxR4dMu1LDJ0YUVPjqcm5Vt
2V6WGHXIF5GX8ggTEWlOuVMNQ67IV1vPhcu1gKstfwWvOf/kYH9N7K2MIGlYAo1foim/akAOWkpa
JNjaj9L6UHKKSXiR3r4oybq5cRS1Qo9VZOlvSCVhNEPXKkloOpnZ0yJ2AhNeXjWCIuwKlMT4mHGM
jp2WuD9w638vXsZtAUouabTJMKNxI8SitCMGjR57JvcU1erD4CVqtAfNb+CFYmGtrkp7k+BZsTIi
WAG4jdzZgduxF9nhYlBOHOQjzztotXh+dgvWzvgYlz7OvfiJysieKV8qO7El8sG8JgrpdAMflTs7
whNAgZu2Y0UEwB6ZNmezeE31DHdRW8y2GCgHR3tgJMcNiG92/tBbFGImVynBb2SVtBmlUDUTW0Du
KcTdaBgyGdVpyFm7BaOUp4U3wXXfZVaqLaQCuhXQGoYj9koi6k4TmZOtUW9sAn8t63/VHff/ID2z
PoLUa2fP6khVFtvar5sXE0korO5UPJ7XD/CovaLuBmEPZnnEBzE6AK1C4n8THRSaYHCpUrXoc7Tx
USLOy6PsqLTLnX3padwYYgTf84Z8T0DWzQ2COfkzZyl8oKl+CP8Tte/emXX5Xd1aDFXSPFvYBUbQ
tm1UAW+TmRc9BWEwHkIX2cZrgX6/jjnBz8nCcQOb0vtu4cgujfhGTtn+BaVJ1kUY3jqQtkxBlrWy
xy8AMi/vjyWPnVefs379zW/KhlaQEqaPd2sfv9YIPeABOwxd0lBBBXKNjbztuoIieAnRM6TrBJk+
87OFu8gzfHfiWQo4npggfnEiia2g4lR1M/yy8Bg1dpT2+GafvMPNbXY8r1XLKmUhz0augW9KApJH
zbsNrCKAnGB9oAqvdhRsvWwVN2rWSzMpdPiNZl9mWWuExa8Ux6z5ZItaEcJ3DoiLPqZVFT6Kz5fB
8EvAfvobpnq4xusRT/inz8JFp0+PRmyzLLn9bdFzrXNttk7xsqUzp+urGqADla09aShSH0h4/sFL
9gSHYO3NZagQo9VSJzAaln/lTizHVhXhPCqK/UFqD5WLa2OHuJuDXksY+wGTaoAf9wTmVCBVTutq
nXHjEqVVd+IfirEcQjkNJnlF1USHe2GNz4blc2zuZMwatx53iS1MB7XBN+JxRsIFaBzeAQnBExHy
6Ff6h5S5p6bTD4nsH5X8tERuLrtDxBPZSe1nPn9gd2rt/3A4XXoVpzceTkiEsuY44opjD8bnTHht
7PF+Q7vdjpRQ6vT7wBpPMW56cGsSqZ94m/luqYt+QKZe3wc3/pgIRR7LNKmkcg+BnhQKNuQ5pL05
we8KXBFPYNO6plVP+3oljLUG9D8hzQAdBHKh3dyrJdD5izDNzVzJzqWE6gdlb1ajLnFYYV64A9FV
tPKhtnfrKJqpgNwWy4iQ1KZlLdgK9aB80bWNT8GvFgrY1BLKm8I90lIv1HUsNMn2SAqfvpCM/ZWN
FI6/8DTkj89fVt3xebXhBiFLT53aUwCgV3lOKq9LzBvv11/DJEGVvr7qrEi8zLH1gCC56C9hOGum
Lyi3efGhVVsQPHXnWDGEqrKQhK4Pec5tZyqO2zQds8QqK32j93xVGCIt6cQPIhWjbWhKTdRjIrcr
tkwNWfmHGkeROPWayWQ6a5jKOeXLpcXGsl0dyXVoXFRniGnGArXmKDjuCc07LTeW/k9/ootwEcaI
pDrD4O1Vr/8crGUsJU+jld4eXPaddxOGMa/uh5qa+bAgz2GDIJdWFgFS8C3pU+qEum5j6tFpEly8
A+/KY16E66GpDgzFadmTqBBQc6Ksp0sm9jV7JpW8ITDskkK4/WQEyRMQdIArOEjttEiZkTpLTBYp
0AB88ubXm8pMqsGy33u7XWUBrzHTo9/sthNsYHE6rzcj2RvnhM57wa7UCGolOyJUPAR6TeibeSyt
d1a6gJVFf1Jrtn1XCqYoK0MJChPCmq0BLJllFEMrn8OBZDCEnCYC32wdy2HCpgyXBeyZrK2pLQwq
xWeRDGpwvbeuNtpxDaB/bQHUbzii2QQCtdIhf7cVrCaOU+MScu+7vJLDrdb3Awbmwp12FZQnQ1yB
bvh4nRqz/erriHQ30G4iNKu/rB7qo22WS7wqghI2gRBe59JHlHsHDR+O9H7DLWMd5I0W8r8HIKpl
bcJTMpi31c0pnpRvlENXG3R985mw2pY3WmffAxEFKKPLAS/OcxphuD9r8BZ6+UNXIyKdgHyC4I3b
5bO4fNkdAobrjDInuvSF/TJh5cYkuqQ0wr57vR6UXQzwelBB4cUqzDt/z1w4VhBzBF1lvCqQWoUT
bRxhQncm317kpJEBg4GxUaDobJB99GH8ZkL6KCSj9RdLn6qt+6enhJn6DlmEinpb+AC0n05lmOLO
HeUD9A8/bbPIj/9I/qjO/xu1WNipNp/IbKnTzKq7eB8g+8zvnL+cZ8tNHiIN1KCokAo6aCtN7Ldc
gaQ2e6VBamg8O2NnfoDbF/8RlC1rb9dAHoJj6VunDOAfgeR6CT5KoyPpBTyKUEE0+8GNkcmolW+7
Hur76W570jWQvkAD9C9ILd2PJOs6qD1QcRA44j94EKIEIR09fFzwcOeJ6MN0l56W2NOMHHasUN4F
RI8DfAb0GZceZZ7Px5llrW3UptZABHOAti2NdSXQ+p5cAEV9sQJt8sq3BukOmq3BtAuAVwEm+EON
CnK9QzvbWtEQNkx8HRfXelQrjXv9Z/0wbhZwI7wTB5/05Q815SjbHZ/hLVToQYe0GJ54X0Dz+iDE
/bx7Dre2ALc0pwI6f7CdiqRfhRL883LIEpT4ohwmdDBmqMLtKP3F1/IfHbs9QWA1ZGb4bOjemzUq
HlBhV/wEzJ6N0SI4ojghqgo5E64KTNOAmxWyWFegxFmuLb5HMMqLrD7C2UA4ONzjOX2JQbYh+AaS
yIu7OP5vyvbfr/7PPPmhsYk9JLAoood+iLwPs8xwDLTvuQygfSQHsoiG7WFxPTVWjj8YeIs7grbK
N9clE2lf0PEBAKBWGA0PGCfkvrLKGclNQ0PEirKCWZvmc7aNIrVq8xPsVmuUylAkuIiQNBmgbGL+
qF9bZonT5p5OkExdhyUGgqrG+aEyV2wYKQ5xQ278ZKlvwrk0IjpEcXQ/+1BKdhTBT9kNvi3bKYZU
q6ihSVKGbVSAlr4gp1mPaoRDqbgDDiZPVLUx/XpUkNZLLY28qAdKb9fjdQFPwSFn3tG3308+C8tf
se+CTspRfr5C3tgfmllQmHFpPI5qymgp1rDDndc2Mxz1IKkjO1yMG+PheUGZCIVieuOoKft3MpDQ
+bsEp2lIgAAYOJsRKTl4GJTLvh+CkZbPA6ohGsjPg5F+4XIuWlJQ151G4326Fm3rsz8vGaVIF0Ro
hkihX+ptbmvUqTeerKndYRaRSMb9zn7tL4JoRoa9bw6Ak2yH7jYbO+j4X1RkY0XRpJT14qj2EmCu
CFvdHrFAoA1POLYoTIDbOzLwSDocmJILxc7whLTWFrOCYV8zSV7PlMOu1jYkVoOsn+6lw+Fgw/cj
JJ29gypQJn6VbmTHEZ4CmQ8oIAI+46wpZ9b+UOxwDU+1OsiSMWRMhEn0PyI8L96c4wKt/nSce1Ko
PMpG+5Y0V7BF9ooKwnVTZgmFaTzt1IgLdssrwL+rP0opTTT9/yAtc1g9gAUx8H8uYKfz5NoTU4mm
r8cU00RJrp2ONuYXoFWGpN1GYTIqxiWF+h9ywh8MVKdGuyKu4MBQO72pX4UqfmWh/qwgi11m5JmH
/z8ExUHFXc5IZFZKWkgqZPo78ek3i7RafQIV3ngCsf+wErD7kBG7fexEq5W7fdLTREV7qE7gIZ8e
sdWTdZtMjWghgm9p2jxmC7eyJ6eTyD5hKC1i/w0BK62VIGovIiPGDMy/iuvxKCvoWoJ4HcDa7Tna
izsGkKivYqcbdvncEZRL0CvK828x8ba8W11BdsUnqczzZiojJgPN7HIPTIKx7+olhdxMjjCWDt/k
Hk/f3lyKDUGQAZb2KRtUEel93BT+SEMhaCPlp3QtSxtDgDrYyoDXmwM04iLqSc/rKpmlrgz13vmS
ofACTOu2KcxF439vJow+zedbqx3593fxA9IoQIBPK4mZt2pfn7NjoDjH8zwuIFewEKbx9ecY3DLU
qMf3brjyS0QWWSyn4lNaAOJwNDeNIxyGemr7Us8/wI084fee6aJm+OfS25jugrOy9XH7Ne+KItzE
NKeHA9070cg9KCz7KcagSA+56wD1smlOOqGiULkyyTwdYUrGyYmOHqVT0oQVpuFdvmswbFtzKsDt
WpMl1+28Yvba28pV+ia+gL93DpcgSyRVsCrBhhOpI1Qgjqh7riI+hBAim3NAdQjnLimRIeAmad8s
k7XhxYlatRZPEybyBDN1i7cshWJNkiRlVTlo6LBbmtbdU6PagZcu57xJVGGc9bXlFIr+B0YWMdK1
MKwL7rjcAZiuiUIdSRBsIXaAxtJU6qEP1wQVbOaHJWipvmuDDqJzTJZWqKrq7ojA18I4Q2qQbt6L
Mg/Gissv1dEIyeSJBlmaOI/5e65ZRv4o0W2DUythN5VTRxf5I60NPNaGx9pKtqj+hN9L7LAQKJfA
9bOjWTJew76tPgRdI0+5v5EE8J8zFJEtdo/R6zL0RC+6HxirIyQcuqhn/ZTTjtU+x5v1ztQ7YurO
NHw6IW6epWnoxKCp2W2IpdHCxNBFXwhYEis0Xt6q17FucoqbsBlL10A2ywm0nfFNG440ZlrZ3I95
MqkuE9KXlvGQo7nj+qlvULP6ojKy2uDIdbb7PCGDuddSze2FSdaHw5NIHV4JbLBr87yKe2uXs7hU
FLtjtpNd1H+DGuqsPzvFfcea+jYjBCHnwaEnkXYTbfR3a0V2RJ5A2ts0V+yLLRTtFt2sHX3UMSXv
jnUHip7ik/2afuelcUrMrAvccR1DklUKfHbx7uhfs9LkV8acy5mBDFbJmubh8izkbMj+DTSK9gMf
CINhifzgq08hKKgHKd08tW2yA3f8YM09eQ/acAQ+yGsbRZLixM04u1MBQwCNufm9D/vnMobYH2NM
PzYJh2x0Q8fFZzSxD+1sXYkVVTcOCnXtljDVH1J4oVp5BmW3cWSeFLd2NFISG65btVp6vh63VHHO
1I5KCunxbtM9jOzYIj70EES6aqiq4SZ9J5DRH0fKUsgUxTNX9Tsnyytz0SDb19aBKPI5o0kvJFHR
mR9jeBsTMKjPSPrtaUX/cLAVigJkfZVC+r7eOEnBm+9R6+WfSYObtbHjcX6zN7KJzRDHI2CyXpCl
Ealaff5RX2EYEhNfR7hkx3PFTSSwa1y1I5D7ev6Y8n7BfOYYkZGy84186kTvPKUQYOlmcX3CbzxS
Y8Pw3fgY6tTeNUX+jsK4t2Sb3lyJ66MeoUL5oO3tyB+FCGWrzc29/YEV19EeT8O1L8iOpVBLdl1I
AYxKtNvTUepUA+rPPrPeiaBCyS+uWbHnonIs02fZlP5hWxDKn6+n6ZcAHQavUdSM8WWSKsOD6D8S
VORQrLx1/53FYTiGC8Il0NnG+oFtHFvLrNd5JmZSRW8O5pxeOn1oOx37ER9g38oXTJ5A5w7mOEUU
mQ+Aqz4jT7AK7/JyAvdJy0qzkI7wcW223HqsC5tSUUTxvy8PieoKVAOQHwbFKC54YjgGUFarXc59
z0zBspJpIWXHWN6lgK+loH3ZJfL4PhNQQTGZeEtNyuF/m7mEP6s+GxOt/IkhCxfo6K5vQtyNY7Lz
hs/im+1V94RVVh+7QQTy932A8toCgTnZs8ZNrWbDnXqRQThm91RE+Hl8/BZt13/zfhvLkw9fe9Yp
OLhdbRT4/GkusncKE9kohZvkIZjwZX0ZoNDIpFU+Vsj6f1WN6lYE03wdoJ10OrTvlgW4dPu5Urqf
M3LsSQtVnIUlKhyGhuPmwA7dhF903hVfeDBIVgugr5DKawMe28T8HSW2DEASwlj5AeBsYC9kld6N
/LRb18v8ViUQlS6yU0IF9/9YWQv/U3bB7wEZFFlx1g4k9KZDitztCUYxkHCPiwOk4bQuN32G/Gwm
IPOF3SWxbX02XTys4wBZ6QesEhsBJG8gtJZa+RBCKkkSjxQqrxrPaCSaP0qyQ83eio73NM38EKCw
7Qdny5vD1aCnKh6/Uet8kDUQfNxnGwtgs99gq34MQD7/dhGwoxlQ14//o3UUNrGU2VDk4Cu0jNeS
HRkprBlt2OoI759scwVAJYwhxGStxl9n8wntlyw/51a4ptqq+g3nFTxwca4WTyQYrWnbAHA0WEAK
pIsK+eF4MQcOPZJumvco38D49JBrTcg86Sg7R6APXb8TcWJ5aP/HeyE5p/f49JL/C6LjpVwZuYVV
m8Auho5orx/7h0nHi8eEmsrKZSNjy1UF/jkrtfX52IbFeS2k19JX3Pn9IbSgFJx1sNEQyLVcZH41
jA5TwX+ftgeABq6/nPGCyFL/iJO2+BRAUTXOSQDw2bseJ5Jw1s/trr6Av72xhLGoohdQQHDVojCd
RBrwcAKoOeNimF8ZfyDTAvywdhuDp+LiFLKgs+Cfh9aRLR4fyaWQYWbFkn886Qee3Fw92Tys8U6w
mBHMg87VDubKmBwKC9x1UsOo/hRNd548YPaLKnCin6GfjwKMYiy2+r6ClNBEzXZ2ZJ4C3j+ZuAu+
xehyQZ5t546YyycUeoX9aKxf51oK31C615+K3476ZircBMafi6CqT8xNd3ig7gVCCckcvu0Nqx5e
VivqWJFm+1nlyUydbVfVomPU/0k853fgM1Eh8hxOP9wD+UnUs3TtvrYd41Vx83Qlt/GimhwHMocF
dNgoyS3KRp6fTaScmPFQROHVU3JJhzYKAAkzbbmV1NnIx75DetEUMoRpX//E+52GhewglJyezGJ2
jGiA1DK001ff4hUkxq36fdwWLU/74V6d8OjejhJMFY1wFnIo34xR2QtNgBNSIBYWirNirw+OUfIU
5j13w0OuVj2nB0UI8GZXj6weQWQTn6m+ERrL5vZfpFYYOje49NOisbuiiTrUHx+zyRYCDy+aDUbM
mcHmfeQ+E2UqTM9soed+3PpaPaHbk2iUe9/Bo2RXlAoDqf31l032A1x+34vCu9JicxxqJKMUQ0iF
aupAh2jKNCe7cGt4Q4mjtxfMHHNveHD7ycxrhr5ns5ysRjYDDhH8CuYs5Eb7pi9zmwKY/kH9HGjO
8+cWQSdSSbiUtX82ypY0WNzaAZdsQbmjmfOy9JeqGuezcDa7TSSjYjkx4eWSsYeurCmn33dOLDBs
Be5GrNdPCnwppaqUlWqV0S/Wh6yHv0HdbWMU5vJEHvaJr6wnxdQnCB27AmrXUvhEl39/dVEcPPGD
Hw9NgPSoPu6QQDVim3gnQ9SKyZvZwTgN5gyPaxD3FwEitzmwYVFZ34C9LRerVGJ9u9WRz2dwzB51
+jhnKDOz51MTVoVeeLWiTLA9OSOjd9K3otWTI/rq2YoV3H4tlOH5IQw8jjWxI3ORpMpoIS+1+K3d
kwsFT1rqCvp1lxDoToCkAoftzS6p6cAd11KpJJCLSPQCb+UvNIFKT/ASI7mt7JNTN58yoL4eH8LG
E2pq1NEQzbkEEaab24bGPaMRYSQx5i7BXxNYY9lLZ119L3KMl2J0eJLFmhPMr6zaHM5AUooJf198
dhUtR/lpCj9owed7uPOidtvSHdN17k/B6Ckhw1FcORlAHs3rqAU0WplfOkFUE7Zx2vEBoKUJM45h
FMaCAiObn9j/h20GWP5k3Dzym6k+xGmlZxpPimxIMgMLVKaoj+08XQfuBZHGhXwmllh9x6j/Oc9T
XEfv1yl92czlCYOi1pryijFG5+Fk5VudHMYeJCQnDoUzZfctfcWKXw5JQMtDjgFf+qLcWWu+c8hj
nTt+YYVMD/p8OGgxgNoWwmKTnu5px2vzP22d77zpt2z0j93jk2dx08YuGQgA586eh8jfNJgnIf8k
Iij8uNNme2tDhpZ4Xr8N59HPSUjhH1I5UTUNh0cpm/NWwJ+FTO3qCRMwY+clprLdvOYO2t+Tnrjx
5yyPS3QcW4grI+L1oIf/iOnKV/rs3/8YyPINXOV885vFJ161/Ow2MEWzvhkqLMu0CP3g866Npt0t
Ub67CCuPxlBjr2gPNN9if/oK/coGI2Y9w/dNjzyKifA4XszgIzxh3TMksarK9sXKafGH5GSiBESd
ly0qdNcpd6yWL07QOPQUeQQnVXcUMtsvNknuVKP6btgSH+yTSs68MHvVo13gb1kGGso2FzIVHX/j
otqHIJSq2aXG9uY74hr1sRUKTNWcksecUWckNu+eJuBBapQvYyqgo6jKHTMtgntxSt2BXPtumsxb
ljomtg/Fbw6m3o5EK40KnWf5Vw574vOPkSbl6uvr+x0QCy08E45FIEPy0WkdfmrI4LDugZlnPTM3
BalV+4ZGlNgXDTrZZakYuv7Wa3SE5qaFLrAv97k5safaaFwZcBUTo0HthVyYHuwhGYoOkhG4yM9z
Y+sXAAK9JQm2sy1YNpz4uId2+IC/IW13uzaFObpkCq9WB1WKk+arrx9vmL9snJ1DbNXNsPyBc6cp
J/BhG2in1K9CLCmvbI8i29e8sxVwt8IIbfbxoe3zw0EsjBRE37ZhJiSjaYfQo/YMtZ/IOHQOYwNB
TdOl1qYV3vfMRQZ1iYeHZ94Paf+hLO3n7NWOspzErcsZ4VbrOgAsFS0v+5+RjDgPJlHJvFDkeXiF
d8e1mClq5MqdyqEdtlDy+wq5xMux63F2p0tJ3f4V5EQpBHqUmIHwgEBPQxZ5itwzkm6y5U+BY8QN
EaFD2tLRVzYtcJ8lCujLi2RjqRGkDjkMvfcKgaKYYc6o/kXiUuAHJ4WLtzWc9lVu1+W3XQ0eUGSc
z2yAY1OVOukJuCs8LXiUDf6AMdhKDCAkGU0VsOmaP9ucJLH0nxpQGsb+nFOBbqkLhPZEWj3SMUx9
dq3fSxl3iHCemNRG5b6Ac1ZFZqvgY/vsoR3UlWs55LU5IthoK6i4U9FqrbihULxyIJ/FkWJ6DfMy
War9wCFwraTqKuURWYUpS/jbyX3aPcXXbjvIPiAqOYhL4PcmBIGQYxlP1lvau2A7Xgs7fnZiptMX
dRNfbIQJ+2Tkca0zIriFgj/BGahJt5TMLrtYlizwXNGeLrVQCNAo1lFwtA1t7myz2jImQgXvMJ/l
LMsRThR67J3JzuPJo4BIewtncs7JPGb/Sz1McA0DljLUdyHqrv5AH9DNMTkPlmh4jrrGFXBq844X
2Uz3J+QVqzMKXq7AK7/GQtLK5de9VGvmhC0MLknY/rOktFP3DZElVgQu+J2IbOSdTLdqIdZveUzA
jK9T7oSI66Ke1P06Cc+RC0MGjw52L+s0WL8d4Cjdq6r7NlkkB1FDcWUhCoGXZg5i3HClkTVbit7b
mKW1FGuXawReg76JWNPV0elEKteQvHN6y7eVG11hxqhED1HijtCDb4hoQSzTw/VK8RIcmAlDmsIl
yrZrAADg+YYDIu8l1h8sTINQEoHoWPolhOZFtXewEot6VDoDW3VWlr7dZyAvWe+0ULGOw2z4ml12
EWZqgXlEVHmJxyOqcmfFElHhSqKU99H7tN7+H6IOFe2/jGOmG6EhU9cb40a5Cpsd0DlInl39ainK
3SimCYFCTygy0EdsUEapORmSziffc4+hpZ0ID14HdMtIQ9EFg89w0dYdrU5oTWuRF53Jpqsxu5ay
8pI1B9VdDDDshcxFiJWEs2xiwkPIH/iaNhUWMYnqSjUyLxzDTaGr2UYNR8yOfhZPer8RNUVLgpjm
tjSgjfWLN9e2gMkGzdBzh/i87GDgw1hKW1YLk5Gj50XvdbXTkWcezi/95iRfU9wG/c7wAWU8xPKN
tR5G8aKk4T1nRKlNJ6+aJdDTu2S5tPrywgvcTmXvSJBtja9wCDhQG/Eux95ZbHyUqwF0XEHTxsml
7GLL+m8sRAKROlj63yNMP3t+jFgyo6u4zPa8DxEkS6DAc0iQtputIObQGX3ppHwQ1vmPM82we880
NkgSK0Pz+EPOhQVgb0MSxkB/NH9mrc6ndhnfGaDJFzg080DtjW5L9iCHm/zuIQ50Jaa9U6DrpWf7
yYQIC+RugDxXa1hTLIEl5s+FKTDpd3vL4BqEx8N4rv01gjJHfNhZ8p9ld1JH9nosKaj4ywhWIOMx
mAO0Xn5LFYdVMi6a3awjOA4I18IGpnHbGHT76pdFwZfZmgXaVQspTW9UOqYLpSosZEMq8afRf7BL
kC2PcOQXfC6vAwFMhTJjIFOPQJ/RPnXFChQET8Vn3hAz80+Q6t3a3+0Orc9cx3358pnTD382hihK
1rgvZoT2RoDbm1MU2jaoE1WmldE+DlevqKGaN+IW8iylDEA8as6FPcgtYkGTrImYV0zXotrZxC20
ASlR6/S1HOa4dyhdcWLg8Th3FPD3DcO+X17x7wl/0Po1nYeZyTYdybhZQ3dxw4A2nZOVMYDk68X0
zwihrqaZCUEArt4wOBba+TtEPcZNEOo7naLaKeyGqUBJtDsxFjDiJuYPizxcLGp2jJXE6BgGzjf1
QOo3YIhrVqfD12EPYCJuunvu3mkFDKfOwREuhLaBK0cc8S7vlyNQMWkSQKJEtZydOj+03OM1fk/Y
TqUJf9rV6BNhetPj6wHJnXQKgeU4/ThxXr5kuzTOB/SZqsmGzG3CKsUziMrYe2Bh9u52bT192wFG
mBYWWe17ngrPCs34guIDha+Z4VUO0HKNPLmLdPJ8UZW0PjU9r701mtMyAoMFpOJZmIfPOvXAodAG
IMUHYRQZPXXCdOsQoais4dK6Yq4GZImmCL5dpj7yHkPK4LE3LOBSoKbXTwMrCyRcA69wrJAHYkph
p7BpHM2xgEgTDtS/8l8UZj1PZevSnnhVTmckELIoVqDMR8Ia2byVhyPYy5w91J+PlnJ1QNGb9dHt
0YHnWljC21Hj5B817jGojL2MPoMiypPH1Wdk9w/9H3jIQpKYOPK+cC6CEQFY5bRKuu9Bi57JI3X9
J2DeuDFJRaF4yLqg1rySr+HMVL3nEIOwFrXU7oC8YJrPq6fyN78vplDf/sXf4iyT3SZsFVczfYh8
dJCLK3Bs9W7fUBxzaaqSUMfdX1K16ToZJVFoh4py8e3iGv17sxbYPrFCWH6LNkWLtLgaWI4c9WBN
D1yGa3FF666Nmhl/DVjv4Zq4aZnP3z09R7Na43JQ2e5W41OH3IRT0On5rLzv+U3qY7g6RAucRfWP
IUhGSb+pQ/F7EP6qBBFca8G5/qXw8hfcDjQXvqIiJaOK8aJ4xMauUTiMVZNA+ubaLfUO1Qh1QbtN
X4bpUz9CFzqTUEieHvHiaP1U9+j/JbiWiutSi1NBrFe9ftRsuWT4FOb/SiojWyB+QZ4PeMz3ZbJj
LkLvxLpt5L6QDKXdqiaSTVdvvs6HlL6S2Dkj8DYVFqTyM/IHYTN084EbMuaKUZHAXQ+tbPbgqlJ/
o7ecQ7YUUifvQlRsEtivRBi6ky+uxogMtZvd0wDZnzpTUqioz2+iq6iwU6BthI+VOJ6I8ajsPuMc
j0uHMEzWq0qrDh3KeoFFWvPjycwnchGXHZSMzCggrWrFs5KLTQpw1Fm7tcURNI2HxFNTc7tFBnbb
r9GeHoaJ/MdXBAsNbYnxGHtMCpv1Yyr4Qr30I2ntgHoi6t7549f8KhXDZU+114xhPPl1WS9IDKrf
jj7+i106zCaYZtlFLTfhTzI8TtbIkrFnl7K0stWlzvoQGlSJbNNgDOXPpaOnfwd6OsM5ievjE5OX
hzogo73dSMpd3Uc3LixhRmJrJmloISK9wyHivdI9Ejf9Zw77FogwS/g4/UksxOEwNv+92MfEsQn5
3btl4XlI2DzcmcYO5htwP1mFq12sdNTJ47IMCmIpMGHFJiEYNTYkJgnvnN/tqMP/JziJzCPZQ6MY
ZRBaojeqBcZ1IsCTUDPOX81IHHSDKbdshLSBbr8m9mpOvmgCnyJwushbCcJvCEGlFteTq77SLfyS
JZNm5NSLLQ1z62BXjEkpngZ/fE9gWFfSqAMA/nz4laNCzYziXl0taj5aKqSHwW/XhKEj5d8d57aS
TqDR0tymKtbktpiRWjybPk7rdaqWX4Vn9fZnCwHrVZF0AdzWMkMzdG+QkV+yb0X0+Hq0uHZsTqM/
dprBDFA/F5dko+YuRYdNrZ8sYXPTuhJL74vEBS7bhHa7EDF+NWCbZad3o2V09uoVesvHROJSdy8/
gpY0f/mv30T4JZWAlhHJRAXKPTDUCWqqT4igre3tu7gkgfZwojaQgQUNmavGlS1crr9Gz53o8c4i
O53ytYpFpMSayRVlCYSVFVtGLwfq00XxIIcqh2fffral716VltolQoqQLveBOUL6pMvBhF40WP+g
CVRNMWgRxXgLJUp1AeRrnl5/YxoTdlaCn+XL9k+5eA2BWWmZC3UiQU5UySd8TuVRcL+s2LoUM/8U
SpCy6AKunLZNcnQftPMOozmI0ESuAe8AGP+Zb0hc7zpNSrQvQGJYBvRgAYiwv9kFLBfj+RfZXlKK
ZmXej88L7j73f+D2fVyfdSqPeO/dS2hENHebQgKS6/PQBExVZ8P+adAEL6yr/tWYKJBWKjBjPCPF
4/UKpxGDu9PGYMy3/i2I20ycIHqU1CZd6iwqehB2z5Cvsz4pT60SR2N6oPoVXLMgM8jFoj9hyMKq
+4BU5kk6i15CB3NFdNJ0ywvakwnbWW2p1rRE0wa4MT+vLlU0LHqkQdMiyjVWHihLhMGx6SDcGcQU
QuL5HEBznZOfIAMC0ZVwwj4WTY0cUkaI4WMFhU+T02DReRmQ4Fh3+9zy4hjjec5lEt9mpTgGdtve
8eL4AheP8ccK3rI+jg+kBy0dolsIi2kMl0zf+SwgbcTpUAn9KTSCcRKs8RqXU1+lxozSxy/rXcD5
BguL9eeJ5vyuZO4HRWFs8v/kP10iqbAZsKvWVq1ml2RU+nNxSa4GOsrhucuzSwizvIZGG5Lkjgow
VJqZw/sH2ONi6s9YJlydGBo7RWVCOZSGVmU3Az/hDmwry4+EQXnx7SjRetJ4TG4GbhzVn6h98pyL
a8O2s3WFRM7Yocp/65sCe/PHgjLU4QT+FgcFSufUiXXHJciF6M90IUW2H84y5SC873yuy9peIEbC
mSKWC5F4Lj7eRFC4WS+Y79HuuqO3LBDtRLvDPReLbcRIzdJpBf+H1KbzPe0bcXA6TvlMIdHrwLXE
GG72McCuHyd2eA62WI6wvKmNMFkXITPqZrmUaBNydAqWyxPs1HHNbDox8d4ethpL4ZUdd+Hx8mgg
DnMq8cMLIM0jbJGKfdkw96YCB0wvMx/Af0m4DBDkhOmwwKhBdLc8y0xYTruiv43Kj0St3OpnyCDK
FYxSE085IeOLRF40JFn51vRa1i6tJPc0UcNyGRSmANuDkRNmVVpaMJ3r+h0NNzogVBRKKKfet5Hf
bVLV/FQAtA0i+Xs7FvtkvJfle1zpqeS6Salq9a32K52L1P8qkfDogrFvdDZK1AOaHbj549dv5syR
GKuYpLU6ddSZFOBm3oucq8NnC68zPQxaXElVeiT2+O1PNVDhPCugzY7iZYPKUpL71oOZ4sPLfZxe
InMTWPXNCHlWG49rEC6BdBq8HRIcqTUU+FpF1eO0O1ET/93rQmI3yzncjV9ld/dzcnLB3PyTX3zA
JPZfjQxLjYBqlmagJteOtFvUisLvlivHkJkSbur5letRmSxq+zRTsOTY86SX2v3vvtDH3YqdLVdb
uR9LsbgvXPPlMb1+JdWg4PSm9S0mG7TzNqplX53tyGppxEMJlHM1+g0CyauJE1YDcxxVD/6Nir9G
S1IZBK74FZgFHtkxxq9U7800hQrGZJJeKVOH7mSB3VlNGrym3+vsg2i4QGB1YK11zx+bSYNJzGHy
2QkSOL7DciTxUcd9yVF+7Ad2T20AWAgYcsy5AByOCQu3X2wLEWJyF2EGoFKidYC1jITk9o45hIhp
3yi2EeFYd+psWrsdP92oT7W7eGM0k03LOeo/5bcwEvESHD2YdvnZUtMTLFwxj8SB0umjmdJGLwpG
3EWItNOsn92V0n7qiQJ0NSAo17Ble59gfd1nF2j9DpPXk9NUdU7zTFy4grCRDSqgl8P2yhHMhlRR
RpvMcynM21JtQsN0x/mxM5uw2mlV2nEMBvbs6sr0p91ItrZ/ZWDkSHTBTvVKHca7KLPghNBRk5Pp
xUUqODThArYNV5dppZi3gpgGmJxW4qRsoMlIvUTVWW40/l6pIttwSHM4jMW6BnHfXWuAy6k3RMMj
/U7mmfx7tW7rcVhVBCBIM/rS2C5gAPGuclIOUYNVQSirwEbDszcNylDKoIyV55FI/Zep2wgwK61Y
6ZlC8L45HoF07mPlhep5VLFpmeACuvib87rbECAMii90rHcpbyB53KGujobpNgd6AYV6e7aHOOSP
o0kT5rKzWFMjMg9PNIHyg7L3tNrY73+CRwCHp3Q6CXSWu94q7mJt0MzvzI4TOutS0ym7pFKAckcX
WTh8MI/k1OCr0PHhmrx2wgNVasnuec57DvVkbPSauYRwAPPBFUgF3Lj4EecyGQSxINhlrX7USsqD
hNmGLYbOuRAUpI3PzyN5a232RnxeHcFDbj8HFqpIAvI3f9/EhlIxLJeiIZvwPNoeLhwMfPlXEa8r
jptc00cSVPNYD36JP7Boe6IURE1xfC9fZkibiPOq1Tpic++JrG2Eqex9gpfzdl+F9WiDOtQ2gYKn
h/b1NEzWZhvC7eVhHvUMFca0CGGbYaAPazVcyWvzhdPYstSlZZB1lKA/+K8PomYWcdkUwYHcARE6
EwrTKosi1bZLVilMISi+JOd3bVoeS9l8jFmN5RDwYpEqlPpqnCmk2Waey1QYxn5okaEjYNJr1LxB
otEmI+RwzyiPzgG3EM567COAmy1iVr6uR9Pq1N/1O6UJyUPWk13zh0p1jgs36X/EwEwckhJj13p1
F+POyvsEsdC+YuF5i7cfGKrhh8kD2LGL+K3q8OoNjVtd5WRXdeYRpE0x42BKBFXo1jDub02d7hk8
2Hu9e4M5vlPna2gbVVlXjZ035De+9no7LE9nGrs4jlERh+qcj0FjUzuwefZd45bFQseUQwLrnW4e
lfwq75VRg8sA+g2+LSrAYzGmJ6Fxppz0pzDWi11yUsOAXuZY1dTmulf05we3Yx/7xGwYvf5d+h8a
WtB+47vSh/MclV729jMMFZxkjRaIXSD8dz5bj2/u7q35S3GBvuvalt3ejdqiUUENSQkbvSG7lCSQ
p3TZXQJRBsGoAAtkU5FVjm6wjAe07TCrZqNFmSHHjzHHVCz2jtK3TirJUGhhBr9c/3GZ04lQkR/6
NMcGeh6tD/h+FBXHtdrUS1kMd6oUe7yZfScoIhtNCGKsjZNPIAF1m3ccuu7EdvDSiW16iJZLur2Q
7yDwyGrtE+YMPg0pfzoh/AhELKtCft+EBZMBCUxLMMgVLxKWIdpdPcC8IVJQ20IJ2UbKqOL6C4l0
Kobydz1U0avVbJx203OjzwZ3TfmuwJtL/7exwd8Zp/fqjAdf+T585np73hEUZbtNG7Q8kTafSACW
HFuMKot49UhjCS1noMV6ToyE1RZZkGrQ9lemMwwiVfdvOTFegjdN22baYWD5yAJcdHcF1dXeoYpL
jgl2RO57rzMoqiSbLTYitWvy9dVYe7ET8Vq8qRhgyB9mjbIZwanIgEfPQJ5ZUrV6uqm8SvXma29M
YlrYgJVqcr4SHiI2s/28kaWkV3Q0y5JboioRLb5A8HUz52yRcTHdX7l8tfK2HQxeVCqtFju4LokP
8srTm/85UKYrtmJXlNi/xv82PtaBaUg1rVVuZDZNK0y6w/LVAnsGYb24PRbRmwMaRdLSGliWog9C
C3SL1qtoa7oyn/rZZzZoKfbXPl8LW3fu1oBWiwOT9RLPF77VBGqBLFbyKXzdaqCxhr13lLvqselw
sIFWS4z40MjP+bTWKSvf4mL914Bwc079oP74e3ntb3lzZLCsz96TwVjbYlUNJur0Zj10zpSvZ4xo
2tVVGff8E1RKwp+9rjDPtzXhKnUhRJlkVW3+eSRKfjwvqcoTZiBDkJ9KdqbYnsp9J6DxHcZfrwJi
OWVvilzeyKCsuRvUTF1YWMQjtVSifX2ieEq7WM8pKoXutwcWdI/RiWF/FuCqiFzALESdYDGyxj3w
k8QdiliZMuP90pHkyhJ/0CBv0GTdno6M1kMEjcUE6GfLKxtcNoLLHX/y3dBeteZCK3Lj9l85d74q
02+tVgWQFHwYLdXdcC4pbVhr4OSdywKnkFK9YYabrtzDX5vgOIi//yQ5J4hRUSMihgh2uOhHZhQN
fB1yB6ZKKIuTaSjmsdcGiEThUXSD3dzqH7kx7WxJ441sxBpOoNLUF1RYKcwfqZHIMcHHrkPHiKD5
GXGIu+SxX6gJUgrAzcnTrhL9jIrR9LW/z2l5h8C0G5VapmQqu9U6du2dM1ppSph4/Tm/NxMkdF4x
vJI0kN0Yfbi336yLs3ACR5NVBpPl0Yph0/6ACJLeDJbjbVxUp8L4N9cVcY/CDTZ1lwxxUfOMs6SU
5/rYWmhl7rVnl7uqCImQ1S7dD1DDhkq9tvC072UVTFIFVYoCxImigzEMGxA/0afO1EmikVra9bvs
xGCLVk72tP/7mK20d+O9kQn+MiCC0SQxxijkULD0f7u3ApylZjZLD26V3oRWYUJqJjj5QwnWUQQz
b0aa57O1rTuiIw+6yxVguu4Q1vNWqpOHvQAD29EI6VcZHKP8XemULZgMXlEK+S+gYPx2rB/vcUnN
b/b12MU/B/mFmtmufPHnuxbs1NLNsdUCe31zUWK7xhluIOBjIWa8siwKP3TbD+bQY7CqoCEr9lIx
URpJ7hSVTU6WZ5m8l6oczgtDYeb8Cqb1SrD/N00sXGr8eZyvv7SbEs++qf0WRTtigMIjed9Ci2bW
GpnWmLp5OA1MaRG33//r/5kj/QDOckXiM4u/52kLDbf8yX9WRgVphQWNkU7TOaT4Ax6qwIv+U4gI
kv90i0uGW6W7tK32oUQfSNmS/+9A9TLJ/2EVnflJB6rHhyU/4Zt2IWh8HIX2hbbEGqFT1B98odBX
RXMuLdWE7/X1gT2Ewcm+oLQFIAjrMlkzdV+C+EMA53fADxMrcRlakU+NBk3gGnxfn4BgySULgoR9
jTGznBLdej3A18EoDsaiHMeWGp0LdZsXEmW6cL2Lvtr5NXKqMhyPf6wx1JW8cD7nSS6vsLiQtroA
KsqrWLQEPRp0SI65ODaV8D6+UmpgdveRNb1F2ZM8q0No9QfDrouL8PxaXiC/cuFTRyCgrbIvQYNb
vGhSWGLQTOKzRfCtiB4ITc8WmI72SvCr7HhkXxyWbXRyJhFzC4HIGbIcUHU9m9OFXiXIvvdA5KiE
w67xkmBdy1Eulj6DbyTDHkrYaZxKdJe8AE23jdc+G02mGu6vBHZSgkHpss1jcVC/vkEhW/VZFj+l
9Lsx8opRaDwOdszbDEfpUsWe7E6OUUC9GMpuOsoRB5PTfrncv/KghzxV90shYwBgYMA0SmIbYIjA
uYi02FI2E2d4PJ+av3oZ+sp/5BkTsxWNLWu+pxNe9fRezQqKPi86Ajj9Hj5lQ+H5pTid1wEFhgEB
GamsR4XawBBiR/PLsOCOHX7W4yxfeKVxOg7HLTPxVWfuUkGRakKHCQtpLx4B9Ez/SGwAZfJGWYlo
yG2NGPyJsKqCzx9D94Pg5n4cgQrvne1OtHu2q8shBgg08b/o3TuI7MjyaFMD4JcB/TA8X7PgtKrc
YCUv0fV/9n67GBEKnNE5h3fOyS13DI04JEhLXXCWwCzIiSE1yKeJ6xKt31RFUpNGX4A+1FP2pjCd
FSWgcjb7aO/7YyvmxOOnfCsHCAlpkTJzlKi97UvtwLuWeJ/wRsbxFUvyDsWdrKWUbN8EofQygdbR
g0c/7fdZyFV4PH7QhY6NHSOKrXS+Gx4wuyILWHmhEvOfnXL3f+7spBVO34VbJh/FkBkRN9r8jUKo
VTGUQLizPtYgGq3SulORsQonCT23txbPYJCVH3IbQnp/dnP2KbIRdZr5FdP7a+TMPkqxAwDHhvGi
ddhTnbHoKg+IU18fvo6o7ICrwbRnm83YDwuuzOcKeImHjcAu36oC4Q9xINvVIiIWyg2u4dQ8G32Q
6RFxwBi0SLBoIxOwqO9PlZXyrVssU+YF/EsbX7WQMyLabrb2MLEAQKtSBC3Bd8kPcnwjwOYF6Exi
NWevdIVKf7GQHWSx1R3wNAE+U+9SN8lfRdfCAVIxglleZfTf/FTLT8Mh6kxGb9ZY4ghaL82lCf6S
AbrqDG77sSBwVdgrGMX62fstDoYmRsUt0b449q7aQxjlZx2pw/c/iEEX0GF5ap9kK1hfAdrqhoqE
nzdMIfIDmL5nCXYruzId5sTOQTmRvq53SEeOnJgSIJxmOyAl6nYOR9LtYk6CJa4agTnjCJ5/i4JA
r8nZg9xfmIT+Oc0pijZLhMmoYQkjIL+vrtKQX3nj2p/cLtyvGPRH3yZba2Yawr6HlFWTdPafE3t0
dlK5Oy05xW4VpcN4lZpy7xB/AExEUTb1wXMYlUoLHQplBVKUMUoVolviR0VsGdKCcUNGDn/iae14
8JHp7nAnf+9V7d+/qilNLFS4ANM2/EFi6XLB2hVoKNaa8oSaTl6VHboAyVDNlyH5/u3Wo7QukgmU
rLz0O+2GjsvXwlHEM6BoMQZb4gC+NGfXvjTW1CNZAyEbcZ3fgd66eKjRCpwEjybUK1A4Ht46kDaL
OSBVaGkExARnnik5WNOYYIvWNEjuy3SGj9dhyTUQF3O+8bU3yzrnpRPS1NQYOyTAaQ7/iSCxcnq9
bBXjDwVuar/FRDo+qY8T/yCD1R4+yh68bT2YFYHIiNHx/LD7pOrtCt4JAfYzBeDnelUuSxfxMbsM
SycPbtHX+MoV39JgDplXpNOefaCs4xf75a+KPrTKpsm425Ir2TRxGV8YFCD11uWbsJKJi8tbufe5
p0X7Go7kcZbHpHN78BC4BmCsOW/YXmfMU100SIl49tbHQZYtG3mi6seqhJ+Trxv/5LQnGs7vra8D
uiNPw0QCJC3bw68mRHb0G8mKIehq3rg1LdWM46uanpOpUkSaJ4auYBB3EhLLWLhUF6RXzt5Q7EwI
XCUb81jrJ0E2LrR6aionhUpPcjnRUYzIRE1b+8aybeVkjIC/mGsvnD2ZoYb2KAcJglU6wH8wUqoX
3JxkWEyxDE/yCky01JEYaqaX09zxyDeWL7VpsmMDNvsvychuYZ0a56ReyOmaNZw3cgIsEkrtjKHb
puSHaSY52h6CIIWJnFmcRMcTSXhtduPYXVllVFdvRcEIYewHgFjRvFDkxVGvrUaQvfWCWJ4qpJ5t
71eq/2o5oDje2BdP2G8BUVJxKxECT6kSmk0WVyXYHajhnU89q3d/QB2qyihNvDRs8UejP/h64aE6
9/guJQ6aCbAIcN1NtwI0nxUGCN8mn7il/FH63Od3iy8trerXDcSLtgLaSm6e5cMYpY4HHOzoGEqY
K3wtec6+2OayHaKUGnU9aGSwMtZegXV1i8l5dNPQZXgMafBbp8ciVStjlxus+C7R4hk1l+B9fxOP
bLPYdgkpEpG6Jxq5fQc4DbmA1dNnmb3tUp6yT8/WO6E03emnWD5Cgdp+N+M0gSDl0gp14KodvuKx
WzBGXBeYJr9Y/qfOzj3W3Zrq1tS4flGu+qh9EJIDy9YaTfxxMatoCFRAAUp100O2UyWBsQvips94
AqLr/TAw5d33p/aMbWJ8/2wWYUw6QNP4kZrpyzII/8ojaUKJs2IFcnyVCLRJbH6aEJnoT5OHccqk
dq1IRtOX4q8Djb56q0KltCCZd+0PP/sFlvZlqk2cq87mP9txkmr7C+uvuGGtuYuaGLMhFgiUHRej
jiNmFnc1ukrxHcPOD2v+qwGxgCwzi75goP0/g9Bma/4VEg4U753yx4kmvUPWi8RaH8YTAu8tdFrY
AXRJhca+cwitTUNZNMjr2xju+HxP40iWFFbN+QFGMLXv7017R7tVJNLWo5JD77J/KlYrGOpJZh1z
DA08nmsLqV3M02hpe2MPKiJSVegxNv2p+8MME5xxlk0WbZoSqQ8f22c5dM2Z4qJv3FCwCEV19GYE
PuStSYMlv4t0dulxYsdQyrHmSptPYg7gInaUgeqEqjKZVmC9sQ9PF36hI+esQ732/U1cnkBWOwRb
2eWNQy2MLsy/bL5OsjlOZesRKCPTsK4E/F6TRWU4DY+8K/0bCkYgoXRsxMCuw3J+o0MlL1kD0O0C
0dLLUQ17/7ZgOOzX5O/mPEoe7YNZpGkTCzBvtDLKHBxIktEL74nzuEwroTVjqPnOdRu0+6vwnxm+
26LmmnMasw/WnVnvCeM+hNiJSN6SkDWwfEo5VF1F+Y0qxl9Ob371U+DTmNGk5vZDa4zB5bgGR5zc
oqT3pdOUQaPyh+rYgqOz5fJv0kTePLSIbfR2wG1qi3ElqRW11accbpkHwnbDm7wGQE9hYePSjZbe
mwLUNzHFk9KaQKLdeQU2FjBgB5BMtV8ZmsdWNCfbCtvJHe3Vl+ajS14VLir9FrMmVT9BRVdesWf4
rwsjUXdZA3NiXdVxcv18pm6y/KKJ5ym8czrQILoScA9CpD5j/T4h9uTySch5ToEuIke0Yk4+Ltg7
ZJICC3UnLNnkjBqRSsz9bK6S6cH1OLJiGK5DUwj+OlU2WAZom/ni4+fIpcx3LNEUtIU4db2SI+aO
MpnjJ35J53Dn7b2qjoDD/6+4Qsk6piSU/3LTB0jIwr2Yyxo7orWCESfZQHTJ09IOxGgr0KsBIGwC
VwJBjSu4NPF3FUIRvRSwlzAQpza4YwOdi/MNS3VF1M6VUhvjazSPBpkfiqWM64ps5jhATkUo1syb
S4reLnbIa6VYaRKQtRVTlfibJOxf/AZnXmI8QOw8iMYi6CshuTiuc9ekka5sRMQTPItu+8E25xNU
pBCKx620lWJ5iJSVClLk2ocflogfpEz+9HXcVl3utADXC3ysiHtK6hhPlGYzycpzi3JM+jnt7MjS
naPKEARhGCDDmxtw+4FgCAZ8XSRJ+4rac/AmrTkcs52Le90c/67fTtz2qnuwyKaaziH/RbltQAvo
O8pPtdWesvr3I3seDyX0FdeGGjxJ0PEOxTAwJ4kqLuge+OV8774meoH9jpsbqP2IrWTChcAGe1gg
aqSusIPt/5KjA5QHw7N0eS3vXPk2nwlmt+L/6R9PR4p49xGfu9uvuGsPej9q6V+5pXqbJraM2cfy
/ctiF/Vb7mmsDn0cIJV660SvvnRVsdi04IrHXUl0CosV018xrEwKqrhcLOxoz/TSfgiDqx28I41+
nAxS/CcTIKTz3/ywxj7GP568WVOU/ZLkuoIk1sATgqix0GEkejVl0WUdlzkg3mnDhLNN32rL9Ipw
i7sYNehPeUjSM/MJT4uGszkrv1RBholvQsO1Yuq5xqW5xbOE6D0sNul61wSEbFnC4B/5WgYA918W
fJRls7MZ5mP1Qoobcb2T1YOpQ4kABxwZvZUMSfBHoHKlGsNK65i/Vz3Oa+3IGDGQgm1lHYp/GLKo
LW5eiTnw6ocNTiLM5ns3ia7AEFc7lRg0g4JJgztdtBuBuWZvrNV7xNEGgrsl/ZC7rsX7Lh1vR90K
qDgoFG6ogXRtO2trcFgsahPwzBhhY5q+3xNErjeMLs86l6gAxPMXdHjynouTet3tgzkTffZtSrmh
nklfBT1L2OR/cwcbNCgkH0uuWJ/IEooPF7UQSlyTiG6hTKtyYwluPFiEEA+vNnj3Z6TCujVFFgUr
jOWiVDDzBxbCM8NGivajsZQvTEOz8OkDN212B4xqV5IMSlKzbABcYFvKLUyFTGo3W1envkCz9FIe
xt2kEA2ADevo7S4EsbFwstAetTE801K0BMmN8difOhknvfCMmjBgsLdbQpVWw7gv3RhgI6rcfOku
mTrvePr6romqVlbe8OH1gb66u4zHWp9YoLUABxVmYNSbSprLL0Q2qJehqbaXBVZfwSjTb7UZ7Q/m
Q+Vk7zDgfgByRdxVNtSPN6Gumv1Qtb2kHhVZnPHWoRv/1Xml1/X1aKYpyrL8Flsa2VcCFTI1v58X
D+9YgOkpY6kdS4hQU5JmQG13nz6bnNYKMksgHUz2DsISpqRJA0wqF+zIiyDXwbTZq//OqeMGF65C
gkXhcgB2CCALF29ri552AxN+YWpnKHmEzD8yc7zTmgKEUb3spjb/EOzw8qsXceQhY8QHtY2PdDLx
tXksphWQ0Z9a1dEHligWHg1PGI9Mu4nJlO6mwRSi/AEtMjGupBbwN6gNglTQouBTy3gT87TN9PcY
MYzX8YH/pm7SygKD6eCSlM4NwFEz4rTuvnyJozdn1ldI4FngMouwUN99CMRZOpdFe2u+zfeU6uJy
Ivc9S7HOksBPnL6c0XESy+tJ+CiH6UBkyZVOMmubBXtDRG9l/DzPrlxKFeHCD8ehOOWX0czZLXCf
de/LIXZgAS6n52nrUqily1D8JYtM8NUU+6+tTqNEsPIDBUrEEC1GwA06miYedRSN9tVhJl1EuI1H
qYKn26UkDxNmzCbmLJf4B/GqZrwwGf4MbstaRmRF3t3de8h+ED4ocAsti20j2g0Bmt+3+zkDAKKj
wu90DiZ02CV34H3+M68j98h32Xfx7c393U4GMmZPhG0fLnz2amrBvaltJYqjw+mS0WJ/xWKkmv9E
4OySGPyGD4m9XAC/2ZzL0lsPOHViZWgANSwSOq6A4TvyfGSzLw5IEKl1Edv8k5yGqV0+byfoFkPk
SmneOF4MnoI5A3mX7JmpvaEsJPAu90QTLIkgK5mgDw2aevHH18gMRUvkcluSjkABWyRpRWN79yjM
5OPB/mxro/ewCYX82NCH5vW/gatIZ0OL1s5fWIF8K3dEsARfnIO5OdrXFcnDc6HfuBjIm3wlQkVN
XXwppvSNMsDQeeR9K7XaoY0YUXBcBNyCRLkaOveZVrhwhGN/NO3ogFIvhmP+rrezYsOwwfT2gpOb
lHPVdck9jCDw46YVZ5jPpcvi4+HBlw2hFcblAxWKeHQssMbQXqnV4I/nIJONeUqC4R32YEDT4+Pm
r16f2IGnjFAKgYXZKdLMJRg/FfAae3Anp1lPCHJiGWOpfNBZ0urq5Pu89/PbTj9MJ+0wowWTl/03
gSEBtpSXF1R2IZvAg1jTUwovZ7BY22RxqjISkVkzhX+YcR42UpsrvsSmM4CMuV8BD0sapf1MERF3
dyv0p2fx4XVfzzKsnQv3td9X0KKIOj7lz+0dtjMEo4+umpeq4sUEfcHdc/6D87vFvUo1z2Igk7aR
ER/cG6B5gYQLgV4H6GgjbENvSuZbppeCgtZR+2fWA4y2FNAsRYzdngzgMryZ/aZNg8yr7qz5ecdf
dzNuvrEkMfdCEygXXsv8akTtF0BekjDYh5JIgIztDtmorXenvFGmejuHx0O/+ubd2crbtjqcxeD0
lR6yHB2e9oXV53dUDJKKhiLiPfDxh1G6c+eT+VAhZ6mc0WgFiK4txN6nNHGBssnoenpXnv5IojJM
1phPa8h/H6ZxD5HRXIvt+04FpEP9BdyVeI+lS2VjmrZ+smh1r24INbNxH6HhUI5DzbKEzGUzG34Q
AanTamn5Ni+sgllFgVZzdgz8V/bhvMViJTF55YcSlMWqSNHYAMVkgJwHZtJXakvXSXp4rSjjYQHB
VcAk/oj04TyhpXoNOyisHRHPQ6/ivAKD5hyQ4LogZzsFpb2jwLER8z+p0/98QvtLZCodgJM0KtMo
Pd+RmLLcHM1co1hQfJt9KUT3uXSlzxwnCVOq5HZaxseck2bVTIYr4BuqXuufkLz/CchdlP5FvLpj
H22HcQQUeXe8knSxVZ+wca7ohA9l0NkmdLYifo9JCEELt3a1c6vKZpU7q7BwveGDuHks93r4NjtL
XiOSTnSvNfcZblgmTrsQ3FUPN/vOf/ughzO2w4HxqalMGcfMt0JUCbJp/+4NTdS6JotkfIXLOkxu
J8TMCCQLsHpQ7fQoWd4kYWTQ5lkJS+/prH/+Mwqv+FKH2bL1NmVqIV3ClBTObP9gvQOH71eSRmQo
WZlt/cDefTo+YUE3xEagfZv9o47IFI2ogpJAxmmssdVMqx3bhPXab/z3ClLLsYZmvv2oH9r/v7Us
xHzskU31I9qJVVGLZa81ce3QW1qiN1aFzdPYnmU9QwZbtPS5v9bT7xqi+XW+ht5sCAJU4HqXz5hT
5IV0G9PEJsIcTRsfLPCzmd4QmLF3aw5OePe8trT+B22H5wiB+MB6YhLCbfKOI31X9tZYflyWHkNg
2vEdAxs/HFOBIXIaUPoXsWfkAtVyGZeX3mwcIcuaIQMVXzbIpNcM8BnmdK3MkK5NW7Ulp5Az8POT
xUKLKLb6KEtgAUwQLCSIJq6QarP2h3VMVFsSESjKstkJJxz3n4RHkSuUFQKRfXZ9PXVNGs2ODOzw
YMOTiamrDw0Da5ZEl33ionaYYfMaXfVFUypNWifZvPCYIgk8a/ONf5bPxggbtAYL7WKlyd71iMII
hT7PdZKp7un2aG0tpdg46DAqKz4PBF+ERJ8jjzOhSzhJ15SkEcpQ5esjZVla5z2LFw+xgzkaapgm
FYb1kJZkawXcHOFaQGFtOJqq+6DlNic3S+aiIBkI4qsvKEXbZdxi6x45ANjEvnhdwmNysr5FKruS
CQPadjXnXZNq9phMiMYgZ08Ukv0BvvCjRzFmJZsAx0GPfgSCaBujaEgExMOBV2cupT1698919N4X
0eXPUph3q5DX099bGLbCXuXHzLDfs4T2qiefhbjUg0G0/EBz99sMRluvLLzADZWyqotiZEnSSvBV
Lu5rRkTC1/ycLR8PE5hGO6KdJj4dirCoVBoMvEpF6tPa3noj3BhgLxuzdAGgy5R65RXN2ZMetQQ2
EVBETeh0TAjx0BOviCLlPjFVgb9oZKsJdlJ+t8gp8+1p+7gMzB5k8X/7rjJ2McZwI8/UaA2X6OhM
PfX4VpW6nT+LuyFv7OeRlkgEC4l7+G7pxv5qbHD3e1vj/pLxN6j/DpBscE3qRldS21pMFjkXyIsZ
1rscZSl3YhKUA7n9j9cf33LlAuYB+N6vUvpG82hArt1ssHgMoFKTFDoLj81+BZ4WyFlZq00XjT5m
oUud2gyHgOtAZoealu3NxZzLD3zyVnz70Bv4dIcou45Mrq+uZZWP7KP9scJW9R5+19w2dJktokyt
qiwpnD4McSCqlQnNVxldGgqVHuU1SI8Yp5LioF/NLSh7ITsnYJqrKgoQtx8+qGE4oTnELji3Lk+s
uwbFeYyceI1rr9qQsnQfWsifar4uF9EoDGDByAa3J41HTI+F0aT9iGGkp9Vk0vfOyy9QgFs4G/kh
aR1kvtAOObE81iC8W+Gy/sesIwTR20hzw0RxH1czYG52UN/um6xfcM55B8Qlrn63S2u4mC7/laiY
wP5DXk6ouF6j5Ep/sjhNHzo4Kki4jiUkmsdEtCGIXQ/e9NhA5l9JzYaVMIpNkaodaW01rsCZIzdW
bICv6n+Ipq4GdpZfbvSXXW+PW2AVpA83379IOVPpmCNUBc68Dyo/CL+1hQJx23zhHWGJu8pPxsS5
pJoMj0t54N5c7m1sfdR1fbabUIM33e75WaszdBxO3+heruYZ9Mw0Eb3zTFSyyV1ZzJqpPxqTiTlF
C3zDx00SFRUa8UEhiWKQt5mXVGebkHlsWVqh2S5x7of1coPT8zeDHwuKVv7K3i6ZCjsNwa/YmeWs
rvdDSAEMjV9sCGPUp6sSTt8/xYehODVYGpkvxHajAkCtkkILfr4ACCkuinNiPTycyaWkBNuAl+BZ
xVKHauKVxJRUIt8Jjl991ZutSQaK0Dxls171RG7NOjWE9Fv4mKpENPXVYNQTQDZcHKxdm+dqIYoX
qp8BBeKUrhtyUBT1U+YQtFVfhy1CwuZVnymwv5Eh5oPf2TC2Sxs21H4PE5fK00RgeRg03iz5nXtU
pWfvRhrPqECXAouS/1INxL54fHkQEkIdY1eJJcS7KujSbBbcVMNo26d/Nn7/lRshULbcUAt+9OGW
VGxYne0KAb2XqzkWw0xmVpbKiVpLT8UAjQVzG2Ktd9F28yNM/DpKEE2TRH8HDEh4lqpjx0BMuFfl
X1mNSZWevx1SAVPA9M1kPwllxM8hFhiuY6PMEiKuhbJ8k8ygnGKEgR4PbHY9ympMVhZCVVX+EisK
ceMBJa3JnhtlF351LyfEdu8K4iN5pc3CDaIBy1NuduYV1bPlVnxkKhiAhlEfON62Q9SD6zgvoWZQ
cYcol+n9WSuyDfe9/XfG2KNptwxZwVrUPY1gX1NbqFoJ2Tz5Akc/D4TXqRByeomp1+3Cu1kcYcv9
W0czfO1dx8fBCf0KRVHVOq80hLsv6yyMR7jk4kE57JD/VK2Z7NsF1MW7iF6flFgLWp56mlyIUFsE
yVXsjsuA8pbFJ7sGpnNQfXXMNcdMBH+ZSudDGZykryaDDO/2Njcvcv9eAYqQsOfO07TVuSeq5ttt
yZ5bPTUh3diD3n6BJAMVb0AtVSt3yswsahNFoWn/EAOSLYuE0e/bnN//GCzna5t3Y9Iuydn4zVks
CzPPqFB2W3C9Up0D1YOjbP7lSCjxosNRSjc6KChb00Ni1Pprh3kyBi/0brLkjDGAt2nWVSWwEgh/
oQU2CifzZFIAwv1MbDcIvt8Hbdb95JXNMeiSMbCtlLw5Gnz/1lTHI5EndlCIp2r9fxvdICwWTXao
kT1DDZtRLrNB0SWzSo70NaF4Q53gudxqyNkH0bic4b/gKfIh/1FeBM0j87IqCuoNjerBFYvgufl1
07sSe/b23DTli+DOBGNp0O4+egXFLZANeZCCGxKovabH5ryfw3Zg1gnP5rC8muI0dVUMy19wN7Hu
XqC0cVzCsoyGxjyBhpcG4fFW4JGLEFzWXhiSZEQxSoT8xDdo8FTdytetkMJnW9cihl9vxCEeKM7u
/5ONt9+JPZmd+KkZwpU6iU5JQcSuanOwM2w/0ACZGQk2R3Lw2wwuNH6+uKxTLvUykly4STygMMVQ
B7LWkiSpxuJGeySa2wB9pVGcjOYholOK3S97AJlwolzBdq8X3mr8BlmnJElgArZLtAwT753+Wkds
iXNpVZQSfS/V9Kg018td5lbgvBXZH7dutWp8QQyy99g+gCBkQWf4mYw26xnV9Mc/V+gn1D+FTGMM
y2U4bsML3szUJgtWQ/FZDpnrzGPOibzZkubD/Q5LWYCKN2iAf5EUuU16UOvK7Kb1DNsv7ugQ5zhx
QLTLGzxl+U3nsRsZAvv1hJk72fUrzbklHA5YaEf7asYn52aUsrCaZoiq5rWW7shIFu0vxNCfmks7
N2P9MYgXURLpT3EqycldJzjYVj0pwGOAh5/XNa+Smf8AC3pc2vvm+S5I0EUBZWIHYgJtBypgOspy
BRG0y/Vl8BMR9YQXaGRwdXCOYgd1Fq9q1mtFglia6VvM7YgWirYf9Ufe1dqAmTQsDQVh7bBfzOGE
yIxu7+iYV2qGZPVfYtMeRsUGBO7Je70Tr9wgpswZp4z2DpDMaSKil32+PxDDxyKbs+Ctjh2AAVWA
jea08secc37Ol/GNRPYKAtn2wLhXrgSyRI/D0/8+QVj3ohVh/5GcxG5nkugN7hz2t3RjeSh11mSl
gkwbJM8Y3P1D5PoJUSqGiYaonO9NYD+SO7UsHuuyrkud1jXP2dmDq2Hv9HVbSMOKhwUu13lJ1wcO
ca0kpYxpi2Hi6PAdwWcLKEZlYpIN6Ko4sJQ0/QnnHpa1bWhLhLHxyaf0ba+oW3BjPcUcLmXBGFOe
/+dETWGIWTYtJntjBkq5DA3cmlxcljWiLAoCTJqLzuQPYTNI+6egE7CJ/ZKg6H1iFF0nevJFKPfp
Z1P3T7NXj373suvqHzzeqJzbhkQrhxNkFwS9V6EmtHrsKarU9RFD1B59sPL4o7jY8wPZG1Puq+ol
qfKXdsly+KI0J5tNGwh5Sq/3lqQtvpXbOsZAtcJ7Hhr+XXMDJ/jPK1cqoaYni/Tw+C/RYTLLa3nB
L3Nv5FLjJMJhi02Yfri/5MWgRRe9A0hfmYoRfNXhd54BZmFsTpvi92Xg8aVeQCLJ7yZAtTtzQp15
7OdLJR5SqjB+bznrm+5fWz5FsR/8NwaYrSjPfzNT3ScKN23BMUJw2IY8c6v3crsi36rhC3hIWePT
Re0sonWYRbpDIer3MF6GChn0Xz4m+tv4hl+z7iBHoTCF7WptWR9u7ewkfGv6PPN2ilEgnlsuWmC8
Rkn5uQagFDIu/SoWD8rylSJ6gQZT1y7sY8HlwGJYT3jiteFe79L3HVSsyH+hLy1UM2GOnbAyAMyf
GMTxuBCtfaaSWx5w507ftX97AfA4vlgkJzoVkSmQNigmLskTV07PhqnDqSM7PYj2t9ALkC6s2QDR
xmU4Jb7egfegtnb2Z4l9c/LrJAFO7aV79r/oNNWQO8vx5R2p1NtxKb0/jOcgHSNGktHJWUfLhPEq
eJofufguj2yRtp0GC0xnPOfGSE5cdWkjiHAIGTpUKnbob0cOcEH7HzYcaHRic6cxtRPiUCpXy/BE
oJ6ceyeuZQo3ZRc/tDDd8KVi8V+C0cSmLfgL0mNV6+DrOjTlIXdMVlU45jXU2BoikZCT3ybEiBFL
J7tqtLszq2CoVRp2PN4ZegL7L8avwW4IcNgIHmTyujaGdZZGraoJQRb9hs2KRiVYn0kagWak+1OD
v/D/16RYT4zBVuetzJVzcyWVUIke4Tp4DtSoEY08nZxOB2C9nRmj8iyh9ZjWGcqSPKzbuK/O1ZYb
IA0p2mM/EO03fz5gqPUmcqq8up3IFrYA2c8PHo9cYkhy5rAGtFdRzwAdUJIVNbigUOjtYHctn7aN
entlqFQIw1PzvOXfRsGBJXGrsRUFm178sQN+Hyp/2AOzdUmxCe1sav70/eHSfCrZoZK47xtxO3Co
f+wLiSebqP05g8hYX8Y+7+SHi1TV2FXun6qSCTLOzRpHbgPMSKl/8FMw9niunUuATxeFlCgp67v1
6TcWjWLokp0rJba76aRzOVECKhodOWM0fiWvCoJbTMgf2Fym9Kn+ziwY+5Y8czfO7fLORmrCutx9
6bQgI8FpB2IpmEqz89yCOTHK3lFshKMVi4D9S01bLgNDT2go2FKU8UxCoU3kkuCqsYGj/AHRxOjP
nuJEeBVc66g7IYlaeL5Jj8N/es1Q36hYcjji181mVJ0U++TAeCovmD2/J3CHUcJVjVe5k3k3uPiR
mwwwoL2pzkMulLqEFh+uZil1nw1UXy6p7t2T5NmBw4YKKQABHttbMBY828ujmwfaDNlnUmIk5W1z
CD4FBMewPtJXMldqnX5a6KvDL2idSaXNSUj0h/XLJu6BFPzcVgUxHOscckV0PTy7kljDtmvKlMw5
E4wumhqwMHGHw96QCTkPLiwUyQoiR/HTqt8GxU78h+8ANH5pEQD4/9wBbxlO2DQW4Uz2HcHIKESd
1XV7aFZsJOJR9Eb/zhYUn+CtNTRc32QwQTEtn2GGd2hiR2pIhnJ8IFo4woMqJwHOP+O7Izt1nD3g
6jq6PpqbSd31rgmxvBtrG2LR+eHikntsRTjFhH7TW4SXayoUH4fFKUF2r5fJ8MXby1A4TfDhhra1
fSq4vMV3j1LvesAY0LzeW4zyHuGycVCDJ4OuLzmGC+K3tEGPYjL9AfAcfcfVLleRULb6YDz1B5Ar
rRVEAi0zj3//KyiTiqv169vYmK/jo2olsgLtOlOwgZqCrF4a6VvXdmCMq7wOpDZ0hkFBZ2owBFbW
G3yFGFWUyjrtbk7Pog2xEZCSZ81p0olP3MuhP3IHhZYLFb9xKV+Y/1U2Kgx9JBUGOUPQKdzno/7m
jOCGyVFpNOeitELBw6kzqnU/jLrN8e0KvPrRSknYeQ1SCpznD5fPcG02p2w/FCES5+ZScSQf5Ffd
VK46pL2Fv3woIfNFtPnP6pKPLeIeb1bWfj7THuExGKPqiRWRCX7T7sR4DXIUZ8arNtzM5ZBByzbK
+I61oIcoswqFhHeNlhxsrqojuBD9L2tm0Ietq9oCp3nfShtNA4pWpx7y6h2LRcWgH9v4o+bTCScQ
2wUUfcBF49gc8o5OmfeY3rthC51RTDMf5eRM3e2XO17BQPx+QmU7Dwd6YLRaximv+G/AbHm3r1f6
0L3tWmJ0gMz/wEKQuWJxN0aCAQdUMOi9wX2CUxtDIL8rATgHTRdBHSgYsNJny5ZjMfc/JavDby+o
bREsKKMhRqaVNRMewG0R+6Sujo0Ez3ql4pRMawV5LwGEu9hCHmZwGvLDuYUJwhzVCLlrhXq51UKt
sB2ws3KOuZicmpbJxSSiJ2VByf7D2LSn5Xy63cTNpBTTcnqDBGslZ9cO33v9pwNotdo0G7uJIxhe
sSsUshFuZdWtEu2rYC7gSp9oiG+9+y+ckPbXpGb+q6yUN3Qws3yDm8tWCMappvVnPEVdhpRhujem
6IHtv6b8HFfNgbXfvkwbEfhU+aUvxWCYaBd6JyIoidk9Kqfg2D0qYlwccv3uDfma65KGeIhqixVH
UBQPzCvcHV0P8LwbyHuqGH+z2PsrN9ftbCDds6pl1OwY15/Pafe/zK1E6FUWUD/na8yjEB7UPOUo
y6Hb8jw3nXA7OqKO7/U+ioiQ1ZgLb/p4MqigNCLuFDJXPAqcAo0DQzMAHwQmR7XjOk854IqzQMZF
h3YUtRvo+kgI7h5Lps8Admw94xKc+/1WFdbj+m65Zmy1vv0Fu/5eUtiOH0osgWOQJRKQb8cKQWsO
roAuE4V7TOrBR09iLrz8ehkSNZxFULrqh0cdUHyJtt8e3N2suYdRF114zUyQ6V3VYxOUNYWPITKZ
zEoB5f3ouI5cskyaEGDSXpA8bdHdMVkMpoOy1Txnu3SKxoIxvBwy8VMvcdEQeDXjKjK8PByspItq
KlAdNirU39IaFEFLFo+Snjpy3X9NVd3p11UdL7CmTp/ug/Ol4IvhQFEdFNuboLtK1KWK0txtV0xH
XzzBzyoc40FnPQr2QVJNrkAgn+GYo6grYqoh6u3uXF8FIqUvj7mm85Su/VckEJx19GVfHaXq6yEu
mAEcrUn/TCb8KbSvIP433z1VNCxQZkDjdXAE/7DCgVFTLE8VqdBuD+qd+iHrePcaX/gIxE3TjEl4
L3VQFRtaOfcwTyu4Wi3ZoCcG9eJ1JoqHt45GZUILLGq+x8z6FZWdYWGRe6SaHItbS24+s8dy79TP
0ifkK4OiPQxjllXPDB5BdtMB5Q88htm48eWlFxm+uGpVsgZPEg9LZsnrdp+bwnUrrRlbMZy/qJK8
SaSldVhKYfVZBlqu+d2qKV6nIQj9x3IgxFI9SzFx35lpT+dKV6oA8P7BHbgW9+LlrSg2H9vHipUo
oMLICkTBwn/CUh5aPyd5FjaSCAJnb2Dw7/KRIgJIOx9a96aS7NludP/ljlOS02iC+DskzUWYRKGq
xDDqGoySoC2Xu5g37gmcjibSxYF5xwMtK0lQTeiKcdk7omD8x74JEyCrphXLi/E73UL+aKxxT1VF
bGXghZoLJ1NVL+L4t6WwK9G11sefcmnKSowminoBzLgNkEyfvEG7MsbiHrsYdBDUtL40Ykxw5RKQ
S90LvI4WoWT8kStOa/A0TYBSkzZ9wdebGf4/IpcDAJZIZ9fEBGVFMqZHWGnSG6/GdIFkKEoOAj+g
AXQTr+qk9MFYF6r7RAXb8vS7qs24oj2araCawzDg2m8n3VFjH1nrG0hCsZK8eE149nrL0CfjaVxr
lXTjWybRsBsBwrbn6lwI0P8xQFgHWy+h4VPVBcq/ZnRNdlZA475caxLZjIQr+nDZFyExhJsM7Pme
UetOtLV1WjOavXz/IdxsiB+vrTSukevcoijB3juEjhLZTN8DrZn2L3KxYEGjIrtHwssZC+8XZRAE
7jab3lWTX3l9MnVi40Xvl8rnZ8Yj9J4eI+PQSzg/zTN74HmTF84Za5UBW+9wxuXwV7y0IvuPAMNb
ed0gKOulYZx+yBzxPX37JAkm4tHNyZLYLC7Na3R3mWaA9jStDRK5YPXUA2lWDKHiY76/EhmDKAZ0
43lYB+oNLZNheeAnM4Czt6jAL7AVJQeYnsk1nSkgYcYor3z683FKz+g1kaJ8Lk329gcAfSeDWehY
4fX5MxD9WD3l48JPIq2aM7Ag8VkbXDRlKA8QHczUurhyrNFd9CXaSV1itKPlOtIIC2XI62gY3QxI
XxSrpzxqP3kRL+nlUPtuj4t/eHRYFzsJnEgbRtUe7N7ZqucoQRIL5PxJx6dwphV4iIap+gJ7ZvHr
i27xOEampxMZ1SdZISWVPa20qlFK3+8rAiEjpqZKb8CFptdzIZgGQrWA8w4P4keKDiy8QiinC68i
74bHLqUz35Uj12wtwRdp5/lA4IVz+ZkVDml72ZR5r4mIdS0+grRC6Kmooi2cA6ZBQpbjwefyOysn
XhpACc30vlgPvW1SrYLP+3z7JRtc9ZUxaPRHaKxpcXnY/UzzgHuMLi6svTT/+7z2zQjaXYkBw0W5
Ukx28bBsE5UVLJb8Efk5ngemHODXPsw80UqEEVG+DoNImBgxKPuzHoAd8tPjPq2ivZjEoR2ddBaf
m3WD3G9ahID4xwPK6j7MDjPEeCVoCi6zfobNr0UX/x9GwXv/Ku4A4Rja9/BvBlvV6Gk4WR5w4eSk
uLCy+Y8WywNGJYPgWd8tkQi33ltuNPWdfkh22U1CfIX0F5UjyKuALyGPTrlbZnwaUn74HZgTmLXL
NaPrMEfGlkEXVeNAKsFFyzaCKvMYrMzPhrZA2fo+FInpB3OtPav7IKKLL0/iBnMTNpwVuxwHgkhS
37xCYjLKKVDU9+yS18Fq/pnxE/cUw+JSxaQJW+rYBsLbngwcaWfuf3rig99ZWaKgCcYK90A9GOU7
wnl7E7xuqjBPS4ijYtPjmpoerNt9rPq/MOiaRgcCXixcDH0eVq6S3t8xwH+rrQrjN4ZHvSDyMKsx
rdCDkMju6qN3jF46FQw8EBpE4XQGdsDxYjmzRdpXnoQEs7uXkX7ORpfHw9PMfoWGdTRDI+qFUk8P
NIC2AMgRJfK96e7ecVQ4un/hCKzgncsAv/ZzMtlRu4u9geElQOSxMSL54AADq0NA/XlDO6aXyjUG
kD3trPIDYAem2gdQPqkfd3atg+fSFA2N94RhwsL63fgMMIXjH86zlY74e0/dQER+kGlxDp/BQVma
cI6zg1bEpyBGYXUHlzROtaF5/mvhQa5c8VEtJ8o5+hNJKJ6jSmgz/8S8YU1zQt/RtiYyh8raQ3fe
8c6npgBIL6LftsY9qECQ3lX+v5E6t/rc24OrcN1sW1bEFw0/25Po5Ji8Ubgx7Ib2knTkPPKTj4q9
Hhsn1pybMjkBgRSK+fKGPPHnPw0YniU2WzMU5h5/MfbePzd+OQFUCnlKgcZaTa9Pel79FALjq0Ro
g7n8iqD23zb+dhlIt/GbCbuoeiemC2zkFt0aHNDZ0KXWi4/zZnU42QBNe8UdANLajmxQctOakdJD
YElU9fNGlaGIQ1jqM782zToDsBy7O2jEosl/GsEbqWr7FtQ5TfmOKyl2DKcIbM7SvRoTlBOBZzmo
ExROQ+JbYCA3qAA+jJw8Wr1z5NKspv59k+8/DhWYhxHOiFu5/KELmGjdkERG5nCc1veoy6PsP6EO
+/i1BSkLdjFTIEHda9A+2RQSuzR3pBiEb4yH9EZo0fwSnv6dQueHehNJosa2ub6HBYWEuTaEaUO3
NS20uBQPpoVlhQcXVfAMPa1g4+EmkMPpYsIIbYQrOQEZhmjurzm/aozp+uiVzg5V5ZWoxWhiGaQP
e34H89oYN65GnuWHuWAByEcHPIUvLliEt/wyuep5A3uMs+811d9Z6hOaJgI6/cWETBzI9R+KmfEU
Cg5qpPUQsDrsQoO+OoBiiN0nzB6kgIY1HF8gbtciGAJ0RWVBz+hIgfR9mnDrZV+Bje/gf84kcrKN
Od8HfbA96LKjFTLFo6qiU1V/bD9AFe6nqLi90tfDSFElWiE740JLtmtXim9IZ8KDGZRqpo2ftwOs
BlLDftQXKY9t1F1Sed/kO0/QlnPCOnRk8GE+6ZFWrEUKvLPkbnpfQr62YkoE0mpp2mdKLXjGI8hQ
cVd3AqKS/SLgsS0D1lMGk88UeyxKpP41+FCozu19KyALkX+8BLdXnCC9GTfRx4oZaWy9aKllEl5/
RsF+8noidICU+sYU7DkdFdEq3lC8c1K3Zz/kE8Bs0sJ3+BA5oBFtmdG9rxc0hY0jE/OLgqpjNC+o
M2tQ9i59cR37PXUHCdESYz88Vhggax4+JW9MxH7v7rC3JqKImC6YER+7/uRvX5sWRmU2qVo767yN
as/tkCcbX/5O52HW5iWxCug+nCh944vgnwHv1J5WaPZIQHKs0AD/dkQwfKFpVfFsotnQia7U2z+q
YS7YKVAaOJVG/tSHRDaDh+SvZGWdzdMl48GchBdTRvv0RUli/t7/zMMn4zR805Xqzxl3qRY3X9QS
4vNIBpQLNBogd6dJeDTQAvSbqMIyTYTgl09LXIpnJxhnnCoP8TIgurp5R2ROeZIzEFI4AtLDykQ5
J32QzGOF3OqhCTIei4qei+ary7rGoE/D7YdYK4StIsZ4b+9W1Tr3rt81CScqms9cRU+3WNmi0bNc
kizhgzJclFX5FvpRRE1SManNlX92X43BKUZpKtbzgcsb48tpV+XcWm9vaJu6+09LUC+FcgLltTYl
uTnAgVJkyhB5ioIYcJk06li/QnJK5KjKHh7xkQ3Whwll5oUGJRgqsXW0K9SCufx6q8IAIfaNwK6A
tKr1bLfq4vNNoEBn2EzDslFP+c0kIZLmbVKE83+hSUfxBg0sly9bjN0pw37uTdudofTyHm1oIsNe
r+YkG0nbKoRXEY27ub5QA2Dr2LrFnjgxRzTlr2hC413Ll6FkYlf4iT848IGSG7EpwqhFl72ee7TD
FPc93PgiqiahkSHXeiiAGGaeZ+pPXXMVqjUCN8XHhotg/PtHPZ9HPoo/xUoJLAHY2Agp7POeAGdN
O4U9R532xQ97oVThsQ3g2OqCQnxrJYLIFhMZLaQ6QabHM7DZ3IyefoL/Q7krZ9sMEJgcBhcvnrie
zWh5XczN/TnBj3RDxgBYljTQpQx0u4LejVt909dzbwLI+RD2i0UX1e8snyZYaO9I8mTNPzBvHUcZ
TErSljwUpaa58V01NFdUNB3EbJQnzW8aLpQ5V3RHDQ4rv+cvc+YXEDHEcK+lkreLnSiHyD+gH3KS
Ij0w2MQinzZ1qDos8hEFSNLli2uK/swHCtzBt3mEdiS9nuauy7ri0uGmv1X8xyNtCPrEt/Euljt/
hlvFbT7uUeOYGmnxXXTDJHGOf1igtq5qrO8ryZUXXWoFGcgSl4cp8AU7vk/blocGKxr72ibYAmC3
K0LeuHh+TO6jT35BBNyQL5LV4RdvhBVF+3GEFYQlFPthGZ+bRdvWcVl+9xf0oKhCnVXc23Ehta9g
5KtvbqhkUm2KZPiu3evKBh/SfDyw5ymdZVYe/rX4S0T7RtSsAbZi04S7kD4LHFtLXTicCbVH2R8s
vG/o5fcdVmUa/yZyf2By5KMPyyA/+b8ggBbnZ/RY4sLEQ0C5WYa/R3ap6WI1RYdlPR3ijyR+F+UR
ywupuoy0GloWMqtHvgPZuPtMKPN1ihVLF4wHzoxVlna99K0BU5STKoMyKANfDpS/QNsBYJmXG0Qk
jW8eatHwdbmX5obMhXqh+1NCZ5quGGOPlxORpUQGM+bVsv60Hh3QcK4kTA0FvHU24kVFHaqn+5Du
sJYqjilwWuXYefQ2/Vmu95m21oX8Y33t9BkfcEAkih4UCZ0zg+xErOfvQTYvy/5118El7Y4aopyJ
OgHG+wc58nLSualuPOq8YI3tYb+VLdI4oKthsoMgI/z9oW8U8Eld6PSqj29UYCGdcb5q3/rqU/Nk
+JdvQ8v5+mGWNUissYpA4KHL0yYomrsgTPT6fRgIgLCO3liUwNJw5a5nzVIom8VARQDCCNvtNlnI
A8r3BKLgLc9dWLXswsQcgA2rBmy1UxiNnfGmwH9gBGesDLDuR2h25FhBk2hubIXsoRfZb5Kns5qF
MMG+jaENN/xDC8K2yhJyJVsJpVPYXTOkLaqfNY9PqEUC+h38JBJqUDxwAEnosVjEcg26RZ3DZiPY
OhBSazMz7rSjMsjrJb5kqLe2axscYPAt27E/QOM1i9+xBPABg0MJKyxS2bLG5zE9Vo/XGWYhCB5+
qSCxsQ1M/qdIYhR/IJlEFT1uBDZwP3JyYc4IUpG9lqBgGtTU4Xtb9RpuCJ4dL9feZJD2DzzFlJwB
23Vow3Tew4yZLIyeCFrEgMxDOfIwW4g0EBiegfdtjVqFvnZ2FFZ8aVr4lZzKt/mRleBz9fMxoc2b
GSxWV6CS3KwVtlstmdE0eb8R6j6FTdAgiN2x2pIaHOtJhoXqqNlkNWY87vGU9vPbn9KGqe4I5ydm
s/UUCnmsCrYt+ATUyyPEIHUTnNLdcBMymUy4YWzi0QhZpeb/9Vxk52ihiXS9WROgPg0LHRXUbg/d
zjPBXisRNA3ALKxryNTmT1mLzyGav6NzIgqYstxM8SHcW3KcjpEa3K1q1/C+WvVsRuf79x72ne/q
xIl9l71ITZ7EkTgRFyCURZAUs8m1ACVFp9343wHgNcN7jtw4qXaVTrrdDUpYb4HQoJ/eMdAdo3xv
xCS5099Wy54mNuADI+osZsSTJ7HKPUNyq1rrOoLH6i7je+J7JUBy2TZ7cmwpaPb3ZSN2L3GOL0L8
n/c9Ix4koDxLhXRvkBXTu694m03ilpW1C0bl532EXOuTadTRz+HfvZMla1wLACkr4Z4KeVQXF989
bBtMYufaTW269z3ONDeeRDAxu/ZQeBr72g9mtWAo0wl0FX740sPTDG/Gw1QAS36Fxyh5rZRh3IGv
xfUJo+UnLIuqVPDTiapb4TknZZdwR4+qMF1AdJNrj6jgZ8y7+mCLf7rFpqhmVcJLUpysAzjSnkvU
gNpVj6Ze7f8C7L38btpe+dhdQw+4OFXoXQcIuGD+ebEFRk/Tuuc9WILVd7XaV2G/aPn2Z8fh0f3C
1HG6viXW+2Kgejeidxa/wONBgB9oozTLSURrrlEt/XwWrklDasD5KBQugIMMq7rw67Evq4WtpA5+
jE5lga677OKC9pn8Wpwh7W3tCsOy0vRXbKJ7CzVfA7lq9e9ssoLby5mA/aeqZfzjDwUWDK+/bxih
lMtVY9CB+yUldMCXTtDUjIsf9sdQMGOVvk3FKq6xVuKLi1u44TKpM6O+4yPxopYg5IAl52eXLnDB
YKojWg4jNIaHneEVIMhj6epon5OohumkfqmEzmyXcJt301OZdosykh2gnCQnsvVWayu37qNh6gtp
deM3tVvr0lgLL2vqPEDJsGiFRfjqK2hODlI2O7ElDKW5huyOsybhc5RwrPlI/EbFbYtee1MZTTIZ
K3L+WzeTZ7DiBane0XvXGHmjex2/O5I7P65b8C2g96YeftU5xkZ71bgWClb966HUIUDjQ3qk/1b4
TA4w8Gly9/1QgED1xbdgLouS0Otk3t2XNYE4QKIT+66VCk5ZtwtLI4b+O1iA96XQvdSbyyt4zruM
Kl5JK81QurFy83t+jTs1EOr1R/w8X7QphWgU/XKgERjI/LrbqvZoyIKhHK2Tsy6nwVRnA9Oe8FCE
rOZeFP3hWEb85osCdBlTJoIcmv9FGknCq/XPOX6b1ungDXKrgvGqaK60CUqO8JNFmhD8hq0ZV2PN
+zOqr6ZKILFjEu7sIPhw+P88O42JgcN6K00CrQzs9ghyeKQDJtPzPHdYr7LwG/HBk9s9IFaku6m5
zOkv+z714J34QcoZI6gkontL8/5GG1doAdL7FSygsQmzrnfrru44ePiRFROONFjhUq9xYLL0m9sj
bM1FrhKFgA3gjQF+O9I39dG91uQUC1+m0D5/18X+Z5aYPkb6mfR6hhTpD+Ycp77h8da9+6lcsOod
S4TD8OzDLlHbSqKXmQ8xhQ/r24S6E6VsRwE3jpJzgv7iEMMbf+Gmm0d+DxBkvfMr9zSSNYXk9ov1
IMbZOY8zTSPg9Cds97wERl2SocOKfSuEn7wpPZ3YCT48Q/6/xAYgtyhsaCvQuVpgZTyb6obSbg1x
thLwhfoYtpaPyfLkhEH/LbxaRq/kx9RtFNHjNeuQxMeYDg81ZKtYzyVaHWbz0dg94swz2Xk3MdXi
xj6Kx+n0eyWhhizxBOcYIdPjpL8QlifGmcirzH6cAztAplYiD20zLm/DvaLkSA8H/w2Dfga554nB
XdyDrxi7yiXy01v4K/56NUI9z/nap3qESCRc7Sf5P5RY/KH3EHI23KJTjA9oKaQgoYYF5Uf7fvnU
lNDUp4lsG3hkwxmJeiuFOQIQicEFO/B7iD/COk3Kp9xBWdhatHal7R8ptdYSXXa7cf+sNoCaByTF
LyoKvo/g9wW8YnxK3B8BI0ksvA1PsZMllIUFn6Orzzv7UIUtqppbBbgGuh00DjnOHy0heuEZ6P1U
0Sew5bDtsPFXPGtisi1YSE76fJKyHCn6s5tnI2YlCj4r0v7HUYZV84SneR3dfiXodYP54gYL+X9Q
eJgcxri+WNyrakzqiHN88n5YZ+nFiUF11z/hsCto/7bT9TGK79k4/amGzAVhX9RvHOH/SxE6RsHp
N8G/iy/eEt3pxYbtlXS3dU8mnXCPYdMPK3+8lX4nFrJrSQZ0Uv+PQMlk0aO5HoT9U4Yyh/CrYvzm
cnlgiK3xUZrzwy7m31GsjAehZSmF2x6N5Y9Ao19HCFCxXpWv53aHm7xxoVOaroeLlxc8Jf/9xxOt
qSby9xFVsf7YwTGRpxvgFGeObYJ1xD/w1ulcA1lL4nawsfYyIxQFh8Cm0I9YApcsRCgL0oyMGln3
plkgiq7aGiPO7hP787vDEmfq7kPdIyLbMoCMlmLBlSbxBlu3QOvOLwF4UtSPWwbARczQJwHSj1Wt
osHx0v0/NQJoRoSC8uN63BvQOx0cgnvaZ3OXoYmtuuHf8qn7404rWlEq0sF9juMN/XpAeBCcyjp1
ZlQjG06tzVOoStfgdIDRvqojxnUDqECBr+Hl1SP2Y0ZnZp85WwDhde3kLN6U4EPdoGkysAx4NN81
1nus0/k3CeQgiCyy0slQpnpcSxSq2jbxjXGt1eVTu8QBJZO7yaNHgAEi2L7Oze5eU3I58wN9riX7
MtTR2AJnhU1mYFEQ/xsW6KpDFovkyYEsMtDbQpq6DKoOH6hvPaM4YlrsYgC9aZiI5A9u9Ot0AC6L
hKqZUuAOL1varG1vMp9pXZNa4gDPPLwz1HpnNifpQIS+apH017UqbHpYHddEdIeDavTj2hwDevh7
xUlMQ7IzfGnjNG5Axr0M78bxKtVdQFsKPW6V16l8p5LZcWBAK5A35EonUKdp/6JJvgErWKHa1PzB
yavQaAMgiU/9JQjnGRQmupnqgKcWqVvgS0QoGcVjdmpte1pQSHRFuxrZqiFv2+VS5fbYN8RKSmII
kGX9mfGrs5pfJnzaJ+lk/SXex9gZHID5EVHlI5r5+5Bq5nqpm28LaGuN6t8NnP+Jvf9A1YB+f7+r
sVsOj6liMz2l2wqNHWSvy+Jh7wfgxEoCZf+tvuhaBKZ04R7Wyr9bUzPw+xltAbzLWeRtVHQF0JAv
kZZWsJcaX8pivO45zKkL0bLjoqXqxVxwEvMhHeDYyccyGob+KHMNSjKBJVCB60LAPDABluDdvYY8
DUjgUmUJAnyzVD1RLP/IXN+IHnB0g21JMnyiaLV8gRddpQ6u/Z813q26IOiEOAG3ul6jZw3kFqAR
UZ5F8v8we6ekiLEtjI+ZzoS9PQxNM92ywFhNuLgzms93YKipbNS19RmV0Mz0VMVoCHRu4V3MMN+b
ZA7qiapMkVwTpkQ04OjDNr7y1/9YxYkRe9Gh/3c8q3gdH6xsPND5xcAkejxedy6azq2J7JvLlGIK
wHquLDYIrjAHxDY/nUJrlmIjBvZcKjia4ei8s0clJidy5BpGliZNJOAJgaGo6vYz0NLSfu0ghpB5
SmkEgts1fCZUCQ3brMwHR/hJrDz6LSIvTz+lklODwriG0E8/l8XgpmxjkV/9JOW1vUm+wre4pRom
/u+1cmII8PVcl7GQ7RT3FVvdjZepWN3dM+8GBiwHc53fUC+ZidtwELiQ38LE5b5h98MoZzntUpgL
atSgzo2Xaryhdc0hUlcQHDwZfICTkyV9BZ/jrGFQaZHCEV1feZ/sjNICPlYILTi1k3HvUSVoIFsE
yqc8h/JttV0h/CnWNy1PHzBoEfrJ3263NSy3f6szQnnOLAlejy2yLurum+LlN9E2b6YoushRutNz
mVDFcM72J5Fki9O4TTFz+aPocll0pQniGpquJmook/aM7fkFKN27tB5b2w0YDl70Q/r9DamHl6hs
vI2H9KAP3aNkdngo6aPK0Q/Edf0jv1I6/jflo3/hN7ZKBXv4a+M/Eebc0VuUdhj7sXOr5DTR+Lqd
GthyXWdk7HAiTOqJK0DR1F8FUvR7K2RPlW+ZfGNGYRZthYzVuwVJkGKgtREgEU1TyMKkX/33NOYx
LuLcPxireKyrbdcFqqAy38XcDJL0i9s+ctjlgPFEOXe9bo7l6uhP0qaj++9IE28MzWT7mqOPkMmI
i1Bf+jFhgfno8qaB6kEwkdFz3cGGzS6LphrYcKI4BQIHdVyJLJG+gW2gBVV46e2oFCpfekYd0n1M
qzlbQxnj8QYOapp86arKkQKL8vBC8dGsBjGdXcUoavkwgP7kOvXkaE0cIaT4lHGsilgFRWAAX/7j
zAPLZUHXmunGtvVHxER5kkFJ4KsYZ9p9nJl4RvZgo8TgQrGPKbrTpHFVesIHgiftM0DvwcrsuOhj
BfLByLW3B1vaaE4ecp6LIR35e4C6KTKMtfGa9z/LW05ovtAAzWvCYTkY7gz4bWc4dDiOMEcf2jb4
Khbk+DbMf0qYT0gAc0fytxlyarqs6mN3z6IYj7JCzPLlzcmCsxx4atkhUUaNoFkN/AK1jXPYQzZN
BDP1epv9YiX46xCYd8btmqsgspQicv2hA+iD1LQNpxaDHdySizzCRaq0AQT7GMej9hmykNRV5YzV
UdAWJNSW0lbSmlI+8KU8YDLc6nGZakVCyaUlerxTbR6ny8qh4OwR391a6/1Gv2qvIcp9BRQIvRiq
SafYGMXCmso42xBpUJsV3yCTNNjSbCsV3LNsy44srVnlKNTZe3Pqp8AIvus/+RpEuIvarbm4g353
C7+r0BYvn7F1XT0CmUwVTlIVnQfz9STcjP0HZEV+U/WWe6Fn39RzAoBWWdlfY5gUhc2X8SiFUQvP
LhHN48/AbGO/Y3NXIuuJyOx4iKF2lwmDJ64sALqacbOuCx75TAlJu+JXe8VRIlv8jdGVwwERQxNx
4TxVclO9GYIiYPbe4oOChMDO9mw3UBcgn96JFg8xf0rN3lCmu3MCRZwn8Yl3p80orbupOwNW5Y48
y1wNGQNUtJm7SZyr7CvU0HTaDbHDqCfireVziitdE5A3lhIhAHX7m7qwuGE10YZGxdDKMsKGtOUm
++mijSQp/mnRaUZfk4p5LiQrvKy0e9qrOhT42rlgaDFcaPDWnY1uQP0ucWLH84Y/giFl/0JfpXSe
4CNkuAtEuEtUHzJIw5qxCkbJSlm6k0/C6ZNEQ8yxDdBBSNiGYbi/gbnvEFXFhzgMeJ2tP/z7DPrA
l95tgjcZXd8nPbWJTcunsfDN0c4pG/u63ss2985GkSh5u16dA8Vlbe3tuIqYJC/2lQ1qZr+Zevf9
mKieFPDn5JkTBdB62on10ybAs2wcMiMqlzOvoER01DmrakLCmIPxUids3eShfimM00Q4XcLIqdrD
BRErXPB4twWFGmyzPKmckqGX3IhIG3T3+U8OIU8cDaQQV3vLyPSyhvzcZWUr9WUuwhVwIpbHMSE2
F+K7wr60Gftb7JEfui/IPPXBIihpSjZYKGzD/WldK84U5oyh5eW9Rmr7VkpnIzxCBxmo2xm2qX84
k0nxJFXWNarnFML8Pjng5Fcysbn07tnz6pLZtEc9hv8eDZIXkHBsiWngLogr5uKo7vjcJLC9iLZA
1S0p7bSevTveEnVesLGwDLB7IhYHVMiA0NJNaPl5J44SlEi/G4f21Sjhc/+kyaslJ/lQYXo4Sf4M
W4ymLbYTNTY6YMRu1nWSro5KLh+8vr2Kso9iyzs+41W7/QA51NZSMTwhT2LwDDeOsXQ72X0lkuf2
YhvpHJBIpiLgzNyl0Rwr9vc7TaRreGZt+kYGIBaxExAaKX0k+o2gN2phxnHdhU36aCE4TuvHK/8L
Zngkm3SiUQPs4iMJFa8OPDc+oya6qHGO5P23f1HUSPJ80JeBzJQbiEjxH20sxELT3S/2yixm+vL8
laqANy7dBwC8A4T1xWwTCvF/etjRWtzstx+A9VZpK5gWbMGFLoy4inj5PrbZoaJulVrpeuhrmXvY
fMv584oJI6o2ETHV7jGstb3OGq7olDX6IQrO5Mmd+PqllXzCp4Pyyq8AIv1ZcYwSu9LJF7Vw5UI/
9K4FgGKAHF2z73wKwK7CdeTpv/fREINVocgb8hzkfXn8tcyzwYZmFv60WfJklEM6FAAZSHmWlPXj
deqmO08aTXdEazKzIIzoPrSHYEwLDB5f3tIpVeI0dzb1vPYIYBuAFks9DXthH49N4gKilm4PmQtq
RPEUEMfcu6d5MMDFbNgullyY7A99BcpnFtkkgYPx1nSin4QBXmG/npa9hpMixs/Tg4Jnoqgmci0r
U/mTwRPSOnonrzd1DqYA94hPUIG6La5ePK55l6HwMR76N3j91AjuYnOaTaAqxDuy1m+LvdNvCVdc
IyWoFi+/gaS75IDPgTI0KIsvK5G8Xk/FufjySUS0qrEAMREEVjIbanfOoo42elET6FcokPCeFdS4
Cp0mvOoUs7qSRiJjpPn3YhsBlSy0Zhm4FneSWpiIr9jmhMq7HeLURdmgr9V8phcAtocN/SvSN1qd
lMT27Xi+/Xj5Hx7eCB0QFX5As7TafscyMhbncR+PcdS/KVHLTdgNXXYVRTg+mIOeu5gG3TvGNyWv
G/ojIbG7inR2uBBfJcBGZGmWlsZhErXzWlrjXLEbVmUD2Mef+oy+vPjGBwj8R0KcUOtO8fT8VTw3
lLg1fW9uhWo8x5mB5/p7upe7n1hiDX/f8eHCkeMHCIHgACLdinB9/YCnbfGeepbSwR6QbN88KRfq
K8XWMoCOy1/5Mls0NM7Ruiu43ejTPiaIqVuUKN27qhwLpXJWsuEyaojdSmiDzbpCv8XPYxlpMa5L
me8FRC2NRZeobSye8AuFW+3nWhAlXGnmfcC9kZatmXE14XQ+ev3PXO/omD1LV6ZVpzTpmAdrEUxW
35+A/vF5+n+FsoxHFdeNhmPwtxxabPZgZLIj4DBRzabUSk0s8iMQJahOu7DT67+PIlamzRLz6ah2
v+U5pPAYv/8g9mIsQPCbwrtQHG7dUWLX+rn9zS8HKlKMKWOnLqp8aHcvx87WyobTQLlipF91LrK+
AR3AuWMKzghiMqXtEFlCEUoX+U+SbKvjvpEg/rb/5etAACgaF5rAXVmBwHUqJPNNgfa8ucOU1nGq
b6uZATU8WrMSG8Qc5wQX5khkgRTD0E9W/OXiXj1NT7DXC3ekOH3k6vSMk5uNnO/LhBy+2gtVN8KO
iYnVZnyp/1LwgcSa38uEr5lRAuJwEfQsaiamv2Mk35VsTV0+g6HELJSFBwDXfjxLWW7HSnE9szQK
lx5YTv0bOd+757ag77y7byJcMqBpr31/QUx0F/UWLy1R5kTXSIcMmdJ0oQYn0Nd7IYc8QqeD77zZ
AZRkdJM92JBxuxNTfWVS3XavOtcNWSn1UgcIiJefpzxU5BpMX0QFiL2jD2W/Rq4bFTxMo/1PzpYG
VAYBkvXVr0rNgr6zHKtuQl65n02Fq7biK9GPZMlvMI+SvJFJdcuHYgpl0J2d+SDKrB1yEtl4PKC5
1B9r9gBSPd/WFTsbG7AUKjYj11Ol6OgyyW619Kfdf7iuq9teNeAkpvTDR/wfbh3IBOpmlXzAVugc
cG+dya+Wkik+NazHZLp5+fHUo6Q8St2xm7PiBLKMxYBQeE+xUZJwvBaolWLvBSIYZnI09rA+baK1
3hXFatvo8EmMuMlWErJLLCd7Ui+TMcaCclrwjTg967L1oAkGWtGS3xDV/HzzO4QkRZScZ7+ME8Lf
WOmoSF2Ka3dQMjnz/h7pA6Fdq4WCn4kSHiRxoGntSd1E/2sV5osWiLrjixm7BkQcZYB4gFUGcBZr
lg8dXBLQn00jhxxJnXcNaI8uSrY2/bU4TbLA7trr4TLDiRV9wK6IqGFJ6UwItnhXFFZkMnh3/0rl
+rGTra9cQujuJtJflHcojBzodNf5nbiV8oyJLDHz5eadyAfwIFpCWrKlA/5GtqNCCqT12Su9lSoT
oKwF0HnpHwlJ3StXpHubXcNnRSTpcv8KE3wN05h4eXOVidqGpZuH2lBXd/yQB5vtwAUdx808tv9m
RUBEpfuJcZoZetltXyvMnQASiJ+i5HbXrzTT1yjFlrwTmv9C8Otf0kr9ffi/VEfCyWR7uaUaIi1U
rd4u0WEA6kLe4vKsNtKahimHIsnxa2ir9DyhIOjbRlnv89mnwQXGLf5klAeY5fu9BpLlzzqlMfYi
2qXiZNJK0wnSx37Y2qqm9AK+ee8DdTcKgiaAkma9aaT5x5DofWQzcLCuiSHVnNKLYS2Vnjf4mC1Z
CSM5qYhe2gR8HlRr15jCs1buz12YqFciycL1OCYVk+AupsZbIcov8lR5U9T6htYP4rCt7W4FrU10
xrhIeD/qHu147mOI/kA0MEJFiw91MALXfxTgoaHctvqr8xUe8UVeUwLS2J1shTisDznPQGeDpA6d
JjF3VFGBnIU9mERH2ZthrTbUT4wLA/njVrvALKdbsrFBgwDMCHnIOrXyU9HAB4QsmbgKAmVZ9AdR
m8R7/6OG+doYnnrWAd03gsTtOIJvKJgX5SCeY1K+bcooz18M4Qp6m5c+lve1KGDJVoX5EAqV9hiz
QOObzMJWYK2FVkh56+tLZ5mvTwaGvoTONAoJF8i5hH2ZHPw7x4ktD3pivsSCUcReanGbJFt8Cpun
7lakOvyCWD5Xfx9h0nsFUfDFSUvXJUIt2PIryzvGFbEQaoHuhpR+ld3kZsLMe752U/i7ArO/SHjR
Dft1eu+JJ3Gj8DSai88HoIWN6zllHD0zkLhDik68Y3in5gSVF5IMGGlMBAX74g7dECJa9ZZkKWsS
x9RQ/5bDbhHlzMR2SQXmDQBFtr4A505vJPjiZeZeYFMpaFJEVUBulcwi6y82pTFgDfyXsKjFNnhw
S+R01BSuHSEfnElskskUMZpsKz6Hvk8/sRxKkE2bxUE6aLEJisKWEFBkNwrk5rlRTluFMderZV50
FU2ptDBv8jNP9cQrIjkkWiuDKobso2vJXcBmtsvhVdY6pEWwDXHNydmUz9VePzx9+JrnZQuxswuE
bQDwdUqqQis55gPcSjCWNfp9ZCCgCsKfOX5Lv67MFvnEa1d7BLMPaI43oLyWRx7FGfvNKiaQ14FO
0QrQyoGko858ZO2nUUe7EV9HKDPYGRd+LKBvbaer0kzd9sYjFtknf9atY3xTM0sNCs2ZGEdhqhZv
TsRU+DTRFXIXkTPXh/KkfAt5kcaaPlPSpMtT20uAebomm+3AJxwbkQfjnUcdfDNvQ7b+82W/YQg9
e1f4uZ4kp7OEjWduSUnUxfqL+fUHG9LJtZt7Xc8YE7H8uLtdBVnYCEcAxlWviWCZ8cvSjTA3WWWM
qPDM0RJUyYkzzqrNpXAue1m6WT2eZctc3Ixn/COqo2jnTCOZFw+AsBHHpMttc3T0m07qYw7PhHNL
UoHx/VRih10FcxWR12j5FriRdfm1drbNU1//T0xWXfrFxGj3ZePYbrHRxntLJ6T1yKOnP/jaJmBP
gaBBWRF8EZqTTOwEOe+0WvQessJ5BaKkkzfR5mltJWxVJp7qYjvzWwPEqX+bw3nlFmZowAmcRvK5
CuvbVjJJkpQlwL697NYjd3pDetYkyaRv01/vtd66lnwjPLrbOo8eLH+ENyxBsIsbACM0c8ungj9d
GUS9f4qHITQi2xQYncver/4TsXCgOrUhAJ1QEwQ/IWQJUQAvbhLVbUFYFx0Z5z7ifWfWpDldYitF
+09QpI/EKzKi8mHkhQFCn6AC+OiZISyLpBKwf+6B2bzdtuBQq1HKnu/KJEH5bFMzuy5HN4/W1Vz1
Dk5wD0koKzpAteu+CYdoC8uNzFtQQZyLJOgk5F0fWyQBl59qy/vMR1/jy4+SybzCPKN5gHaZFUKA
j1wgBgoRXJzNTHAyKw5+1xP3m2QoF77jd9Vrv1OYPuGUWX68ndNf8AvgYW2cGybYYZFUqRkeF4Pp
Nki5O4gQ108R5AWZ/HhYmC7EgMInFUIA4uKjbkGYTFNK90LNjipuyjGTRUpkCymF0STQXqK+hTX/
mZZwXEPh/bBOyz/BFULYIsaKhtHHWShCAuGpQoAI4AFdjYg5laN8Mq2BbUnYDstz+7A+5KT9b/nf
bnidKuF7Ljp6MQTzAJx2tahznQKhpztxi3pjcZ/QeUM+MApr0Z3L8qJa7/PrZWgWRyG50ogLmBOh
r77RWVVDbX1cjRg+FHGHSdyz0EUiGvkzpE5m1OGNfH0bbevDfjNbB/3DlXruyuAkupHZe/GJA/qf
pmDBHRHy4fnDQpBtCCUz9A32qQTXUjGmh7IyCj2RXB0bKNNJiCLq6r8MiAEhtpTvxT5C0zDRRmd1
nnOhl+k+iIyGb5pWiHA83jgjaxbYTbIlAn+8zTx4rrjETHlZSI5i1M8xlMzxYImAbnv+id6mexId
oAPNb+TbRpV5URJ1MXcRdxUOEIp/DvpbEaVvoK8ol53g2eqldn7CYnNO0/HpDGHrQ86iVvmf8j3e
KkF3TGW7JfoF2lHo4vT5v9vvLyMJ9GC5dsw4hz9c1imuEOV7A6wS9U/JmLzX2EPe2JZKYwsvS6AD
1o1VivyKGIJCcy4xAy/OzANkDw9Zjfs6c3DwoFnf8HE5+tXfNXjEIsg/UD5VjvjI5DLNWC5vlcpC
sOfvVJJ3DTH7oW4dZnwz+VgFmGxYF8NmbfRIljb8pAMULRlNi1r/SmzBaU313vcJW1ZFLwPQFSYX
ks5zlwAEcKxWWzOsq7u8diFnlHeUafy7936Bmd2SMS+3YWZF/bRS5r7r2idn63Qo9ErXe86R2NEO
gVQFaW4THDUBY35GkEiuFqTzSBHOB1w3hAkTl0jKUlCVWEuwfkyJchrLn/bJ+W3sMMn0IqSOF3ph
YPJiQDZhCvrHpAvxd5fDqRNWYufhcI0xOv5MFkWf9RQCuujYIhW6HcNzTU9jnGXDDpZbu6JcYyQ4
6HZNkdLTnN0eUblm+z3Lo30YJD8o40zpPF9i8FvZ1HFJbjh4iisTlArsMfmA0aqQhkJyjos76ddm
FdzzSrBCcPwBtw6sCCfZv8z+CUpaFq5ZZtL3trAzd1Q/jLGjojKwsUX0NJz15XC7j5GKReug0+RW
Mk5pD+4SPcAEZ6Pky9HPGBSBpl6ew7EOlB/UR1tZbYoBbGg5uxDpHLQXRwd5KnYMacY5tta+68dy
g2pQ5kmYaAs537E8Giqap38s4eBdnlhhcO2sI/TIVadNwWvoz1YAqO/ZQHXtjz3ET4BV8eihqChV
ZIHcNK9wQvwNLy93qC7eRW2gyVQozFokRTPStbdOxRCsTMRjrY8suKCb9mWK7XUjufw37yopuYPr
MZ+HsZjRCPloLBw4UGjCDh2tha9i3bcAN5c0ubXLXRK3wGTrSKFt7ZqpC1EqPj/y5X3qpzCXRLb6
cM3Zjp3qCamzoafdxvoe5W6HYXtQxG6MclNIRr1M2HmUzuTq9WVqfdZfPv05yrxZwtT5gZWNqAmu
VQOKEBn+wd3ZxAoO8SJqsmTD+cyKJOvgBzsI4OSWujznbYkZuqz9+HdjOqRlsQVrv0qNC1m/bonS
iLCRziFtXyIHKD/dOGfNS+o6rq0bsht4c5a3CVl8u8kTzJs6asIDfNRxecPI8Pxq9qVs5ELXqkFL
39s8OsU2gzsUAW33XB6CYzlkeJhG9UIna4CLjXlxCQ8qyFbeiP+xfwrB7NeoXV4ZjPHfy1Q8JGfE
9cDJ3PXzYCXJ1WHqCCdiDxlEtKM3CX2hlreFsphdfvFSG6dIhDb4YMpHnT11t83ez5cEYaL6hC4s
io/D1pJpWtF6XjZibQAHe5qjjWET4DxaKfAkA4B6OXxuZc/BxHGme0a/u5knMzArv3jmM0wvoECe
XrNuigf4jlHh0r6shp+k3R5PI4wqWdhWwJ5XytO/tm1kMKiOJh1hIEepxJ7Uq8/TT3wQMEzSAKLb
BZbd6sR+tBk9QIKcLLkGZNDt95JvA4kl2ev3CbjzkVvJ8irr9IPb3YljIj0nf0eUOJPc6zgfMv4g
FeBv+2zA4SbpeBDPMP0bCJA99NEZURAtZyzZq1XnMmafNZggMmEYi5UT9veoel2U6a/+3SRYmnTq
pP0pKGWa8Ey6rS/DQ6KDjd5omaFrSWVI07/25gBjUtdZmPY8P2fIQPbqwIKOibj3l+ZfZxtCgTsN
TjXnPg9MJbXmdaHYtWoJ56zn2FN8Gp+XsHMiV1W+BWYpfkbvL1LQCJ0OP/0WF2BYVfnsGz8TFlWy
7uTSZt+u8u14M3KSTir+7g6U3OBhqAUcORRm8/ly/wkA9wIdr66YX3SXpmGw9j/9puC+6Q/UzAQx
xEXCIqd5ZJ4tQwC2xJpsFH3D8BmsulyUvoMVsl4zA15et38Ngs2vY507E8qJ5BDQ0QE11NJcU1Ra
+d4mb53ANenFSqRD0RR9JXHwLC/A1brpHfUTg6Y16Y/KLVDuQmzoNBGn3IDsaIraiNCRoUb15uWE
JPkwm5fCy6lKQZlzDBSzOUAXqX069pC6aPml3+RU5GFef9yMUfqd9BQSLzr+ui2RQ03kpAgiz2lN
Ks+DOOBuZ8SEsQzy1we35WYcFCffIko0lXQTliZNxVKO+O41+xlcADzhlNk6qgoMUlqJ7yc9vwyl
W6uft8t3tzCq9b6hk+wa6hImRMsRrdGZpyRyyO6eq3LKBhThpa2OEMt5+EfvKS5yEOmPpVkjEpb1
JZKKecUVaPEuS8OGL/6cIWlVpG6MWDrJQGQZ0hkN2KpdY79d/tm3uXRjNXSYZqS4i4HP66Fe6MX0
y7aZp3uMjF6zIZu1weqbmz+APmKJomkBgDUNOG+NV8qjWd1bXp2V0iAY6SlP4KeXYtJBrelQnzPI
iJbzIz71o1p5M8H1Nx8BmmYruavs3947pkecUQ2kNkkkysU/FmAoX0+4zysRXLMmlq8kt/sDxEUv
YwNzlOGo2ZCw7wN+YpW0UkfIgkez65iHK8PalnN64KzRIE9NBxI2bFjYVAaFL0WcWWtIgP9NUygg
Ug5uPu07xfE6SCZTE6kDCGB4b+XBdHSoqOAT49Ii9lRwB1Z2Ui2WOEwg7UbN+e+aulNxDvH3CFgs
1bFePueJqWplw584BtoXNgqOxJZ7+OkQ8lAE5hVXiAoTu78maH/pS5Q66C2So+IFfS2vTDxoDt0N
cWIY+5JWfIm6ooUMsA2kOi2sYCFZt+qwJEID1kKYcqSrPuMJVCPf+WqGpahjCuDLP7zjhHZ9QCzl
KIdiUGToYsYz0pSuDz8x3kEyXDduOt4/Glv3YJ7io4HiX25AgxIC59/CDrM1t15tq8aotZ+95hRT
1To9SoiK13hMAV4FF9nGCrkhhzGj8sSnT6bnnfeo/vqzSHIyhtJQIkO9HR2OLHunTXnlI6naB2YA
4RkiV/5UrkQHJlOeKa/yeoH5+QwekMhguC7RQmuFIOPQmkS2l4xy0Mq0nNAh8Ovl3ly6RA6duHea
Nn9GGugUIInBMpXUcwysElAH04jLIGXJbEzDSMMpg4jz1E9vyeDu1cJth2GdrXkbyLO79apYXb1a
khNYzp3Xb/6/HHgZYY/R4tEU4YpGZ7ACuKaLhkxfnXI5+uk4FdnymZqKeJoXjyjID484vK4zMIDX
N4rAjAzpuV/UpClNip/nVAEsJotu/s3Ruk8k6yM2C2ywkq9RTeNQDi1DbiYQ9SZqGUtRgLlM9tnF
fPcrDKEQV84tizRLT6ClWZ2CrG5udDAHJkf8IG3fT+wQdkLu7obmsVyfejtzrNoiZLBUz61UUXyF
y5jWdEpPWkYTyKE7cI38xDWxcfsg6s+i2hyFgJt7JXVBTbWjrv9Wc56DaTLD4PaeSZa0YHCWnbjM
gAM3jlQIUWhByvxiT369qjjpF+iReE2ow9/knLt7oJH+dHqFi7LuUYnwGyqgTw1652ZtmT2iEmxI
bEnSX3dbe1yLf5V05IjZ28izmcVUh9fY3dwT62AY5o5s0ZBLRtn5jt9eLfFrmtN/0mz7TYvI0o8b
OcGeFYNyH0L69tNQ9YhfAFDumdMs0zW576DX9MyeXWpfNPS8qXLH1dm7fIHe+47JZ/Pl2IIrjeB7
LnxAD8CFcj76ZC5Ui/UnMoH3vdo+QWbPNiMQtBqlJ6goF8ia7stksQuYy7aXLEBhSxWh8SzbHcdH
yohqC0NRxvFh+O4vqTLs0SLUeZd+naTeS5BS2vy3hSGf7aEkUsvKYY6cPB9H9lzny9ZPTdtun+L0
UUGM4La6L/wACDJ0ief88mxrGbsnr/LtITm+RI/M4L0+FJ0lR5QkHjT7EZOWv3TiYQPTnv/oSAe6
kq+QxRSITvVa9EHQlHuZLMdjSWXbPtn4e9yLlqad4TGlSnQbdQ39jykP1v7duUtjDPAYIO47e2sm
PvsYLJ2EezcMD/CZU2VElOWS8vICrQFTQ1+5jTogOr+V0B/dNpUBctmnh3QdqqPKB/dyAKs5nKLd
WtCau0Yd+/yWBCHPPps/B6c8MwfBxJLOmj5XjyEtm/teVvzBfOOqVZPyEo8E9OZCpOV8JyO+8r/P
7/itqeRtPMaN4VTAUkxkpLAoDbBSQLQqsiimY/62QTGTl95/3K2GsXEvVZUhOl+aQtQwwSEnxD+r
m941bbgQH4W0zYFets6YVU6TAcgZ4+khpyM5c1vCSoTMYuegFf9eH1Pn6bCUhRD5v0rAYOFHa5z9
kE7THGpCMHXw4tPvvouUi7fP/ZUlW4IjCoamrU2F1JkiEcDWrJBicppVi5bbtGY63KO5U3NtqVdh
/qKG6P4L6MsVnfsDO7POLTdeDrPFVDTGbLt+YJKruDsSDgs/0XE04CEpRdIs+kMJIsQl8+XpK3WB
0cRCQQ27P0cQwngLArKYH7lxVRbz81RhLnZKN330rG+3jZIh+4EwDSwDbHXZQIcutAWVtadVWQsV
/qFIWSATcXKkDKQ/1IXwZKrpThVAnGfa9Xx2F5ZqSjVFdllUZQ2iX0gDy3vp16a/joad4kL/E4z5
2qp5dd5yuM6R9jEUWmXATy66PZX1ujEZFiR0ai4GZ+6nkXrpbuqWv+w4pNASpmxWi+RULRKfB7s2
sDg8J3y+FEGjk5lqtBsZTCec08tqSf6Z7ky8BklrEXu74YUAiDdWk+HYD6qx/lMopuAsaiWN2Sl8
MTWTX6vZSa9x07w+ou3zZQMbLbt50hpw5wL3IddY8sgLFqfvcB5L0AjRwhbAdVMTnjBL9HJyxW0m
d0BQKSlFJtldbS1ou+BbTDl9/ybk0qEKuFt9tWRowoM1K8ppvmlZEbugTlWhb/2BOe09Tj2kfHck
8kYPR+bizDeD6xyZCAEHEhjNZP5Jc9IkHAUYDWHlyiM0VZHKNVLTkXovMF4blDuAMb6qFZwv53Z4
PiY8NbGFRZAGVvGGzkL51zSnwjXIGg+puIS8uT+vQzE1R/d0+SUeC3eCxaoJ4FxjhdZLDqzJ0w0d
vBQb2mFneNAVCT4KWj/zNlT6P45lRY+x1qK/ozRD9LQC2LFTUzFR08D6iAAZ0BFMBjXfw80+3r7w
r3yMMi/J8WaVwyUx3NQdENF8hXJ00AmKqyzgK7czZUjtk1mWmyzIIf9ErsKWOJE2+numJbKwxw5U
eemTJuvnk2tAqcr3Xosj+8WLoT1b63hxEEFuxeyy3y6EGQDJHeeOiuIyg05D0Y4GH/ciHJNzKtqE
7a0DP92GQa2OPzErJnsEDvvFQjpgED748EEW86QMeRL7iS1luUwnHeMXeuf0JMSOlUGyWHK5bUqi
XEEGUQeKDVvuAFbcm71grmc66AIGRBLQMy1jIlZrvVhzN2T6HJIh7ukqIM5cPGXgjCKBi1sNo4k9
vuGqH8IuH0R6ZlYUGH7NSTn2IeozAjReX5Ld+iCXhUWiIYr5QWReJ9pPpwhQD86IM2pekLT48JzT
ORCkUvtlhlVlx5Nl0bWl+wqxf7pbWzqVBrbNmbnQyk/L6TakCm2qeRdJorB3Ze0Wrvn7gw2FD7zm
814D6PK6uKHiRzoCUiYG2t6xYSk+M0X9x7I34Ivnqdvxg9lGlcSJQ6lA6HaqIqqrg3laeVsDAtuG
dx0LFETUSdDGBGXJF/vjDV1jBMi6P1qzF0LlA/ABXhB5BMs27dLqLZya+phdbqkqgI1qdtXlk8UG
kcnHmX/hKmEK59zM4XWCAHLm6JTnl5toFuKGFjT0PxlNRgm3n8pTaI7GLK17SiOeojSePo4H6+dg
Zz510Sr5GnGqVHwjLDnsaPcE2VjONdJ0CWN+Ci+sIwfGG6vFbenjxWVzwK/J6B6IKtijooSbdhhG
MjGeIEV90r2X+v+wxU5tK5soCb/os8A2ZHZwrOJVF+Js2oVyvVT+YV17tWaC918DRgW1EqMMYEMd
lsv1N27Xt2byuFNRbo5sR3KIyybOuaMEnrkzhEHYbOGqbGpGDgsGsp7NnfJzfaHc8YWbAIzHyNWf
GE6NhGD/wH2bfFwgpdK5j5y/wn9NJZSFgKqZvJ29HjZu4cGb8o4iUNjBP//RmJUBrdsCpsjiyDt1
jZrpjgS+N0OX+/xPmAo+g/1r+FzHWg+AP1RYyV0P0zjdbRSdLs14P1Pfb/9xDj/bQGu7HowfTqU/
7OwK9gIdNU1pIuvpzV6/lT/YN8bESeYVCoyCv/mBaTxKiZvi8SJqmodKw9rp4+pWsVfc/FDtkup4
y8HEj2/m+otR6kQYrA9ag6f0vauvOXzUHuGGgYAglA+y9Tx6S15oRFguxCEcYI+pQ0Hnz1sVFo2h
LKnsMU/t8G72fyFFtcihu9Cl5AgmQA235BmB7nlsO5mzenJk6ZbFv9tSvILotz2NhOKl+LWXRMBt
5Sbzd6gqkHVZHVqxPj+dxTy4SuBap0j6We/LNhxm0b1qhIYOWAVz55jKopD79eeJfTyUzeJdjYE8
nY1O+/4u7iohaIIwDfoheDwpRY1X5Cw5dRcr28fjZFO0TnZq35lRusGlYkdbSCQywKWKcLSHq2qP
9HF5VShdvOQIhq/KVnWvdSvNvnqoMVO2FFYyB1iejQJ2jqH9pU1onGELCegZNzJdcuCsULYF6PiS
bkivz1E5CEw3wn54hL9/0yPOM62wjUk+bXwD0UIVpv/W6oT+y9TEe1r5ZP7VERPwe7K62Mxb9xqa
nWHOZsoLWcYH5w/gVD7KyF4Z+eGHHJMuN+C1tzIJrqjVKQjhkNGdwfHlujw0WdZCJK0UhtZmc60w
Fpxoqn9oRWwfCCvMS3FuAOF2z/KK8r1PPFWHrxw3RkVvI5ouyT69FTQIBbTD8VJnc2TCtPJKUggB
kB5OBGQp7O5z/W3bAISk4E5gLoYmDWvCr7fYPHxEnf9pv8HfcWB8yLdqEJQhGQbx5lZwrnHb3ri8
pw/PQi9PdW2I8lRMqaaJEqEvnGQbqUoOtVX0Xxm72pay1H5GNWSQJux/ObEFQGgQ4qe2WaoJrIH/
Af4uOE9+VPROhGOWhd0mNlbmrAMlUM+MWOmkH84ksrrAJDk83d/jdA/7ZMlsOzqAttOGLBFW/4fN
nIbYinjeT8UzQ1WdICOjnSU3HgB8m5p1ApXqQjK0mAHkb3oAmshuSVci8U2iBrF0vJmKxEoW+o2F
efm/3pZ9mZzR17HALB/7ahAdXygMsaiTTMecuOR7pyuuSQIpLPohRtuGMAMeoevhZswyoCrYfVTF
B4xP4mkQ/b1Bq3BbXDpnZ54wlHRY8YMGTO4Xzl5QlgHpOq7Tus6q4i5NHWxAhgpSbD5xPQ1z/o4x
H5KpBOdfkHh8yKkXDG+S7sJ1WvobJXsjkMYIb1KbbnlJmHTRPmwc2154gj6oVmZup62WNdpQOyHF
Nuqr0XfXTqWG+/aZekpEM+Y43mXa0mx169OKaoGnXx1l+DTFGc+MeFsIeXqIqB4kjKfMYq2gXHiA
n5w/MayuClwRmOzEPq9418O5bgOcyCmoobHMtqDSIdFxDIMT6j177LeAmWkTRK83pG79rP6rspln
yH7P3Xz3B6jGfSs3YQVLsjEl3fwU3QkNzrqv7H2FGNv6VAWHiQldMijrfFkEGG5YSSlRTekSE7vQ
uy1P0FyUzGTLVIQdyqwRUl6el3Pz+/NyoO9/nSocUXSX5+RMJgklQE04mIKWLe1Pca8bMtlwbX3/
9s+2tTmQe2qhID91cs/nUFGMteFIqbxOR9/Ww7d4N3OuH8Gpt4tg38iQx6L0QINl9yyrMKI+tvqo
F67FwWrDDfYzRZfse1CfHd+LDkvvWyvRo0Pqti8LBRrlGmSd7VQSmZm3xA8J3pLW6Hr+zHuGLTB0
JMsV5g08j5iAiStILWjm/Sf6Vyrvw1SBPibQiMnwPOXdUK0Naz4O4eJvPCD9+cgfOtSaoQ6cSmAm
jETgdaLaFKD5skTwcu2yBkoFOE87EZ3aqp/AL3cEQ1VQDrRQe+rdzciH1gk6oMMcOG/9jsy/zPPo
ZBkHHa8Egi4KD+nKTV20Ecw1sqlbzgx3ioyHtZMYXFsytzHAPHhCpEtA4VI+vZu2XCrtVKUGYMZb
eWtmmD4JFkGt4PEff9nALvkW5Mq/Yl4E44KZ2pygx81TS4YNMh8YFVq4U+TEgFZ6580rS+kgFdAf
HeyY/JcVCHvQ/yWtvbB/plaJogA6+Y2lwGqZP7bI7P9DmDlyfixpgt/+kXhtVufefYINJN8nTkqU
WRDJo4DHgRA2iRgpx9YXfpFZ8rdtrQBnZ8C9sc/sXaPF2iVKGuOilll2i9HdMUJMhGjkbCd9plEJ
4mSjvGGo+uZksHRIJYZWpgC++2Nn/9R7B0XCyRE8pTo1oaN5KexpXnRuSAM2R1e00qjZcBkaSqZE
SFoLhU2c8ghMDP2aqwt2kNaZ9F7JfAQ2UCiaB15J220A1VP+FtA4qBuvdYlLLtnRedJsLRxaTbf3
+iZgByvfXJmDZVX5BLfVE4LOc8dl1334mWhb8EeqP/ba54z7MNWU0BkjxyTbaxs+8Fs/TZI9FusH
1xiKnCtu3p1+4R/ZUzje0dbl11mvSq3LwndAnf6UAZLixCifvBBh7O9NV4p+RFVzb8rYr9+rE8+N
Sv1ZTw+7slgcZ655w6a33xP2hnz0+hPLNSsrrRXUsXZXqfZFpkua2MTLyGeBthzLkNC/Rm12TlZc
ZPQzWukkiRx2lfUNZlLcaDzbblFLJM3kX9qO1zOqCLnBAIZaVFXS1jVH3Ess9BPS1eN1UJ87wwpQ
DM0rEpxD1/LOMT2X4h7Nti/rWO89hApC5bR1PZV1LbZsm/PcgRxiFnTucfKL9GmqIyW7/szwKAQ1
K4AOtteY0QPLKcoR2VnssA+bBPi1PmmFVyf0pt3W695Y4aSaAMSm2SpORULhGgqrTPiXHFC3Ejxk
c/TcYqIpexAXp1EnGleA5aonrRtwKAFyihewmQw0hEnihzMbTt+ulBR1THaP9ik2uf9bV4aEIM5v
3dn6vTATH55K3rd5nGWkS+Xm8tSsxnFNSo6PSGq3GkBD9k0DAhUbmpzq5s7Is88UL8TXhyiIOZ6m
C7YeU4A83xjrFTU9yzafconKp5kghndWeodHl8/vxUqZNbktw3Uc+f7Z+HqQzy3aCIDYHRl/Wp4+
qZ9B7jO5QrRXie0eWd5MpW/amBJ16h44cjDs7TU3Lk11YPDl6o36I9bzNwJwm7cTuOPQGSbC8FOR
fSouSQoULn0qmqbHurNJvO8Z11s991ug+Aj50k/a+BZmjk7YrKQc8g6oUjmD+QZa58Fma5O0odZn
YQMDWDkd0V5fYnc5YYK4BFKwAhOrqfwi/0TdlMTw/Lwz3KonqOw31kgu4Q8qgy4takjd+q8r0uVO
+2RGGICj/zh/sgnPQqgy59MMVix0LeCfcCFmIYXItcYontuEgBXhBnAZLRQP1jJrk6outPaIZDc2
mEAdP/E0BA5DZ4bIJ6yuMItJQAS220lfFU0sMWL2+JDzUrm+5a1E2VJYTSCR/K77UBCAUo+l6p6Z
XMynxzLfKNpNkmPwJybfuwlHPJF3JKl5JCpHasoBwzYnZDCVNh40XQF3UTZ0V9EHjNTOKBA+CtJw
b53SCYdyxmL/8HppsIBpM5XKTOPbQ84+P1UazGuikB7u7NWOan2oglrK86988W5xKiyLUMTAGIqM
oSZXK56v1bVM8pBHfVuVWQXkeGnJnSHoC9sIlbLfIrOuA30JudY56Roxn60oFf7E3UIeb6iOnIxk
eBFgdbfJmAVooGt+Ur4qS5COA6bBP0S28OUULLN5wntv0x+VaDWVRG2oKJ3KaoiDKdthX89Cyp6V
I7dgeE973QCwSojHiHn6pFKiWukKq4fabcYvBS2vGh6pbOrA6H6t3Btvxhc944WR2waU2RrCvfS4
anjLDqjDI4kGYPC0flCvfAkVU3QzymwjuXLnQq/aHReykOOTDdCPJ3sxVd9/og6Pp8RonQe8WSG6
TLbaIbbZWRnVQaN2uGD/wuaqfazwFibFAGt1f0ipvqpp/JuQDMxblf5pbLj4T4ZreDlgoS8s0v+h
wb/obHiwVmqJ1bNUywlN3Km97Y48EMWmVUJCM2yrSEBLt9BGzQtGlGUMkeTshdnd2Oxw/tosE3Ne
Jt/0BPQ9/RnexiMz04zy4SWL/BTQChQwcfYthPc1K6lhYny7CPXxrOdgwWin1IYA11Vhu7nAU3wl
scc7ClpeunUBoU9b9zeYpuhyEZwzO+hERB3CqGTygsPKEPfKl6JuJBv0UXsjc7MKPXwG7T3tV9VX
Fzb2vSPxL2a9iX7TjXrS3Uvq02e4M6RA8JMurYRHXy8iBzDW3sGyg669XxPdOnA699ELf3U6L5DL
W4FKi7Po09ycc+fklUBGd80PzHxqu2s5jF+IJmFAL1t6dK7jPV82QGPdG340vxRH3xN9QVvrkIdw
DgBsbK3vrJ87V/f2pclKto4bdNJWx6W20tC4l4mv1YS3zWH1Vx63PYX9xdOeRpgGJBh618qv92yh
yVSMN5N19dnR2mYKUEjihqXcCISyBfcG5R94zCq9NGuXhqCmE6WR4Ac9MVzNIppDlCxinTmPZcFR
AJo8y5yU9MQIt8jVEvVnpaCs+oCFzKSBBP5hhFZxrpmaVWFAcduBdoX+HLIZ0+hNY48JQSzdSLFB
ZHOM9agpIQD4mWRM0g4OjfkBSYL2OfJGxr7M/b1Fgk/QRXw1k5Z7yQqwEOKnWZw9UBacoUsJNhee
pZK3enQsO4uPii+gq/g8QviXWhq676YvbdV4+xMOxFctWO4E7k0a5Gi6TDp+4tw8Mlm2TI2bT4pn
3kF+HsNYwiPEepzp9gYDrO1PMaBiXTSTutzt1UXJQ2UXCZKV3xJ7lcy31A5NAac18jODHUNAe7HU
adIiIHSeHhPMhMTxfVJXu4mWKR8XJpYhaXvEbHbLFlhPfG7D0OUSBBE7quUN/Ft4u1xtwNORyXiV
ztTD3Hg9tHbqym573TWQTwCbchFeNKbT/koKK/71t20/VCSmdYSJmLS7vZsBuObXUaoOj6J6r53V
ZWh5R5lJRVVxlKxzciX2WzJEDnqxZ2VCjd22iSDgPkx76j3FQuOFqppPAjLJsaepgzFotV/OHoQY
P6CyHLGSiacQXoegNj4sb+ltw9tFp9TbSoX4eKuJBkkbPGWy+90OMb4/358Lt4NhDV4jyp1YlokR
5V4bGc9zqOaf7RrMM6gBiOOui++tDZOHEP4TVjYmKA+bwXRMAaCJsshEbffeAH4V77sv9TaYbyeU
7lH4wOKsm7qSwZitK7TPrUtVzFB4qM1xcWNt5izMN9VxMXPyq4v0Qx/nVw4UOAFsexTw64w0qgqe
YdWhqovO1Zk8B7OFl2vb42NkzJXco5S7NL3DFsv6pA4yA7ZPXDG/o59yF/VPBt7ep1TqwLnshmE+
m68ldt3BvjAy6Hz1G4I+DwXPHMm6+ARmslrBJ07vHzRxvlcBqK19zm8Y1Dr6Ou5aPiSnnjaCF3UZ
zeVlKMoAV83gDD4ngM/JaYEsGHggble/4sJ+0YKlSrmAr9Pzvz9owMHBeH1Isk30aFobyimg9UsE
E5OUBLd4nuLLx4wmAU8ZyWPd+xE+LljpGX7DJSSkmuMm+h9/qayYjMvHEkR0fEoDiz/MxkUrh4/Y
Y9knxz3zgXek+j0IQNxTai34cDAU25xTVbDifCRBLK7Uyv97WGnm/YuXsPiLo0ygXllJEMITm6Om
PqGbDKmx8OvBXjK8k6UieZhsDOnHBhtZdkn9GYZC7iotR0SPW1A+rciNrEf35ArS1YakmJfBeEP/
QLSDrF7VfMqtts7mtUB9jSkIermd+OkbCqeemA4jaLhPNRWWyfR8TK5AWK20Dx4T48KxaYRH0zfV
V7veFA+4sYov/BbFslahddxJ37ArVr3icG4GwoT1G6esuydd5nGeCY6vSObSAnKRaULDDkRKW+Pd
t0peD2AL5tFp9kfEIISevnUz9XWb9aZZvpcjVl07Gkd1m0R6xdWGI0UCTkotlYe4vQ2Luz7c1G8q
FjZhbXyNwx8KjJAeFGWF4gcAVW8uZosvqq5y+JSjZe4KX+/nf2mftqZVkYAPX/jV0nJvYvDq4seD
NJZmfy8kJNazZAhi8xITWK9RyyN2+3CTkURjPs3I9uoYAV2Sp32yccGOca5mC9UGW1hFr1Gw8AW+
qwyxdvbdXBUkTdxsiTbsSfATgTv/MTGoNUA0UogRCt0E72I4H3H8C4co0OoslQfzdUqs3cV7sPVu
sS/TjEKMSZ9oHUkPuDtaVdff42xaWR59A/STWTgDc9nHiYO3vjrb1M2W+Ji1LTg6sCQg+doBqt/X
6WHNfJ3DRYsKQt6NFsA5j3B3+JUTn+3CLNDzmYinCdjIN88b7fL9VB1Xxuv6vth8eSPF0WMwCxFF
FYJxrRd93U0Jg+bpi9YdHtRj9kg089IJD1d3eDHnm3vOm9pF1es5JgSmtekaPJ3ZXCStr6vZli73
UG0Cc1DTM9wLX+sknhD6Cw2sruazYVvYOE1a9NnWACRk6RcvkhYUXWm4f7QCbYrJv1ztNTkLyLLS
EmhOi8enKsFDBxDCCBDPzxYyEZdzwpmRCA/+qDWzip6Qf4FIpJIB1tsd+Tkqszy8q8kz7baredUP
MurHN/NKIWUqVC4KO12fbJ9bN7y8Ol9aucZ0YgH8UyVqxjBTUf+Hd6GhO0PQ537S/BR7Q9rU+GVM
QU/Mmh95dlmiCHNBHLC8EV9kHG5CNmF0Ecg5sjpM4SQXt6q2X//YgmIHGNZXRFsOuqKlS0z7N+eA
l3Ln26X2Dr6GedY3jOyoCl2MFMOO83jcYz+mjxapnruK/fT/35qVob/xT7GwFC58uIs1J/c/FN9X
e6PIHKBHMJ0AWDeQtt3f+PgdiV8utBTVHUrrdDkYxd6UawNKCBS954jC4DRfc1XSeOuag3+H1WJc
1jZQCgN5y0wIhfLgH1QTgdFXcfpJQ2QAFwkYNjKnfS0Bh9rGMfUkEe7NodrFrqEVCQt+HHViIo2s
eEtpZR5jsxGNCq7WvBtQnjJZZEF7HplieXRdstZRTSZlAVwkqi/rOmsfX1LMDtANWcYnukcfqqJq
3GDgjxZCo2VKR9dXwDN2EoAxtuxn1SZ0cfM+j6c/9dELLKrDwo750Dn/HHzeRK9L6zXURQW16fwh
xrxTw5Vl+hn3R+2bzGh67pUU/EYOlM+06/E4h63iToF6oqTzMJzvd4MpoJCJ1Aku3ub43dhL7klA
pM4qRo5fV/gqC1rqLKcqouVIo84pwVvDsL7OblnEnbSbvL2onmrJfcQgKZvVQrglj7jWMHGcy/hZ
AkaDUCIEX9AJVpSrkbNhWapYSggSDWf8eBIT5umu1hOqdexRbWK99LCyMywukry8tslFFQ+6metW
SJoM81c8Dv3jF5VEiUoLWIMRfWFldx8OlgxHhq3H+YbNbGuicgrVX1SQYR3YVPIto7WjHmoQnD3H
qAbdMqyaGUvkdBaBtXkaqbHD51Xrlks+Wyb9bio9d9NxPpxYnK2HL7KAOsJ871gwSLInvA8HiCvD
HmYZxqSn7M2osUvThqRSu3vucjHmO3TwbC3J7fKkV/Cgl/2pE3VqE7tQE8AY8CQNxzMAZN8Zeg4v
sg/9ews0/9LbWZES2WZ+YpvLKvTvCm7+5Okrqr41mTiv0nFbkT3CDdPYnRKtFlBMsEP7b34unTbF
NDOwHFzQUniD07hBKEuhy4SdG/QO0gH+TgsH/SaOOT2cybQhyx0RUZ9KirCyN9Ep4L/1/N9TgrKk
L6zaGJ+250xkcTdYJKn8xQkcoB4QRxti1BreQkMPrLmxe9tZu0vD7z5RhaKi7RkKpMMqZzJfFjxh
xro6MgzssHkGh2x2AFWm6VvB/zFp6PeF1IVZX/WuU5v+gAepOhpeoQWkVv5StVZb/ZomPiZM03A7
TuBpL88ystHUaB03EQ6ko4MtJMGl7wJHgTQ+//bitWpt9LjbxnskO3Y6y3Ik+TkbCM3VpjMp3n0V
YsoCD6z9DqopUl8BjshVu4OeM2wmVONSqSFVe4F8AM5PFj8OF2Pkq43sxqT40E26QCpXwEUZUjyB
P8r5PtFd+10dri29R0/RnWfXfhFEkYVa7pW6QoZ6tIxa8KXWe6+gZ/TbZiQVeAN67JSjbnqvUu0U
BBP0dcSd6Z5v9ZmJ/JhEHX4zxHhL+k4EgP/bZsZ4KUnJcOmJvPF02OhlzMstfHUMpcF3TzPUs9Qb
ZBt6Jo8xgqhrCJ9BuZnmJQ2Cbv+ROtdlf13W1kTfcG4FqCZDIemw4Re09gL3yTmy1fkxqYcQTSKi
j3rc+Rf4jKNwxLO7OLJ3D7BXJ0nQrF0ZI5AQEcHfoIdkvqpMPJWbABdTbkWqmc2T6T7vBAfDBtKi
mj7SvZ2VoXsW6kc0MjIU7q/2uEvCaU3Ao8X0dSm5UC0iZVM01DWJuSyzxUkJIerB+R5fwmQUFP7P
UwxAJK8uZvH9WsRGOy3GRTJ80DSWg9WrOLWofUGQxd0WP8rR4GDFfg9McfQWvZVVZPqisGLewftN
cBI6wMQrQ1HUcjaZkITkpsfHlsB4R30FSMqDeJj9Z7nlXfNG+9uWrwqtk0fJiZrTEiRpO+9e8I4i
bn2sURkxKr7KkiDK6oWzjt0gg/WmAdntN9vshYYmnhrEXLucCMQuZY6cN1zIgkK6L3at4n5bthvW
FhpnvwHuq2t1OFsgfdrOC4bZmQmMKFr9dyl72MT34o7q3GybvkQsJE3ocGIOLryHXIVzXc5M0upL
gIE/OxKAvXaL2tYTByjS0Rcxnous5qWj0igdk7uyWfAaIthsdKY+oY2tNwJVXm5GKtISBrTkNVwl
TOhjr+FlDgLRoN4EemIWnU2Di5AaEd8i6sV/uQdHgK8TQ6bN/nCU8z7HhsIblUdifaue0LO7Kke+
8TRuHWPGlmGOkch4GOW6d+RA4Yhsr1SM02nf2o+eb79Q/M7PJKphjMwo86CYgp2j4TC//gxSqV7L
WhSySGrc4iigBSt4r6hBcLKyXFscVvBk7LbdaIuxpmZqxyHJfO+ma4LkSltN6PgzUr4Vn5UBAQMn
vu9TEXdD9tDtUdwgLdiIFfnfMx/upjGSzhruBr6OPYGZAJnD3/+Qa+pwCzHuNllfczamenkImQtp
fh0BT2bN2PQSEX4eP9Oog14YmwIZbzbDL7CN7av2PrynUe+sRLdfncIjwXX3I2YFoqhPI1Pe/16H
ab2OJeYnvrraUN//ljMv0vFViqesXnEK32iTmstOFBiqTnMcebWTtWqHpMrEAT04qeKvy20BceX+
+V/3e3GhIuSGWI21iubMoleW8qFfjHOqavdPXg2i3pXeutpdfc6UJl933vBZAuNQPGE32x2fckZH
xWl5IQP89HMznJd8121mVj9xooK/yuxk7dcd98JjHntjRVCGClzc2iGF909SL97jJknu5v57VNga
SxWURftl7z0kxhnPEgHkLF77/z/n7LjRV9qhSu8MAEbfarNzEW4NwZ2NqdVDhLQNEAEiSTRGVhXs
MrUuKmZ6ml/Y7m3nQCmjNww3iOLvZRDudInH/fhOB1JIkiyd/oVZkKk+4ASjECOKseAECviEszbI
sBqR7Qj76iV7VspL8aJ6YCs1Ay5VpGI11WAd17hfLXoxj/DFnkxaDVIE/Y1qYcKro1z2rmQfVQPs
8xZrOfJt80EGcM8OAlKpc99B8oFt68nDJm5jJVsBSysvvncort9mkwslpD8EynJT0Fc7YOaYaQeK
0fjC4UQMqejFDPLChwDJrldVkDiLYmhrtBMMnNPhPWiraP52CzEca1y9k6tUx+fvd3kdDiAo1uE+
GAzDAND5DYWvJ9XXqS0cTpq6Tcaulw8QcDMJNJ6RWF2fKFFNykMoH1B2DFGZiCFkkPppjuFPyihv
OOtNBthDXx5QnCApRFEWCI7gMKgTaBf5PMpnS2zYMbGKNWBA5WEeVJADYT16L7jd5E9oYPPe2Zk1
Kw2OVV/xS7qUJLgWkOWBKact9d1qvm5Xo6/E9Jusm3X8dpwOAWWqMeJamv/BCabvtcFn/98LVgtx
7LhF0J+LQKYifXvtj0WJwr8Czx00fhQW6DXNCP41G22vC4cX7ymB1lTpGe9LSmah9CTHw+xuG5pc
Mfwkw1Q8BE1/0CmnGGR0ycD8XgodQrP3RlBMzE+HxKj5rxYvbDFPDLUcW8+h2YtJ/3bBSTH5shRf
63MVQ9gvEwkxkmDBTHTY7cwBC582jxq5Z2r/uxLzCw/5VCHQK1OdGAyqFz1+vLQVc4wA4qJuwME8
ffDcoDexy8XcQNaE8M28Q3Rxo+N6+8lYEj3jZlm8xIpBqifuAgkXMs8YZ/sFslCR2lpMoy/t8NNI
O+b0hjA8kKIlnYaHyXn8O6lP+mIZJ5f+BiQtOxcD0T8nmF6cDouOZbp+DEMRH0PVKf8hxnDba6mK
j2/PCLrOhLQh40KM/b/uxxJDIDtmPxZG2NII1f5w+h6srV6uHvCN7a+IYi05bw7woRC2AFFiDgY/
egGBpdMBhyd4H3ra7uDx/duTRSi7VxOFWyXKlMTY0rPprv9ck6P3yo3RulQl08Ay/4szJ3eHyRnD
2QWfarVtTVJD0BCdhfFHfrF8+wYDonBUGbgVUrHwkYg2VM0fdy18X/H+EgOhGH7ukTdqxTapkPZ0
UvavbxQb6JC+VvpocQzdUGD4KB/IEwBNLUWP4OyVXxoq5VX3I7VdVlbbpVS7AglTXesuMAOOH2z7
M68KS62ZjxQxNDTLgzMdg1+f5epndXlrNeEhl5EKFjhfJK9puPVBZ49XoarcMyB823saMfAET3HA
CQIcLHESMH68VHKO8xJ2HesHFs3HuppLT2ox6P9fGUDl02+d6wYV0euQAZIdZNmmw399i/s+7wWy
eXt0EUqa6Sj3SVnAYSS917V8/IT6ESD4tkSkYafuTmhO4TWWL3czEmbuULUIFVCspyJ3PSgKM4PX
ECnxNAHqtKIhK2rjkCsxzUelBIOjQfPBJvKS4vLW8mRDe8Jq7mnyreYb94j3NadIyWL+Cn3ozJp1
64IRBi6R0dia0xiYg2sWUZKqrtrZRU5SFGCj0dFAL3r9teVuMqka707tWG655vWOWxpyRMT/pHoP
RpBz9o7cwYzcHEHKjDVzi6MCrgaViIThtXuKJleMecz0/3VQT/cFZ8kUh5cFvMW1o1VZXGNowmfI
/UT51NXfSeczAZVI4fyhhbqJqqpSik+ZUbb5A/15U8OdsveodXL8QoTtBBnLAM9gcL3udQqtKQ/r
tzHiilpSFtuxOYrg09Ct9zYvXJL9PIOJyz4plc5fwxEGdt+YYHItsSsvjS7GfaRETka+ZJMr99gH
LCeBv5fRK+/XkN7WxgjyJcBskXfm87EYf+of5eBRxRVMzcSXfK+wfotr5gF/FgJ7tCbPYE0K1B8V
aU9cF4oy59dtHAeOyB6jL1KIQCqOJ1H1lAGyQkWLsnSpVC/zenDzFZGq38uomFqr86Qzfmuv4wqY
8gnsMCNlIpnpWXkATwWJzbybVzoynKhbX744H9Y/rqID4Hd5K9PS9fhSgbgFiiPQar5+NRNEIBNc
jnzTmsm4QpmEe22ViGJQl/5IQArrCIv8JaI1p13OAgAq2E2UiMkHD3cr+IzaDu6tMLVJkJ/WPE9J
C6v6dHlzkyOBnKiumgfFNMiEZlqUtOcSA4vkj5KwYpzLlx68dQb6ENW7jMzSytd3RsXkqijiwxNl
ODzr47cjRQ9gCgRpRDnsTXkyToZpS0I2Bf4eUPZhgA2zSAyWiu9m5Pifydn/ZQQHmLAjgdqccUKW
hBN9YASuHE/FM1SC6ay9i1dx0DDz8+oozHhs+oML6t4wVMKgwyUYsLElTAIN1pONYZ/IZKc6CoGF
8o7QwwZeFWvkfaj3r2SuopVwrJVzzouX8Z6AxNgZiSGSZSMhlBxGO0aq2G29kqdmcDtv1yh1oiza
NEp7FV6/mZSYj9nTN+d5SkQ7zc44U4aJ2eIsa+FfZri2PgPtjJm10bxctpqegq979IM5uJ6EPctM
FAEdHRNFM5y8U4PsZ3yJKeAWOML/jT6agTZQHKyxgBasw0untV1G7XFa5vHKmipzxxAv+S9L679q
owgeposjX8UWSNHzn+0SnX9dw4X0BinjNgh+er7dFNCE0S3TK5yVGI9Xj9v3Tn/gI8tysJP/vo9L
6yYQq7d9GC8VWGQOdavu8EQsEk3V6yDfu2UfYVaz+UQDqiFF8Fi/7mZRCdFbGpYQuCz0iCgb+ie6
140JeV4e+Y8UFvGaC94zKPxL7s8vzYiW/MSD+NovMq6EhseX/5k8fwlW8sm/VgvKDn7dC4X3wEbE
rYdiRPJc+1qKI4PWNsaEC/Uhnl1fyiiBwMiAq4gLcIUAZfAoLwYr5BfK9jcIiwcMcPDGKYKGRUxP
ZhWgoLtikAf29707NroLTDdbh5ehqYBqnqHgDJ3iXyye9aaUU7VF6NdafglhGPCJW6dceONYtjI0
ikHkCdrKmSuMyT3Obyw1qpp3+LOO3SmNsuojnbds/iIpUqVoxE4wBWM5SmIVmpy4DdkQfN3QfEx9
9Id2Hn4c596B2Ec486YZ6cR4OP9OeFHILoil1ZkD3LgPl+1Jd+Tph6PpkVELtO8AMDQEnpXhC2gT
kJNvAjcbxs6wr7UeVYzFk3o47LCxjU/ikVerXp/Qy/uusHFBFqRoe4yAuuQo6Z3aTl8YDk+xocdJ
9NQmCotSlHkN1W1sG6yCAb/UF78SSHmruNW0/tmcrse9Adpy6MiZLF/ZlDXlD4Mn50p0b6TJf8/1
514Dh/rjoA4xWP/OYRdJ/uEdGUoBVgzpkZZNadX6oqriAIQT3DPPRYM5X+7Wc6cICZUaPWM15FM8
hKsRBqdiO2IdhaOOHqfR99nZYL/ojQUUGXR6QtMW2P4wo5JfwdH4zQw901yyPdqKGahpoVXCd1Mx
BQcU08GeOiYpreWNMhWMQjX2SQAS2V4r2DtjCrLRJYAoKk5MH6gPYSLSSwUZGgocnuuuaEXykBEr
R0VdqNJsVnE6AULh+SiVxhCvMAW0ELvSu68Aki7yTM1SOCXFQyjd8Oj0Cm4dYuL0C4vgR0o4rsrj
KYzloOCjlCk2jVOXmXFinmpWwhiZmWKvCGnyO1ZgLMQF5JsHhAJqW51F75GTFnsqA94E0qezmBUc
l8QXr8PlTJZ29gTlBd1w7w85bqeJDxsWZuSUjPvJ3dsyK/5KsuDrXVsmTkQmwbYviOPa6s/qael+
3HzcxOpfTTIDaXqsuOYNGxk4m22wTdiKITdhGMhgkzQ7fvamdCBM6PFU0/O0dxbCDCJ8X0borU1h
vSha8irxq+qQsJhMP2vHoicYSjo2NcGlZmkLjOnz2d1HrYbz9j3vUO5CcCaol1taQCkKqBDDktH6
OdQ1ugNl9Py002q2vi+553F5mUyzpEaXpiMpwaqaAOc4sJt+5fz1hUdSHKG0s7WbP01rpVfw6gC1
2ZXX/JOYWdwuRB4aDbO4p+XO6IqrgtbZfPax7bsydza1Cl6/6d8iACnwOpdi7BNKAJJNiebtXGpy
H06okVGXxLTSC/uzIRnLuI8a5uA6XnlA4PVWbTjGLUep9cE0Q29qBJ04BwGdMusxrNxX0ji1TcgV
4SdDmzYCRAzBHwB1N0uslt2t+IRubdBqJKCHmhl19HoCo/SCuNo/E3Y+Ta5YLkDFzSc3978GqlMa
0lfPuN63zPbV7z4ktcMV7nXDL0gGnjdo3EhzuflRmNRI9fgNpSjf1dmrQzl/iOXWnRpgDrNWTqsz
AkSBaRkpsot5tzLiXRgDUKnp1a+5cgq7AAr3wJg8LKMr3mr53hWI8J/qSnTGtURJqjOqqn8+rdhy
oN2Le9jTdgDVdryNa8mqZTut4o1QFkno/gJuOQQJIGX//98Yw62VNnLcj7m3B0LX+9xm4Bf8uEt9
B0T0HzQiquKyJfAhIqaLObzeZUDBE4JbDiCF1y3UKltPk2wruTZOPC4tywx9paE/eO+QsnkV3gFG
KYedyImH6c2YV1Sc3B/E+NJrMGKnfE2JXnjTfPX2Sr1AApgfHsRGF8s8G3Dpa2+ciJ0INgSjF1Ue
S5v6fnAC+C/5h+MJPV/HQuUbUb48DEuerSRUPKtdmFfPBdYZx5t179CAydFr9cIOV+0mWf7vBtiD
rYd4LVRfPUPzdd6EkX1v8Bl72MsKc3IVSPAm138ECFzaoxGDS9RG0R408PhBStvOTONpKNMCzEhD
qioke80HD1PNajhTW+1dGFlj+Y/vVfLBOHPprGDx23RL1bInyLGwBPGcVd210TQ4BbXty+osG7g9
DVuLRzufa2vLtrq6Et4KU3Vc0MMGnNqY2ziT0jRSxIS3b8oVbyiWselX7IonN2uORVifUdVHslpo
XEdj3Waacc8W9Uk+FF5B68z5BP7rmBCUHIckxEusrPnS0+85u6WuPRFnwZk3n60QpZOG1Gnh9QQS
7h2dAlSIyTp/mK4bSjDRpcU8I9R34t1J4QM2cUt63TKPb+GwK2ZBT+fNDuWEVIkhicId2F7GAsS+
BS7OZ1yHgh9jzO2cfnkUEjmI8CJjbI+B4nJhEtZdI2Umo7xJdVeawZa+4iZVvlGgCRZb9b1cfhOX
vRg2p2W3RbNp/MiBJ7bxQ8m3APk/5CkKSix2jlEbX3f0rs6D5YAzbnvUJFTZ/eLuOYLeGhnLLqJW
/iUpfrZRtsLdTpvI/7yqD/thYmLRFwBNJPsS/mxq45srrnY0Xdxa802Jpiuwtk1ZMqRwOOXceDNY
nImpKoHLD1mmzcqsMUB9Q37cKS7TiLPxW3QF4Rsl/ZSssoTLbDLhm9y/WvFfY6zv1toWe5CZd/00
DfZvYSCgnRPbL7joYxZqaFOEEE71CwqNZtSPmvp1+5ZDqu2sePuQySJ2MYSIwzXKr2VyQfYAyqO5
rb8yoKMVoO56MUP/SPbU4LC23YxpEvBogm0D9E6eXOXMZ9Zhe0XKYEhUHBambzmwx3hu3f1ptI7r
dDwyQyO11Y1B1pm6P26Hl/yt7PnUnlH/bbEvi5ghvbjgZ8I5rMTKgJvQO97bWyC3U3hlSkBcV4Cr
MxfNMRIAt/jcoWmWzgrt6ULx1I2p7z7SMWy1MrJT+0QXFz+OzWte6ei6gJBpwX3F2xf5Q/BLPdMt
6n5dqV5PAZ2fkVrbCCiQz+7gmYTLmT3Vh3rKxJrTZLH4pzl27sEzwnNqT2gHgTOswSCroeiUmfx1
fFZH70Whu4t3D3TTc2QaIDP3qG8/zR2T08fDe38d3EdqL1Vb4Hl/ut5I8qaOUVhRn6pGAS2nl1ck
e7/0TH49f34VcZVb8g4PW/6TAUwAL160S8l4pgqJ7gcAcGvt01L78OTwhE/jg49DxaVfVuUQuu8f
CiS9IqzyHHILh+ByUjG9UwbEcof/pE4O/QhYB7JtWX6VI/M/ffBub+6Ln4zRgJWLjyuIqChqbYXh
nj2W0bv9EOGvmdERim75zMDQxs6Qek7XIiz8C2yZctWjnoaSBTIq3v9EEOp1Q337/XSYfSgNdEAM
Lp7WxWbf2kjO8aL80p03UGG34smzK6l33TMbKcfyr6XosQJA+/uwEV7X9gZ6kHGyiE0n6jY7eLq4
TUo43DY/+PS1R293ogjRCXN6qscMSNriaccqz/vdD3EZ0Gm9+lsDlxK2TyuItTc/RNUn0il8ctWy
FAvRQpwvKSTEuasfWnLtN53OZPxXwer+dQsWEzj1xfrxTVJSwyHQsZxVR3OECT5pl9+kJBog4uwR
ej+HLqFdTB/kah+cEWws9FFeZmRKlNzqucv7j0P3J5Jw+cBcc5xaLu0Do86rHZBBLZqW6Pd12J7e
UQI2w2wefOY4ZrMnTrtR0xZYG1D9VKI0/z+4fB7S0T6eFWlxP0CpzvqR5syCQycu3x52C8WmaCZu
GWxtGKCkI/r8sXpWPc9e/0kiZb2ls7XBJmI9JPhHoUboE2p3fcrddTxbN3KkjQQwtUXTq5DMEjmF
13tLbgvPxIRZeVURu2QfXyCYxfm+uQNATYBz6LBYyrRuyaWtVHccwXSVRjisyJ4+X8vwA9EcS4/d
+FLdu4zUX4FU3ry1EpS9M2WjypOT7rwTTGR+nux0QT5glykmzEwLIXI2UCXvx+pPlNLADYaUPJMD
FoKBpE2BUBWpBJ2bED/oALyTiGAZGcYcloFmNGX03v1Tvj11GZIAIwrfYELSZnUsXYDfO4loztGw
E7vM/cE/P9Y1xAakCA4XpWvI7jU/1gJzNM4K+chpSuFyu00QADay4myGkBkTam845h9fztFih5N1
RVgpnsaH8H8rTpPAOuO44lYgbSFvb7atzgVpWWMca3A+CqRQPC5DHNNUF7i3Yi0eS16k4SzD8cVQ
rxC5x2sR6wiEbO6QkeSUQLRnL1URlqFxVwYYuBOmOXTFuxspgpU2FyP6vw7oAAsVRTbxtPsmwxxH
/z8e1LUigSi36FZiarHYOU+pJ9frrb1ArT2lF2V7GKPTAvzvWa+BKY7zzeaCePv/Z3wmbYn6nQtH
s5UYID+etFxw1EpV65WyZT0WrdyriNBFt2OpABehArFzkei4H1g1VAnZQfEjZxZ5pCybaPez+GMB
KWE0E6kAdAo/zhykL8XN6yLJSDiqcxL3vDIFx9uHekaWyDjip3fmGo+Wz02XEFsUytbmGzMwJH+q
dq2/S1LDFm4qBIa0Mg/PH4lkECIjZVodsU5Cge9UQvxOrEyTibcJjsiAgQniF7F4WIQ9VC/+0cY1
+uVr/wkex08TpRrtvrtDvfb9oADwLjHJPgBat9R7eXYuC6pE+Gl/ZhY3kufkPNdNaYoJEOUWOGd0
/uKW2eIMz2QZoJRJUX98GjeT3UQOfHlfAU7S5XtFU3g31kEOYxYr/WxlvjgAB6h9a+A5dLK9LoD9
O48vRW+kWFHSK62/hyFDFVGM/3AUQnEO18rMaxeZMPwL5JmxlvLZyOJQZ2KMtbLPU2nUw4U2HAfX
rqJxfKSNosZun1JF0pakdyE9cyozXYxKYHR7J9h7GUKQfVuoBV8HGs0LNI0WEeSqJRRT1r3ZSHud
URV01Zqgm6uwsydukU6xHOzyWin/sOZwSpJt3f4w7fioDjEsaeH08KKkznSxpKYwXmCR5ssCoHpf
6gPCuZUQwktR4Mk1FD4OUvrs3umNM7v4vLeIjeNzDkGcTfAmiaoyRDe5annl53NrC4hoYtissZWU
/Ge0IFDTl8Ms7TsVq2uOZhsNwYEy7eZDKI4ew2i0icxMfypp9v3m2N+PGNxUR5cZ+yRpgL5RNjY0
i0wjC/armNuRHV0u399iEzTmxn5ma4IHIkLjIUpcR5yPyIOFe/GacZ5Dr+GMvsQdJWnPnfxyo8GJ
ZAy2cd5YJjZ2FtTHSfjp7grMXVW1V4pxigVAR8Qs8ewQo/IEsn7EMyMib3/aMbmbaB6LKvDSdjXB
VICGH6xCHzPtkJbyULDaBTGXoHZJYKGb66Ml7IpA/CVht4b76is0lbD+S95P7//EOvkSoaGI9f6i
eM98xaBqQBjsmy59GTPLRQhzMdg1dARmVINGiSLggBXcaUN6uu63XeSUMs/nKxRc3I6w9jfibVv2
6bdSN2LHHpGmcMCjptN8r69KBXzBjn9+JgwYdIOXsRNl2Jsytk1IXu7ZUFghmy++P88op7B7JuAF
+d+XZaPXxQ6BTa1t8coG4QLpX4ElClJZxXkDkX+IfCGkLzC8yV35Ay11XRDjlzTz2m8YgRE7SvcZ
/MURjFle/5X/Rri3/cx3qfaumMgESkhKy6/3TbtULrL8PfW6LbIZKxVr7iF1LF3BGexZX2jSBDzc
5VP2nboPjl71QgRqXKqveaGfgSuc9FAvq6ag848u99LFpA9G0OUSkx7L8cEZpBB7zgSIr76pWb9L
j/IBNMobwtGayFcNDmaV1FWEEi2E0/JeSfWnw6mU4jUAm+JxbeVvQx6NwOgu7qPSIyt1dc3nyOt4
rmT+j7aA1P39wr0tBHNJcqOZcuLA9oUC44fyRmeLHWnpWKQET0waK3gmpZjvqecV4GcetkrlLm4K
tCWGq1CS8f8MRXRh5ZCU3Q+udhChj4nSYoW+nZmwx51tbkiXSJ7rpL/nL1K1sqUM8cxArKNvHBLL
nYWHNdDeiB0CnE02NaBkWc7nltP4/QrPudHfdzRcTA395a3nJjY9lwOvon/fTh2xVZJBjZC6hu2x
XsbmpQP7jcztWQXqNJ5zMnIr9mTWY4xqjBX6iF6q5CdLjVrkmcN4cvxeOptqxzpqmrNUy0pUdf/r
jnyJ0yknkgIAzoEN+ivoC/Rx+rOLuQE49HaI57kCpt16tyQRtYsa0poSWOQeENa04cFgVWoWsN8M
zKFLhdN9NTUVlztnFYfw/5B1h2LlqbQ87/Y4xiLyjWGyCM6Z8IYFq+phvvQWsasRSK5t7fzF5DHc
RuXcbZB/hc4G2rVHks7sOUYPtMkVbNd03GtTKdiVennE+BO6dNMKxGAmeVDeQ9uMTMMl3AOwSefX
6WKbg5EdM1bqlyKyOIoRTMtC3pu3pwpvy0RE/WNs6qvc7xd3ad+EQaLg/Ty2tFuxbgiQJzGWm5N4
ST80SYsM9EQ/RA+8yb0MYFnWXAHOV4uFEQrcpvNoUWU2Pc2QGFRqIydv3Qub7UORGFEE7qHaoDn5
UiF4jl9jhIO0soCiHrMbB/3/aBfxMXhx7IZ7oWHkc4N/7D5XS8p6QEbWKQS6niRcwjfvbhjbdVVi
yFE4cpcPQQ8tFFRCFgKC0asCsfsVkQqlO1TbZ8Q1Tk4XZHDpBst91IxhD8MpAH0Y2HwyT8XcHplW
rZizfjZ5drGMFtZ23KOOotDShrgvljXCYEgTvQPOX0IBtOP3Msa2gJAVaHYBcdHiVaMklThKh4Ta
aNwO1mE/eYLsBCdsH91TRqCLuWDBg3vzD1R4Zv9IkZmfUJNizXlm2JeUsrAEDm7V325C2ayhDFx7
DFyQbKkUfcOsnGpGqyxyKFHcJ2q8GmLNa+KO02J74nGIDqwciwB3UJ7HHWh0JbR0AFNMBwq9hAgB
rDJgl64g1hCywR/KNkIeUgoHefiCebaDNp/46tohEr+okS7xKMn1Pc51F/KVX6xwtQioAtpGuhBI
CYtXiKAwqOYfzmTse5tXJO/+g5LZlCohFm0GfOdjkioEsa5HxQ9sKohQuPFo3w3HNGU5xfP7wgRu
ruC41lZoiVtBtiWuaO+KmcDUOYpr/MkEnP2huxSbPl09Vve2UJWW7DZrenS5viKhaOhiKpQDrodk
er6a2VN0B3f3rrHgTU1+ulgPJyupNc8ZL1rqVqvk4o9HkUayOoucKu6FpuRKWyxGy5X+z0GGQoPL
kAImOFzCc0i8iVKYQoo98jrnoxeDK7ImnK2KfN1pdUO18osz4NGe3IvA1KaOXsgYlkp5qkgIw7uX
+9EGDkgHRZ9um/j36/0qR6RgM+/gnla0if9uI9yu+X0+F+w+dh0AH2ywt4/PY/Mw8QUE+m2jJ3by
X9TrGw44OJYIaKBrpflN6ITYeZv01rP7U1YR1Hzem2uljCXkDvaa1MuxKx6gyH49ceC/TvZbC1D6
XewfGesGb9xmssH18Rv4NNXBmX2EWbNP7Ib/Itgp0EF6pAuI3Siqi69kT2jdw9QEUQbHvce+TyKD
VmXBupNhEdRK6Knqr28WcNn0h9sdmVbJF7LpA3D0SC0v/P6eXOHh5N8ODu/boUpE9Msfx+GfABlt
dn5ImsDEc92IJ9FZQxQfvXdUlbtiwzvoXMJXSbFGtSbJut+lVmHeB5xCAgz4ztrmfYrcGOtzI9au
zL1WUbWc71tvIScNCJe0M7LMkgnjWKd9k6EavUEL/rtyXrhKpR6+5xzfHouP+msG6jbkjAKCKfQd
rdBxoEK1Psjx1NN/aKrSQxNz0QvPfo3bbqU9INGW0K4ICzdchlzFdJoBK/CxJizgDxFxGO/v/XdZ
3mmXm0nqwBfyJ13+KgHEFGQ48Bx+4yFt1ptlvrO1/A4XoJJZ0dR5j/th6/vECiCZo6yw6baF4jFe
CQuj/0URD8KkAXzvABott2ze9HigCItYcTUXOOJuI64ghQZd1viqqFXasqgFpa3CFtASQ6u141TB
7TdfRYT9n11jcyaLyBHCoSY3RDdAcf1k/FZGk9mdUTNSiyGrSdjQiM2f2jr4iIGbJVqjqk6fIswI
5zhVHhBAdDyESMI3x3mQucYngLrb5G8WrSBxsiNyBI01zIsbtTFjQV/rqaoR7YIs3MfBdz//f0X0
bW4eNCFxeHiskYcaimjjF6110MwLPwY/NmLLzJtCYZzSeUNhkV0bdJ7LAT+RCwmsYZ9mHQ2K4kiK
LCebNI5BXD7W4Z3RfkZ2VZBOEJnevLBMFz89Ci/vh/4HE3Avnob9XMxm16w3uXf+Fs70DBrR3C2S
30r0tPPBXp0aK74ldSC+L91DfBP2WDmWM+w12lhmNC1mIQsubSk7LaG/ZVYOgqcbHYdyLfs0WVcx
SmweQap1i6ksji8eSVcttbGcXzJjvCd93SgF7ZZ2VrCt9ElUCaNsc47Dmsq6elU2f9RXLfJ0j80k
f758GUtsrwtKFbKXx8PhPYFSbcQK6YvI2gjT5e+ZsPw++I5yR64p1QjfRlYKFaNDHlx3SwjZiBnj
Ni75TgVj7bzGqXY075UGlgjdtf9e9etPOsj2VwOa3KWUtbcNeoJN6/Qi5jHaObqEqiMGOxv7vsa7
7YsBtDAl9Bczp4Zt4dKYvY2TtJpwvp5q5KbImSPtrVh1330tEyVtsbfP8agaeQ5djxJ5aeFFip2b
jJ3m8mY5gRg4khd0Y4RXO/nx5wNDHozrkl96FRpprwMi4w56NezCyAjR1u6WXtN0CvQS5E26wtNE
a/SkXrZXDEzUh7x9079fXV1xFCbaXppQbtAwSF4CI1YmocvXmBohjpHugAFjIiooKoPTezvHUjeq
Mbhzsz8cRbZRrgAmHbEdzG72NOO7B/rsiySNQ1QlV8E56bpi63sAZrRLGbw9zl2e7gpui5eOcGUr
W5tQ9vDOAjB9OoDo7nZkosd1X+mDhQaUmcFzXe5+D8v043c3NwmZMvdnI1Ajtql3H/tJ76xZdYUH
d3ScFVfOg3sjz79AUHx19y/dmPaQMDHs8KRheTq1G8jJnsN/3GSL026P/7EbQ5tJBPhG6S0bVdHA
TWdDHsnPqPUOmnpJCSGCq1cTLezdLY0aQe/oWCZaimVHjgaR2jXDp2Exk544BIunAppQVU5oppwa
9TXk4H/3knkFy6513IzFLVnCBNHELa//jNA3wYOCBGC8mmn0Ykjc73JsjD7vSofVGn91BiYqDAR9
wWKO0sgdXL53TLdawrhjEwlNyfE14S1WHNBjb0RIUOxaDZN0WM1wnfJcioHp5RunWSv/QgmGjNrS
6kd54RLNXVoFJg7i4hkPWeMUA2gm+AJ+9Vx9EUtnAT0ftlypHvQ9Q3kyFLkYx+CdY59/0cfpPbms
mj6N4198v+Cizwx9BVeJmvh04orWPW+XExyu0SsaiCNUvZ/FGOKWkA1JqUNRhCY7d2lMiLOc3kdA
XUH3uitmli3QOSFVLjMc+YLxKqpHArBjOq6m6P1Kmp2L6S4TlUyTfbXtDW/8CRlw8J0Z/rnJqNos
LgKmNh53gGTtBSWPZxuGFwcAKIOaYRcYI6XH99yvFXRod0R4Nv7bJczJBePmEn7MXTK60ogjedqw
ggJ5+tNPxd7L5bB5j+j46wHQPmVl6FuTGBozNkw+oDPqzjh35Mw2oJ7VmxDQdYmSqj653Fjex71w
IbEoU0Ckf2f/xVHIyXA4e/QDn6S+ooW1TC8cDeQmNLks8Wb11NHIapUl5kBwcRlieULzu4DeJm6f
oCPmUbEEMSfOG09nYPJY80iXZHSAFlOtQhwBOj7p2ajz8H+ZCkJltBgPsas81RdpM4AreazGV184
XTKZjwu6y6pUm9/3+IQHzXlG3bzsve7+q0nrso6ZkZS25i+b3Iyk894tDq6Mwn9UDDGRTIgAl9FZ
fiSTdvGdiQoiCI5OvrDDOmCn9CV39HoESuSLi9Xjsns3V1dw0rJfUzsniU7Ffu+NnNiekcdKRGYK
ipYYY4Sa7JU1otWRYa4GvsAohf9fHe/Gy/vr1fpbxdEPv6+hwhue83J9t6JMFcsfDhxA5g8bg91H
frpYhxm6zU5JBfL6T6gl1CrfezBwj8XGrcLKXSoDFkZC3zSHv7y8OWOpBP+kv38GHZ4PXVvAf0Wt
UD5dMQ5gIzo0Zc7KIyTPlxztGummsacWKDraf2vjGPGrqfiydK+4q4hRoLDFjaJ3XcwMhM9O2IUx
t7f2XCn2celKVm/uWlhi+JJlegp7uPeLgb//hjI1zn2l59OxqqarfM+cMGAXwsQ4si/BHwO5NhoL
eLiwiazhlfsfWi+Au5UdYxFClMidj8O/wo7MaQ7sEzJwqDnFz3T9br9hAmk2GjOYJdbB4GSQooVZ
MTIujYJVqpbOqBKObdhulNOrVDWqkUYbtNXa2ssqh9JieEb/l/IEGZxtBmRdf/jLBsXuSj6O9I5L
eoNDKNajRgmAVthMhOC14fCBwGsGVqSoWBg0aMIIDmSktQP2RDXUBQ0+C2Ez9PEwkXO1xoikD54w
ZQ15sUt9oexwJM+/QgcxKLPNnaoVSJARQ/2Q6udZ+GR3iYmLVHi7WPy5aeglnRPgsMSzeO3Xb5xa
5i7tKJcSMFkQVOUGjlervru21kKlocMP8PgApiTy9rFcZeIISSPbpKfTJwDTgA9A8dv4Wnc9fltQ
9Spf3Lb+SEpYhfy+6uMDy1bh2wfMy2JP93FfrJSL1CMlUOC/d6NgGPTmLkS3Xzyj7Gu+G/LJQ04B
06GJ7WklKZ4/bpRtZadrDQX+brnPdu1SO4GJmrbA5KElUH5TAK8ZbkKLLRrR/vZ+7HYzNTr6oatG
RxFjydVPZtvgCn7I9QUkotMRaq5UjemdkA7+I2DtIgL8kiw1KlXYJzhmah/P9QGBsYFkBKpQm8T+
19yAa4oWibef3gE5mfgG0GfyhWYY9cDSVhMkCEAuQ/UjYP8NrlKYuVEU2vyHt38jCMfl2/TQ6kIP
U8kwynccYJlC8oPwjqNgKeIyYeDjk5G1cLglmmm7++0YoIFPz9F9GXz9V9G2x3BfC64LIJf78944
rVhcq0RouhkpPXTkeNV9IjC+3tfroPVLC3jY9upWUMaRk6H3H51/AbpZ7yop0p3zrPndadpFkDGR
sHtcQX30M+R3oy4XaaoQ+4hqrhpaBozQ23HFn37Tdcicgi6vud8Fh0geWVCYqMg5z+eMyxxbwOTd
8vlGFVwKhfhwzOOt3k4UXEa4wOrB2lm3EjCdchu9rwEwc9acl5YBF4MQXRJyHq3EMJVKjW4RPigL
a5nBG2yn9MJC0EivjqVB4+F6V/OZ3Tl2gVV8ei1ovdujPBcqccQHt6tHLtagWX1l3FX544kzcbzJ
/y9H/46Sujsw1wFKnlp2OpBZCzqDeO5WGjR7PYN/GtV9wRAKyKQgR9sHwMQcc/NOmRlV4dTMNIax
VA75eP72MRIUYu5ZXde/eoGxDv1bpsFrpp4QUsXDcBlpVWej9gMHK5ujfldPzfHYsBbj0bANk5Lv
+Gdx5PKGWGxjlK0E/9/adNDwlTLeb7vlLs3XNoh3eMqS91IwrAfpEgdtsP8FXDNvU10zfWXYRABO
YQqgPoBxFauNvZDZlx9zxVzPEQdIiPRrK+Dg8pmCevPOQmVdD+UuVGGT0wG8i11xXdej6xxxGUnH
E0jSZ/yhfRrNy7cyCcn9p9kBFLuq7PqSoIea1jDzxoNyXA5X97Hgpu1vyv4g/RblceFgV5siF6Wk
euDR37YWWcNkRjpxlU2V7eBINJK6LAdvFpjzkkH7eVL12hQet8PA4qIGYJPCSYiNXaKd8/+3caKL
NkM9hVmoc8wQZoeXVBAddQ51gG8PBsyzOWs0ZRCq4ILn1UgHNbu33Ez1Gt8EnuFIwJibgrm1rCEk
lH6fJzsBrr7Cx21er2WxjqArfNghd2xhS/b45FMKrqly7d2AtA/HM+VyOKZ0iNDU1SU8dniVImmC
Jfy6r9lkzifNx5HwWTxUZ0b4R2tM/qegkFXON2ixGaYD/c3Li3oJVaW2Igg/73z5GdPTAdAkGhfo
AhKNGHqLzA9bP+nO2vsY8CKOsid/ZXsk1FwzmU2NWuZbTHbi2Dyqy4Qnuz3jLgNtlSvAlSIV+n7Z
knUcD55CilO0W9kVDg3exRTRuxQspn/BICe4NZITkKGSwvoMXrSolF3ZcyoP7yGBrXfoXATJHvtH
zco481N4VFdwc84Ghru07ih3KVHLEjhT+FbLuDiKn/XtbLuDP1jfssYzP15PndLDBsvCcJz7CRRj
CeqXwfF06TWPmtSJsosXvs8G/yDmpxyQIFOTH3PSViZFPVvvC4gXt9SHBkDQq6DyM3qYwXpiryDD
SXsG4xFuH+ckgWDJ0meBQ77QSuwPUKcHXj1pBDgRSl2CrPnEsV+ov9RFKlE2gp5zFTXmZnpnBwqp
TwRhEN+BQ141/hq6vj1CPksRJHzWQFBPkAJkJN02GtrlGvVYd6XScQG91ckrvUAupAf78vkS7GtY
7ljRaTc363FPMkSF53lNJVCmBJ0kMl80/SXYCVZl9qTGSZUwSBUu9fmQnB7qX9Q5e3dPME2AVibm
gzeW5nP36ODOu/d+wmgi3/gVUm88Yf4Gutum+mIPn842JC3r41xZM4+pk0ZPvvx2AI+0DuII02PB
QU7FKLjrDksPLUNVtPOVxTUXRczLMSgSqvbpy0Wjvxg5soUCei+K9VyAStb8d9bnbWQi7UCtI3Zo
9rn3I3Oxp8qGfguo66ivpwsfLnZ1qRn+falKPvChJnJurhA2qok8t8GEKny7UW8BitVgTkpx0PtA
8bhGU+DmGxyCqlmr/EPVi+0RxpDy6riywvxBsIyPXXAx5cucQPbeBixwOFHCC/J38GslsnwqQFr8
sVVRcG20qnfA8gduCpXDTTWA2hHLQVyV1vp9g9eO1oHbRid3PS/900iFB/2scmugcC/QlXGEl/Iq
ZFOn4SsUHunqj0MWq7m+AZc7UswNHxVXft6rGA1pfDpket7qZEeGNiyxg66MuTNQBeMGBI9IBMMJ
KL393AoYN9T7O4w4cPieJLAtf9hEgT7OkTeeogCFoQhd8yfvijGC+1Qx/4BkZbZRX7DsGewEbDiN
ftUGCZdoVdBzTxRTvS6aqqKsBwQaPglGW49c84eVMzdd9Yv4RvzlGwp1ycCvb29dU8eElICkiVlI
Cww7k2VCuVFRokorfOVP4AjKABR6jVKErdM0ukyo9eMeS2IJcgcmljfo7yE7xzQc6ZyDExrBMICg
PuaBXDJzIb1y0/Tf1BAuaHTSYwFPXbk34YP8Xf4emSuFFAjp6BHaA5CEKXdLea06NC9/+E57BKfH
YPRqQ+RtDmgjYsnvrJwZGKnNlH7q0jksjkxQb6LLdXESAiRdO1lomn7WBaidhWeGvy6ERU6gSMza
pUJm1F+Cqk0JA+DWIFnQSpo5rLm0jkgOip+Nzu6T+DCRskOUjzebC/AlccIWLYjqKfj/q3XCHivu
Q1zoPVb+L7V8Ld7HUMwuUKREy0UkMMk0kqYH4Mi1y+OLMS9AfPnwsXPo+7GLbVHCPXoxYJOariLn
peOt7KN0tbdCS0SAQeuoOwnKCGpFY+CGJhsMruHo77pFzF8jSlJHLbW23sRqYGtO47f95trvN95j
cV84RhzSRHZnJZj5XbrQ1jM/7wRwdBcAwLrdydNODgtC9d1TZ8a8cdRRnQYKkF4FpYpHrdZvSCJF
ThH2/4TVwmxrmyLRKdNQcYHaFMkOvP41AV46/j0ci8iHGg1pnscd9NikRvZ5rUw0PDDS+vCrY9QH
7mLrE4MJWbtBaaCT2FScaSAOd/WFQkh3H7Qu/Pd2cSOeYq1gJgw0+KbOzlkUUNlO9IM7rNLHCfci
TMcmfiMDhtCGz5nJMzG3d5ktyVpEG7nbQDbER5FkHqmub8KHt2s4zpji4z8MDMMmZHnIZl+tsBft
+aNeRQFHGywUwskFYMRUF7yCBZ7hQ6qoBS8asUmBLP0CCY/66kOIq/9dWyZqVZBE0saF3FYIBRZS
4HSSNpqET5D9+ws+w5wSOJt2vYuVa7lan2k2Pv9zqy4rfLL1HxWg6twaq3fliaRsW8aU5ZxmOgwo
Dq9O2v3hHwdGQRWedNcLAql08m+wJsX6gD2C2Ccu3Hn1hLcUgkqSt6N5SPHvqgzolTMuuLWo8Bam
jm7yr0pbe+DuaZQTN7ZeJxL25n0vpMr4wDGLqVfNRQk/x9pbUnXfvgJjg7fic4Vij78FNE5WTonf
TzpkgMdr3RMz/NAshDacomoEGhyTlcNM08NmuGlbWYELfX9pNXPWSRsambBwofbyFqoJgJDdTBdT
T+dKCLeB38kqIMI4KaAELlIAesWDdZzlXgAd0fmsVW/nYCfutMpeuwXw92xQqKiFFRjqzX/akcjd
pwGuiDha+pDdb9Oe3jJZHgKDb0qypMxmtw75uil4DTr5sgtlDpQ/2VhU6K7vpQUo/M23tLWkueWN
YaNu3xpmShfNm7HnldEdhitlkj3ysNF5ehlQayc0fuJ/ALk83iOqglkWaNCht9Q1gCqJdvPsW2pW
8S/z9rD9vSYCMgtILhU9nLX0uQyoegs4eRzch71F0F9KZsEvoie3PTYEAPN13UINrzMNkBqVoFA3
GY/6uNuwrzsX3duo3V+i+lfaosVk1NWfBB6f6ugS8lDetljidAsRS6r+fLb5dQIGylXt9J3Ti5Pm
TpnwryBOPaAQw1NQwCeV4HhnkceHlKHY8+VBwlF4XZfFb/fvnL9w8RrTQ89hvA/SpE37k1NDtP3G
UVYxo3t+jk/Y7hgFNvIJ8rTxELxiUJpqkuWaiyMkqrnvJeYnlBWxKLQePHSXyGtl7MHgcC17vfxU
ZXyo5WYVeK9MvudVK945k1IvdhAXuIwxjQqi26Sa5zCZ+JLuDhNbXvX7CDbliR+PkDbC2KqXyFEj
T/iwjW0QJZtgLYFUuY8eTD9jFRZI+3EoCm1GrHLHlonpMuEBwp/KcympUcDvG8/LUJh83s3d6ZzH
Ed4dB8noz8W6O7RFpwKWC34VHtEpxkj/doGeqFzJLmzAsPIK3xnhU89qk7BITvMo1+fdbvKs7Abu
x49oZ1WED0wsZqjxhFzEtxDmhw9FjAxPD0SMiXNO0aOzoIUN2/S2AameJcDiCh51kIcZzRppwe9R
iSORddDpPA0jmCRuThILNLPZ4yteJwRGoBZPb4EN0QS5zAcXU4huy+yuC/V6xTnMq/hbl5yKYvQN
hIuNIZLdxie84tKzJfUhs5Gu7laDrHnYQdnFf9Fo7KAENXN3kp45NN6zsF/Q95yr2POYTuFaw6xX
x8Wy5bUmM/LbFDq9QzNaHZ1t5ohmAaUjej2NAVJUOt3Fcp3h7kM+CF2RyN+NK8rwAqYVTQWY/3lA
Rwrb3aZVswuGqx4OexyMO+modGDQq/dIFhVpiARrymXQzuuGkyIKNHFB8QoTViKLCdrBrWPYI3rL
pjaYdL+ADKCUluvvODSzwpaqeWnnwmQfuq8flIl0R0oK+wD0sJMeatSrq3Z19A1sFLKXU4isf5JA
Dm6RV204+FngUwVFFu6iLhgc1aQ9mma0qSwUJNUOIbK+Ysm8YJBkV/w8gYIokhwJ0TnJEeDL99JN
eHfeF874YrNqGyALg/a9mOZYgIWzQ+SRYbs1NqgTZySlvkne4OEUI8iLPmtGimEvxYCiIvyO6Jko
D5QGLja3DKZuUyLchNsIPecHUAvqgkYJGTbC0qxW9lnwteDxtvKQg07zWKxFDNFFQLCPVx8zx6fB
LGKj12XGnDLBdLsOsubvSqt0LwyQWWeV4W4VuBrYje/ClzHjbKIN1hp1x6hGw43NvAcchbCZKKe8
duQ9D/BR0oa061s7zMuyg87vF27xdT872MgWTL7zwYAJMrk0hLJ5J/4JlUEBtksRav1zH1OIblot
DRCdhtEgZndpZFP2GnKaBHo08g0R1MVHUhIMPN3QZzfRLAQjhFG7ZHj0f18mhvcBEDiobzeuZcs7
J5xpjY1n/KVuqrKD/GCK5liLMrxFuTLW3Do2kAtFmKcrq2y+IIuEEh+yrmmLYmhRqSmKrVMH6UDf
cs1kW8+cnXK/cMKSuCigwJL3wECVVYiR2GEQjLlkBwYds9uuShnTVgMdOKa+lZKmR4q3IMWGzyLq
nXezzz53HAvb1mtlbaEq7gjTZ7P/Pk3YNCzvM65UX8jgfc6cjS7vflgBJ2+PrN5+1ug/kZndrlir
/pU5lYb2XYWirPo1sjb9cA7o3arTabqv37sCG3WVORG3riRD/DmekM86RoO//GUsd3PSiJxadf4h
z2pGeIO8w22H4Kn4DDXN/071DISk5pxs81hcu5VqO9+99VJnXjYGrMTPzNf5ESkj2E8l5VcIP+LO
Jt/zS2s+2/HsyIGa3Bg7TsvOyk9Y7DGzT0HaowSW6RvnV4cVh20hTMn8B4Mo5RxXdBMPEFFUOIqS
XbbpNxTigEGWAcT/OtdoCVquzemZLneg3Tv4tjT795wwCHADoLmeSob1fCvtwJoQUj7sNna42WIo
sQirpYX3GXM8SiK+bJ13gDNJcLyUiycOLrrmgJARbkf98W40OKwT+PwtDzXIKfCtTFoEoX6DYCIB
TzT2LUVwIXCfbKHxpV/Nk9dgpdrzNlrV/m6OBritl+h5nkEC/dJ2oAG3rxUcZSLQR3Lb0ApJ76Nw
AVl9ExUvUsdxEfxKfzmkAMEJXtmrKwpLIdT3MsRGDynzHJJO62WY+bH9Hjw6+3I4l+6fMGA+BuHu
V/UKgaS6Ojf4fMmTOsZKr6Hipva/FKieCIfjfLFoWmgBI4HqTQ4oyq/a81UO92EWgzlYAZkiMUtO
KIC4jr2s0+HlWAQbNNuBhwe4vw7ANb79Whsf8uQQ6dxB5sN1TMriT8MozCXpP2Ue4jt1Jfd79wVI
2fmnsEABOYbgnWTpE/HgtgDJXHK740dF9qepPRhguhKYzN8vHMteLQS0wgwCpcTcTg9RaPlmPyQJ
yoWnjAVYfkuk3FVVAggkPWjEEVyus+lsvKwjCzCzgbXD5OMjMt/9uZy46a74BYsm5Tmhdl7xtdjj
pRIdhfWNAKqBHgxObLqFGt8wXy7BjM8SsPzHxvIqY+H8l3cBv8LE7EVhyLFmYWY+AfIX0gkKD37D
KG3FvtKMK0CqpEvZc5XOuG5MAGa1tQkP4h08ekF2CXeGr9sChukaRwYMDW7RF41ygdDx9hCz7mYu
C/KT3/tajgSk0BIvLTzVY7h7mSu7tzLdIZj5YPnzc/xaXRQtE3IXxCFgH9ssUuu1AE9kRNXHpiom
lEc/SSt21QTD5D3tAjPNPu3vJF2l004UmrGqUZoOrjiPcxh3eQFuBprkvFpgl0Tw9FN2adWZvgtE
QzmE+DDu/N0stTdpEYoaPmVroDqbVxWEHvrtzx/wn88i837ebqxKSymcZeNJstksAlJGhT/wcZ0s
EXyZfNUL76RNeIdq/5ZoepF5w5Hx7Pj3zN0vqOZd7MsiclAwAOmfK/gzv0vIQbuI6jOdHTOuRx79
WT74M2E68dtdVw+jrPMGT7XWEGKoNSbZs7KysX45r56Q+y1ZWE5tIcoZnj/Ep+cbySLA8XTSyw4/
am6mMSRAnCdn2Q/njHhijnZPtArE+zG5VQ3hdNlJdDtNs1vHEYt80r05cE+JLKIbTUkUkku/uSGN
8FVO8W/yG0WsoNCTdM/toimUn1p81LiN02hD5IURFT63cB/rurt2Nrh8qcWAKzxXbj5Rx5l41YYB
+TbEni6D1tVIpYVhQ3Fum3cNI7GYZ1C5kLwaqRz8Bxoe+BB5QMFNUvErTWKJ5eumUOktnkxRgXHH
zx9LycR4Y+bHzqvgd2no6Xe6SvssNWHZKhUZTHa9k5gm3HrFBct9yppI4Pkecndh3zVkq3a1Xvrb
jeMh6qSrmAM5uxXifx2LgXSPSJQ6tLIkNZl2mduuydCnml3/U+pOt/RPgzjXyPC0EDJDSL45TckH
1WWb7OK885TK9po9a/LRR0ZjSbvCWgjHWiAWOnB17ox2YzGSBsFp1F+j2ZGK0ptaFMWv/JGyyqmU
mC8M8w8F6un9cgdwrex03a8zY3AAUnpdgdKLWIkFUX6wqvwfgKarQtaeFFimQkf75aHu5gmpv+LP
LpNR3xiIUb0oQaBiZa+Uue/sFigUO1nlWjb2SF4Yph+JL+g+pJ0SZJq4s/pJnqYNpaVU3FhNxUYl
PU5l+z1gjQYGbH1g5Ieof50C28stn340K2O183ISasZXZE6+rqVtgCE58pUeRQb19XL7sNarklAf
E6g4RChtBT24NgZvM6OM9CgBDhaJ6jE4N0ChTbmTA4HFWUY6bXxiXqKfIjN9vwPeNFcVmAQrxw3g
YxJVsM4XdTvW8m5bnLpEiCo9zd7KqM5GxWqb05BA5LjcaFuPKjzMEXBRlhQLVn/fv69Tm+JcJV9S
QNrU1KA2JrcEx4eopFcvu5hzeCpRiAvezBGqoyYsNQVBF1Zuq7fONCoA4QiLErXqoRTnmpuX+FQ+
VRqZVnQBF4ZNSsW6ormXs+FQfHVk0J+vcI9A4LWwjDbrF3F2mp6UFaZhtJKHLYFn0KYtWdo1scGO
yapK6rm4roz9LyJcxb78v0pNOS389oAwxwQrXEnmF6hp5bYYtmLGsMWS6eveuOZVFgp3JiuOQwaX
GANNalMBRn2XhDkM28B4DLBOPQu3t6IBZO7ywmcwRf0h0IvKI+C+B7JqlqWy7g/GSbx19GiCAYMI
VqxJhLfuXy6FfEKmLrwNb9tsOvw/6s23KpMwCC4XP7Rgh0D1ebyOFeEXOmbBIo1+ft0I/YDWp3/A
zZGN+mnDbm1JVIbCA8XWvD7J8o17ZVRBANdG85dEyuryJILWaaK1lP7f9dsT4j7XAKoLmfeX23m4
/34yEt88am7jpyYI0V3jNyN92cJQOk7SE5DIjqm8/dUgbubAMxofofSvLvtvy93AcEQylrdFjDgh
qWZSs3+k7KRFxiAtUc/ojDro4sHi3tfooI0VfxD8fcyYCXo//vLzFz8T7y6hS1Fe9JMWxApI1j39
a+vpBXf2KWIN5JNZKRA9ii7XhWpxVNTrrMAUPcfmkPNAmmG6n7ZRGYk65MJbD1oGvy6aXCz3p4wj
IGVWeQHlShM2ggGVcQKbTBw2DQBlwT6g9cg7Ph/5lpzyHGxC8UshcIYBFHFYUQq17XScSfcbX6gC
ldRdMLInl9U2+NT9Z0ArZFCZ0CvkV1FVjlLxuXZPKoWPna4wWy9XTuqpUQaXKQUtFIKbRli+tzYt
c/P8FChL96Jp5HTCezje58PzlaeGHHao6xggovK7c/TPXK/S4CaIKqkwkKwMVGon9wdK7mHp3nRw
3IApA/Cg/qkBkMA46YhxeL2jS/hrS6X3Mu4T0DBCt+FSOdjhOAZnjozQOR+jdqRqQWeIi4rHRCmq
6XaWjQA5MScWSx07Ftgl+tXciScli8AbWnRlkLwG2FfQ0qzJ2pStlaQNcJQ0nMrgDVwA3f4U3bBE
9jXcRpzj6QcZ40l+OJc1Oojzixf/88izlMpFa3HVGVXCGe7s81FiL9QzHZC0ZOuvCjW0zQZjPzHn
dBw5W8U2X3a2zZh8YjUYTTnyOKGjmmBoGVv0g10nOpyd2FZ2ir8WL91jQUo60zcpWdgerOT0BZVQ
IbhILsNN+kHx++6Y5JlA5Yjd8rcO7hmmN0CIveG3iB5tx9g/xxq8L+9Tnuw4WhkYtwv4tvpI6xLG
BeG/bxWStzOYwWANts8LTzFyPwGG70tP1MeAGW/WZu4+ms7+7I6CWdBsn6FPYlEQ6MWZe7G524L/
oi2569qW4FVa/wktRlvFoJK7+Eg9OrDtBpRW46MzQg/8BSDapDXp2zIUzYcMIBayALZFMSWL5T0m
jfgGF0y5ZclmInS3nLgl6ZdfVa4QAWAgl1ZuiHHmayc9d8PtBBbN2yvgoZfQR13h+RmQH1CM93UO
hUsRYs72Y+QL0/KnK6H9+IrHP/2e+iicV4b8NN/+SdqKNeqL+qx7XmNTsg7cDuxxPIRzftze7ZTL
wTgs5XRcK2f6EDx8dRVJGQ5sJIT122QccJt4Yts146BzJkMyHIogTN4iqSzkWUUyXJYTbbKDAX+p
8gZZSvFfwJdn1tfIXhx1oGrs2XE+AI9l6lZeKIF+LLfwkz4nzxqgTuIjM/ZHohT5nFTrKwALI2pW
YwcLH+60bhfvVkVA7aks+lia4uOcrFLP6xgKFra16mn97KLVODVwYIWNz8z0qXaNn9RxgbOKjl0Q
MbmvgdDq9+AV012u6rPWtVJLGKX14bYMKANL0cqnKXInzraonTN0KsuXDOa1DMYXeGyKvYC05HTT
KKtivlU6J4hKrdY322SKDvjCDu0H9pjErYvoP9Hq0M5/dv4aH7kt15sPcyXZM5KT94/5dAkEpYYo
wsadYIrSYUbST0ONZjrbObYg7qrRzGbeUp7ZcPzHQ184zFWXo8YpTmvBoGvDgZKvXZ78eqPLt/Qj
RVFoHdJtbdblj/YnNxMy1VA/bi6T9sAnHxQEdaxzPK1+PcGFvC7CDpUkalfuO59Niis4SEsOpZdo
LQ3OcCYJ7OEgzwheyvCiJ5SdBH0PaHBfucev0VwyfQzfCW9IIRlpN3mX4I4y2teL1rcA27KyG8az
44o2p59XgOiiF5/WqjGSpfboU3nIvG4P0MSmhPqnVTnpveSPS8er/m9shPpNuLBcNuseVBuS+P1L
bBAVSdDcad65IgfBWhZKBR4wLA2BuQ5U3kFu2IMVOnUyc/Awf4Js16bFt2UgrMjJaQ7chzgPXqU/
TCMiyZfRBIYENJooDCVTr5LjJRjKaAN/pMdND+GrZ1lMDp39HXoe7lnLynS0JoWZw7Wn87LNonkc
3VHPVXYQKsJ6wQy61UAnD+qtBvyQx3QXiI9hxdughFy7+ljj7BKeZ4pNAZfzOu5vulqQ/IE4jBr7
rJAEskwrqiuomOzGz2+XCTZVbIcF7g2ln2eMzWYPcym6U5HCnn2e4ZdqXiLjrX60PZn4fossVhmX
LpFyNohSVKm5p6tqHeWXXfNRLqa5FZYBMbauJRD+e5DcdwdquufWadng0iYcqlzcf5wvLiU+bk8B
Oo+4qPLRIErIZuY4gIhO7D36Cqc/hE/Whh7MM85GSecpwt44XyGAqy4bdpdAoBBVvYHEKk/T4Htr
DJnLFpvygu2arNpbl2eUPE8ee581RmsNsdgvB1cMTyBz56cUuiFixmhfGVczr0KtDPzsz+nWYWl0
qqaKC07yvJbIjntouQZEqe+wGRcwYX9uS93HcfilTEcKq6AnhKaZCvM5//3KOUydHA+C9mb4oDTB
auhe4wbZZCfN/ELlTwN3Tto4S8oHBE8LPB17SH8ijt8kqkzEixIq96Ip/lFsfihOzqfSI25xOmk/
pggeKEp461cwfHHbEkwkYV8kCoW1DxMrayIUdWowS/ggO5D9xUAuSQy1OrzL6K85JOwI5TBDSCxm
nJz1jBD9LjWgB8VfKJHpu1o+hbwImiIhSPmT8NVByMckSzWBm68qsmdQVIfcTp9qjKuuueXVTk54
+T0FwA89IHlP877HCnWpYcmQC5e/8TKaN3Wl6hdEtH4/x1oKfeedfI6lo0cFTtv/D1X7VXDCK3Mu
fDjnitwTGiP3ReTrtnSm8DT5v3hsSCbAvBhmCEvKIN4kxwMgrxZEbwj30cHx1x83wYEeQnMMOXm7
0OpnCEijHwu3KYSdVIZa69XSZO9MLLpNZkPQECWIhK/W5sjwk4OkQj9Tx77gPE6CShMf5X7ZvJrc
uKnHVOCrSz8snMrmHiXhz+JwiQoVk2W6fZNpbxm3FnSCHf7qr44a0ku38Wdzu6DWqic67E+0Gj7i
cPl+WfVXH1VoZT4MnQj3JrBak9Dj6Pe6CGGHQaz1T5A+wKbPD6g5xEhUuWwMpZwVsjIMKtsG0M4M
TysMvLytY7r0CJK3uFA3MASAUOLE2Kl7739uAnmg+dEt9O+qXtSmHbVmH4uck+LRbzB7cE5kvYHi
spYvbX58MTx+cDx2j+FUFGIz0tgWXBpNGi1vOHurqnQvrPORVQMr+NKv5k/rJjtx5RqA9LUdhIvf
KNdD8nmeN5DzszNsemvXLcnuSlkce8MIcruWbzao1iiEvq252x2kprTUC17rsG9fImxS2tKfV5/C
V2nzUG8zynL3zGoCM4Z75LbvdAQTuYclOS+5jFT6VnGB0Ipc8xqte7zOlu8vy0FjHu8EwiT1dx2P
AyZWbulCPEqd1VkVKxdYVwZQO5oD6k23yKzlIy3qM4sMVEolj8R++WcOfQ4MRwg7vH4hpzin0huX
L06xHS+VjNQJV7bCKqSZPjuM73jRHp+QbpH0ynYerroMReBEzwvcR5zPxZs1xCRpZHiPwHIV0gtS
xJ+aCgN43gS6ZtvvJdEPVat4rNakeznaBVaVRjBpryOY6KRYPm/Bsm6sYJBOniumem6UBaGZoGe4
UIP4tFnCFEEv9ZopBxQZxemyI6lVs66Hz/8YNWHk8obFKeS98UkXuJFZlMRMj42e0sfNMwzE4duM
qyZuTvFDeXV7IcNH59eYMi5ay5xCNF0kSRHf3p/gZDik3XZadsdgTc/qiwwy3YTF1gH3gOVQ9tUt
0rDjM1AMOg9/+VMVJBEvjIYrsMQg6/R5EM1PRVbx5duF2XaG5bZ+fJGHYyTp02apiaijjAFDjxOy
ENUEnmWMKrNMLbLsCu8AxG1B53l0aDSXrmJbtHOat/LE+Fgg9751UHdW+2eXCtrSKkeRSFAxEVDr
K92MZ/bHQ7HcKky6PI/IE6H4oGaoumqcIcg8Ufs2SueT8rh0K4lqrReJY0SK1d1M3qkUUpJd3Anl
lkkW0F1gQAhaCHHBs8TPH4IGRoePnc3yGDV+6hhRTfQ8dI+rX9TRDu8m6RUrKgXqCxNBeB8V59Cg
WK/07CyjVjGjMSDuaHe4FG+OzMldPAmRhdr1OcPUuBB7xjc19c8A3dywndwXV0lCl1XDo66c7Avy
xCp3AHIt2oHzrW8J7EUa1Tak8oCckOCCrYu5yotp1/sg+bEip6Ytsqk+aNv51Tr2Bugjt9Ca50Zq
F/6uOpmOaZLTRyq0dt+9vBwUT2L1JkHiUltMn9laZP4HyYtk56XJE4YwhCyWIgWMxNcFrbZkYnTj
x3z0vXwU8aMu5jcF5roG3vLjFPUKk9f0ECgon2xFugi1vDav9Ku4obmsOKac7kGLLomwUNlH50yT
2TLhYgWx8NkhDPIV8KgC4i9jeV2Tmlvbm3xYOGw1pjEFUDuzm09i9UrW5B0ZsnYBevMSd/tqrBfY
KODcEt/GCADgXzsjOz7puYKIXvHOviYqfWSoHY3QuUD1VGsZVT+e6wqG6+CP42bMICB45zQ6SrGe
29X2n+WXuUTu3rqhJgZ6Rc9ysgNpDbNAlf1MQMwzPyh7qfdyigrUANzzQLUhxwv/zTsuFIypjBCt
ljP0fS62SApO/QTRqA9OGEbKX7jn+DRLAvuGXQ8UaqcEsnWqd0sMpNEF50mFjFomNKBuaEGLNbda
HKk/ebAUUWsu7NoE9ztb5Fw+OvMxpPXJspPB1WkZ24aiPHTEjM1A3uuSKO4ymyhU9d5s6TJnmP0B
rCCV4tEpc3NM+ISP/Jc21FvvvcLsw8J5SzF2afwVmDCwq2aAA09ZQVBvB2YuQOd+/P50o9QuyO7/
/s8ajZ1xYyIvT3qqp+UQaUCLb5f0R/eIpVYwX5xBUQcqIxSoRQZLmlahV0v+cgL8AHkysaouGdrn
Fj0kTE9wB6vo56uJ/+F3PxTvCskrqQk3AwvZtBJJOor1gBiWH0RoB3/tWqmgNVzAY7u5+V/Cd0pg
oPN/qp83SKCTeHcWFjo6grMh94Oi3xwKPEp65lNi3AaUbz6LoN2NpypYEq4DVc552usX9q4B+oUj
aCi4RwFGa31kEdvwusjlOevTkRoZoT8wb3AAnMzEkQNsUzvjI4HMEh0V4PGdPZ1FNDV+ovY8nbon
iE8UFFkzySCkgpdZ/vmPezhBCebM/Snjb21XmGQ7j/a2pMf1+UpiRCPInLMbEX19TVSqLVG+Eick
ARyKkGIdJFmN+G2VyE1fWpx5QvuowP4BdFhQfBQ7pXDfhnwDSQJUHULZWDXR0Hy9m297VxJzbmgR
BuIGS2m+3T2wHOu36mhptGFZZalzw2Z3eacd8ct6HEhBnPA+8cMZYWKGeV0CuB4+5ozbtdGtYjYm
QXlwPGS43qNb7iJ/AeqPWMIQqB9qsBKXjufRMN2Dj/G4zWnKDFkKWKvfjaHwUZ4SdLtBzKkwvCF1
oHL6tngFb3NkvgCjVo85Op6+LRS33SKut8m8EppKyWByiqvHJtOjMrnxy/i9jdc4Z/vooMRa+nhL
L5UW4u1rx+SVRgEoU0QZDtGx2DvaqXOKfqS6BAmfJbOA8mgHJrBI2AHiehavKBJ78mbie5lF5mAN
gE5Sq2sRuEuFjBpKQfvLoVVJx0d/9eX12kj6IByIcEsFTcarPKpB46QDTuQIH3z5RpPMXo+MHJEE
yqZohPU8rCgno8MAlvkYvK5T92wYhbw8wpEQGwGQUh9D/MNuTJO+Gm0MHmN3I06pU6zI0Boxwcck
wkZWTGI1Gw0SuBnOioU7+vhBBj+p6QfLnpzS4Llvh61KejsBfekNVREvEhJVtIQj7Au4LybXGJ4E
gJtNrA4LRhM/lGNWAgk8JV3MD5froS/qkEng7p4RuNU2ngnWP5PelnAq0J7p2l7bP1hf0CsSvX5g
IFSqZooYybSDaLuAPrK/xkhB53yIDfvrCeL+suY4ZeOHya4AxU9QDjWYRDZADzgzgFiSV61qRy53
N91z3nGzzGTc2oO78lyhBhG8DB488tXJ1OMMvHUpzNK4y5+mp74SZW9Zu+/HGv8Jb/Gv0PGj8qaL
5RAonjqDxg+0ttbggH458fUqa+CSPKWAWSbMhE182uFpBai5paDwqBu91aeMnMej2W96ndoFDin2
NvrRGhQPWKadICCS0TFFtxrGhTGbFlh834Ods794Ox7sLllB0s2B0+xgB1wZ7WPH4c/xOtvZILdn
5pKGMTFyz5BALGryow+GHKmnYArKoF91fE16prxYJY3nz0TJMO75yqKxXDAUR6RrBYEzrJI/gLu/
6MoiVPKvi/9QaLDVBgQQMOk/GKTMpP04N7SsqsN+M+vaZfbOkUzNpCfUmsEMOc0882eY9W+mdRTC
zEqsO8p4vYDFISAN+XNGoa/tzlkRcO4bmLHwRd34eRK408FeUclO+0dL94TEe3aUkq9idNub3HFG
U5X1Yrb6u+n0FSAc4VbUIxDvWiKoulP09GU5XR9Q5K4KF5RdCZBFcC+0esys+gn3jO0Gg90ej/VM
tuJoarTtVJvhCbx98mS3fWglBkaLnr5qD8v9FU6IkxR5kjYe79LP6jyEBydX0FygQzlFm/E3xMt4
lsagcSWQqz5Y9SW6uN//Eal4hXd76ZlMrRdog9xxQrf4HOwoCIGA94+lMV0Q5g+mUpHDWEyAoltb
Lh5Fg36QP85FHfcOCvscDYguJtFkz7NskflkXfZahunbRc6d1w4BbjTeavyM3h1TyvaO+sMSOafI
cp6nxpr5kpO1LQ2Wto3Yt7WbaHe/AuYcjaN6BuDW6OVgvSHz57wpRV/hIV4foz/T1zozqLciuwPL
JaCZUT6H4j68X/Ht063P6JqnteFGQoLkq1kNeXJV8EGIly0w5nhDnqMChZtY8OUj0Z+QfrI95g02
6TqZyAbRGiDT/NoPpBY8bdqeFw7qeOjosgV2qsmqbZyU+DWtuYSndat7+BAmEQlyqNGF3Pvz2MLH
SLtqBFypxrXCtPs+ZyFR1B8RfgirCxlL6dEvVYltr/TzarWjnEh7WexGNz62JwvCuTWbzhNMPVyQ
x4PM8OYLUin0AbHdl9oTJsHfP6Z9aWihMaj7HQhf3LUEGPMF16Gqcuw6SYNFom0XB0gziOMoO2v2
UtepM6O3mUCnD25IP71bT+AVhD9M9N6FbS9B+GVVM7u6ub6BYlrwUvNWlBK+WM+IMZoeG/OjAb1V
xhlEITBohrA9U3woRIfRGtxFgt1w0FpzdmZHAVwovK9aQch5yQchVcNMmlUPXBIecKdFJpjU7Qp2
V9KlS1gDCZAC5CGp0q6kxD5mI6HRdXbe1LzWFq7tEjJLb/QpJeum2asnzFMKRBHZDZUpZ0gerzvl
ciiwyASVm87x36dsZJ43R0ARMxWNG1APSCgzMVB3JWEiR9IyiicG5Uq2BEyZrk0NAxxJp1cr+AhP
oc8PKQbBCjHG4ogBFlGTItq4fDAPeWIZPzbEqQakW5HrqX3d8l2iHylSWw538ozuzXZYpgwOaKF8
cr1jk7eiYyEMmJHMrrr7i55ArDAPnf2KIRxxFlb1vpk1oqLeAOb1FB5E9IHg80li4IXGag6BoXbb
y/4E5Ya27+ItGCmg/lR6aST/bQ/4WUA9h+HDHwD6yVD5qq1WHHXoumby791NlxPwdC/z+n3+1v9V
PH60ubQpEenTHe3eXTHl898hnD1VPnCd4UyKwZRvLiWDpS88NAsFmyTRx3UOTzeHQmyJwlmr8uSS
Z7wFcvssE9A7c9RlSlzZlSAFLmqXG5oifIg3MEO8rQ09XEcyKBJNTrfEzx1JCB0OObqRW+IU2tF7
HxVPwgT9VVGurL9gW8Dx+jXOVAwtxcz8dTT6r5WR6/ZLQdgyptMk8Sk4iZU3gtuzi2V7ZS2V4e94
NVwFycIFXNcc315dA0daqKBqDIAMZPZGG43RVZUz9wdgQlGLMrEDq3hRYG1OyQzXe0J8kZ4KaYa4
OREFefVxSIVITBZP93kr/MdkCgYD1FmYP8LZZYiu31LgE3VLrXtnWHGnwVLol0FFtQadm+sypNUJ
doyM+acXI6VfpDWdv2oHSHy1e/tPAZaen9k/KghQep4bQiKnM4SKxaLzCLae8JxnlsGsuf/i1j9j
p5exUOX+IYkJdI06kXXSkSsouEACoRSTAo1ehIBjuqV9vR/6XdU2ZSqNvRk+akdnnYKCBz/zLl34
ZevxJhW8GsQiRlH46jL+7cLvDK4eEH74U0qZu93FvM4G9xDRU2CGNrRVQquOHPTE3SkPUZWvtLgQ
nF5e44w8S0rb6QNhIkKbv3omlT4xVcRuFP+LTcQuvDu3/nljqqQYq8qSXAY2ofId9YDjPoJ9eroC
0om7w2m7Bul08+c21r55VuRI4ajLetLQ6dEqYEuNj4oQ1JMdQqee2mf+bzegFlFzHkeclC/Fl3l3
/Q9Bz+975UNF1rvmLLH5BIy0xj0qwlw7X+P533UJhYNxpx1JsbKVMdClgK4fnIBqoiyOhMBBcew2
nRn9UMcXlDt6tih5IRw8fd+Cx5vxc4Qv7w1zWw2he5EEMWclwMbyBhP9szeY4DFQ1buATAg1T01A
cgpHDri+7d6RYuXrXGmuo1IlvYrzPxfYjLGKvBn9ggfuAEVewm4J9ytqEXW2jNCL7BjpjmaF19Ps
YPc9DkluXldu3z7+e0XZB4F5dh8jA8ITO8H5JI7jlU7u2L9lBisX8bvJ644rV51KjiYNZ7wjT7/H
+yWrXW4J9lpTcXyE0VAj7gjC8SY+HGWs90uDsparZlkKsFnwsXsh4RibgO1ewaVJX/x5493h80wH
rf7aDPQoTNH0puNhY/ma68kYR3tfTeP4fi3ZkPms6nIapTr9eLwnDxPOylBteZycl0iFjBZDvHbK
epyRalgui7gPUe4+GV4/VMvYJRkp1v3eVhO8OBiJi+dQ65Z4jgJINPg2WTN1pqjmd9GHvHEf21kS
driFIBM+afdYjcXHNIyhyALERYfyE2eUy1jud6eqpP974w7aRRcJkuKWC8wlmCwpxPt3rr8VRFWN
2sVDsCs6mkIu3LuBRZ3omDNsFNgmz/C06kV8YwXXZ4MYU927g0Ry1CIrfEo3933AFkbXwBf1TqpG
PuL+1oDzQMLo0NrmXORhZmPGh74UnTa6gCZSmLTEHftheNyvWm+Iwqf2FBPhIOU0p67nmwTMOcRD
kzjTOvMS2wonyrm5Az1okkuJLlKXOpAQOA+/4Npw1TQ0NDz0AiYHPDFJElMocpBix6hBWJo5OiUl
YJgeQjFoc5hqvakB2A4ICVuFEhmPXaMnh2AVpKCdq2pDrfmIUjsCfS0bER6XP0SaqOxTR8B2dZT+
UooFbphYWYx/hHqUdAjMRu3kAw7B+McAluq3d5mkS3KIGNQ+LbrYdf4vfwzV8AAqfYc7jrdVSdVX
4hoSUp8/Kh4IF5iYxk+JBfMBRGH/0E5dBqYdO1+qTTstIPPntPiHTCBEa0sTBJBfqyDPdWEUR2sA
Runc4rY9500Z6KthffxuS6J7VVs/sEiubWsbtmQIbxw9eUGGrly2aSjW8GvrsF8kzt6ixkcbcS7Y
dUCgh54mN1VGwTxtgfMdPQ+E+9BjJp7s5IW70WtPSSWHXoTUAlR/1sjarR5ihlR1Md/ZF1h9bEC0
jdf0MMBFPW18nD8wKZVIeUFgoDhMimbrlmbp/oWwVPC8hmt4cADFnfRIHXPxxQQKxlW/Hi6P6Ry2
kb7Pl+Jdpzc8cFZOYLMQbbUKAWVJWB9T+Ru5iJJJbBZXQrYwrYvwGA9/NaSEaxc8pzVcf9gRuvdy
mptsd7X/mwMw6rl+s7zKa6zur9eGwGgrjcHJ6NlzJRf8G9wH77QzzP9/IowpFe8/crpQPIb8fOSO
UuuRpR2XgKSzTB++JntM6pfxaX9rp2NLU+Q78pLxOohFtMyQvdetK1jfwe8tMpl7MIxwdyMBWyOY
m8S60hMKfe5/woKEBNa1yoPR4fQLnrDeGiogYANzn99tI3bJ0RBs7+HkcmdMAEWQoh2yrkLYKNHb
3Wo9A8qaXJW+3AnphFGYuaj0qjUWO2ar6FHeXfJJK2WXjrPs0Qc/zzgGj/Eyvv4CDBttM7ypZ2SO
SQTlHhaUwxnIhZyRl5X6lhjQ9FTJV3p+6K3kYlXmtfGbMxSmjwxmQPBr8lmi3Zwao6Y+PD10AJcp
a5D7m7xYIvx+wJpIaQ3mty2KHgC0AWheqGmMFunfCmmUMQ2jmDVf0jNi/L1fLGbz9ivGQIeU48PK
kAkT7bhTK1jsZhZ1iqflePJw7qLuGDRvegl4rM5JsgXxe0AKYylB6h3G/k+W/3auKHOK0U52HTOo
XIFgQRVq0/4UUsDhd9P9UB+0BOWU+bUmRdpSXg4nPOgMetB9pYO4ORnBbHv0v4E1LrIPUT9Fe0W2
g90AXnRQq6zCicEyKFMbeLjU2QrK6OevYy439vBOCQuwd0R9gaNmnFKq80fLNzqXn818BW5SXZM0
6JVqSwv4MG9ceqByeZMZqKgC2ig5bFetdIMESMarzMky9dxG/vI8I1X7PNtsUv+FRCyEs0S0WOky
wx8WIcGfUelzv66hZeZ329eYfpeX+WqTxRnXCB7N6LrgtUgxbMI38Z6fET4b5HLb616+Ko/83eD6
syj3fKIRbkcKkrEH1hAo0h6p5DNfwOG5BSplLSQSougHjbwvDR/0GceZpsrzKTUxL/459PkYCJgr
q7dGTwu5P3oyxCoCEAXKs0bjMKEpJ6hzLJzJMYj/0rnEqAhc+BqHKIrHWuaBmVlRoJ/Tm91lDxOW
1Bc1zDrug58Jya3hNRBrAD8wKqq56FC0eAxAUedIRXpzQ8tohQjfne0pok7WkK6oNjuuYUewrhsj
AZaGS8tK9a6AljWA1huhPNW9EV6xxqpLLCO1PAYRv0eX+U92gqmxBaifcaCivSf0jDvvvB6qjWtW
qGUqRZdJcBQsAryrhaJLpQIWqY5D1JEw2wd5gQtFObW/BQgHiipfpK4vDFHfbMbnHk8DJDYENePs
5/HDPkqYmEI23Nqfxpgtsg7Qm/A7KHh6Rwe53pOgd1JmvtjlO6pxieHaAj6NWsWno0kXwGJJilmN
/OhgfxRJfiuSzL8wWH/7/rpZlJkSDUaLJT+kDv+99vMNO8vl6jIX0CRngqoSDW1bJez9+IOSZPHD
Cxe8WLFuOutY/Is2nyzKgC4cvhIVig7U3o8z4if7PZZ7T4LjEj0wmW9PXvp6g2rEiN8C0E5pipAi
I1OqMhlNkaTO6Xhkarb2RXtOCrcuvndCh/WgM3JFIduHpmIagSPRLOC0Riz/ye8Dfr5e+fd4QLBN
vlQS0NSzXPsJccEJdWOCc7mHn7Mzc5UAvHfbI7gBhi85QH+/+ruw918k0jNgZWjumlIOIbdUUr5h
NK8mw+4oVszMIQKBUW2DG8+OfySXiCBqEEuHdzku6pO4DvabKWMyuT4ENo6LCYofl5xDG0SvJR1Y
lNnUPo/wdVNHEB91No1UGVX9FWwIt1MTwo3J/LL4/xUMk8Uo5hPEDR9pBIEAYT0XJSE0T1MaWuE0
3uS/PE44+sPOfxFEgjJNTk51HzaXSNWByCIIN8IIo751QZ8h9sG7nwEm9b3yKQYTCJx0uRGwBo8+
AWL6kJ1y3gLh3Y/3bBPkivnMeyn8K63xzyLVQa8+nBDgkmB5CQ0pThPpenyAnjvraOaYNRFe5vkN
w9KUVCXs5wclsSNH6Aw9aTfv/XuPkS0NcxXF61S/OXMUOIskZ+L6JbnRb3jpDbsgOx3gaLT0LIWu
BX2Dc+Cck54qJyYDunXlqm1Wj/Otw4mw5/Da8pq0x24x9uHqEWxml5Vpf11l1wa//R1CtbSQ8FjP
TDJEsuVpXm7kC4jjxACYgSZWJssqr1n6nRA/09FQvJER2GGqXqqocj+kCh/0AFz2ioWhcelRaUaD
V+AX/RmTOjRLeRcz9d4cK9ML96EnRcA9WGag4iuYbmYZEB50VpNiaXxgzVDT9jaf7zOHfJCgwBOC
P4Odj3TqWWNnt5aT5Gf2FnJORzPE0HSQI/r54DFLfoLNfUaKvd3vreDlCbGmECaRTUnpvm8KgDNZ
z2PlCKpEWMs8BxP8K6aAf/Z3z7lh8qZ/9Ykl6UE+hDDCR3noRm2cjiOZhELuN2qPqA8IdZ3Jlk27
M/OGqjBjgClQtd/1ivoNgYFigDn1BODx4/INTmiH5XvZiUKZgN7ESssk/IczDvLprtyCPZajamjK
j2GmFigrgI36s8cAR08Xg/JNPNENc4/ORJjdv2HcYnKMHsbzzLjY7BSwMYxYap4n6VnP44eP3Z0p
RjR3WY8ebGY1xfw1R3GhgQ/dT47SIck4BBGSj/zpEsfQeTXb6KfwdFL7WpoHtuW+Ec2iVBjnVzh9
kD8Oye5QS7wo7mDntA4+j1kWTiFOaGBdAm9RFScTopEs28KB8IAnsq1wETsWA3YmAeGsgtZPqkKk
SeTRMdRC8uuIEqaQAruXubTFsxIGH/YNKLijuqjx+4SU9IxzgCBIzEs3ywM+2CUi4sKsFOXbd6CD
clazYfA2uKQwuV/Ib+5ip/VfjvBUtm+7Msht81UYYeAqcm2Yslgrss8drUQXu28Ehs53CklNv3rM
6pOQvZpMA6mZVAYnum7zcDO5ePLuc+rcejDLo3wU/3Uas3G+zohRVEFGrvE2bT049W22u+ZHt6BQ
/Gd343QgXdUjashpo8Sj6gaBAPOSfDpJHhbu2wwI+LGycvQa5bA8iQ3JHJ+TN6BXQ8nHd2QBIWtz
qUr3TuPgfQwIak0a4rqZCGOIlDAdI/mP7gs1pBMAXZNUtpBQBj+obWR7Y93fKPK9iPwja2tBGuz3
yevwdVDPUJpM+0yXWFomLCyrtIX9TE9wBdyF+TW8/vFJ7goU/wWGtuBXNAr4MtCyH8X9deIPmIRq
v86sUptDFY0vSAH/fhgeZAArzyXCRsK92Vk1xHrNBWu29oRwZqRNaWwDi1nnDVo0pzuv59xJI7P+
+asZYOWgO1h6mI+ox/6cCQLSZuuRNxVPe5BFYd8Mntl2bJYKzVtzcG1qEG3VTV4YEigNWLzzgQFK
PjO2Nqj3D5qPG+wnw5rXvKODkWZCvtDH5cQJOkNWr+j9DYRsi7qmdcPaC+r5D42Q5YajUrBY78Nu
1Uo5Z6EYteznw3k5OEdjJZlo2Khc9Dm5WAjaUB87vV+izyccU+LgpNuuXNQcivcfTTugtE3RpC4e
zmtJG6xbGCFgAmtxDoahg+O2PAlqOkSkrS0hoxaYhLuO2xEsUiNjSDD31QiBZXL1QCJirmHImfO5
Z/DfcRTnp8ngXcGaRGjbylpyq7AYBEJeMhrmnqVt/8CgXHesK1pZeHvJEhpo2OBFMJwQyXtzpbtq
UD6exOizEvwZI2kqyam0WOr+ujsNSNVLFgYdzgVSS5KgRbc1M63hfQtut7nwOfUBTNedRIvEh12L
116EExGXF2feZNIwo+vCWcX+Axw5dan6WL/JTqOVfSl0fHrAU+2KZpmM8lYjpAd+5KmZzafc85/B
DQYrQcjvWs3qJddPDqGGSt/qGXF8Wcbg9jDckwUtzmOWbH1tRr0CsECwEJVeqmwwWgDqkODKAoDY
7Uj2miWZeQF4Qkv9pQOP/XOU+r06BSdP/8ZcpSNER4gp88GwDM7ERhroaAGvACS92+4P86Hm2RxV
NcCGsbsFxX5AF4v3qnGSMOLjXVH1OUpDsdN+MowoV9ua/fuH3aD7kgByxSyjyUK58R3lP9hXYQOF
H+7mS3JBqNdnHuUpGeJ6WUNYoqzu16OB2tDRq9N9Tu+PAMULQsdIlHat9Evz7ohOAnHb3dfZ3i6J
U6X8CDjkCUR8sxkF+n/P5yxKGt+CRJAS46Uh5I6TciZc6aJEgi/X11gL8n6gJZX4HoHM3/oFqh4I
GteybMiBFCY9meDFfLkRyqzN4eFGVmzu56EzCTg9eCm3v5nbXB+ce908GypXjHYCg6xqaJPf4Njm
LU46WZwoWofinQ/Bh43ji2eYM7IEee1tSAX/+DBV9MLvS6S2ZbeCwFUJehe+riF0pmgcWTKSrNsB
+EVLYA6hGG/zsarm38AMA6NcALWi475ysFsWZqgWO+itAG3m1TXcF7Io6JiCkLokOC2JW55YqRT7
byNiCEhEn+9afu/5JKCWQKZMtjCuka9E7XKOoUFVgpHMu/LCu/v+L7ukjh1AyjA4Jtsj+64qxO94
lh8Hz1hOxUR4AyEK6K7V/ALwnSUlOttQZ6y8QZV7gDQPd32j0BRdK3H5Jn2z9QCgZ7s/juFqwyOZ
W94k8A/BaC1xFuRmL46hWKf76eFShw2SLiv/+XnMwTyXbKEuKruo9KXal4zogzbftYRbovyeA5/C
mr/YSWLpzU066iw0ox0Xf42g7fARxJO1Fyo4Qltm5WtD0pxwUVheL/+XBdZoUgGV1x97pFann/he
op8gXpgCTIZKyyxP12rJkMCzhbtLMAzfw6DVSA66jmNBCrdvGPN9CO14WyN4SRRohYyPxAoVI5F6
YyUcQEfpVc8sL9foo0L5D514z+B5v7fkGUlkOyQdOse+AxlS/HMR2hPCc/4B4Glpk9xpefELkRja
nm+2tgyGTc3fG59GnCaVW2Jkigbiw/Glwvo2tRrOv6qFL1wj4J/pfAel3MLMOkV/tLRI4GfIXHy0
LLUlA+ETdBnD92nshcmqdQ82h9/bIjAi5IBc6qOtitim8/jLNnpsDLROiGZR4cB1fgfb/zh1/cOw
sGgOCLiJKiLNySxuTnAGT7N5Lo6i7J532PFv1Z7BNUN/o1Y3D5fO8yz8KVI51dv7LBEL2lbSOFq3
MavDR6NNag8tzwznSOtqX22iBVVJHH4bGk/7AsVpztSIdQylNzYIB0Vq4tCyyQ0jTLsEOCJBILMy
nCSJVK94tcC3+b0YA+ofHYzqBvW5KvGvxSsIRyl4rsdAFwv+RJLxxwTkWWqIM2FPVY1B8X8ytj28
GoiD8Mtc4E0pqET3/+t5+7UuR/HDlGI5k3T2MucddIrz0vv+k+WEutfxp2zzTle1s+oI7DKBGn5x
bMZqezxEtdvjC203kMealTyaoRKgYEAg15RY6BwCSp8Iqbtabvsyf6udjKx9xOnk8br3X2qCeE7T
0K/Et8ygyZjfR1wCR+0fegi8H6TUCA38jdu8zP+N619sJw0sM+ar7/qVqU6KzqYAIj4PC7fqBISO
h3+2MK11iermp9kG2Gv+OhRPV7aDhn2h4SUPvuzwDSo3sibY2LBxZqYU9a6URE38UVqyKgnBNjxW
IaqWd173L+IoxGM0A1mZ2XkU1iqx0AJSmus+BwPDeDlBJNTr558PFtT5mZky/a0r+RBIzNmkzdRs
WYf5A6sKyoTrZp6YrOM87OeOG38jcoai48+wW48Jc7aLxfUYkEWjU9+zfH8qqY7jFHy79QbCj3/P
6WTx3YUO3eTxvx+XWcJ+zehujuwba9CmUb6i2V7ily/LLnz2Q6K0MyuanBqwsV2VGkfCmdn5JT9c
0uNd0EIEnY0NeymrAqueIalw+8gi6h19wXWvRxs/x3r4q+X1Prme+wZsKDq7KeRhbGEXXh3RLSSS
H52O7/GCSJpl3FnG78T7Ga+Vf3OMSwI7dg/KnScohv4v5osoDZKvqJgImMTWVTizhg7u/Tqj5zk6
obFnNc8wrEawYt2d9r/J56q1bAEAmHEonWkYWUtsW7VWlL0xWqkczINcr6WRooOYiywGbjQyCFva
6Qn6u1K5SQhzYPuswKwisrXnHlOAoQstis40lr7tJr/xbRGaWv3LuP2RDrmSSwBfIi+L+IbRMbar
RGZf7AsJx1gBzH+8ShmNWxmKky25T6ZxdTurPr/EdEZXWtCQr2bBhi8kU2vZcq4EWGFaNpDXqC9E
ljFMjNBPnmPGWwbX2DPN3eU7Jo6G8K5DpHJuyPBAAvF1bHjchirKYkYceu+juuGaqZhSjViivhTC
gyY3uWkph9rpTz/NN3Emi9itNc1sRV5VAdQLEjAGrUhNJIHHbgfbnOiVt/PfKpHO+ewZ2NNhyR+C
HurFbaOi0xjtEFctXpN3nrgwdCcSaQw2FYc+7Ou9rCe5jolbnSpbS4QMJ7yNkjXcM8hKMfL26Gyr
HOnRoo5KKHf/CwbvfSiWMGMdyBu60+IpD6sWOX7PArt06GwHiP8ToA1CbtyXFrTjbiUZgA8nmOaK
xzT/DCrCI+/N7593/W5/8feEvaR1lXoF5lEcRoELvCZkP+YUhy5N1iDjsg5DAnqJATrCM8ogeV7N
/iODzUEKmySDJ5Q+bfyX4mqt+55+W1cU8ib+A72Nm+waoyvq5pwDaTxWIqg3MsBUJf5fmJ4+VSzO
YwZSSY0dFiv6vGn9fT5OL2wp/jzfLlKJU4xsZyEDA2Mnd9A66v4+MCLjEK24xaIINBgSCaqAwmS3
sftXfKWBuQOks6KZJipf+anNnMalkDItTrFm3AK3WBlRN18fxlPMimns+XgkszmmTs0lPDKkx2wa
p6V3CASfaKmex3TKz0zVtl66Mi9Zg8dtX1tT0iGorXoWj9/GWXVudOjouggJCfPfjlkat6nxgXSX
afcFUMuSUQFWQ8Em6zX5Rx2vXk1E846WYkNidrsbjUiM/uYV0Dj2eJ7IJ/zHNgfX5Lb9DUatVDzY
IUdsQ6ErNgQCPiUXfoXKBRuOAFh3ikKiY9bBgoTd4VbJxwX4AHsEPLGCKEEtf4nuMqZzkTx1W0hv
fPY8cQfmXv2aHOnpv0XKA4B4MVSc0KJ5ropVeqckwb8GNrWpRGIA9KE+3Zry+Eko/PgdQdWABUa+
m+4f+sSb7StradY9+Hz5gG6gS3Q5/8BzfElg8irAfFXSH7lcR5QHXx5vOEbK4ZCW9mwIoKBcMpoB
+ahq26lu48caIjA/tR1BMx32N35ucGkLEYo8cqN1oOFG4Wg7zWxcUCxyhxqBXLY8/k2orVbqljU/
GKFjfbG+SoWh12VbAr473Fte6m6V8g+SJI9NqTHPsbMxVJhF5QY+Y/4CaqxxNLryQNYfVZdoDiNw
fUsrR5nUG3VuSk+4VV8rMXu2S5fYsNnbxYnsALYjKJ/N8hdd8XTRColfN2YKK2O4KdSs0tgbDZLT
WAhJMrEaQqgkXzDU0syi2YrQeW7ExwGXz1s1qJ99N4qZb21//nPPjnGFhRCvhYLXA1aHNO+Bsi+S
rlUG5DRSdumOB+BU7gd7nqCWEbLR0L6QpuMCE0fVzPw1TyV6IH99mIC5h/p8KDMEmZq8yE/bMcwJ
o1aawiQYcn/8VS9Xlzd2iTOVbbaxLTnqFANYd9nit57mnMc6RSL0Y4jEZhRxj6UGcrH0GjZgg/xN
8nNqteuy9/aBQR8MnEo1SnIsBTk5qOxxraAtM6hxtLr8IZadLNYMBXna6zJadnNtv/HXIjnGZa9x
IIV5KjidxmYhPpCUv9TDgtrjD08qV9VBrYo06x3JGLNaUlJR0SrNpViH8OkS4TG2Ja25EwIBs2M/
qcg/yH1bB9PZTCSd/KtCpemXEh3+ajjZutop8RmgC+8PDxs0YWHS75HKC92ktrLqDS3UT2daLwEx
aUco9ii+FLjc+ha6/p1JXDyQMyRM3roL/gsCWGKmmTuM6xsHazSZbB4bt6ODY9UcKFZYqAl6Lpej
NJ6MNGIJHu+8tRhC674GhzpVXiYxk+6Vngr7YNs8udgD5F2cJGlfgTI3jBcoFr3KUH8vpR0f1XJF
SNHMzZGDuKbDcxwBL7u8XSK0xnS2CpE89EpmbChNnSxoQKwjr+ywa08bwmjcaTIDyvgracbKFVY8
KxXUUOG1RDxeajJKArndEZhMumguZ39cVBdH0ziHAbm+LJYODLSMOs4fF78GBazfwAtlvvX6IeY1
XeKar5lysXg6i7HrPtFpelBD2ROxEhv6tpsRiVAvCBoGiJE0mbhYg7+lEJv42Jvr4fmq/A+rTNxr
HL+vSXCUCX4FxDMbaPJNfFmq3KN4VdZBwwo2KIKnQ3hN9PbfkEYiLH6qYH+V255/36iRJ3/3Xp7Q
LK9YwI6cJRhd5IbAqCVRfCJJ0S8XWCti9AnssljM/sX3kFZmQW/Uf/dgDm6MZvMDXeRke09rGpE/
y4yzyITohdnAQSpfa68akOjJMzgjzUCa+PzYeByAclYgykJ8AKRl3HDK60cJaXWzVmwaxzqa1sz4
ibpnLq8964rdX51cSSW61gB69v4z2dmVjnTrgRMR8S03Z1Ag7WjLeoTBNkaMbwYPo15YQhTk2Pnv
HXBGkHpuQ3RxabyX1gaOAlHCgqCmis01WWU652Z+8ZnAOSikHPy2KxTeUJJGOkF8Y7dVIPE6mBdU
u+t9CW5gddMGhH1WBsitt01rJL1vavQpYJwv5hkYkaUHRJj7gQpRhgbJzWYcSzXortNREcO2OWnw
1SUtgopWzWappqSjG6DYsfqeude61zSQlNnia8g0nG0JgPgWRymLpjrR1ujb2M1V7gNKanLJZWrF
w6AkeoTH1/8AgbeDI1a33SxNpHbwti7n0YO6Ew28qexIiKYQX/8VzEtZz5lkMgKPlSZJ4UFVbGix
v/KNSeaj4+3uxfUnTTDmeXC/W2tZw6pGQ3qdjkLOhtdtc3GMMOks8qFgUR70urS8re7pqmQk30ej
YD3u9Mo1U3laZljCnevPk6N3YrZSxT6CgYRq9Thoqcu30ZluqMaevoE2h8cJEmvM9FrY0J5pPc1b
9dAMGvukjbx2RaWdim2XAIKUpf+Fw9gjA8zPcoJ0ZJ1eSk0RbLMPvGNr4un3Mhsc7HQmsdsCEoIR
/r4nNpUc42mv9ZJTrXFYJdcqsgpL+t0WVdsgJ8zse5Ptuk6l7MzHqEIc2Qj5Mlh0v/DGE84+itPD
Pxqt7yi2Ax9PXeALp2KUwjeGpG1t96Kxc/KAWHsgbH3IT3r0aR3H57y1G3R2imFckhHMB2CFtI1h
oTVrRP1fltREmOxVLCHABNJm14ulW1ytvNsPbHxW8YfwtcIM+okF2ASQW1aKwV2VSZiPxnlIAzSM
yPFtqAbHjeEEkIE97HJhbrFYr+4uw4ayzrugNGnG/Nbzz51b+ZACTXeaq3QDILxkjjoK1MH/cSD5
2qFotFGLe6zSAuLDh3JMi2WeUDj3hMKlrYmglteWVZyndS/9+QBPt9spLCcZAD7ZXSitPOUZcL48
0SS8vJxXSqGTdrfUM84i29fzcd0+Mbr/RF7/Em4nel0+cf90/dFkDe9k1Z11MU19MjHhRRxvIHlW
dFzMzTK3i5r9/GCuwPLjjH+uvbxwnFzvS6owgrpe6dPhqRLs2lXdzKXKqpJNMmjQVBYFAEP3BN3C
bWTatNp+luDIK+Myxs9DNDqg0QSis3DskdLcJbNwOQRxkRMTqPWM7MJQQ4ArMkDxlc5ohaHtl7aC
tLXCk2T5deuVuq7FAS1wLIMmJ5gr5UBWBmZIz36lcMlb9gAv4AaEuIgmn2dyz6Glv6IxihwjHmNj
5Q5lqcZvUUhp0S9wTt/RTo6O5t245JZHKk3+OQZHSQuZ0fMqC1aZcZXmoDteEcKW6XkBU/Lkg5EL
OTs5ayT68RSd1EDJmJ82Z51ZH8FW5UQvtn+fOQbCMh3IxLoNnFBM+7e4zXHQ7JVYgukfwc8Mbrzq
88AkO9t1EhIlzAmi89KBRqL/sWMRnWYezKfBnrv0Di+FKSn3j0cW85pbOY0lHJ+3+V5yE5OwvF5m
2D9i9uSJ8u4j1B2iwsf6mf1IX1VmJRdTTiRCLeqk2OrK8LqqDO966o+8TPRpMO9903ipU7kr5Flw
j5I0XXlEYGYwiJwR+79pvjUAkaZCTun4ICIKvvbMLkBOxwg1UTUNpV7sW7+XOM/4fzuEZyjEkoj+
3wpMoFSexjYZnjiga7G7S4+gbo4EF2Bx2LhBmyKFBzm83BiHDXUGZnRKi2a10mKRfjAJQ5BSaFF5
nP/UwQCAY7WxcwlavWAWyYIOcI85e0CQAAiL+/Qx4pEttGP8FveShmZK2AtY23oBm4Er/v67fIZE
QEcnukoNVaKH52H2HDC8lyBj7nak8nyuZ99XInrD8tY1ufvMrCAZELDZUdRkz5x20wduYRWo5dcD
LYt5QnkUl+JCBjDG+T67LnWOtTGoyZRWdiSsr9RgbM6IwuZvOo22FMxjN5GeXvqvtqT4zx0IbolK
kw0jwVQYfJgMFsZnQA5nUTzPFuId0e6bUs7292V4NXM+TcSWdpZce9T45VPUANIqxDxJnZAqFGak
8RoPA3VQR8zYYKqWmMroqxUpprmLHNZvH8srvnB03JrD+EmiCblLSI/VjOJtuFtA9wg6Kwh6VLRv
TOa8M7cSnluzPn4zhtVNmH2BjTz9WfRKUh+1oCXMPhPU4QLRw/MdK1nqz+1PeO5biuowTMl5PPlm
NCoBIbHeZ/S6XHiybsktAIHxBtQBXhRjAvcBCuqq56xjFFYPIsJgbTLDdELqjFraX95c1Uv1Q3Ir
k8/FZid2Wt1YPQEVlOc0UN85CXsF1cVngF72m4u0SoexgUDBN22X2QOSm4V5OQzcFhr1SrGGiLl5
4yg6nZt+H0xEg2+YR4BQB85W0l5qNvZretOhmukeY4DdzUlUHxsPbLtl9xPZ6zG92FSzdJe/vn1Y
ZdTo9uGePhCD+R1tFhWXW8Zn/u8pObQ2Yviwdwyi1dP7VX/LISs+X8vLDGL2p2KqryE3+9gk1dbb
tmom61skTgMEu7fVJ/oBKQY7tU69dNPKo/AlQan8dPLkm4f/wkFclEHdKZvSQdWucMAq1opKaYka
nNobz+CVS5ftPsguESFwRa+lqRLWWnDMLFd4jU++usvMXI4JL6K11aGhseZEHcG4D7zKWCFT3zmZ
MONxlDrC0cilKt15YPtiUf/04wLvCAoTBpxg709OwBRFkW3jcYNRr7OwV9uXEsQzPaT4whRjpg0x
kzHl7Pwq6OsNqZV5hqVfYJxvSxPJcWtMe/hIdfQ+mw06/6jNpC6nPmKRUd4A2C/R4cEjpRAHWnOQ
psMFcFc0LcsYFzetEJ+nh76wfPulmnrWm2nEbWTOjIlGAOx2ROw17S79XTeNcfU6WPNAQ2/YC8lg
7xQUnC9mW5AtR8h7FCduEg9XbgjKXausJAIZTRtakWa69BMXno/QBYyys0BJves1a8hETIwXIXL+
uihp2C6jeYUd9TGUPwza24f36g7NCi3ONW6EGi5LX6A6uCojT+A1+DGpEdIAYq1F0tCrvCGQhWIn
SG5bmIOQpCFnLaOsxz2Pa+hK97rYI4/Lbc0Ui+q/f4XhTNh1g3xU3ovHQpt74E2es3sJ+3qN2Z65
0fenqm8BW/HS1BnrvAYiQAlkZEkeUVe2oRGQ25w6btcqUxMCqcUbc9CsBsE+8W8XTvc6tWnovfBp
YBLVKQ0lJk2D1MsFcihg9vrvfVcQEVH8FXA1C7+4pSj7FUjtfPe1FNKIvjfWrB7GiYvyGLZU9sF2
a+Ib+Lmv1eOIqMO3UwqEmA9g2E4Ff826owfhHm8YdgkoogxKI6DCOaAevPHQ0tMEBkppn7+zlwG5
BMlWfPF9mX9dWY7UwjQMW/4fXo0c9O10zNYEWi+ALmKpiA/ExUVSztJ5OTGCFGlO5P9V42+rATru
gHyp9zBgWLyGPzk/9ENCWaY5mE9yhoVAUSNcUcIdWL6Mf7bzNUw3k5tsCLQpujjMLl1/0KFpX3w+
iqfQU/K6Svj+85GxTeTkcM9gQBH8vZCadunUp4/qNGv5vkx1Girevs9dVmMP9HNDsytNTNBA9xUE
e+ut/LAKCOTVZIinX74MNA9opMKhnG6GhHw5PyVB/Zom3L4yLnjD6MNKVYoEwsI5QIFlMHRVuQaj
2+9Li9p0gphk3ZavWxYM2qpvFQjiDPUehOD2RG7rtPHTcyfCccN1DHuQbgLFlt+v0ibRZgNTbvJy
+uT3ynf6WgDIl3rgvbnfiYDJILYOxoaVh7iMT7t8eaDhvNqF1FQ9sxTOnGhkR9mrhH4VfFRVsl5N
V9ObyndRv+lDBCowaAelcveTA/E/Pckalf9ckN/GCMVY00JafkTsiH6YrHBEpzK4OkswjUqs9L8U
ILed13wqEkFF6fTCF0R3erWBF28/qZW/RSOBEgg5V8F9o5vElubvUgP/rUz929yRzBreLyYzRK8F
CwNY5dOMKLCm0KDBBSlHK1Oz5Lli1RQGpezT0fdsIUI5nTkWAFVledgKbpYKnyfYEy2VrojVVb1k
ZmjlD0gyibiIl0v6tpHgm+806t5iG/2mqXU+gl5aBiV5rWyVODoVVM2zf/pNWJDXTAkvRNDAvRUL
ZTXGlQRjmnYr7V9KxAeKhiDYulLkgMGoBGxS0fP0yrjH8YxdG5eFMmHb8zHcQuZdoTDlSxx67GCA
nrLWYKBqfiuS5GwU5Qz/ee+h3qasBLY43GnIdCHQ4W3t6pChhMYUpOLQeED6mAc0CdyRrElccjX9
KZ+UCobE6iPjoEx+CxSUB1El/Ks9kssF3mcwNhKt2SXL6ZUE700VEazbcVi7AHc8lJQ1kJOX+bwP
dVX412Y+ICL1W59kalDiQmS5dT5mSr13yg8l1Er87JmwktI08840ChDKQgMVLgfYnjHTaWOb8pFA
mebvLc8vhlGIM0xgXfLLI9aqmrypcGdtanrlWOG7AHjIfVltwZWtJzYrCzxbc0zVD+RFmmNS5Fgm
gMz1M1UWaWoldZ++uZmwjd0auitEyLJtWy+MQKvCognPNrbuGaGBgYA4mSFcyoELVXWI9ThQ0tyX
kP2O82sip39ulgV0d+Y3SFPoyfRv9lBZjHWkLJFH9PbN7rxKd/R+bz4HsY+zmdwrf8HJjYUsNVlr
sXZ22Q5CjwawT6MWyXq3rpwZF1YfFmloxr7xK3XXENOmMAUBX3HNBzSbmxQZq/konvBGejNyfG5t
KAupXAiEihvgFFVvG94IUdyS3Qum97bUyRuEVsYvWhCaXlFJR77DKlFbSd2WP4IGdKO501pmNeRG
KbKS/aPvoOb9Tv/A9dU6MvAPHlv7b2LyxcQxBXrYQ7SA/V/ojWCNB2oQRk88ROcA2xDnCJ3Adh0v
ywVUTaNGtn1LTZmTzxutbLmhow9D6MLQ6E+kDuf96fJh6YDrAPLtNGTrfaH+Y6VYsGGxSapCOH1W
zLduLuRZc7ZILUAVgO/xFQSzVIqtOhD/oVObKY6psrVXC5QWoSkG1nDiCmDNx63kXQwWZpTZLVgy
Yyji/f+6AcJbnK64rcr5JE/Q0rDAryLVibXUk7pZfDU56NhrNe072IcezVjXdADnEAGij1S7fVau
n73iRgP6f976TMr6pIcps1U+eL+qOo29ATVYAgbB0ks3lb0VsVNOdYf0VNdDKIjcB3VH6h9YTdEK
8lf+W4Wtrtc5bNZvk4lXOwfDHaU3ZZSRm5oHaheahi7W5g6oGzg7eDCyv8JALQCrLncLQqhjh2Tg
W1Hdh531nh59O9OYQv04ydJvWWaW+Se2yK+OPimoI/RBor+Vg4o3A8qdzlO+58nlx3w1GPbgYv3T
DU5S6R776AtDrOVz3wUIBp2D2H4ueoxQ5hUNHi58OxcXn6PEj9ztuOz9Ru/RC++vWFpzioGeXQwq
BtsRiMlrAjwXaNBTOOcg1NajE7vK3CK2SrEwNuRjACI1GhnNPH//+eWk4iJhvkHRj/BbeTYwIA4P
kkwZMGpQfgRSYYZKYN8AWBAKcmPjteoEkT1r14EPLBa4gozjX/EIMpqv3sqer54L+vaB6J135Mfz
lRMjeomcRFSIJJoqfTQwOt9sl/67ag3cIpjxh79LF74/AZTqOV29gNj0F5lQh/FU9x+s0bLOWPYa
ZrX7iA6IuvSA+ftw8zmWytzDL6MTk1ovu3T2mwLcR68Xe7Rv7ATIgf9omASihVmXoaeikNgvWnz7
J/DuTbeQsMDGk/cQkFLeciViiMMkixShVugR21yMQpedVVf5AIuv/0UZ9kMkH2Mhc4+mH58GUYnH
m0Ne/nWQ8F0pCVZsOL/JXc2Yaw6SLSgMKEr65ZfVVXt4MGQN3W0UvenVIy3fdGeurVZaWFd4GPvu
iUe4E1nWKPG4uNWcYUOehSo+3oMVtLo0/XHPn4CGpqok8BEdAuXce2GycIUL+gQGoA0iYCnyFJIE
6H0bzBxXiFJDexDkXVV0273aWY9SYptSRP0DTi45IDtaUu4ggb80ONcCqrS1kOpQMoCxNkzU+ZI9
zVvsvmf1CwQ+zx8SSlYHD6dAxbYKEmrnXAOK6n23dFevmkBxiUs3MQ/zYZ2OQ153DyN+J2FRJFOk
i2WM1HBiJeO/IukM1KTZr9/zuTBNDX55aoQn3kDnUGkz3Njky5zuT8o+UiBQFPSz3Q9eTJ3SJq3y
fwHlLlQaSIekU/rRdgnhAB6fxkYEYvQkFB/nEdI39Qq/ujROhe3Bjlee3q9A+tEu2anFES4AlIi3
eM5LrC1YP0xSEGkFZakMdJgt2e0uXSVcMZX/OYIyzwNhvC3Jdk1LnwOaLUmR1BWMHzN5W7hXqIwG
NTZ6kgjoLOmfiOoGONII6RykX0G5rYoZpwrGUVQjnvFZKADgnFYqWZOP5EYlNhKtNhFsLYW4l5Q4
LWsGDMpGISWB4ALo8CSC47VS/uOPaoieuXG4dIChRM4SCKfEhI4Zmh2pHET1KyjR6D6F8eKnE31k
RtLj0sOnGmMzWfRJK+iwcvuAy78NwQ3uXeIXgs5L/cPNmMU1qWHrq9gq2OvegbMfPcqXXCS6M1qV
X5EBrWKoY5YsMwHUIq2LUNXcUIkLDWcEu1dzd01nO8UW1XpAvo+62v3V+x6lwS8ccuvVpmnL4Jat
JhTlySN2HMzRz4FodiCGpvZHYUg5GsCY+flqHvMrre2jYrpHTTVa0edHgjuFsztNpR5bN+Wq0Lgj
K/0fvtXXHqnXvr1mGYNjWwYVpDCiFTJuwq1T23pnFEEeDimCktXx7auZovBF818ZYMGK1U8BODUg
PBnw6V2B4JsOaeFYJVMP9nDHhJY4ZeDAQocrWutPYOTvgoNBuMqaxz0KZWVFHp4Q7oAQleSGHqsB
aOglnJs2A571fdNO3Esrj4eZIM31b/vruqapJNp3zs4BxA0mEQRy6/zLQPazNSzvVf1FdnpM5Rhz
q2AMX3P/65iiscsrrhmyZr0DmRxyzLOnPQq/FBBQ7+eNkdOJ4/RuwU+ty5PbQ3Urqys/a0sNXtD9
Kk7MBqrQijF2TH6WNWCZ72/EO1MLkk24uiClrpwQAkLQO/qfOl7SlSqrPskxbuw8egy6RvzyV64p
jGrYVNvV2IXFIgGOXLkqArASj0YBd8gP8rSk7duMxVIQQ9vzW7Ejz//nrxd+X4sOV+WuVgQXklDs
0fkKgoTH6cld3CGS4SfnywUeP8bCx3h0N96VGKzQR397KUKPuuEc950OxDE2keexCZUYv6m3bqmR
N2OUi4BrR38JHmIgwnO0v43D7ly9Z26xHk7DBMBKC5Tw6drm9e+Paf/j/+eT7WpYwKy1vL/VXp+7
53VKWUL6gkTnE8mjZR3vNXrywb5xcUcVjEYQKIpkRbvzeEmO/FjFYVEw1V60xBjWB9d8a+R00qqO
9yo5bLb5DdtLDq/uGVw3NuMGHVgqo3BEAAI3ipnxPdHxTAuGxlUwSqUHLUjCiAAPj0xrr+LFlJCK
OWSOQwOoJiCmeLM1WV1W9er5RQnZd0TLGYqRba1xcJUMtNDVDRLRRZHLZWO9p0uw1ysR+3uqENJn
EqZN+pg5v49TXxGTD/FmLxnT84XENWwJb6Zc2DettpwKgvISwgVWbrdNsRWNt+GZ23r4uh/+Frc1
miYoLCF5UQKaMDLl3cq8+4wUWzSb/+7JGB5tj4KSDrFj0sohV/vsTfA7tWOqefoRmw7GPxrheAY9
xArW14CMNypN1OedTojpvFOr5mFZ/cJ4BW3j5OmKZmf+veM9NhBcNkmLfhSDsz9IdUoGYn9nWnV1
Kyhu+rpjT3fLrbSflTd6SO0jEz9/+Akk1zOpUUpTRvgDtyB9NhoAzjOBLnl5WmqVRPW89Q+YTSSF
HQop4RtwQqh3K7JZszUDXFaj3+STZ1w52esl8VYwMAgYr21U+mg9rL/C5V21wGP7j+btLm9Wqoh+
GcHBV6k+x6aCwi7frelEAjK5ZVsUK+PTRkFMjk3HXPH44VDMYwKYFT6ihPGgrbgfONiACkBkh9aj
BYOBeEWOqYH78ln67yVmyoB+sWfS3yejMbS7NdxcqnZKLFKnCNjfq5XU685/mTfQUDueGx5ir6r0
wF3IYR+TgfRo7CMKEYtSizKv1tIa/5rdm6kLRcK9wwcUvhmGJn8fS95Iuf52N/+b9rJW/2plcvbw
f7oBydekZSVRZL4VQBqoChsX+hi1AYQZMBhEDIybYF7uRKzJH70Sp76zKMQBu+eagxA9C6PCzO2w
0r8Ow90O6u++afGyOQjiQpEXwAVzKSYXBfBOncCkIxLG5rH+7cYp7qQhx4RKujbc35ieWjslcIM2
4x8DS0WxxCQftIO2QFmi1KmpJDm5krlAYEgiWN84osxwKdK4DLjoj98gR9VeRFy9rPM2VnQ+/epf
t6IGbU4k4XJ3rmcew8FwWZwbPix8fT3yYpISgbJ9HFcCXRW6erc+B2rCRUV8RD5ouzTw17GUE58s
9QxihTVYa+/DWHMe0AmtYLryDwokEUozenv/+yv5ktamYWxQXVvAA+TLlfOjZUqvQAnw5ZMw1VP4
tDdgyz7/IUyrIajtB9mBz9mxw9kglb4/aR/nmcHn1OnslKVfVPv/hIvmI6RZDdi0245GddBaY9O8
t6FSYzrkQBQUhv+EMTQrkA5xB8A4GdszLEoGO50S07j9wvl7PycyMzkU2g3t8iSAwkSYvHjG5agT
A/xUfdcvSWfRV2DVYbJgxQkK+XMgvXFdL9A/vXo83d7l+NPIp1fpMlDg8sYS3Vsjt/xv8twlmzAw
tRh5fF2goWkWwtLC/jA0488t3vN1xIytGhRb+NeRHMeS0vW67B4FNH/v4n7m0n2h+e35Qz52RE4/
zWQuyr4lxuiWEU+ps0jyEgNysVVq5gKKXI2eXXOpn15aWIMwiXEgnb/wpZgCtnQsgjZkfBWZrPd/
WFV4efJpOuxNIkVr0TP2HIiP/VaYpvWHbXr3OMaJi9p/qYkluk3kJiLpr4LttLk3pwqAvKoKi6oC
Gpg81amDguE/YFnjul/vqA5cbOZJc1/R2IoFVW+j/FczjnvH+/XYhMHKtuLPCuY5tTpH7bz6FjG3
4CA0pzqnsabHH+LjbdDzAWM2e3kEQ+Wd+khDsrwbwSWkmOZDCjz///fU3P9FA7a7HltjCfwPCYy9
G65/mLLzbJCV/VLigEc4c6tfo/OfmjYfd5GfrI5I6n0/0lda2RCdW3CbY37UpXcIntyUZL56cNh8
9qIOydkrBwq4BQ2+HRxY50z5Y98nM4PE7my/OtxM2LMW7BrMSrWwxsBqOtNLL6ZDTZ1+Feaw6tBV
Dnx4kE6Fxj0b2L/+EuqJ0d9u7JHV23DEcooVIZpjWTkxpiaSRAZ1RkNbqfEiX2Irsn1nvl5LALob
yNdtHaDZIperST8eYBb6QY11LTZBXqGWtWH9eVA+H999F9F2tNIk1kiGiPHbtEjP8byKP2NlSfKY
vfegKrWwPwbRg755WkGgvRcjyNZULwRzsrgPUlz9HCQpwUU+BQYFBMS9YhP+CgCJwRgNqXol8QC/
RGmjejxqHOwHIaG8/wHav1xrxWeupU9gpPWR5G2qzxtzcXbZYMMgvIitNlnN9uwkpL9dtKZGuvnX
3DuW/BSLRQemK6TBf95rafdB/3o5DpGPhTHqHDThZHN/KJJ5XoPxR+McJC7OGRu9Q9spYYtBqNuY
67bl91jPw4WTMjnCRaQK0UJeOPUemKpl5OyLfbd3nzrU3Kh/aFh5skiqFjNgNj+HQM6TQ6QBQdNE
YhuGS9N5XSobBLHp6QnmgZdfCHhy7nOw4yliXBKBCQtkrndifq7yn9Oh1YIIYR1Sf0HpRxZ31zsd
rkPT40pvmCNf5YAMVrdXJVQozWE88Z6r9hYqQc5feBA2ea1PSCxb+GIchUWCXSoWDvhmbeQQf8LP
MfuI9wOgUbtfURy+LqnIyTfudzJ8QFIFGhcf/b73CKmF+S80AeuT948qDPVvbhhaUPbnMtPB94m9
zBILocGCbKZfNhdPdrPWV6RpyzZnhGIqmT1cMrdjNPRZ6Xcy+71YaA4KjAsTc9Z+SfW9A590G98I
HlLAyKboz32KA0jUj9ImieZ5KCv0WJ+iQlYugUQbpN0DjkcZmjFumWFzp6SHCmflHX4nc3YyYwSO
2qvyKd/FSQhgkQgs4hfOTm/CUX91zX5w1HslTpRiHQrUXl7IxzvsfFdHOk0RjysPg0Kj4PQ/GsFd
vJ+26M/1GC36ICJLrQ/NGvoHGgOjjUUy28/p65Wq44oKziN6WsUdNjONajiFhFI2YzSLa3wYd2/X
sMTmQhiOv1/XOy3RWs+YQ4aoks+Bfs7WvvexN3YocCKhJAbfgW56XOY5mejwtLbKPNZwH2Oh8hTE
Rr2GEzkkaQcH9+gdsgDvsk/mW/A1sNfqH/XtHQ/UubfwCfWlM8ynbIi56/ouPHKFeMSTa20XAbh6
Sdn0BZWckoDMkAvzO8UBI93B/nWnV3n46DGoiHH3iFPcYV+KUGVpGoD1fps/LwoQNeJ7sumMFBbz
9XFhnUWDpm6z9WfHbcPVQYgt/AikSD2Aip+k76mWLXzvUmonU8CE34j3z4D1NP7iGJjMiPoi/kYn
G1IskN1QbhoneuWzm9ePMciBo+IZKAFjtA1fGBUJfF/JwMjcaf3kcFmTS5AzAOIWl+QELZ0RK+z9
54b3SqwZshSb3ELRYhueP09ScmiAIbI5qyTdVPOEjhsT5Wza7csAGbxq2at9wdxemqFn9qs5b7A0
KSrAh/XWr5NL397LOXrTqbzPbS4aIqY15IJ5Kwq4UUsMc/hvbffzqtSMLLYSv6qk9iOX8X5hxrf6
0s6LK93EfKhH2vGsilQqgrhR7mC0sv+U0PLlQxLdfwR3WZ6pdKCx2uELPHlDXoRvZSwVgf0Ldgpl
QDN0AnpZb5t+eAf2Mfvxkee2Os7EEOcwIgXTlKEdBbFW0NK788ugZ+/3DFA4u50MlGXjT6RnbuiX
qxyuROTJExpJoSL6MRCDXDTyO+hqOo2wdjl08v501Xw4rQFqxFvyDsMGV37YN7MpJlTqawUXlsFh
gQ/yekPd9wTFnfYosT6piGD0MLFSSp+IEYgnZCKEujQ4EsS/l2yH/Rj9WQegqrSNx6uS3Sz5TqMJ
1r6N9Bww4m4C43JnPX5pf7yoNVeWIADzd+Xrc5DpC2AXRXYLqdOGEfirmSjwybtcNkDAfVq2yu7H
hX4EFEh1fyGk3d/KMf8u1EvsukJarpPXWAbtVUsSPB2cc8lQpUSCxJHOXJS8p63XvUEtNi3gyc+B
31ToSoGTU7SWf9uzrfQGIY0rvy2Nat3+Gj1uMBpRtVUxsK4PcRl0ygGNtkJjXXn6+DpfhTUwvcOO
tHLSSg7sVZlqPmb4yeWw5jhwiDng2ZTf/jjdL1uRyxJ69lBXAlWFp5Jd14YAaBFgNInaV6tMXg7Z
mt8nkHXaD9SPXUWTn8GrqzN1xx1f0GVOcmglPtly1lpYZYmSBqcaLoFaWjvN6K7wn5sgpx6pc9BZ
NbK0LFY605qD0YFrMAxeIBwetvXSlLa0YWQHacKWhmdrH4adnS2YNrEhj3uf5CSoYrX/2nOfa6dx
7jDi88Al6PQawbIAbWP1Tpdi5g5t6qUD3uVMc6snKYR+/0oAsLWcyKGMiMmHnYLz6ykjGTK9PRk/
R3iP0/tpme3tCZNw+m4bbArohTTPDXbd4F98zEMNhuJuEL3XXmtj0dKv5NOFru4Ws5MgirWXVyDq
c0wLOG/Q84fE/kuvB5E+QFU6DddLzRMDkPPK6DzzL0r2VWwKlfqinmArd0HLV+TiYqV+XHrbXT8f
LYpy/oLgmCWfP8r//mKGQqPiEOuFOxVtDoigyqwgxt819wzugT2oWhW4VqGLo6OcPbpTM1vuYZNs
PA07TzMYDfkoDB74kVi0LLCoP9mEMCevYyb2vhxoMSILsvrXKulmdR3ixpGmZ35oM483HgMiRJWB
CV4T9bg8Pv02f2muRlOt+eysOYvEcrh+CXQ0Ci6J9Qs5ou1YkJGcYP6VH/4mi3tNUDSPy2KElW7R
e3sg2rW0+BOSrKwaADMNij8ZbB6z5uuAcvAeGTIS0CmrQwQm26iQ+E434XEVcwBeuNSD0rTinE9n
cUTD+rN8z7xnhwKK48RaPONB2EmJnfiO6qZC9Ck5BAjeneVtu4Umj9QGJjjlPmA35aXVUxvcuHdf
zw088Vgn0JXuCf8JTpuY2wrDyjLa+uEDmGqiZAZvhfjrTN8KfTAvMvipSN/gJJcGn5g/m4A2tO7r
ErubiRFCQHex6xaXaWA5YIdzawhlRY1fHM4iQ9J4RJqygisMO9eAyFoDaRtfz4DMTdD25cTWs7pu
gLh/7E9tMhtCPXuQR1l8z65GFcwsRSFLmyLa6GoyiNIUOhKtMmw9pU+2NfkP4F5T7MCE51bZuMlC
O4TT5dmpE4AjHeBs+UBHBont6WzzWjv3h0UfV6PFY0v8P4XPfMmaQVW4qVIbTV0TQYOMiblEdODO
/Opf87X6VHvlR/ae+tYVBKnGh8yF/hp+ZHBYQdmRx9Opu7vKbcorZhxxF0+SEBg6jFRNlX5UENM0
iTO8qgOjjxJ6tGpPy3f0NmnXOXbSOeKLqB1gGiOT6BOofVcyRdqWoeso2J6sH3VR775kxrqRK7C9
x7GBjg+QHujQf99OcSmVTyuT/AK2NwAXR8EfvXwT9eKI/+XFAWplbbLpIhI5K/p0DooZ8jeCYLBf
+O52kNLyS2ZtEBBn8tmf56hrE9eSVRTzls8voF9Gr9L2vYZIRcuIjeEe5qlZak5UARnzK+oUPECy
JVymWmwZLy83L8pxpkqYkYN39DwFGAL2qLb+hT6qYuQYML8RDAa5ZsIs2nqaEgHNf6vHqJwSX26s
ckX6BptYaDEwKakqO/9dsVPt0qFhJE11HxqGCIalZVpE4XrFUlP/2F579BGWjd36Ly0TJmJaEv2P
NAuAaNyKbME/lJ4dVW3EBayiZwX1GFJXWhRzdQo4f07TXC3CkGXYbV1j13QamqrdzIUhPEbzuwvf
2E9PMQ86w8dw5UeyeSOULq+GBzjDyyscnFKjefE+LKS2liWcTmXv2aGbRhajBRyobEmYtNJRHNcx
CCKpBOUVE4IGEiSG+NQnm8diQt5KgMcqNaKwPbB76ftBWpWaQkJQ6qese1Mk0st+TPIyV3WzI48a
K5WvWR3ugf5rIPJiPIdsToqsv7D2LEO0v/2FNF07HabNCEetMyxlqwZgbM9bpY+CpdRE+3uw9lP0
9ZmeB0863+ZvV1TYbn/F/qNYabMc5wN0IPQjCE4D1uuBsCmQfSn9dE2GWlNjWHjINfdvBEGIoCMA
oVSE7b2vdwxnVPHweyTGUlJmf548nr+Wv3+tynhC7aePnNkAfnuNQR03alOn5622r7PM4bAdTgD8
pnvnn7fBB0hf6Dgy+wfDPicWZGDT0NMfM7vyro6o13DklpI5a/JvsERH2rqcBYJtlSrSHiv1YipW
Fz9NNvkpSkKtCWcPtF9xUjp18RzpsH/Az80UeaRqDGdNYKiHo1FAezkMa/0EHH7gH1+fUWCuDGHN
TMiiN6h/4X3emsQOwpypMA7AfCHKakpl8vRnIugLx7WsrUMO3XasgSumDNdNcba6R0YboYnswqtw
sL5mzPOmUOSuljzywwDxMfbfkALKqcJmBX+AUUJ5tjOyHPTsnoOuGz3vJlCNxixeRKtqFe3Htcd7
NdgVsIf3jn6w/6MNGadp0VGL2XH789CYYZ4P5r0Zv8oaTUY4vPmhDkduBNNb64EPubRUKtuRP8vV
GH3ohh8iu9EZOmNo5+sKwiFysYbIMdDZIjnQpNkCQw7W0EihuZrjN5fNveyUGkq44dkrKqBw9i4Y
8WNt4azlQXXThW29baeOwJxZCS8gkbSBiUU+UPT56mLZwS1uMOf+byaoFcvKoYSB8N7lbKkybXAP
Tj73hTi8YcsSoqdZZEs4z/MpLJskhJJp06oZcj/bYVzU9KkagTSn8Q5O+2jrNjxBAoyC4qIhe1Ay
Ywxnz95OiWMACc2+cHM52M0LQVrDxgI2W3Aucl4TVbpPe8AcHFlHvlEeks5dCjsJ7O09g/NGO6SF
QsnGNlp+9VCk7gi76ckjDIDab3JU1FKfDoesvMXS2fPdWN6bcMOMGrb3DKa3AVUtFpOzeLCNVHSE
c3aFW2gLxoxySoZT6RsvhkSa1P4h3EVcofsQuQxs+R5mb7uqtwWWwm8U+0tVYvRihiRcUwCTh6y6
euQ23RLvYL5s4VBGH+GZ+WDLLvU6X7XzaRNaVz2RY+TrXYhanmx77BgpBGWcAFVQzj57CqIHspX2
6q/TSW+xLmYUrRYLHmpBAdO4M310/891xQcq6Qnu0VOb3T0yrd6RmvdS2Wenik10ypRmQtjXiFjo
mrSu8FKJxDihlnwYgmGET97YWXDmEkBMj2vr6/P8kew/vaFS8HQEbpMA+mA6GHUaulHIUPZ1wUAz
4zTFW3Usv1DobkhrxCZwAW+lc8c7KlwdWSyz10F1K52BQ3haKHHzMrqss8Q/FLF2+TFqBb3PZAJ3
ZdMDGF8sTxUyHxCeTHYN8olPl+c0d1XlwAy9hMy2+mneVJUhIzrFh7nC4LzRKOJMnYGdMQ9Ut3JI
D38Ye7PK99cKjHOWVgGfU8Nq2zPDdedxhEeOvfOy83heH+GMppagVSh2Ve9GjeK4rHcZdnqSi1QB
U7hIjPLUKRWZo7R4fY3DNJ2FXBTPtflG9g3zrq+9sdSNrntWWSGaj7kXisktHns8tPPy1hQjMZHd
EQkeBMYOoe+nf1XCcDOWJT2RtfULzLg9H3HGNmcx1+cqxCeCbym7d0YvFElxfnR7S0wkuDiJrUEG
JT+mngCSKdLTF9lcJhhogGX2AtmQBNQ7HU7H6XWg+ooi5v8iOuPdmfPRFHXFgf42iwshKeB3CWJ2
WkdEeYBJjfPmQRMZ7BXApg2J/wFVQ5YAeMMe6O12XlO1oCKnWLvJ+d3tsSlf0D00l9LuhyhjTxY4
jSiMG1lgokRZ8YHqSxPEjCo5YnvjEYwem7UEYp5n9N1ki+O/gzSov+CK5kdWDcC8z42d/v9NKCsI
du4XNDJ/Hb1gnNMq9K1AXJ2EI5E58VLD6u/S9gFxjUlyMS73zwidQESPlFchvAmm3oe4XGKE1sqe
uFJXTZYCWP9MV7AuqPeFZKsretohK4f+Bb2vRokXwUwIZdMHNHv1t1vKKtH+webpKXr5RT4iVh5b
X0T7FykelF5XdxlUokqs52RqaDA5+SNwJrTqWATwqF6EFnttqqc0f/Bfi4/mo0US3h8iz7ZiV3sG
DeAeMoO9uUCrJHq+3SmAJdAyQsCu9yVrtCYM6muNnuZ4SD99FDJ2+nBAyNwPpGahddxO9Py2u1JH
Wcih9yrYdKOEEUW1hjI43mVgoQCAREOUCoGXZEYw6+TPpATcwmKPW4b7PrhRG2lsj3Ci/3pNWa92
4/+x2tOUXCI1ziNIP4yY07scebTph5jInssRgWptjLNkgzHctkHcIuSggvoTE1AqoPDEBPS3xAqr
miG6Gqrmi+8oejRqJyFMTfba31P5rOr5l3lXTckv7RxaX6ixm1KpZHscIlfC6B33tFE/LymUD/KK
d0C7MA/AExjM/DmgPo9wdHK1vcbR62Na1isHq8fJ+3wf17tgknUgLLTxLCp39Su/n+DWstOGYNDH
nAVpuex1Hh0wPVsRnToobMv/0T8D86v040xrySIxq0nlmKTBgwnCBW388eU4tsnc00C31zQRPW3L
hx5wBrJqEbb7GbPT84+34TOywKvqv8mvQ2V3dN7UJq1X6Sl0fO/5cQmpmKW+qeOp4pdQpBLoI6lb
3uwa/JEYdSz4mmxhSu467OQYwh201sMjpVZjer6W5XWldzM3UUZJ/Rb4NmPOS4QcOw3k8KFtD8nE
KdQbRSB/VXtQVGM8ktHZw/srhugjCRP3wzpk71IfBlYh9lJ6VHeOLrz6oUgxyS/oJOEyR2R9F1DB
4sf4GHbS2+2TT4AKqsFcwOyDWW/3/2ZGnT8GK2sUzFy8HIB8JaRocNLiMukNz3EU7eIKgHu8LCeD
qI/HcQ2tTo/29l1Oio3CS3hXqMsfHXuByYTipYCgf/dz+Dw22nt0fy5+YzyXz2IJTIN5BFN2TIFG
w0QhYf+tZHu6sXe2gAQejRBhPy2xBT4wZcONd91RZaIJChX4C+POvImTSOl9m6tokty3PrSxc+fA
4SFGEwfapKLCkoN5k/TJmlh3am9JY/hEAT4fjlG5upNzeR/QYTbkKsA0hLXB2Luwzvibdd8K01Hs
kNuqDEC80byvzDtAoRWb/MTU4HQKjlQiCIqwA0wzBoEgOF+rGgQeMZadSD9fhB/U1blHOrsHWgAb
4W03XG8VtRLi17R88nj4HBg1gweTW1tR+Nofa4K2TSGRDFdelLkOyAH8uSc39rSf+P7ilTlaNJM8
bCvgEy1M7stKxhGVl07azdhgPK7+cBLOQfkF8cI//m4P17xXQrCinisUlecGZPDPb65Id+aqy8gK
IkRrc7nkNvvO2hlCRu4T2N7ePWszUmDSjeX9YWQruhzTT12IkAZk2BZxLPjGTFOvjLR+5FSMCf7s
mcms8wlEYuWNGgniv00a4A1XyyevepjK0ONtfdpVC6fQMnj+q/H24RNFaY9t3iiSddpgV1NFgQf1
QDYy1DN4o+ICzPnRPWksfXO6mQEwLaNVOiNy9Xvd5QarJgqHrZy0TNT7YCuiT/hIosLhQmQ7jhrB
4CIp78FxLYxJW8gU/WVxh9hwua3FT+rMWCiAeSGg21ayRbTxY18dFAcBAAerD2zoOYI67LDohWKl
sv4Te/RCkLWxaIB3hrMWHCCLx6wuijSkU+6JKVyYVxzIrZ/0cUhodk2fX9p7HwjBVhZPLktELXCM
tnLJTQsvvvxVgWVM/3yL+1WhbkQKsmuzrT/6jN3bHES3KHO2J/D3Nl3C74l8+svWN6axoW7VU4gc
QzPqJg/frGSENZn8cHECgTaIB4xCUGPShmKiYfEwxwzRURsPx9aSTdmCJf6QqluoqquZgCy9ciwV
xHSF/7wiz96ZtUoZzaFMx76lKTVvwPJ0hMqPd3AqdHPdsInodDvuFyN6fa/O+S4SnWXzac3mXsMB
//v0K8pnsVbryj+c4PjBxvDu2Gok92eeW9SsCKdeCx395JhgCbFQ2/r3cgNU87o+Q67B50l9HIMi
XXOxDiEFirWB2hoArvh6kiajCJ4Wt6Nb3LYt1yyHli5ncAkJzuKGIBmY3xQaV6asKc9yLfFOetiH
1Kjz3bjDT5T4ucbA5DJWXCFNPi7Ue5uZIRdzH6fFl82sG0Igpgo8nMVAETpqyZ+2Lm0+D/pCC6aR
XDba0wbX7HL3RFW0pmQ79i5OwD/Tzkjrn5HbS/HZe3acYuDe8ZOdfn+0w+sO9/psLMF7lxhutcaG
EiREXDZora73QTUoErOejLFYhRj9xtEf5IXI5Y7/pxFkaDb07nlGkdUC6kNKHZsG/gzZuCmm+52l
xm2CD73IK0NN0PwhgjFTd2akwS19ecz4oYz+Jf03Vlye9dejZOCr5dcHgpY3gtcCUKyUFUUKbJ4z
V0zsJsoQyvTiqXPGJfZL2sKbLPH8cQmTJsQZU8sqTitkReG6uU5TefpUolkg9JW3xhUBleaRKdIY
q8MWrpnn/4Qc6ER/KpuEe2alzohasOonY/CNoBmL9wXnTceYsJIeixEmpzvrF4PE1GsMMljkWxDD
LuwwmlEjZa0CS+IzoFxZkOcFnAyQd/HIKzkP7KTlzExeeNRbzM5r7abScguF7aChlgaqSUmYw8Bu
Vm3d8V2RKooC6zOndIqs6dOEFmiuMUY/zTv8HGSn8ebtC2MvXqNp+kTO98wiLr0nnGqYlZ5BcKff
LbR/zyLpn6zZHkDOpli/inGONAy0hBXCs3xT6ihD4LMoxmcMFfLum7xYtvc79KPIH8qcHilTx8/0
7QhsBojd/jQpCIhIAShRDa1je2Sjm83GEemQ46UbdaNMxOAj8x+TEx5n6sAbCcnLqVOBh/w7jaXs
Nm6iD1j7/sdTY8Tv6MvA8GuZBBiJBwSbxcoXY49NrZhbNnZcyi49aFsiurKHYe3xMvz6zmbt29xA
lYQhOYh+5316IH45loQ4+jge2dHR0Gk7hTMkrN8CtmXHv0kOtVHP+fiSsMqoRp4RuXJsZwNf0zlB
J2W4cIt6zyxWYkMvqPHVsvPFIU0p1q2NbLiMoU3DzOVxxFmVR1T8FPy2+gKUsDuqv0j0M2aPYHcW
ls+oTQRaK7v9FM8Ym44G+rNh91jvXyCZVIZl1+RNcYLct1BV0fAw2y6GWepaErPNMj8fRGsrYTTV
23SWBAri+ZlDvI7JsPpXcQj5j1vWVxblJ8GfigRsq3KJuF4+m/UAgumDIxALSNR7+veFMFd/R/Vf
O/5lUS+P4jMaQ4FkAmZgOwwBlR3nLRgtOoIdHTkqQ61zAcOrhbWD9fWsYquHmgOW9haooxktTDlK
Xi3OPv5AgiQSfUobCwFoZa+WmkgwcgE0dNDr3+ZOPFeHNZMmGBp7AZx7a1nG9etCXwKJfo07Pnli
76li36xzK05h//cVjMaqKMKKU2HpeWEOc+H0AQSaPcsV2tks7DuXd7AUo+fSA9tDFzdHxAJdJH99
Vpdegv5KV/7V4OqUwgHZMdzIJuGm9ilC8kYvY23A1QrSjdaFv6kGgnffYJWlgkc71WRc3ao/fHfo
wlsH5tGjj03Py3WdPiUlkMxmF0FFeQJAhg+Vme9N3ffau57lwJ4Ndk+ep2pusgWoQBXDO7pjVyFC
EjM1DQKKijPGFh2BuH62K3iUa9CIhubxh72PRmDKfBCloDAg41l4ZRbZFvvHw3/TnFBVIKJWl4wx
3TLEs2ZK0uhlZa16j/AFtt/prRU53Xj0tCbdlfmoMnDBvP+S4tMc8Tu+L+Zd80IRhWfMpekzzTO4
el2DGmuxxMILrsTHn3vT1uJphkK7WqkG3VTjyFBGTD4DoZan8KCRBPlIX3rYULuzCCtZhVLmnkY2
6YvfuZ7RhQYbENjPrqXRHaWtKMxPpDIGFQHTNM0+IWcYZXeUVIptBOepvuhpmOERVvHt96jAa5vw
VkQ4cfOZ14IWQTdSV5irF5AV7W8UbzPioFNh8yevKunJKLZcVWs0Wx76vfmPPT/k4TM+23i1isTV
I+iD0bMGa3k9tuckXTNpHASkprL8dy6yMhS9Cu1itTyupkluYY1bQLSbtnCrY2eV4TOiRMfhOVez
vom2CDYnSHT+jQewNpj/ZgAsYz+Q9NM5o+cqncnRY3jfS9OtVIQXlgDiQQb+oPzaqVxqRwcDPdw+
Pw92N60SvkHQSO5DVQ4hjawTcIRjmbp/DfXCuQzhceot4yW6M44/QNB74rfUmDTtZFf8RQ8lNi6i
Kw4CKgfJAOt6mpvPPH6/h33syOiyw5lJ/OdLDERITfGUhtyTGHKf2maIP90h9y3jz3dWZy8tR9CD
Fotv5uzLR5nQqtwrMj8VGu7RcgbNvf7ycWVVwBSHye7giMm31NGld13RCtQAdlixKnmlq4iBN43z
thK6WUe8nXUgw3TDwfb58L7R6ei05XtFjL6wllItuwM0458gqWM0XLWNaS36LOYVslkxZDj+LUhq
IoDnZMW2C1o0bhWMdlIipAPyRu98fLexYhGP0kLAtKOd94wPB4tllJOBNlrbcsqCKVLfcnupjLtT
btoedqhDYiJae0wVupyLV2vCpWF1hZkaqk/WtzG39ph04jbPO5cQKEEuf8MCnDIGPGp86wOgy0N3
vB2sXxZQ77B1oa2qARAcW9Qhx0Ktp33D7k0RWmbXK2RASkM/jlRdYm7E4lPmxbRgkZgBUCYsy/X1
uYr9mR8tQZfq98Qthqt4nrLiuMLi1G2CzX0ohKXaH4GXeJ77l92hzRHMkcu/asUcGyigyaC1xwAf
0/RX/vNatXfGM0l6ZuWhkzI0YiB5GQA8ySgNHMHAhC336ROoF5c/9/tIox4dJlPGE7vX3JloQXL3
8Z3EPzRfYxxILkCUH1Y11YNBuutqftqUXZUf3Omrm6TutjBObLlWAa9KQXFl4nbMbjxGybULaOQR
s1D7fJW0ANGit68XM8uZxwMauBlZDtucx4Om7PWzM/Z+Mqsht6fnGSdr//D7ID4RwGFyK4g3tPUm
2wn6gSlS6rrJ9TrxEjLa38sjW8xWeO6ZxPzIuVRO9Is60FiO0Wd+kbcVsThcT6OpFlCaZwlvZBPa
bvsfQV2zY4lfSkecW9M6xpzCGJPl4SmrVot9DcqQCINj4j5iyQGEPKeGLAfJynfdQBeDtUdtsvoH
h68e+0md5R5EapTf4in74e5dP+gyhqno761NJz1X/ztr9jct4Bd/oknM+q62rpMzezNlu4c+xuBC
dqORZfUxjCVPjOgL0Pww0WtDluNhyJDLKFqIGqPj+PXmjYygFHCXqEuO/iOKT+dFw1Bwet2Cfctw
8/XMK0A7TS4BYk+F9jljQkr+0CVdRARe8PrvJ8VfdYxMxp+8NjzE10yxsQewsfzgOY/1OQ9hR4m4
1QYHQsd3FWj0XMNgPK7yXym5svxgtpWowSfSQu7wt416GZjQJAJbINSy1RfNwRhDP0C/Qp8kMv9B
m5aP2EtuTie3p0iQReDY+4fu+/XnkJ/diW32Y0m/IFfiHH92Zd7Ao6Rnn2Xm9bBrKH9apT3XGdD6
t7r8H9zge7TF7TugfFf82mnlowMKG5uhya9OMx12TbuzlbcLIEyt19TgseJDyeSga6TPuZa79nkm
G+t4TopEAtPySZ6I3maieVqhW3WYgu99+9mqeoo48potkwGDEHHo0aY1U187oP78MNEmEfqk/cRT
zXrDt4X4zOFsMzoEpPmSdHB6WQz+ku3J8MWBWFT0wHKNlMFMBnlav1Co9PUGeynE/zpWyVt/hXz4
+ikkbCPEz8fjKscqM63wGnQrxqZ0P75RC1VcTrywOIC/35Et2GHiRLmcS/zcwTEEINzFtt31ct3i
tI0b0+lcu/6EGpkv5XkNlPTaS7urbtiYbxGEwSi/u4coNkD9jt8eua7yDh49ci+n8UD4kVAXSOdv
avERI9CCUk8qDtcXn7kSrRA0P/Jwnsvv9NAikppuTi27fV2ueEfEwssXwi3YIKYIfkCbmC4kcyuf
mwAGhAcsSozwiYidhncXSK72ds+rERUuU/Hmf2kJ8xYim2v/wEKrvIPWj/Ci5QmrzQW7+m5MkIYV
0NPRwwaiAmWKjspTXkDf5z4GYS79ekCcsxq6/R4XnE2pShjxWaPElAsMM/XX7zOIaty/wnH82zWB
yEKhoGrBuX1wYgSV9O3o/mOefcZGOw7Dqz+Dz2SNhl4u+3Pd2GffyN/OyWtx/bG7LOVOQm6vFNrQ
YVp7clGOgh6DAEWqrae9brxMg5c7/6HazRLlgWDaRnFx3P4O2erHiMI9aWtaEfgy+4+2FnDS9/VD
eKQGECASd2Ozm1L51RIxDPujFfzyuxajaz81Gq1RuY3DBkiFy0vu4Ep5ddj9CWOSEJcVAKZype45
POh4D5OE16yigsExyeRZfckDd4+ieajuV/EzvH7XGPbswNm9AadGuUa67wTFhRX6wj84Exekd5ya
IiAEGt2BFYX5aGi1oTRLes7Wxw3rfot/Y2d44czkyeTUlAhGUJW4j+fKhyJtKwmF+PVLxSU3Hig8
r6xelieTuG/QGOmRYQVez0BH2aj8ZiUgE+9CKI65qBfPg9tDnup8ZALCcxZ7BA7nnGCGKJA1pWCA
WpKmVfU5b7TmPsNB1ySHxSCopo83p591S4PsuTxoML8q9oJugcAiHQ3VMf9MeCQNRVTKv8IgxyMt
AeXKE4hYsQ3KtV4CFwXZQwEZnvHMW7vQimUO8TiTc8nJ6/Hzikcs/TkUE0Et/TeX7dHoAfSiFT7j
6K4HlUARQvw1JO8vUf3kM8pPxLYq9FWxXKd/kU8TFHpuSnqVqlyLk0LQJfsT6lw+ZzawugAs33CI
SKBZth6enC2fFLQmz4PnJg/hfcUw0hcK6AFnUYIkvR6HtYjXzVbzfVYPL/7/8z8zbRlcXm2Ki3gm
pqUUDDySMddwXs0qyAAg/vnXqwHx9xbX1BOmL/neve/ArY8dcJpFQe9woCwUVhCfUmsgPSOWIGQS
RPN4PQfWUoDZsd2aLQA2hGhWG1WX22VykMoB0CwgrrpjaAvsxrsIN3OrR/6PsbeMSo8qnn3bYmz3
yhccs/uMAkP6n865hA2+9pBsA44Gix+xwToFI5vDGgi+XaAx/tKXNq7g+eiRpyoL2dHLYT0eQznq
ieTcJHOl3505RNl0iy2FaD2tCQroxaJaDeGffgSsQyyJt6BvPXCWqJzAn61kgbKuCQdBMKgxoWcB
/JVf9c1vrnmE64ESo6bnKrPGbqj3QH6vC/KRM6UWFweC5zGuV5ivzXBuH+Pzdtypx6Iuxfl4+1lm
UtHbLvj4o4lM5uKfVxA4vS7KEd3NJ/NcSrgijYMweI/SXhIyugPCcmm5P03wsmvGitx5tUDCvM/F
D6qVuQ9h/qmap9qcqnLNqVMibJAllaCzearKES25xg14iB1VTPUmi+kbPJqOKEZCvd8uGDJntBC6
lwK/WH9y8np25L/jO3YBsas2j4bYqKHY86csQjCJBWKuToOxeydwDIS4Kt+zgXrGuSIqQw2XHfuo
+yg1AstfOdI85b+I8T6z2ZKxS7HxPIexj8SjtngxRXTmAw0pFC15esrmboZh8nWKbrUp0ArSnydw
Lr8u0bHd61zunVQX0rrVd2om1Os3zJXvvZrb3gYF8zcD3lT70CgsXnkxSQVd51TeVXbrcwpt3EVY
MWoJcp7IJjGYDqgzR+CA18GYWPZxVTlA+q0K0OybVnHE+cu0qplmo7quZZOQCRuiu/DmDLjx71Eu
cBzhZrvv0RXkRYntt8wCyMxCFxbM4W+++o3UQqRxtMhQeduE1adNFRi1QTqZQCsAEZy+bgAnWNWN
mClwwF2dCDGmoSSab/8qPsGhK7bQaqIORwk2vjE0GlVnAqATXeIM47uYC2tLDd9wHjQ5iXPPv4ZR
qtvp4gYuvuTQ0LvLSlFZdwzFlxm7nI8wc4iBRdWCFjo7YzFtU7/k+MRIqxn3TYXLgIZkJvT991xU
mZS3SiECkRqym21+6ZcagXFLqefbgms75NOfjItiVdBl/ExFSUtNk8svACTP6wlKe0sFsf49CG8D
xOQ4d54ktguvOXxqsDyHrxKv28OLvJSa1+FL/kvHpVQJqGFWMD40tmcG2LkXUNklsJIKZeYLKkN8
XrlHXHxcj/RUv5Sg0hDf//8zkigTWzcecdiv9G+v5j9odKL1Dozr92vF42Qq/Kf47995UjBiteNP
AQtGX9YpZfyS5nLuvBUx+GFs9Kg065ipBVZvXq1x48P8TA+hiM42ppmDTpjhEMquROn+X2xQPu69
GvVWKyt5km0/qDtkpYJDOkrUthDTWplOP8kbFNS/vuwjjoAOh67tUKGfHvHrBzZdutKCHnRZAQlr
AQnKfP33b8255hOsi3YOLaHgCVBzuJOHPr9c6uYmW9aroNGeVQ8goRPRAPeGOQ0/QhUJhtEZTyGo
ezLWOKAq17F39/gUFE+it922Y9qEl1db5xASoNACxeatvohbJd/IQaq3rcxCRixG2+HY6AaLB1+2
k7eRBqFOeX3Vgw8Tg0wsrUXdd+/2vv/q1vMBdoysbbfeut03Sh6bZvxq7q/TVqD4/oiYAmD8CKX+
HQ2ZcuBQNcwPHV1bzef4Xlbs9bCmstwo8rn4c6sMrp+XvmgKNgxeMx4jRpN+s2a22Tf6XUFUvTB0
/9nI6gDcJy8tTufAjOVPKWuu15U3LpxUKAHiN6jIqtxx/MT646b7CXuMMjJZ28gPTS5chHunQVr6
2lfIAtjGcBTTxP40FXUtHLGcP/8rwA74ZyNoD2vlEQ8yOamw+peuyc52eHA3gJ31qKmquQGN2ys0
EHLzTv4j+Mev3nK1aPLC1ftfk3XC4ZMrEz/BLtoLywqIceT/e3IcKzn7GHs2tU1S/hU9yzzjsbDf
zuyF/hm5q/huUVgUlRuFip1+fmE41mX3u+e2jVZAH0tmSJngxF77jFDYsbPOY9kOBIURKL4HyeFn
PSJmK+xfUH5KSvruFIsZDtTw+3e3Q9fVQBo0KmsJxIwzF4FhB8sqtMAQul5URbzdU06fULo08xNk
OE4YgEu1cyzxX28R/gaWFx/om4YnDSQLk9gF7yAf1Ipz3UPZZDSftF1TO/DzECm765t0i7NeHGEG
EDp6S5gtuAuFo8ufF9VL1l6glR7WVxgp2sR0qm1RTsjLqOXKlbjNk1ghdX218yBp0Y2SqbVrlC6w
evHC1rfjH98SLjPbSJHkmgS+DqOUElz9icBfm+rAw9W9YDHYNPMIEsKm+7qgQ1Xn4xrfR+yID4HZ
rX6Yh75KGX/aAhwZP8t1O1Un3I224NGe2f3Rz/i+FSVmT/KIMNEd/Hnx8b639M1fS8M/QwLQrmTB
qR9W60HYV2bcr5lLIRDzlbfOmiZ8oHOLhCA6H8uwxZbp+C5YsI67Mo2CFVnqPFle5xRZ0+YO5yu0
rev6Oki3eHPI4zo5JdkHPF7vCTtZy4Vd0CyRi9c4Lo2ErbVXdrH09fDP93FyO14cSdc8dUMucevy
jG7hFOgcRPg6TjFupNPU0+tByRqEmzzbNMSj8uv8NueI9JhMcdJDRLKev2XjGliuC5nQbnB8wMvy
S4I8W9qMc2Xwva757HgDOLRFSm3XwUT2K2MwFoKNJiGu9mLMAcwdMt2ISy2EtJxKFeLiL0VqB0N9
HYnNZAorXOH8Y5PLM0Di8zAi6ItYCcuk/Nf8M5cPTq9AcnxORmA0vThg/GuD6s4IQssFt60lVEKq
XXpdmbvBK3BtbQJuDSjkSrrvqGnWVuHRLZ+WsFiYwlvDNmj4jDy461s2oc/gOOL4LRVvogpqm977
/C12ccxZD8UVEw2M2yxnDSvXVQb5rrpnBEeUg1OsD+dihL/r4bfyKE9Jw08tYdhwS5EbVBQhAmFN
df5q24am8cGOx5vA0s9HA5MuTVn07zGVs5vNVgEc0JeEz+KgOT0NW5dpo7NbnN/jGT4+W4xyQuBb
70JwsJfJSpXtJz+n5Q4I0072Ab6/kCeixegjhtjWF0nZ1VPBghNc79hQmGmoJsakgT0jxLEFfJxE
Mh9cDnFx+Ar998mtXXtQfWTnh79KtryHKp3CGKAPh5sjt7g0AW8HyGROrB9ysQbwgkgRakNBtO7N
+OTCuHGGHjmi56wB6WkFtXo4M1DjZOXlK7u088jnRKI7sn1vt5h4EIzh8MBi9DIGTaFCvcS+o9fd
0p496GG0dUcsCwWPuRE7V8EeAJxS5SWZS/K/+jFA/fhEWSA4i60v4ILZzp/+i9yH4J6/zwacumCl
pPSlP2dlV0BR+v0uK9w4xZBYJVQl2ZW8I5ekm/ERk1xInJFd1oKoPXrIJHnRcpzdSlpJ/MVy+DtL
BW+AHIviltkh6Xka06tzfKCHfEJhoQ5ZcFYR4AF+0o/hIgiA11oNHNuFMyUhLdkxEzHvZZ6fvc5Q
ZL0jBdjM0BOZEA/4GjWHZsX8xuvRggYIu3c2QO9x56vvI6gcfqsDEjnjLxVFKyk24IcbnqLW9/Wg
QRLlhNSotz6QfkXMBjb4Jpob4toTx+5XwZS+E1vZEVdnRbU/0YjuS2wGxNvdOTXKCqcJr+Mcoi7I
lu7apkBLUPwbIUIooOKf9Ed8Q0htAWfRcZ8BHIwGo/cZQ3vp1eMdyk2YdbOBcQdoX5rQq1wE2UV+
2izN4dmBHZ80Rqbw3+PGQeRC4HEWg89kqQWVaqNanDDkx0rZD2pWO2DpXzfSeaWfxXpbt+GFUPB5
38yKD5P72Skk6UBTtFUDTzGHGG/skM1yU7lFkgL5R2siwEJxz4PGEbUsU3AAWXbkea6hk3eunoTE
tKZxIFGXU3YGecTw+4sYpkTh47xqLKJjJqpuRhjItAbO1/3unhGx7ILKWL8uVIq/1akVbWne9qin
BRs8LHvPCeW4JitBsRX5KQ72KWKV3L0ujV443zoHNKp96oyeNis+4ZYeQVLoBlBfq0hxTPTSk3WO
1+6h7edOdtOiGmuyc/aMo6jQgo1v9BLux8IPJvVtpfTof7afL0PD9gHgDPZmZQIPNmsQrccmoa1c
ICbT+MmSGhC4vJ8xY+zguSsx1KE42UVaZzdAaKQbZ2Z5YFYptukFF6Dsnz+YWJ2liDOCvx9NBuQh
VA/38fkdcl4Y1yLzLIZmvqc11EnQh1a48NrO6JhYLSzBxjyeVsKQFEUPS1p74bAgVHY3HHZf19AS
LakTCN0VF9UOIOaqLAJ8C2OQgR2PDz75MCOCAVr4ZuSxQGMUMuexM/qvlf4+fiN/5VvFfjaO/4lC
kTcDkmxYEbz64uydQaDAEbmDlkJg0hrp7EyssutmI8Uq2VSKrHQ2YwLeH4rZCsADWi7qwOTDFVcX
wfpXl+oQYKaDqJxX2d6/CnwI3jF+1I5yF7wHwACJ5HwQfthqW0n8NSkpH5ojB8KwWQEEXF/IeqVB
Nf1EeVZbivAtQQyrO/MhEK6NzO6wTcFFTRqGe/rQp4BTO6ix7QQXWnKpgsIQdElI8AY+WkCYRqsF
gKC33NuvChTySutEsRknHG/XUAmllMsg2Of5NnQxmHHhNU/vlxCFe78LLscZdu//1ISmLEoxOQNb
yV6g2feVlvLjHjfTkyk7+kuNYHmNtpTmH61v10wARrcBmVHwOQyHM152nmGbH9zU01aTSBANL0q3
z3xXcyPG54E96GyPZ5Kk0spNwOYDr1m5PK0zux+2NlZ0pirkZqDhEj49QPs2QLIvi9s8r8IHeKBX
ani5xhM4vKwYD/WsPNRckULbTTIAgmLSPNnvyfgFfBXDnu+a8R58LZlKBGjlAnWUWmqhT8XGGynv
umbwK/M8unD5A3FgWEIymN6mipJCGBYByD/YKeSSb4q5cPjL71NjoFiuIyuo3szsYKUFbUnBdbpX
H6er+sc7dGIrcyL0CNF6Kvzw2H9G3FAtVaZY93wq/7WTwJR7Yj9U7bgzYx06EI2Cccw4QIPIRoRt
+fiFQzuSAg/BXKlxdXQn/9u2lCxasjGbeJUOBe0pQFt0ok6SzBExPF1/a3eT18PQeisnYNjfQY/4
H4p7dt4ovFo1ugfw7sRrg9m8eqs7oOWuIjgjcXC0zEGUDyjgluBdlv2VyRiJqEbyiNDJQM1maAri
FQGUaYrCqt2DHgrOnc6RSE/vwF5uWpxmMRa4bo9TfIc3P7ETbtWIdBlEJI9uBG9kquKZ4g9Mkq7G
SI0vrdFF3mK2+GNroVfvFIXXuGWVLof1Q1W7pncfqWNQq+0dNCXOJS4wp93z5aXZfbkQP0XDJ47L
lyhDhSjcUrB/wY1pRmidsPtt9IOqX26eVPlikF6wJeGjDQPTiWQJ7m1n3RYN73n2Ps5tFWn+x6GQ
xGwxgd0t93sm6WcOv9dx9oDxIRUpeWTPlJGKPpdbdT7Hf2OBJuJA3xLmRq9vJqfwSYIpVlr6xilm
gs/NLwq8PUdaDexFLsMln0Kzdh59B/PE9Jg+6PKpDGG6a1y6iD9fkH+hqGPzL/cQSKWoJFHDSC43
HvOxZza4gQLKIctSuz4RB72+JnnqfaMaEE/ljKjR8tFcKFLWcI9LfC0LshlAaCA9NKqSSoCzhBqI
3P6mYJXvclCqd3TltU3xDgrKdhEWxZHOM8MvTLbllSpOZPe26apGBnCnJfK8zcO/VcCilZmRcMoq
v2iZHJr7He9uYQtcsydVHo0aWdSdvDrmoNmB+yHXqNGUZbqgyKD6TABMqBOO/VHxM+uvKILFp4IX
6I7rpEGyWmCOh+nyqzsJBA+r1TREdg/ApAxmKYgfwcf4S/xpniERMjH5cLPhOz3XI0Lj7oOQGYvY
zTX30Qmy52giekNyFBqLPq13rhXdWAO1pG8wXSpH+EhY9vKVEBWKFbrCnxbbi7xlI3zwKNptj2w4
7bVxXeet2xoRTg09mpUUN42Ka/T24756gAE+jJDTqi7nFqfaMokYuCC8Ab4PyGkW3fRt3oczXYzD
hIp4KT3klQPmFADNOBFgqgm/CP8dQsAoHoHFIBHpB5vKrZnTTLlk6cGSz9I/9Vf6maPufCVdpRkJ
2mgAYAG7VMlKsfAWw5Z4fv48C3TMc+FPdspmiSXZVwUeY77YDiCaKOcGZBGiNrEJPPSBLJB3DEs+
TrG21/b/UbfyW2En+ohcaYUyrmdjqVATkmT7QQHKbjSHY0WfXFmQSi47EPNp4yfw25SR0G4WdeON
93ZHH0KHD+D1m9iZ/uyjUAInZp7UFTwKnH6I/5tqOsgM66ZN6Q9PuMJnB4ObmOQaCT9wKi+H7cV0
79EakSAPbFmklm9YoQMRB01NiaJgjnvILeK9k8hIon03cMV92gXv1DLpvbHLyL89E0tVYR89zrMC
4GVfEa96S6bf79xGf3XZV0X8pDsfIJirdonyQonVV8E1P3FJ6gcnkT8c+vK7y66oPGUlKhWLAVQY
UPE95SwTAQbgA2NMqNG1OZ9XoTp9EamfujjqmNvZOLWElLGoPRQDdyQgiR/5eItYH+S080+He04V
ejL+nXnebTUNTutSNDkO8FNWNnJNyu/TlOPWaQeyRoAKBarHxEOHoX/nf+z/O6XvYDZtXmVNX18K
iTZGy4bheGP28rMO+GyOJn0rzyLs4FRSHJz03usW0OlxOls3GO0ksuDu8SpP1MlxPGdipf9SZk6F
Z6W8fuRzwpOMVikSWpwxS67JYThqP8AP/eXuxOvjTHyVC7VOtfKWTlyMm9u3QTm5FldoiE9OV6BH
UFT0PkZ8w4Thsp02MdY6prwFH+8wZnfNurAVaOMwd/jl5kxkLL4KVBGR4ke9eQ6Wqd8SHvTIfK7h
c9yGw01lEkOgO4oXrMfxIhlAqubgwyb4+0UxKwCeVTKNv5VdIH/0q0lqaKw4fmbsnqtGTAAQCozB
CVj9PQcMXFJ2mfgdlTYn22lungUdGr0vX0JGha1GNe9/CSuw3oxkPgVhk5JH+dabja4hkMrkgqqD
tpv78RolsTSSAA2R6bwebl0Lx+j7R11/DbDZknspSSjtrU/5T+2Ain+U2gO3slmdUfFl3lq8uf5i
HBiVi8/RkURQJKIONwo6ozIC/sTNS4CO0zAmXwF7e0JOPolejgGaoHUxj3h5cbGIW2yeVXSb9Kw+
03XmJVLZVFHODhFNmyHX1dRfthFZUG4xr9/UwzXiU+ztO8i83XNzvjFFlhDhNlQFJCpYkeYkv9Xz
9fMDrU30PKInYwnhcWOWx7xOQNPNAdj0fZmFz7pC3Z6KmPU1kqVP518RYMtxqTcddsZooJMBUfPQ
NGeRBNuG65qcnNfBz6aRncZtSBv3LFErRdqCTzEg6hJ+gnR91WjSWdyqqE2HGLPHS7MiiEMMT2Vq
0vC3GxeF8UivLBwI3s11Vlq36TnG/qJzLXQSZOH80Ej6mbXyN3Gl25mPUiSLr2nt5JMccllh9P1L
c0rbgW4HhccLYb/xwMVnmlZSwCIv2JzluX/j9l38hkndmJEBFLloJ+0T32hbPG6j/VbUsgc1qlTh
dLem6LkmbCGdM67t/fTsp6nGBJU6XS4SAovNapbqQGnaBPhPWnJsleAbP4uWV9626DRFqH4g4x/N
0whRMjXfsBkR6x0mMlEUGnrRJxwdIAGKL8HM05LJcAB0IUNEgfOKeQl5d0vC4HpbeKpS5GN6L3c7
DOA0wg1qdKyscyJEfUv0WGxgwMuR78RaVY+o6HgjYfZOmCnrjii2HYjFFYmsZhew/HO6XUP13Axd
vf6CSCaLP7ytkJdgM3rKuWAyzqXZtdm8Xh6nDsy3kK2ISzF+g/0Su/m3H3dJfdZU2WWWwRTx4p9i
Q44v/KsG/gBKXHhCxwKZnH4/x/YeG5TrAj+Jl2sM4XbVrlngS2TYs9D3X4Ctdlg1z54mJluSbiA3
xfmMiRv6eWFe1CIfld3RqMFyNwllmbumuploHbHnd+EdYXymAWfxQTxFwFNORR748BeM+WlDdINf
w/SaIhmHy8yJMXjcUqxVjSs0ZNkob4tgYLNLej8fClRxXct2uBgh6EASEOvHarjmJvtje6FK1RWe
4D8Q9Vpz33drnu7V/8OloDauNOhO6pKUhBKoYcdH402d8e98TObuIQu2rrdBIe9SdLwPFGv0NNMK
4W/Nl5bLJ/rFnVgIcyCD6dkBB7mcf9XshoE3cJUB5FtLIkyM/Jse27rbz33MQsbPWLB+cc8vd9IA
fbkHkIHIzJBAm+LkE7+OUUl9H61AXf5tFO+ohGchi/jxPGDLOZrZAjwfV7zaK8oox7f46/NypDXV
neNTL7ZhB0JHAk+zfZ+YXghF16S6SCT1t3YYW8tRBERhbMJ/QSgR6J406a3NKhLBGsp1fT+jgfIp
5UCf54Iz/6GpJ+72lVms5CkItvB7slJvYmI6kEPB0MSjSy1eBJEE9EpuMYF1RstX/4Q/N+iRyWrw
8IWMoJX8gx00lNmt8A3SB0VzkxTqYV1pTbFMmdV9jBSgzleuBA1huCX0h7lF7Fx70Xv+5SMNz4Pv
/Rg77nMhS0kSPTKM+iFr7W+x+mK8iJCwjhIAQMsNqnIyh79Aw4neFDwwA/5I6PoluM0m90lu+4Ss
oLNxiC7TVRzfJqPZFRezspNsplpJ4sEK+ejgfiNza6CzpCWufbJrEvef4xQonICJTpPzoU83hUyj
/dAOQtBtl6l/ta6buvId5nKXG/joFk1udWskExtzfL+Ox6ZUczh3k415cvAhjjdfvDtrLH1TeWzV
r2FUw6Sx+3LmRNFP8l+zEz9fc/3ZYTOrjfBKbWOuNEjPtltJKbt1Ty3HWta+VYCnI7JXxCB9N/8c
j+I4355adUtfk4EXPWzhmXLY+9++A1lk/UCZ4pEtQQkZsrJ9hceKK/ubDmHZ4YzSxPL3jIg52q3Q
zoQ9ULAvQiENTG1vuBB9E7wVPW0yMQM35niqlId3RBUMEqMLoV3McC5MKzMVxPDckwZq2jZkPMaD
SjvdjMLpq8+K/G4gVMQ7qMSqpFAlpRn6/cjhVKTGFv1iQElIaLjDLRREY8tTn43dtlyj2oyT0119
18azNHdc7Ziw5oLplDQEmDENH5Uil7I65DH5oiD/y3/UgVEIpLxgndrCZ/7QDQ1JLO1xd6ShVO82
CY1wSfZ90nERtQ50ASuT2ZJaMfY444eMpT7U+IdaoZwmr7WgTyMxUDuiNVu+Z7z/vdzwWrqO3fNe
kcxWdR/tsEMS0kOHmGepw3vLJTm8wz6KRhDPhClcXcRwumLW/u+W42KsNoqeyUWoxUkw0fgjAiJv
81ZOXkH9jbAAvuSyABRwFoHBI6JkfPitWN2yoltMM4zNWRThPvIAu04HqWFk9ZwNEx069Xjsn/Bv
lozuNuguOtKCnIhIoF1N+5YxjkF0INy+HveUmcKjLkdBeA/hB/XWVs/k/LvsncLoTeS8060DbTvS
bq/YDn8fwpY1exnVb3owixjztJf7GkGyv+pKQ1uOia4mUcrEGiXK5PO83disB0d4WzWazn8yZe42
DwWSuk+y7WFzCSVlhVbFWpcbqBYXUcqKmP41Zdf9clAz881muCcB873cZEnh2SHqZ4kWn40WaIUg
8l4FHztKNioNQexSASBpwsuYEy+FLdI6SfBShQ9gy1ywsqUo2N7r6JqvNJwTy4jnnKim4V/j3q9z
RNzo9owCSrmSOY8dR08h0FwZHzG1PNFt/mcbyknKrnv2WRzkVQkP9++AF1ZjNdk4Ps9GXvJYf521
pfOOnFDwRMIUHWQv1q3p2BZd7QWzqqhS6CPnXsjeyjHdNwtFWzuk1ayBBWRdZHSBvP8GOMiFOV8l
6BDIjz5t0RhF4VFtYyAcHKN/JbC9tzkTXazfCGkG8hldd9BwpIVdREIhHY6U2yVyg2Pq3bUuSEUY
ItwKJNTv6pvIa+TJTAeTovbFDRuKr2wR72FZdfKz0Fqm2aKx1yDf53BwVmQekqqmg4TLq2cRzySs
ctfzcwDd8K/2RwFx2cfu6b87Z8zcVuDOVTt81swEnym6L5l+MJyPeJJvxbTF8XWZK3cgjZKcZqpv
Z6pXsgpcTkMnqhFxZTW0eTOm+Nx1HPQSSBnKy47VkiA6tv/MsAW9Z0LRaq8BNj1F2/bB/5IDSfWR
K34Uml++M/rDPqSnpaMbItPN+W5t9C0szE8Hgu0ERxwGHLOi3ohCeN2W3G3akbj6tSJMtKxAMf9Q
1xSgdEACTLOPHXecSKRZ7Ov9wcO8nTFwskcqMWi0Awr3nJd4mCUja9apdUqLHPEzyj4rovnI3ZmY
VtjlisdHHZ/gyqkSpOUOvz9R05UP8uJSJVYb/7GLNXVRYI8Dv4yIFViGBx+7amQHERjovJ/vT3+D
kd4GTaA59CvtcMMHYqtTdAStCPbASEBDVa8Er/Ufp0WNb/EA3OAOxMWA6Wr4rD3YQa8ebdHs7iqy
NvsRanc3FyelFrZ3niDgQP4TCRt8GsPwyAG1SbqJILEP/FGcM8v7MnCKZXIOobJARZ0EgCeRqRLR
WgckTx/ZGq66xxwW7p6c5lIz9jJ8DhOTJ/2WGnOwVqx1NQr8fKjXXUAYXibObGmhUqj27Lpp1el1
XYiNDCN63RzUKSbJAiIXP61+b9n2ypfVrVHf3140otRziGmPIEEXfdD/41PDljCiXMljN7Q6RAmx
ehDZo+4UzZLkes/zOKJEWKLYQY5AERU5WroG/V64d5WTBF9dBeADyERP14thOzo//AW7UsHstpsA
z7AfB+n5j+9vnMQsRxzo1zTrrio8sVBuZW9Aj7qT3GJj74l6GDTKqTtdhmQYShme6bQR1ySkVf6A
vPVYTqPCGk8Z4JJXpUVjxd/2tsLL8YmEpI2jLB+NXFqLGionr6DpLOWMRYzgzJFYsuiE5Kzjt8tX
dLEWo2R5D4DGEZaLwJd5G7a9EgtVVovSB/8N64cvM5s9NGVvZ+7jigCBdXwRoYr4gohfvXgx5Of3
VCyFwaPVpEtRs5JWydtjgeE33Q4I4GJDswOfby294HUdD+t10VCLK8LdaXCsCCGsbEFJlGhedvoT
yrfbJ9+IdIU+MmkRoYbQkrnpsLG52OqQwc+gBgCH+p8lKxscbxLBlAL/8HeBIOX1jWgSLNp9WbCQ
wkxeU31uiJsTvUNZoOE3QKy1d+axea2xdxXcJzMj1eofb0VzzSQH/6c8xerUQXv3qEt6Xf97PQAt
ISXM0M/nkSB71uI3wvQZBeHBGRQK0Y+MOTkSk/ARu2KFShCcuSJBKRYQqJMghAzBZzZyUi6Balza
mWEAk3GY/VxQOTONgGnqWNdzNdJKMx6zhGq3PScXmsW8h28EqkVhM7Yw7CjJJPXlYlVJX5JioGxs
Qyup0NvMdcvagtT88pnvARpqt44llak/zX4Br0vjzbKQe+OtA34PCwA+9ZQfoWbXjJWEHyJL7hES
dYvKkRcFNZ+IMERefpxYH9C4CLDwKsMmY0piTjilpmqMI99XY1I5ciCJBGx2BwDod9MA1axWVkXo
EOLXldXk3XMgKchpAaVbH2t5BxCfOUosx0JBpdqd+gp04e8sNRaUSjCyaUNI8wYfUXRTbHecXaRb
g/uIhRvl9AFxIGpb6CgQi0V4QqObgDRxP1XQvIAAKb2bBeX1HR2llwdH4YfPtF7ZzIvO3VZD45yF
RpEBdHWAVTt4Z+iCRF70vYbq4Ffx6dBpAGN7pF4FXQH107F7TIxYmoQlZ1/8gwbZnJCxSOyJMZvE
KtGMfrJbED8hVPDvQgcv80+qaj44G00zRBdxZX03ObCmLceSPhWDZfaqHo1LCSfaHt13hIHAel9Z
TvdN4APUfXyfn6y+1NLv0jR7obVLZscR2Lp6PPjWswNOnYu2YHk/vdcbKtZ9R9BpZCzNsgNVA4Hz
leSJZYx0oqxZr7hf4kOiCSDDyylel9DhnKkfXLs+tRjERDinYIT+CxKZXxxLvC/c08vus7ZgRv1n
yNYPn+fd0tGfZH9haMZfKZfq2NRu6evXfNNUG4t1DbOIid5JimgAFsJ5inNqULcHk9l3l1O6Jgg/
AHyjBHZEG9BKlYoPMaIVvPtUE7+iJUjhX0mYq7bOLyiG6ixDpXiQhtIEIguk622gnNOgbWlZtyU6
LckbdYoN7n+UP418r7jfMG7mgyEVhSuS3CrwvdxFMBxb91oX7Qs+Q6pX8P14XAiWAlQMgKDY/pBL
CXp15nFkVJOuosaaF5dODG0SjABYLSzCDgCz5NjLZ7GbbYNZO6MF3odXZu6hsxWjoc8U3hj1YM7B
3o/x7FnALDIpHYx+hXSPC/Lszo877KO1YWJCDJZN9PpE2zNPkzCCbK8L/pMEV2p+nLJCCyeqVNbf
ZJstDpGOCllpTbrn15WnI0hRgEe/OrwwM6RXo5k4zl7kn+yvaZsrNLEw/3vCBNjALeEzTjZp4SsI
udsRdwhMfhu2ASbQYF6J1WwGnRye8h3BN1nJ9ibZ2YANrDPotnWZ4E4fQ972BsGkGsu6ZxcUk6WT
tnfUQORwp22DyKB5w7ztkMKbbzGvD8x0X/DW7Q4Q6YoO9+bdaWrlrE29e0Q+s3fUD8L3+B2OKy9A
SToRg/3cgxHr52KghU3sK5Y8wBMJeAA9muMUE1bNDDXLTHloalTlyn1lHJtVDynM2/eN1/c8SYnU
lE2FEhHDDTMgR1rTq0pwgDK880J78gVMDpvI/h9Vp1+IXeM758OVtVb2acphgJGzeEezlRPN2ppc
g+VcZfk3SuNId6E/CaT16L5fcZ3f6pAFwPMp1ScT5Cd2b+O3BtTYhkxTkcT1si8fTQ3z6gcwPh/L
CIyXkPDpaVdt2SDP8o+U9LbJgNHrv9ja1lTQXSx4ij6RGTuDbccpc1xTuv+Zf6SXLz8hnMk3X6/t
XEmP9AJ7fIPHg2UGAxzUDaHqtr5qbBvnOgs5fY+OXhHEzs0/eigNO6vQ18APhVeDocwEmRNjUT0v
18fYEvV14M8Mz9HYJdhLJ+A8rLr2TMjoyJQkK7WWViNVHYt15P3dBpyesRaiLOzJaDVOJoYqkf1F
sKPJzyLETZ67vEVoEJKX+eXC++jTuZWTETjVBzKkeWJCrmEDmq+C0Gps6FOXdi0/r9H0oY6sx6cw
ltDUn06BmqWxhYocuOZZtxTcBq6GEC+5u54JfDEnD13dmD+hJgAFTePwYi/gTbgX6wzzkKee5jFK
EJUbl8XeCWA8zuS0hz78cvUTYS0jreDP0GA3nQAmuzFM239SVUJaDXaZAwwIqmx9AMPD5MnnGisf
GrO4ntLpbMh0czb5ukUEBpeqzgojSxeFm45k+9rqjj3q2ApWOXd12lpQE31OMb97lq7EappT8qJN
mwxIXcSMYSdetp3EYMpBJZrLBFvnlZDLRtZQs/SnAFOO28roPxajXLnMF2UAiAVQtsoRipp76l7w
JxuiMO/IjC5jtp/7eqbqgOprBi03K93RcV/k3fkkkZHRlQH9I11QGYIMAEpt4zJkjhE0qvXeH7Kh
hLf46627k7zl6khvSccvnAm12c/F7T6JhzQ757A5W64yzIgodpSk883aZARxXQrrQroByKetwR+K
JRXD9w6XNIKYHXVhaojct4NCORsTP1gBKhLYsnWCw64HNTaR0Tzp8OmOLamSp6UKBoZZcMNeek7z
Fww8Bm3bGfKQDOz3di8nIFvQ2ml5vltWTX8vqowB27qRUaYldInIeIO5NdDor19MJiAgQNYw+3vZ
8ysDqfQHHwMtTSNhUOy06eY7Q2D7PUmnSLjotzRWiyg9IMA920g+ocB/4lB3lowAVCE32oa3tRi0
EFI1UjsjjzyQ1DF4RjWzxJ28B+iSORc3tZIom6UaPP6gZfbo/Lk3XjG3iGyWacoOF/EiEsl3aKQp
Exq2gB+GxGeFKODsT+Q6EgqSwtvsry7bTYa/fyVhRF2DYNI4mNOATTLd9YGSVogS7nlkCGgTS9ht
6XWaS0ehOb2TOjxEwg0LaCPVSSzqCy9r0eORJ843rVVdjM+i/C8Jv2PSOstMr9Q1kTpuQ/4CdPay
OJZA0ZekyhmDxsci7MGGVx9pJO2aeqHtreuqUNF43QFForbDGDIJz4B1WkYfehtLt59S131sHLWa
5ZUgwzno7UEHrIjz6Tty0vrOYxcdEHEPNRgtZWx9PA8HbFm3l+rwyezZUEFKLe0XqlMFA0vTN34J
kHidCUeXbtl4DqDcZvbeMmMsS2XWTSyQymuVIR4ci4a6IZg7WzFYTQGSnV6MvlDMSxZgpPYUHEpw
v9Hc16TwU42I89N1YeHw9HTgVFhANx1n8fPpIjWbWbA5AxSrmYv9xFgeCpN56z+95NKzIbXEQhlZ
OEeJu0AiWzYeCVb+o8+MW9d6Mm2IkJQAcNKwMxVtAM9ohALhQOjPFdAXNVNwjNztIdWV6nOJ0DzQ
bKbtEfzHup24/wZSoDdmq6jEbeIH64vVNsn+yGWJyEELqmxlBSqnmP7Ai7AJcYL1gOSdaaObcBkm
HSDNGOpAL+vKzNq1nZ1gZWQrP+jynTUHYhDscXiGdr6qv9AQ7ubJ2gJ7UDQ1MV8EeSLntsXj1kl0
vv3Fgou06cnmLXWSebP9hCyEiycuk2PXYIs7j/KJB12+nO/1jvxKlrqgGlr/C4lILYB6r29Xg3AR
iaHBqRj7EQgwk/cVNqaso3VNXqd998gnj0+x0vgyyWWaladzLqRnVtqgmvrndQqIMWLm1pF2ojgy
AQqJqseX44UyyqBxad3ogBa7FbrVo8xAUGbXGY82Gt1fAjAi9KtVshWiPgkoNZbj9emmaJ6Bc4MV
pkF/vJ9SIYPqIdq1dMFlDyEcIdUufWgdvGqJ1V6A0ad2dZ83IRJvZ7um8y3YAe3kW/YzKYUgJCLq
Tk1HUW/cKhS2NteC09zZHPqssZz7sXJqaUSHSPG8qi384eF63xgtYeVDxE23nshNtKSvGo4tU7qb
+8NRfDMJP4zmF41XFDObqr/ZHNvfVTL0nXDf1PBt49AC5sRQ/kefxBxIzEcceJ7mYGJZXq/p6P0o
LMTmv2/w6vH1VE/Fkgr8BmC20ij5XwZqpKinw5R4kZ6M0CHyz4zs7M3dvVfzZhiF+/N3x00X0tsA
x46pn8PFSib1uUTDNJSHWFzApV62Nwo8ejCYV+/z/G6zgJnFydrUuXsYqs7uwHG+IEUom0WhPajN
Wbtn36AMVBdqjkcNTHls+yg9RmfuAE/kZTSlN980SzpSJ8aVdVhHkWxVworgfleJjU4SIztUwszE
Uc/kUjROTJORnwS23ldT7uUqaEITDs2pOR2e1c55yOxhmj2zowqX1GUAz7GYIE38dDtrxFoAx48i
rCnkn5GNkkdFf/ayjD1ZH9LsVsv3HlPDsqzdjDOWJoxfV9ohcOhxk6/vcZWl2QkqFK6fiEvrzwkf
amJZR9nzM04GlX+6AhOWPheFczCEwGJ7vP1GAtdo7updwg83FKw6KImZUj2vRJ1riVofk68q8J8p
uEK05VlHLmWbZNJQatXvqo99D9NNS0HFqUpWOn/HWKzt0s2ayEP8s4JtscmY3ATP0WD/u+8ycHgi
05/vlPFl+18qfylemsnRj2mxe3LFGMgbBkJ6eWexeX4VknV3F54RW8oFN19mMnMiFR7rOEyhOPla
g5VtR0IHMNZGl0/dgijLLRU+2x0f10EsSqHKIdX3whdcUN+GvaApUFUySFnqdpzBDGEsLBkTucY/
ne+cTNfJcfKEYRi0F4rAOKPC6kDWwjUly7XWmz//Y9HfR4EI0PVw9iuLi++FuheS658P38QBdRDP
Zy09ZgDwqx99aNB7wS0ikaktIyLBclxLJc9SD5SyxPOX8GpeVud6ce2gqlnsu8CMORg0zhtg2a44
jRDzFIRWMjCGKX3fUEoI0axChfHgkVJ+qqnI+TH6UxyhlHA8C+B4CUGkRFp004l29Rc3k7HwbB84
vDtXC2qB+RCsuTXykVYb/FgdVWQdzluBwMNultN8cCL73+KjAXNiRHgD7B8bpywe4sDycfLeR0DG
DhpSIQRAAf+6mJauzFZ51ptWKZ0clfiGaWfSpQ9RjFnBjvYTgersYwffTtUS4PHHM+4gA8+YKJbj
L/EopvM5davcCWTjGw65DdmcF7ul8tDnwuFR9XcFcAxGaA2+cQcnBW0KzZLqFJn2xWYsnrd4OwIx
o/nEeXIc3ZppFgh+yM5g6Dd60Oz3RCnUqWGoGGoXcsXyqOZjrqOjt90bMIWrJGJ4sLAMFU8OpdXh
qZ5PJ5TSCsq3X+ALM5xRqHz4PurPAfsbgN6CG/v8vMrm2/txxDbhpIXdWZuuITeNNGfXham+4IPx
csMtkdVrn8a6yhevhHH4LMFMFdxfjNFSuhmh4XOZGwgnOPSBZa+WumtgSUlnVtc1Ab2nI2SeORug
sGZdibmDIaW5691wcc8M1OVGTtwkMNxbmrVLr+FiPA1kT3VBn5URARwwIBQtZA0Anx1qa4F74rqX
Z7dsVv8xQTo3VaSald0WBVC8mSrTZmVfg8utGZQxtKLfwwCbil42pHec1ybo1BPnaBFd1Z1dDCU2
9EWHhbVRyEK/vPizVy+1fZPbqIJau5nUcJosIVIQRVcdcQGdlfk0UVS+om+rcQIuiZpf3mokWkR/
vCduo/eR82wqqICmMoNVGjXrPpaT3kidNia17TwU5RpUXv1bmhBgDrBBlDkM2H5f+wbPQ71qCCfR
Eotzro3rkrxAVz5wZAWBrYyDJyD4BP0i+SdijUaaMD2xyZ5eAzY//ERaVw2LKcEx/1RE8en90fh+
p2vsoTCCgCwVGChjILl+tOf1cEvtxMiyMHr/jreiOOPwCvxtEIE0bYkA0/2BVV6BqJtGNWK8u3s1
I38HM0UOvQwSP5JGH3GuM12h21ThebhdK1BtLbXTSCI9szguFY1t8s5tz36trsoiPxOVncgaoJGq
E0yjG6qf8brz8KRjFMwL4YJBbk5rIPaQB8/OuKZpa3rQYtj5qIU6jU+6h9qwQd3O9GuXuvYsy4oH
lym/QaaHAdMxA8QpMdqnyEUGJ208/M0sB0Nmd2cTC8qHfvnlcDNE6C6H7fx2JZDksieteyb0Lwjn
xJnj0Aeg51t0rQ41we3l3DWbSjJ4bnRvqxjbj1Ofq5mo0lU9RZj7rp8X21rBrwv5MBYAVgSigRf9
J/z8tf7kXAFNRIuDw5ckFtbjRV8lGmYpGkl/X0bAMt/02E0HzDbdhNPssQG4QL2YIs12Ttvl3gVs
+qBDt+fYCiVp08nGeqpkOhmjnumfRQbZPmoKLnOOUn6U/eMbkbVxsowHRIpiyT4Hfz4f57ZibB0O
/7g8fKVZfnkwCkWq1/HudE8wuftOIW8IC2eqQe81kI1jh668vEoInI+w9FJKoO3GCjgQqPui3WI/
RlNGiAY2vKol1P6zGT11Rp3ZqYeuWV3TpZhiwEjNM0g/9tu5t8V9UktJAQKqUMRXGK8DyWmmIVza
zNF9qItatX+/XNIwys5YGI28LJnfCiu97qolvOhsQVHEyNmOCKAmGbvarJX2sPXYZbbWto5SYvJ/
LsUh1GTbrCD/F9HrdVDELgl2qDECViTw3DxPReitLb0F/lMuB0mlCIyD692zPVAgQgkhm+WwXWBe
jtFPli4FOpdlGGbbbVM2axy3tTzXSR6cVZbW9sfCD+G1BD+R2PhS4/X8QR7v5ps4ajC0yoC+WLMk
HTeyfgf3vyz3Ss4omMWkWCZbazL6XuJpzCdI9aG6PJ6zwWNzp2QnJAbxVo9BWCVnyiRpuVl79AGh
r3rZAROL8G0F9aCpSBI2RUNeFUxq0yvA7K/0prhrKFmKhLtwWUyv/bi4Uab/bAPzUMs+i7aqYZXh
1N0aMlECw9P7xOfnNGzRiqFQmmeanyA5m2HXQbHi5AHF3veAqCp3gbjQQczDfjnZagqCUXqdvX5G
fnPAZW67wzRnedxxLgp/dLTkuUVaqwjJ7VcffItD0ewtmuZ/wiu69c8R14rqIOTSY+Ng0w0zWWqF
eSTlgtbibWkx7/rdZaiIx5OOwFkAzvhHqUU4/8LQYLaqtppHwedT4/Aqy48XkdNPRnuzh7AJXvVJ
ezgSPQr0OTfdIr51YCZMz++J9RlwFlEldfo/6kRNgjP6wF1f6+QgBKzbJBowhyFAnfBosZebKbqf
goNvCWLwBJAyi1+Is7RKx3jO5+ESXM5r4IYm/736KMsoJRrw2oUNabSGSLf+WNwnvtlKF5qFxjmY
+ahA/mGbi0Lye+KhVYjsVLviuULOuUrYuoU4bLekIltrqR1a69UT8MT/mNT85nR1kqJUpEil+DJL
qzOHicuGHtjzErfQpV80DIoZ5zei7EdP7LP3jgA111Lkauv0T/WKZP9WpXRPpDmcCWyrN1iOxz1h
EUIY3Xn5tPWPFxARqMWKxBbZeAwnrnm1OxqurqAxf5rnWVKTVbJRu5bxX57XDMSe45okFoIA8GYF
ew01jRcVLSRy/f9HlhhDjURV4ibTItpa3ab7LErjIcnZSdUlxiJniDB45dEqI7OfsTTRfEwcf6sE
/CTYB6REOSlhjJztzs5A83lNrZFYTlGnxm/+Bnm1Eg5OclNKhvBOIegHdWTxzvl45UJ6Z0bdacr0
FsIwRTEfWV/0o5wR2jP7Hr+mb3SdiFl2gnGzuzjFw7q2DjkxKUFjamKw02mAJ6PIF/C7UjXeRi34
zdREhuixdSiMYunmDbvFpAWpSAldKNxP6vtJ8UM0C4wWk0XbqLs7qm73eeytGV3rHRUUPteq6ADM
uV4m/q+as7zcvdMRiN/k5sJQDc/VZsxdK+b0hosd5PFG1rK2Gzr02TT8hCImLBAWdpmT5rU590RQ
VuL2tGe39sbajTvuYP0ihSAw5skXZOfykaCBItiYGVAgGHo7KhSnx+FE9NkKBjCka9iRGaZJXG60
CfAPugdLUYyns5Y5PuKRuf3iCn4FuNGHmVaCkHlv/XWYWEWkMqYp3xilLpnTejCiZuKNHiTKUXdx
YYYQNJp55g4yddRI2udQ9M9UX1N4wG27CXCnBRuF4PiTqyifSXON/wbds3gk83Q4DkRQZqRYy2oq
DZU7FmZzJJJI1uxZHdW/+cjjpMRARqpSdh/Jvx2W9ekEdAu5xwSjTGg+KsEi7dlfUJxJ7cP5iuPX
vT8CRPEh3VN7cSMG9OdTxP/aeQ8qLT8aIWeEk8dwd5PgpWLw2rl3qN44oMwhszu63QqJk7WwJpQz
AIU6RLlr7qEDXkWTgoyeYngMpmIlW/n2FixTRwpJFkpdPgz7883Li0RSVwPox5yLnVXjKG4yyk3w
LlDu+G/zeBtegjWRtD4MqsrB5hBAqCCPyF3yMawCm4Gl1D0UqO0EryAXuFHhX0/8HrvJQY/Sbxnh
Yb1c4pa4gpjTOapkBNKIvhs71WfdL00ZBevw6v7Jyd9X1OX6BDwfcqqYuKwq6c2Jgo/XwSBVyNFt
yE7kebMcsj36jtQGWyRa+TTl3yhkYUS/g10gsV1uBlV8iGU0+ZwovNm3/rB9e95Qpa4yXQnsEZuF
O/7ogwZfFIZsgAeEKrOf8exdRUuni2W9kvqucl6Qv2RBxPSw8hwWe5X/PfwjKfilivlXSkx+edsV
J7WUjLqsYCxtaHgAyNckNvKuy6H5Xb8RIm80EdyilBdrMf0GH8CTtMMhP0GeMv2Q6jbhCrGUIEOs
TVuMddJsf4aeV12rVknUq7tHiOi3o4ZWWMs7narePY6NVNDSCLN6Kojjccd5sWDmYhvWkurj3DGU
uxw943xqi9cCLz+NYybmY4dT5eSRoYlxPj8ywJRZcrQtaFwnYBZljRwGfm/9u/iS72e6kbH6lXIa
6r01awlFwV42Ns30ri3iu772/iWzY8lrpWSLxrCatUT2OOJxlMnCBYUokcpyFAzUwfAp5gHldZJm
hkbTZVHIN148ji7IHODxJjY0ZiFKX5MednVI4DEUUwIjcqjssKR67O18lpYHL1TcOuezm7rt4XUz
m93k0PojPZ3Vp4/19mhX2ro0Yma45M/gvLgk/m7qzk3Lazx2rFkfG2oIN+THmRyI8RGb/x9+aUmu
wPYd2B9jiWIzRaNELJDYkxQzdF0iDEhhVxhgeXebre4avkemTMQmD2Z8kmLC9J3SNoXvhEiXacTc
zYf4jQwzmHf07UNZFdnrxwBejh40hxrpOHokQ44WZiLVixfMSrFFVIRVTv+R0ivhg6qQJUl+HeyJ
b/HWLj0lnRiaEYFAhf1B/9qkjQF2ETsTHGSbQX2nKaIsgou1bHkejSiTKmJQkVXOhonTlj0DL0b0
M/TcitkKqvc/a8yBGpvVKERHY0hT6EtS5tdupzSSeWY0wvpSLxLYEe9KEQamrzIbKKzlP+o08Ofo
ae0g0Z1Ubp02jB+bFfzScX1DaTn4w3EystTIUNbSZOKHboTO6sOHxjt4E++EXUDjbVWieqS4rTDw
odtkrJ7nMsHlocgA5d39fd+9Q0C74p3COWDphj1a/LaNXsfJAcirV64B/ySAhi3e173y5kJdmqe6
Ol/+TCA8U22yPSttKkgmt2z3pcfXGGtX1llGPadrlb79dGuG/RvPCzE69TVjqq+SB6IVa7oXjyBF
CMnYxp1gYxBHZLx+2F+qckl3FPoaMYQuBhYLaIszwSLqoxwcSg/efKRBunsOvU2839YC3t7CLUs+
RPtIsFMM5r5XEEBwxnQkt/Tbz3aUhyNkcwCyk7ERntgp00RC/ZKXODfBRcmmOeJQJIUlLY8gMDOM
ySUFJY39jkFKlUuybTtca1RYWHCdesMzVBftyhWDs1EZf066NkVnz5RrMF0zkFpLmjO1Gf6qMjuO
ovUyabFFo5sZvjx7izTAxzYOIywBzanjm+QSOEaR9XsywGKsRzLmVusJVH1ZT8Zn3en2ne9pLMHS
R1z6OCtZry5acTZVUS5kxGtY3pLEmIP2FFq/+4q3BX6JibymWARDW2vilhUxQAL383vgBPz/KyYV
kwDBCpzZVXD5fN6LaSOLtGdSEiLk2Dgb7d04x1jdTYnNP4MFa2YacgFbpeBZMpXWiWn1mX8V3TDv
/4RLUn34JwqBa5iWXY+vF2/6eeSZLxIqwD6M/f4/P6pSdVPmX7ObiXPgG3pfEvk38blB8uo+pB+x
CKMVTZyti+DSIGJgqdORedbeQeFAHqpibzcrwBpCQjJ4+jm//4PakFL53B73hwwssv67ngvfsjMj
l4zJF78ceB2EFwjaECfNhrmhAXvP/VdMCDq8TIDcrObKpEWkeOVVA7OSGQhvDwlLRXUX+jzFjoHo
69CzZ6vLzAtkD181BvnzJPzSZOS4EIB95p9v1C+Et9WVV48/1QSmHnJMCbbX2SO47L/WhKeMx6MU
X6RssKwtAo9M3Ye3HkiGTH7dUYE/ocMSF8g1oRXcPLKdhBSeC8rzSB+O10Xnb0RNx4CSopjr7Njm
UrCC/PNmuJ+EWoBOqe0aYbFUVoI1A3xLvs4vnDMZe1DHp+9WIrouYAwp6Py13ukviuYCpogOhQyC
mJ+IGPrGJTbZBrHDWtMWzHdsGpHEV8M0jL22fsDAVEXNcGeulhYKYK1c7XmOo4JAs759uJLhLQ/o
23F1ZzSc+9+GBXrUvmYIlH/iIIX39FhPgvrFeVnx5zE3AehADAKoGUXgqoV1eO8x0lb3+j6hQrYw
b+Wkjxv5Qjys1bcopHTtC1STf7BQD1gFsSAlQayXFx837axxUfJxQo9pGjTE6/FJfIAjSWcIsi2s
DsXTjFOP+tEzE+bwUUjc9I474oYoW5HSZ5VmoZP/ZL/TS6eSJq3LVUlDxJEEKKnMdGwu8m4WnrYd
6vo9n+YPaavk7LHWQTcwawPLLS22SWAJrOXez+1i4ZnztBc+JDuCeUqOtMWCyH+Xcscdm4JdsTvb
Gt20B6SY1nKQfzJL72OWuNFh2ImnCYwRY5EkG2zIAJQqOCnTJmISYoA3SzUWVLdbOmtC2LVngdFw
GA8dHv/GTcYL353a6Qs3ldNIxX+WdJ9T7incCUQklQH+aypqim8SIApAGzblSh8vk7hiV2oynJHM
siSS6nVgGh2i7hirLSi2ocB8Lk/tnAfottP0cyYUpIABkRQsQ6nCWZKMbn1mFE5GXx9zr/aqYrU6
A2MeGHQ55tKxi7bL1CD5HLbu6P19atOOPfTpphn8QRqW7wT6zLQ6szNLn33nBcdQpvvCuxCL0h8k
6gOpsbP1iY/oyvOQw0YjmuVeTLIi+1pW3n8miYgMYkobAqbWJAgxudjE252X6DPjbwXF3CEmg7q+
2k4iwoaiQyyPfMKImbJ78L+e1mJM4DPMji9F+vcZrlXmzr3Ap47DIzELspDiU9XkE/174z+omq3k
UYMQGzL9H4+05M5mznNDBPLqZyMKMuIdzgtq67zcxhSFJo7lPQJy5KAb/SbQYH+m+TAQJtb2CiCc
zGYsF7JlyPAT7s8/LR83D0qbRL9DbilHIhWPPjyXBdfKjgm6oL9tAGsdt32jjl4CTD6s7YU5cTU6
g5QHcTKu7ycQTw6m7xiWzaS0EmjVRtXxsewSgUu1Z0hK42bOVqToUXEjNHpMcnNFcX4SjUIwqD7z
TAqx9WNs8icsygpczEuBvkVbxCZ/4UtDI4APCdmDiD+ibk5fSRCuhzDxGtRwK+M/KkPcXgMFUDSx
2pawuQtW+cqz9RbfU6gnZgxuCOH5EUThs8771M9/W5e0JFV8DJrPVdJFaLd3jbIu9XlvfNt/qjhR
cWOUk/SzHY8F48amO4sOPCp5fXKspzCgt8oXo8W4CWF5Zp1AvvrNWB+AskUif/8kCkC9ucZpymZ6
83Xb7gS3otcV0a5eILBIUtHJZ+2ONUAQqfyyeOzn40HZxa6akbDGWIIi7oUH1x70nO/drjoJAdAU
QRdui8nfgSkdQkNmde32Zy/aBCxN0rOYmbQbeAOPnaljnx4Q/3ybn2nsPgOMrewLzHsCXHSoO67q
W0fr/mteNcZ2B/taT3zeqrcjg1mv/EboLDjlWUL20TRq6rLddWJ0QIZmrkMqH1+VQBvMipjSJqNc
kd4qXy/NdGlC449kkJet9x1m0nCWl0XDj//wekjLBMIP+k/e0nhzWeTtWVkhhTKzq7wl2Wn9bzjd
VDr1wREkE8Q0hd10c07fLAyQOionij3yaB+OXIooKcz/Kuh26xWyzcymvamYjf80ve1kG81e19Uo
922myRaSsmVMltH5cHP3FDnmKXstlLOHBk7AlWvxTct5ZtDHQ1Ft+ysOR1XkpqW0U0kIl8lSzciQ
u8Y+4l+CP0uiqqUNetKHDTsRSLLbZwB9BvWGIT/7TdR3XgkhTn9SPRLjzpDTWnhRRK07VD85RkqD
9uujMMQjzCXiH6wFOK1/mi3Dp2P7aqrvW05tzIx7SMV4xf2jG1J5kXw3uHsvUH5OhCBdyogi4z26
wahUrErG8yHgOpSVZRkvt+3cPKemNkvlT1SxiQMwOMnLLBypZ6kggYAs06PRfFefBdkD4RoXUiRI
RUzRJXD44aP/Fv3b1R+o3P3X1M3jrZYU/4jN0CHtQJxn3aglcOyr1Nm+PHIfHp8Gz8n2+VL+JALR
ZIZGYg9dJWeTyKmKOuo3hZquEVcX+vidUczwHfPqiTRdysgkXD/xxaKNGvhcmkXqt0ILP1yBXBTv
tj0Xb2oSFddmzmRA1FRkBNk/kW3OwKlauNnY02nhCZPXYfqYjzVdI2iYHBkeS0hqAWHHYj6h4pZ4
ODpqaOHUrUWuPzMYf8+8PRf48sNJ+Hib9JVXAPBeK3dGjSh4mQ28nniiuWQhAAWJavmQBNScdkMh
9ZgXgVEnYgKglQEGJ0xE11ra72nB8YaMbnoFITUKUJwAU+8CwDA+TCYM7dRHtncYvuUTSs83uKc5
/OYZUia810pt3xdkTRWaM36cdluJ/zFWDXa39C5mYYNHN4dupk68m64e/v/R713lWs1M/ek2Xbkr
nYD9qDBoukQetYtO4CEp6mHGm4hur0CDfi2crGI3xnYp2HBtIVMnLKlG3vAX3cro5aYG8CGrv0OF
gF8fpE06WIUGpYvBWtNoq8z2MHpytVI0YZ8zuaK0ha9EDtBOU6enMJHyYZdjOantq/pLhvvD4N5h
BgAzrK6xusug3FtvJJn+Y/BVBRphS7SZZOhEPGyaAOa/jazc9PX3GDv55XR/d6lWA0dZdOmhI6j3
I2ZymXoGb3flgk6wTMWKb0FlTB0hv1f/Ag9a2o6w4g+MokYlwg1ufVgvtGcMYuDdDmdv/Zz20c1A
u6eUy9U5LSBCorzP5Xg0BynEIRvGhbSDI3BWUVAPRerMdxjSKgmob4gaYAoosqjofSM5RqmSNLvm
GvmW2q/mwULl5BcUvP6ZT7kiqprnBkvyQ7QlTS6c81+WwmuA9AtsASnBTOWIHycTLVMUrf9U0avw
pR4mu8z2H5xqDwwq/+yP0hiAVqzGs4qoYN3YeNFXkgpxuNWbqj8kjSDZlyVSmJEKnJ9IT1Ok/+Gp
G51Y5KJdXEjgnm2liDFjV5L2miJf7slGzLdWHEelvbIIYepuWE2kUVFzXuU+VDVqjyMXyXQ1xxAg
RJpJHSGzsoGlkVA3AB7goQwECRuT62OuW1bxLpTCacfxfjVhd+TBOazdF9RGzJGfcoqEgSMnKWKT
0tt8sHz0yeWNoUJkaYuyaGl7g//hFAzLBJ2o25xMgTR/bQnIzaRFxovWnN3UEvmwSVu5quLc6q1E
PLqwcg8H3e3xrSh+xbzNmqo/4Hy1Jp0nlAcYGcrsp0wkZAANIarXWRlpGA62yJa3IYlLuDQYLCJS
vizwTFKa9DPiZeRM+N1cFaraIM+wXGZEX7k+djGclR4YmQFTBdDEgtvOP9vOGySqIgEjsb1fw+Xe
EY9rWkPv8X4RZcouDeoDt5P20Xguh7wFxFPViZIlpJPUv+Nx9aXMbD4hmpFtFcWl0/4N8gjUTAKD
5SZpvzoI7S8CDTemg1SPYCo0Y/faOKb0gJeHE6uC+iskElx6o/8OiKWiyjUUNpj+AizAX3yPRmZK
J33m2iio4K9C2i4xnMtRG0Wm/qqCTlWDtBxsCdADsEVpqyezICD1yrq9IFWa4jadvsKSsRmhSolv
U1SGr3QBCxnuKjepVajjQAvVtFr19QpLuCrzbuvzgbPSQKmIaAl5GA3HYQDgm37+uXOEArbtiuTk
bb2d3SWuEd0XvWB/zhzmWKQ0lbtJadBC1mPYdB48CnD0F1L/mDqbzsu7pzU8G9o8uMCL6ojFjmox
RBeJRFBeRC3vZh3l4VW6ma8UGZoAMnfYUHmqHsg5uiHbOBah0BgDi1ianFVpM07YRdS/0Fjgr1Qa
77H6K3UKi17ezKi+jl4VcvOx9IfpYTtz31qMKkdcImCEl7AlhIRw2x3Ocz4nllytfWNHQmyo51Xb
asipFEIRbPqR18aV4/hYpZzLyUS1RE7SLyffHXbQ0Ty0jYzKSMufAEgn8Pobe3KhLExb8JrEoQbh
bdA2Nhy8/V7/gqCwZKVZk2i3BGaOFy3i8hiI7Kq4UMqkmlseAxNlEfd071OFioxI4xq5UovhX9GM
as1hcMcEqMHVbV0B8LpMNIc2zC+ucqRm4/dzuBsWB6lXz/3oGsELWH8Y39R06RcmfX3g3jGcvnxZ
U/blN5o/iGnAakgXVOs2Ebxtj9IQ1I4JP0FnD4BuSW32rP3ovgNCXc4NYzabTJEmIatPqav70GAC
7wwLvVQgUs9pj/gezZxPvXAR8iWZyAm1J9BiwRW2X6BTHt9k8OCuKzjCu7yQSJju21j7L5z1kk0e
XOeT5vU/hzFUzbNPy6+mTkcFUDq4pXK6VcRGAZ8jVnNXzRfLwdC4/9iNk0ix8x3Zaiknqs2eeJPV
wiSk5l08kX7aZIqxJrtc5Azawdm+gNyydDFUM63vKrMkcKbFuGHqVxwTGR09X1V5lUcfQ9ZqTJ1H
jnQycLWuNi4MXsY45AcuksO84sGAQHYj4jAnqhI17iy8PiCn1yZwXg0qvgIFGqBhbuJUSggUwdMu
512YoC5CAH4n0LLrwrM3+mnPWIKKNXVfBqoWFeVRvEQ74KxztR8XKGTEGx2kfgKlVwQeyq01ZfzR
y/uvA1iy7vNRgTqxmFmZeB+yZACLCHQBkqkhh4defJy54j4UiqMq2p0DcKgboQsGCcTWrDKnt5hc
PMoYIGd09BKLlCiRedE0YksIjr19sds1RM7+eRpWXJPooPurT44aAhlWzP1bPo1Jsa3n7fe0KM3S
iUFo0Uppj0Vv4RWaD2JGODYPUwFgsBNmi0R0e2hkV//JzUQvWS/DnWD6c1/f+34DSHb7ibznj9tc
KX0XPn3ZguzBd8gS4kdEwyK9QwNqt+Djey/oLqDcVELNw6dWnfSkvo8iXhzkVCNJqz3hDu3yQbQD
5N/I3QTuCysdFRg9oXqI0VpGBNjRXgSmkuu+N6JfL1Khja4AqWUPiowrVhO0Vo534Qfj6Y3O5Ydv
Cm+Udk7iTBZyXGRbX31+ujal58Zm9XywEyzgUd6a4BFetXy0cz2snAt49jyMC4DI9cvCpKEJa2qG
g8d/UkQHeMJIUFzZq/9EvEl7NSLVBX+hy5U5KAxp8HXONBtpTYBI82pRQR0uvbah7Lb3xiMPZ19n
vpUzJPzAqRDfb5zzmaJs08pyd74PwXarv7tLoHd3cPk75Z33FKik2k7ggDAqW7DyGvGSFe8mPKQ6
4Y9zvxmKPxqDsGdz7uGTu69MNAA7yHfuocQxq4q5cOYexVLDDR4tqFIVQh2q92xHTo7xf1X+0dY5
SAW6bkPcQ72pUBRopFMU7XsaIVH9LD6Rjtlb5DchnEAlZF15Z6xng5IwZlD/suUX5oS9556ZVdhb
8VdwwfJwWPlYSD/YJu4JXD1D4+AaU9VDdxTT4S1Q0yCAH6mVXt2CPDxu9r/hMOStK1BmCjqNUw/G
tKtp8MiSXFzGvroyBFgTDIDq11f9L3JmZgGNq2mAM00YvcyX+FoG1I6Eyb3Tfv7VT+N9gIN2jLox
94fWUHpIv/VJmMJO1VyjybfaOqcWCNDs8DYA9NBiNlF/YtCHc0O7ihe+rHRWOH9eZ6uxi4kXfo/y
eQbw/nK5Yok4LTPcKLvglfMIUrGCKWlK+FE7xZ8qWmiUokUudq2ibibgPuKOOVsYOWCKlx6VNzFq
vPw3Y05n+pYqf2R3onGaXGEm1sTiVicpbY5AqY5vw8JNyHC6dgnU1K9sNzUe++NppLz8TCKqN/Bu
RLwmwKUoSFmZ7uUU83/pR3R6CQLptlBxdNJLk2qXrBYplISg8Ur39k02X1QRCSVic+m638aloeyV
8sSdu1IiPqB3GAWCGMDIDqivNw2RN4QOrODMJvZEEhO16zmWYMZessSN2FTUGvEqYF9aIJyReQwV
aceUOGq9EeirMnUPtvNxE0Vfm0Ger8R2HlTeGFdqwmumhLLcvKaMjR9+bBP+lhFUgfxQjN2q5vLe
hruz52eVmHpsUUbPw0V8H4eHrpfWi+lkLtjuADb340Ji1Les21+V9RtHNkzcKZIKmxy+hTch094M
k3A7hSVakAdv8O2c6w0YPm5iLCqNPJFagbiMsgLkA3J2b7fupGSvHqE8KCjzDh4hRr/KL5QmVJxp
gc8Kvte6AJNB9hUDjZnjthJCMrgYM7mTIw1hSIOpXrlcBfQx5xlViaBJau1cU3Bo+LD3gTM0x0VR
lHek4oXT+vGqTXhAUzwyLK8uUSukn9R25z+8I1cVeAJANZ5EhVcf1Y2tsPWn+dwyYPSvgEtfmlnO
9nR2xMepZB6WZvYsDec6EzOsYPe9p8HNUGFT6tx0y0a/BSyK+uXlGlqVJT3YmIpCSwDvKksVbyVd
BOg0y7BjL4S8zGc7tRyUxVbzTgJ+5954WpT+KRZm7x/wF4JioDdPYerKNGH0w7QiJYVDtHwxH511
W1M5z3ThlT4Dgjq7uCyEmAUzyqCaJx2NhsNNCLJoci5iZmmbgOcCGO4Rz7naMHiKa0aeNQb4aXF5
lmykrxXANod3GxsChK4NvckAeILHAmDISJ2COU8RkM/EFXDWXvbo1a0cMcXe5O6YvY1geIhzI1bY
ZTqOyuz52VIJxHtVU5VPcGteZO/FkKHbsHYRv37sYVfsQ6YcoFGJRd1GO6G9tU6Y5sKYzKor2Xed
ZMlq5kPA5bbKuxN2RA9ATfiw4OFpAgWQ/GV7GqGsRRnn9VRM+ay9MAz3NsDuha3mZTMeyXV0/HD6
5n2Wi7dW3Z7b9mEN1SLZPltzP0RjNM+Pbvg3IoPPMHSCx1cm9Bavx1FKB61YMtxVr2XXtb8uEnnj
KIs5JBWdFFjBYVDBLbM9FYnNeJppEKkQSSaKJK5NoSqZbSI7TZ/ufvk6Lv5G9zjw5UxRvfrCdT29
jdLdq5/xNq2XcGYggs5vBESvyuXWZyPBUUcHcPxpGr8DrGhDFAA+w133a7tjvwgJGEJcYfYaf4L9
CWVh+Q8HlYwKXlFPFgPcj70blnnmogslsXLTlmUkoP6/ROkDiaGwnW0pL8sdAPyC0FVQ9KJ85ntg
eOWOb6gWO5zmX5+wh7z01geOJPzbb5D2QNag4Aw0PUVwALYmwT6pDMAc//5J4fg2So7eLtt2RK5h
8Ewq/KdLeg/RgKijQ9J2OduGIwEA/KIdKDLD4JAwHTW3K2MAQMuTb1rh+b6WwdzFvDLlE0yK04ZF
y07iETTbEy4HJsgw/F86ilqqSXyb+aZipMuq12KHSagMBcf3zkjeyg/ZIGEiIQftcuuvGL4qtwcy
4grtNx5N5CUTGtzRVzFmarSU+zjiqXljJS8EY0st7VkZPTYZFUM08gzSyvANQ14OnZkWkT7bpy0l
pU+f/gXCY99F8A6c5L44Xz0FjGwsxsLQL+iKmQ+FaFcFZ+VtmY1vESXFYF170FoUA0ztQj7kI+9I
cAwt6asWJxMI8vqnvBFIbjccfZJ8af4lo9zhR34/NdGdByjtFcwMe9uaPECRMTb4q8bpOjvgBkgT
yvXcvN8FCKa66B8+xletaJEm3BFOWZZ8yZXmD+N2MLJCIVPGxIFNE0aVJokXv71O0uQajwn1Yncl
eiWdf+rW5JNJ3NRkepB87il9czKJ1lytWKLrkQ4cqls/EAsiVnx5luJrAKM5T+FrV/w2/jLxXykX
YKByKp7Ysk9cTR5edc42oa//Ys31YE1uyxzDR5WmlNOQnwEBJWUOQZgPSk/G/09MnFuVr9Z/wv4m
nqsKe9YsfS/HqXgcOHS7Zfqd0m/Ju6/b4UcO2zZOvZS3EDlR1qBdQNbRIAy3FrtPixRTjMMUfViV
EeHV49qDNRFlIKfMQVyMctkTguT4xp2cgJ7pfpJWItBq0MDo+vb7N2FcfJJHEffuMzpzJvBNuGew
fNe4VpqDXH9tA6GTu3w+0womDR7nCiVh3pK0Mcwg1uCeC7INte1O3Wd6yvDpa2HRAib0P2K4GjMg
xCmxMMEV1Q+aq915qbfey6dsusxO3bv/TsYAXBn4tp7146pMOT4gAoeLKA74kCh95Us9mRtJ8L+0
3om3KdDBxa1zRiMOAq4Iu5xdR/ddbzNxzC3U8tfLWUZa6nTiAWmOq1CCmWvLJ+6g/3P8hvD7CySf
h/QG/NcBt0gEuv+RZowSm8vDmvBztHnJHheggduQ4iSMfWGvtXvSzujtIE/20E9xolgnu5QoUBC1
tVTUQuor3p7XzUC+Rat86U5TIfTStAE7TZiJedqBambTgD9gNV1G5DixxQfcfKeZ0RYSPSNBpmPJ
DgZFBabrd9IqdKuBOzk2JXdoz9mTdyzx8wFzZtjvscbsJs15/DnE0SOiHXsjar/TLad0JfBI6Fpr
wW4o9DvdNn99viRcwMbFKx7HQQMyrW9Xd1bwBIzexu8SzfORqME9WlUisacEPI9zspD5CwY4Ih77
q7uPwSLQv+1aBuChRQi4mDUQgjoZWvWzipj0beAcz5CE4todEuuh5jrI9ZAYjkZFZZzUgTvlcDlb
fc51micuyCHrb6kxcrnIKsLM7Trj8VbE+i3cmafHDB3jRRAKQmronlLOEOocNMvVEda+3taevGK3
ButVdqzW2+Jvw89RKAjMrSyRWo40PXV7oQ+ZmXS5FW4f59XpRfryeORqWrWcaohudt/ji7hmzZQR
dkKyRv8VuMQOEWljw6Vxnlw/x8Yy9fAktHpt+J9h0MmI9u6Gy4+ih8tfR2hSVVh7uzy/h4yiYgZV
iPYhhRHtUejG5JVIKzhp2V1nSmEA380dJjsG4SqDGOHH6qxN6SxZ3nJ96rXR7WxZ79WjZrHEDZu4
JL0N6MDroNduYWYByBYPfuFbseDCdfn3IVFygund6vYGSfu9aDWZip9V6zjQJOTL+XZKOFKV5pxl
GTBu90Q55gA+5/g3xEl5BAZQGLR/j227Ew1fNCN9aAN8EXTDlxRzx++WehXvA6un9gdB4yVx+0VD
kjYnCRZn0YwyLe4kVUW/uj3qKdEImJ+kKbszyu0PwR/IKaKbO7Qnt2nb4BJIGmMjr5X9cJYG68pH
S45TLr+UYnar66RE4Xhb9zFJCGaGyVXS7qLIylGPwXKQdwMn3iM6X2TcaH+QgpN7fbU6p1/Fculj
7WEW+nOaLDnVChBQbAYiqG2JC/Jct+GS9kW9blZgsX68kZz9HgnfoSDSE4RXyy7cK5o2+qf1KT6S
Z4s/COsnX41YkmnCZN4MYjRY88YleAFbbh5XpaR+QIRLBp7cCEbuQj5DY94pLlMAnb1WAHgGL0Tv
gIbkE36+D+XXtseDBCT0R+1ojeHC8tPHJHN4ap+LOR/gZIsQiDxm0TRL9FnFDSzDW3D6Dajl1M14
ol5CXNzOqNI/YEPK+bePnpn47Vg6eZM23Gvv8XqwF44Mhgveuq+xNfcNIRAC+dCWHzRHQAepqTcX
/v/JEegR85E6bA6XB2Z6+/7V8hCdcign5zGe7ye2RyhUvl+wqEJzRIpyavUChHjtSULQU/X+q5fA
1nkrfyDDhWGDPo5z/duxfWAip9nPx8eczVnhN7esmjRKLXuYKS+T59SK9da8nkv5qGuJa2qJ3Xbf
tiZHRH7Sm4yyc+tt9s8D/hjU8zL15Ey2XbmMVozMn6aAaF4V/GPNcqLH55pClczw8NUv6PyNcnJO
gt1iL+nh6AHY+S1J7+a6Q2wShCmXbGagKIumYGp8HffH4ZYvB5hHQ1m/ahx2k6pn195rYd31nLx/
/Y5wqo0d6BDJlLvGpkh6OIh+L1VU0IUhckDXonLsWZ0ZU/dACm/dTLDCEQpqgrNJqi3qVWRlrkkC
cpHN4rMBGC3TwQS6XUCojV1EzMzUbw/ze39itXlLTwwqNKDd2JEVpKJ1TXXm8FuvFLBrqBoNOxw9
DRf/uWds/awDljSw3C56qtWeEPSo+2STXUZYxB3pGVd7YBUoVfnkn6vX4zXm5PgskGHmjqZBc0mI
7H0QDGYU6HtCodnnCMJHVf6nV1Ioqz8LxocxO1pR6qEPaF91Xnk4mFppEFqUJAhrrRNX2zJuqSaI
QKeMeQWChtW/S186ygUU8rGIXWAv9sl4MZq51i3fHANnpqkxnU8AuuF7lGNUUzM4KZ28TUOg6KLf
xVVYlo8+/usK6AuzUWh2f9jahYWUHKU8AqMAnTaVoL8sMplRC1b7MIyEu9pYLtJE8tgxVuLGLwH3
VULRZgWYKhKMC/rPObqU2xsfQuqWwzccZM/RDyX+8WldEsTl0hPFPViSW2m+YROzvpC7wP/XK5Oi
Cx/MQ9UxDNJkm2GVDZk3OWN7nFY1x1GBZp3DcCI/hdJFGmjQ39aZzcXYnwP+UUUXf21djd7fhlae
VCiaGVve4eI/QhKTmUWHKsgIX1Ibb/gonH2KUOpNPOJwvcFMJeSX2jEqUUY15AxYFXCwFPTf0eTF
hMg+lDy2n+GYxSEyHdcTqGCDn7qrFpYI6yea57eMsM8zaTLUlV3cmG7F6ueR2fC7CUtLxsokHbcj
P2Sp3kxhMh6oYrJKuvAAKG/AnI5PM9jesaDBciBWKT0LF1PGqNJb45B7iWWsrvTjGEBR7779DrQb
HJpKdG7ITujVN2lCv1oihW049nPJacxMuqncBiqoRSWP6p3Ctb7ZsDrBVJ4b/5IMAMxwxVUIeMGT
8d73QJ9Qirc46SQEkUD/et71AMQQ09fplvWnQaZmDfq7iCwW26r1x8PuwsIRB4mYJSs9p7QCqptj
2qcJ21Pa918BUPCjgCRQFvcSdVjuuKSLat0IOZlV+83u+UaSvTsiXbB5mWEiGOYSPMe1SJBQQrgQ
SiNAWdh9MrQmHU3t83498nJ8a5MQ0UdXylunNQeJUmryuqpvRbcio3n53hfh2B8gc4duy1pvZf9u
l0NjobKppgg2kXeQOeVSTmQh38m9KxeozN7CRhKAptACvddpl7nbdQ+mckVXbuR9NT7n+SGOCR67
VRQ2LxQp+SoHBHLctnIHAn8moSHqzOcWu+ft0DX8Bq6lF2N4+OIOG3T487q/TQ3Z0KGTyDPSpihr
/fm9HhkWPN2FAqQLcRkMvU7RHprXeLgKgEJRfkD8Q6AR/poa8tc/VDP7tkJ4XQ3ud7BWVvTLJVVZ
7bk4tq3mpFbSZNEVvwM1xPt+7mZfhMyfw77Js+zMOzlQ/FXF8ihYH7FmllsAhaU9tQnz5IY7ShDD
PqhjzIMVRs4mYSF8C6S/bInAnm68Ny+3IPNKecB3j62JGZuOJwebkgH6hco5AmgJYftGa91P1a9z
7SRZTlu+vK7MlLEM+ici+nYkfAs3/mV24LXIMKQeCWcOtp5uy4bx/hKm29sTHzkc/OycjpkDMvyX
UcJd9X6oejI6e78kO9Wmw9sRyr10nflfc2bo+rdSbK4iLakAVwEprr5KvKZRTFw389s0pzgntQId
kXGF4Muy1xPrU24Ua4SdV5Zryoy/o/+P00PtxpxqDYGhy8bPH6zUff+2/HVjwQScqJ2c/j19uOBL
xQ+OXBHGlGwKedoL1xi+D069BhDIeZ6OiE+K/M71leqq2ywWzeaLc5ih26i5lOAoXwp2CB5FNKz1
dqmrNvettyEjWhhUqrLthPspXjB4/wqYX0RIK0L9eK8L8v+Iasv6Czc0WsNRNVFoHbziQE+cPSNJ
C4OqUBGKCzqKCllCUgeeHoxV+/uX5DolVkbg9qaRlIs5NHORsUHFHlwLYJc2VDudeK0BfT35fxJM
E9pC0LWGZ5wgfVViBkyhP65YpZkouC1oJDfqnPh1MxHstlXlyYx2BgcfA7v1ikSTm1tsSEYgS8Ey
7aHTGuVQCBNMOQBpfmYll/intrc4jf9A0s8JS8IKf7ZUXGDY1wiC8RYimCDAvOD8VsFm9f5g/GZJ
/++zygOhsV7nZvGo2s+yivzTlMVXgYGf74WEWxap/lAgDG+Bdm1nC8VP8Ju/U7mFD9V7fEA0DQyS
Wlqe6vi9MA63MrcJM44oqHvBbTHmEL23lqd19dillreSU2Lhr9nlzjVEKA2qfpmWwxxB8IsdlTUM
R20zBpL4QKZVXiGe97Gx7P+aCQLILPRx8lM60tkUbLe6R/mPWe0zInqjMmXgu0FzbSfK0tTFBX/L
NleBxLCVU4hywFoG929e9ElgGij7za4yX/d8DPFJ8BVfjnif833EYg0nqao8YimdV3C3DPXeIaCs
jIE181PPPOBs2m3KfhP9BVUvJ06v0zFPOlbco6Cfo4HtO6XOQNf3EVxdRk5m4cB8Ou1NPBnu9nfq
JG1OCtw3YEAWUd+pivQ+KbB8vduVhuEJhvB8GmjfUj24/IC9qC3HxAE75BU1R2JLXPM4kPS4a6ws
eMqtIXr2mldnX0h418FvKbQVSAGIpYIr8zChWNzvbTtKu1AiZcMEomIoINxHFJzyDOz/MQIhvWQx
boH55lTTd3mbsGpUDvgyVvtFTG8Ro8x+CQjOu8cJ/2RfBiynwxsO+m7sRUYPDpst/95PC1NAj7Zb
N5QnGTzKu8BOl+fKmfj4zA9Fyd6rlsGr31KkFOlQ0iuf42Q/OlFndA533tKeEa0KRJaCkoqKlUj7
q0a0YDf568bNzfH+YybtVaXabUDhMHXiNQghib2Tq0n3OAwW7lV+mXd0GVDPu8zwYiIYVVYlp+Sm
JKrxxRLS/SpOvkget5A9J/KvNnv7sfRlftzSIght4oMJj6colWU5Dob6YdcIfNftMFjffFakbAa8
Ugua2vdjs0xpuOO9RtmuUKxuzL+GoyjdzZG5GKJ/F07BJi8FSf3ETwdGsDor2nmlQvXR9ElDYZRp
57di3nL6XDfIUyS6LXqPL6vvQZdae1j1xrZU3ov7amhrsVxxQe7gW68f07iROt10C29a5yiiOAdN
gj7k12Jd0hZT2OMLBiz4Hz0dXPPye89k2lrx/u1m8efusctOPXo8NTJDtY6+Hv6KnOaKq7Zy2x10
KFLDxxNEQQLgVBrzZojHJY7ncN/3DJGzedWMbrkdG5x5E4CJVCLsNCuerGJqVdJegAUAE23ITjm0
deZTJNCvXml4tPfyCAMVyPjcUHserMQ60DcZ0yNNbbIPlO6kX/wrkDRAZKHycmg4sm1DiwumuiTl
5xV19kxg0b+s57BXjQhb7zPWqoMKQQCRm/IDshyFW8LDIp0d6+s7Oum9jwISf+p//15JpAUj8rgq
CTnchF3FZPbUWlrnAuk/oTlZu2SdSlvMf+ifrhXtDqmT7mEMcMQ93RvwCsUMiE5J5hk42eBhkaC6
gVe609iSYjZV3toPRo3Bm6KICh/HtjWZa4kBsmAjOjCEKKCKnAlLht1NCNw0P9nWBHba02ycyLy5
JbX0abIBMOwOoPKQ5ZUemTMMQz3WX8pOIbR4KMOGaIjwa7NlJPz0zBB8cywcmXWzjzYrhqkE9VBs
81WCkjBJX55DjwY1gaXbY2sAvJggnrIVVElT/U5M4rCbvZIXy40FcB+yUG2+MIWx17D0yz2hTUeX
QmCg42YJH0JgVyblylVEuHp+UXbzxAduOWfhmRPujW1KMpMeR2YN8/b07ERjqE05T3no7SwKfCiS
cuLKGofvodD+mukcWlnepIPIu4wml5BIoUGjuxqvPyb9GpM3pT3V+MhNEI+mYRaLc6hZCEkqIAmj
Gkboe7wHaKPDu+WDNt7UKre2R3hss9G2Q4XCTg9Cpo5BjgtcqZEeLzyhscXBTuPbtntsu7rz3ptB
tSOXEMWXTtrUSsOqK5jzzXUW64HPKrvk+80EVq0J3JVFXbewQpszQ+TjKYlDXrdnC/PveZe81CIO
P6R/kBijzKX/YbTYAgc9LuxZjUTcgVMyH0GtKErkPihye0pamRdeYNVaYGU0ajJYy8T5ls/eplxM
VFuA4FteG/RFmSNjJL7GbG8zk+SavLQ5UtN+oPuv+cXfuvylEP4FCCkweFUARmnEyF79ojV9urFF
e5ZXTT8YkYdsZH9V2lpI4j7a9utFE64hwi0D3TPThjQcVX92qM/36RRjqkvhmOyz5eWkoUk5AqRN
P9HlS1hCA654ygK1j0cLyiy/9GL4v7haPp7ThNWLA4rhF5I3sJFGOLfYBolaZH51QNLQ99PNLX+J
Sx/RmqKAFiw3jrsQE4xygpV0W7nbRZBdVGqvUBTtR6PehXE+RwbOqCcJYmjOELzpRl83FfUaYVQ0
PMoEzcBVUlTPOTx2XgS3CbrcDrzNtjQXkQMjga1V3eokrVuZm857EVf4Fvpl9DMKGa6fTiU7vQJT
sAHZc5K9ss1NPYVND56eAgagOqqaHUlOgQwbA6rsUiFxgmZ/irLfmsc8kJPezJDDGQtfn/O7ATxp
CmVFrWl+kfqpc6NfXNIcJrwP0y6WU6+SiNnpay2khw6S/KAu7sEQfwbJ09JGIx5NwRB0blQCTyhp
mbTmIDsmHmyrgtThw22X8gglKYGlMuIbBGCLjyn83VZ0+aSOJlQfhD3Faj8Zqp96y2I8aBYgXgPT
tNR+AljWsABvXZrmQ6I1/G+62UMTbsKXgANHFOfafJzUNIBsGs4J6odsIDJVOPxO83gYrtVYOlbV
+0vwPMfKyCtQQKJOxTiBzc4PqkWUpbNAOE0hgrGDLAkPRdaPAMv++pUPUPvWolMxPSnr/uoC95PT
kMVBxfzu7VANRtSIsJK12YcQ/1Z9OmZ3WYM3RV8WAkT+m5j0V1blxbiW1qLKdtV2jb6/M9NeIawb
K/WJO9sW5kLLnvJrF/tPc6D31/c2Uhs+0r1hj+GrQD8154pGJQSxlHdhar027m3WBwGQ0rcvOOwA
ASCx3gRP5HKwtywXIR3uc1L6H8i3lZYuZIsr8q8FByU+5eHuW39/evpAZ2qiLxJe3boCqpK3IMMZ
8tOtNjODrDaDnSDBNnyEQFKmucWz8U3QLmxdK9Gy232XJwg/yjzOCIl+ab9Odb+t3e8qe3EJ79Qd
jG2WEuz9rEY+pruyCCEJYzZdNjluK94maw8NvXrwgBLG2d+MGvlBvx2aXI0OBMzv1ODGfToAreak
HuTCjbOrwtLdgUsvWTWyUHUREqtgffEW6rSNUriLZ7+riR1wCWup5As8zBCdSC9bK650/V6WAHWL
HV3YuhayJ8fIfuOBfwO34jyBSAuPqGWXA/5IZiyX+JJ0SGcI0Dx7gqixJ/A/tLuRY1SXwAhQl25i
rDyqi9d/3sSs36UUi0FxVOXnRy0cJaAgnWqYcNblfxn6vfTLfQrx63cg1ic+/eWywJ7bCvChaX8j
BPNmb5EcTphOmpg+xyP6TPp+m2FDSAX4PMUdekx0uAuYV6RVS1K+J2QTjYJF7GIViEaq4Y0hTL1V
zVyqZg8AdmOw1VTbDzv+/2B6ZfQX+QPczZPfpzXQeXyGq7QfEJc/Kl1RLDvwgdP8uYOJl7m0dJVk
fo1610H6o7p+DSguj4dJw1JYuqunsQJCjECcenALDDJrnE0RbqO8oeTn6Vk0HjhY24r6PmGaAoY6
sLyRScRQQBIabrNdMzxRFUqYWFv35hjCM3tKO/l8g0XiSmiInupiyIhmGAIwSIEE8+apRCEyvIvP
W96gVnP3MduiyU8wHXrJ/sqo+Gu240yZG64b3LOpknRS9qLLiYvfOmvAPmgZroAdt27nl3k9KOkA
cAkNYPeX7rtK8hMeJ0DotENHLGjLPMr862CJgjUZn7CT9mFUlxE/7wZ0srlkMp3onClpQfdSbb4n
6wyjt3wrGJPT2sKkGrA/HWsA6C/7N1YdaVXaWKSPkFFxhZBFYYrTQv9ckhYSpJOQTddXNVooC/kK
NC3n6Wxy3AW+r3D/WdKvb46CAsd1lICyqw+kxGyIGzDllWtqFCFIW8UU+XTNUK3mR0KwEgQiswfx
CwtcBLTgt5KjfSxEWK06LxSlG6RvZKJeYhRLmOevyuij4t5r6vOoXPngNwh56tafIgwuONppiH3k
ayd05RldLXo/Su+Lz7RGNjd1SMdsXsRUuneBOO1Y2W4PMei4sA1V6Veb6QdpfT5i+bMNlFU12CAM
+oIIy8/XY6CQeKpVzz3s0AzM1FjNjZNTlVhwj7dj7FPyKw8dn1tQyyrDFAb0j2zIV/8AvzitZZwW
TxVdNnkfBrSJ0im2ThkqBzL2ElNS+oCSzy7kpMTp68AtjydlqeQPZB/F9xOn0MtQO2eI7B8pnJR5
xYmOmRJn6+R26leHWsmMnvGQz/pSCZ/p+1JsuLq7/vHeq8TiRfChgU+LR3GAb/Ag/QjFQfpY35SO
PsXU+llyW/ArinXnWF8TPiUd/zAQABEyj9ck+tSZu3LVkX6oe1nAtxyw5+6ITq1v2t29f9ilO+sO
GcCDkCJfXT9qtRuJ+0KLl4OTQ/xXXMJpRfnfUi5ZP2ojpAMgpvSl361OqB62UsJJvA/gtgd+DKRS
owfpomdPK56gaINtYFoO1+4kaiSha1h17q02W8O0aJVVZM3UElW9BcUfpKNdnnorunTxOtmtpdnD
3ZEj05v2KrB47FixItzfGNWy3UdUpJg9Br4l46C2M//VknHorEihL8ZHQPDnV+hotTtpDOarzpWF
v2aa6QXQBjorsWePbVCAGFUCPFPneDS2zhSL5yEXT/P7pekRbJaPElaqlOxshefr8U5nIQTL77Ii
2UKLBxfwO6+oIl5rCf1CIpcVrHMZwTqGOzsoFRLn6NMRTgJNova7VbuuDqiSQQPy/p3IbK9J6NHi
M+ocXVRSc2Mdzx5XON1Cz5C1qpBp1wI+0ZIHRCc9IzLvuZx1dWO7avbKLlWHsoRJptmIHe44bfzS
xApY2O0w133MLYeY8O+VfrE7Xxuldfr1C8b9bhJTPyVep/DS6zZMMD0XWEyjbLeoKTS+qIx45G/d
1C4koTkhYMxp1a99453XGH9pE2F07eXJqfmsz/ddkGVk50YI4LDi7eN0ENCcNru3HIqzqgiobjl/
gsD4JFtm1QtU9RYB4wUg44z/tnQvCI67z0PqTCPw0Y/8xORwn7D+bQTPoZdNao5h2SIQo8ZjQDp6
RUGqHW7+vs8Xr1vKLZz46CDjaYE/BUz+TcXMMKQW7JTKLisI3FmOzZ49zHZHW2jP+eqtgzQpOGrn
FRfWCt53gIrJnc5wCqln2b7okSphCqj7xjo4do4c7b0UDSlElmUVnFJAmSyqw0pBT+PVoamNLAnu
RCvSSdIG+En4r22gz6ClOMQqWt0ZpasZ7ZDikuCqk4lAg6irXpS58Dn4Px+utAHy0oQlMnPiNAc5
U6hJe2fTP4xKQ+LdtaDyWdQmz72ZqUGpu907MBVWkInHnkJoWxW1ICsBbVLXHNWNypBhn2wHA1W1
h5nryDEa9l4ub6WQtYPn3QotEq90AGrA00/AJZRK1d64FHgTuQTuSiCfCDNeBoomboMYhjRHcZB6
HJa9HJhKT8l9juj9x075Z9RUYRAt0xYzpcXS87aQ8188mp+npLAOpz7ngDvmrit/32ZHIr8Cjapr
H0mOGkd3yGy4OFO7mUNGjOVZuXz3XV6twh+NO1F8gT9K1udCXF1aDG3Vtopw3sug1v7QBYdkKuRf
fJCN4Of3fa+ih5lx1xk2fuFRzhEtnpmAjLux1H0FsMdAiOWSBryVoc/yGb/CM9w18zzhTh2oxBv8
S5C0SdooHoUMDBqVMc2oBWx0+gkZtafAV/njgC0cEnIs0jv4+ZI/+pwBhKXFou5EM5ZMXt9C+BD4
mIQrvNVfNpjKnau4dRoHAQPbQra9rSgoEXP70Ti4eNjUbSxgPeZmNY+LQgwhO4HVk6UKydSGNKh5
h/gEISB5QeA6/htQBhc+98RjK4+XZ/hONs/qQsL02yqwGDyjbxpIDvEQ6kQPlR8ZE3ugX914VeOu
F3UOb1wLCtKKGzd7iJlAPpOlTklkMUqWgDQpku463Brrk9QEnLHd8KNiiiRWi1PJWW5vJPA88z+K
R0YnHR7ejU7okmMFHJBdYnklFRkh1+rTmcFk2VL23qlNAiyhkFOjAxPVLNEGesMUUayZHNvf2lhk
senrNZUtu3G0nzbnuwTez8btHW7CItTsnQf6o/Wda+Df7s/w9zW/3aolQEpTd6eo6JEo1m2a/MzQ
8rF+ffJpcbub6E3NCGxXjIbeg91cDc9IbObByI3AP/lnNpJzvBujSPfVSFipuvNP45McUgfv9DMz
tftahxa2ULxpBqoJPb8eVG1kSsh4qbgP6WsnMPZpd24vtuWVsV3uw1/tQCLUojMMacpE5X87fsWx
0BrwaLXkeotl5k/yHmpfDuG1bbmNoYMzmAYMpceOZFbXW1IAnZouEW9q8W6htwwiKqYhEd0xRpuj
05gqjHfQFOdZG7QV9X9lGbWrSX73SGeg+HMtXNJ1ipDCwIg1oHDyYslbaD/HD7mgWfJ9tbl5P2gW
6vCupPGsAg6m7+UmmSfqe+Qgc7FxUnxsiHh5lLN95b3E+b1XrEPrbWGJxclV9UKiN9r5PjwZAgPi
b6qRqGCOcDGntFbKS2y6g5QQENKZWBmjwFrkhTmpDcXWAd3Z1SMgZ04FOvxJEq2NSqAC4zgiae5z
RUJ/l9l+qokK8P4G1AYcl6y/TRKvPJnVMGnwtB7CXM1SK4LVd6osieCm4RCOXKNjohLCiN3e5I/W
mlsVmSiu4zP4x9FdTvnj6bYTLkTEx4e86WfUFJ7zKq0yYBPG7tbe/tFsosT4L1GpLBm4OfJGQleP
32No6hZT+xFzz/zn10kJgat35Y9ET+OjUbO/s7zyEaSAf56pXj1oWwVqAENwAXosXwpEDDM+FWba
FttvtMYuZgWj2jl0N1RCWYFEKyz8awylKUjOX1/MRyxHWfQ7XB8J8twDNitZV2FQ0QBqUI3qn9c9
X+LBZrDHO8wG9fZVsNOAYpH3BrxJiupSEwSVPwC1Kt6efeEOFioGApeZJFKV2diDnWIk76Wqy9Xo
yp0GCTCtBQrVTfBmtS92jo+BoDAV5lddB9Y/Ei/WeDOxobO8T/nuoEjOZMyMPam+5NeFDo9DfuAZ
7V4Q4JTK6HgyDp1NO7p2X7fyMWAhIpjxnqtCPYrAk4zQyyXnhiowofPIc3hkV+7o0NarAH4zopl1
QAH3exRXWonPSAAZmD4VP9F+24QphXB5U89O600/ukndMGkIYNxwDGHzpRdNbs/qe8oBqn0CsUWu
UrjawyJhDPnqBcoU1iIwdIwJ+WhF4yMrVF3DvURZgzonK5Rwfb4if6KQHGdQ4lCr+ZYH82yph1PQ
EMOHWGbbClYX/nqZjkHlpSh855dGWQYeYEH8E4jbdpJVPqI6+r7LZ8+YrXHPzxciKFj90Cfn91Nc
/qUjmGR3+rZrnLDpRBTX7qKWdDL+M23LHw+c8xri2qrXclh4QXcgQHo49+GKZYRjiHqBeTaGoZZX
pcOdFL1HDJgme56Uq/mGKTyHi2tw5C740E1Nbd1YFocACe/dqL7WPdO8q9CuMnL6haER28cxwUJj
s8yvUbYQpXogqVfFdNDFrYrvrb2PtcU3UXkA3lSvGGHHxz4lhi49E/RdZ4cL6n3C04m1tK28+EN5
O9+9KP9kC+XXfiMhEMsC0Ok7VZrVdd3EeGVajaFhoX8sZRhmQimZUdTrD9qUoHBaLPugAErQsAXX
H76YsmuAVZFdJKv7wQcZESYVOBX5p1im/mXhHXb9NRuk6tLeHa5teaV0n/sK5LF/+QNUXV+U1eFx
XTigKhzNpiRSW0EMvD2z7MX57eFcJ2QH+ZvhHvpAMkefGAkysnzBqa0gb4buKfFQYOCn/OXfKYjJ
kxPcicO/HzapsJ8GY54jSLChWfPRdoQVnQVvppX+ol1J6w2susW/XQdrR42617x7sVS3WY5Xd3KV
LsB7bn9VXwbca3/QmP37JR57Xzzb7HvpniUNlpXPIYCQxr+FDVRHm9VK+kqnNGOLhBKMO2CuLoXv
jck146Zg4UVbfnW+NA3EL05zKLPCjqKe+uuM4XN/SM0x7ePJ/D8K8/cGNPMhmjAZ/C0dVi8MDBfG
yeFQVCsZii78NF2hCpYO43muqy61HbV7e9EYQyPZlRCKHbhqSjMdB9srp025JVjpbkI9rG/xeHTB
Ja3nH7J2pdwngqDqlKnZL9FU8mQ+gBqWkb6RjS57wjhzbZ1FX84zGrS2IVscMd/xqqeiX2iTaSkz
qenU47uVQ7CatP8Sq+Djg8XQ0gRuZ6shLx1tD8MOekJN27yX+1gfHNvDQEZP+jfgNA6PDWjweq3L
LmeRZKTopaHaZhj01+18MltpHiwWbnTrSk9Ep/qBtcVduKX4uFaN2llKjnhVikiWobU2pvit70V6
LoUhIJPG+xCPgvoVafs+WaA7RyV1xnkpD2EKz51vKTiuSR6UXVE1Z9EtVW6mGhKDSEdtc18Mk84p
wIXloo7rMMenC+mp0ljD+9ly6G70SCvl6a9Sl1oT6BHRPs7urTm0LqCGwASTynVzKaZoYTaVwDct
BxHGD8Y54nn3XJDVUK37LjnOTsV9h3agI47a5GY4Vq4NcLmVAyKEDanhp1iOJ9qAdblEtsmJh2Js
KPdE6yGDbqoux9Nb7Mqx4rq4jKxbo+l6j/1q+DacQbpfMCk1CphMlGOV2NMh+m2MnPTG1gsrESf9
eLEFhKwR8eMpM6TRrKbn0v0cbLpgUun1FIEeU5+4IpQbhnzIsLFUgaGwYPz0yDq5ypXM7TfUBDsb
/EKjmHwukrLB0pq4YkINq8b265NcdzNhYqxTERLVuEBKYw+T0QGVU9heSp9sCnYbLm47j2k6Gmc8
032Q7EAeBZ0FwLTnWuyotvUjPScEFj2S9vEnt/JB65TB8bIMhvszeW8te6xDnmyYSgxLbHrgLoFL
LmUBsaOhCa6iQ2dAEXVov5z22NFLpP7X8nDezk77ZjvzwgUm6AkLSxJNezwu48gYE0j+WjUo3llb
+eOYsekXSMxc4lVF76SF3WgUlOzX1B8BiWl/Y08psPsaNHnJGl7X+j91LV2j9tUSA0kZYuo0Rk5L
YMoZjdUrDR1OU7JLSs2NRx1vmm/er5yhwpobY28UdZppBdIuHadI8WsqTufkpPF8MXN/4cTV32R2
cJAmatp0pfEJSAD+uBK2sslsmoERMTkF2klCrBjrVMS8HPVe7BBB5lQ0Bb+yt5ctQOp3H5Flft6z
x8Zy0tBaYXSrfjVUc+Vo9E6S3LYn0tDZ1BelDj0zGnNinWZikqWjxAtxaX9rRyQneDFT08zqRUGK
0hNQ2fYheNWqTC6jxrS71QsN8Irs93RPmMgcKis9sSjEYw4z9cgUlAOnMLu2PW8HBw1GmkTFwIL0
CWwi4YnFlImo1hidAD+xywwYDmFcXV8vxW/+deVJJ3XNpwG4WU6BvgQg/G/4goMqGV88gBMgEs3a
BFMmX+6p5kVrtzHsOu9gi6L0k5lI18Vg/nPoo9kTFt6p6FeInXJx+1SuSAcKFR3h+Wh7jrsNwnJD
IV8qdpHdG2EzGE0usneiIYZW+61AH0ISX/euqKmm8+0elZu+tpzAChvA9pmLvavs3K8TfXaPtZSX
38PaTwkWo9UHdhDnJvNReKRRXcE66qzHemhMoU6I/bvIRNoP3PB0PqIlg50ZMw6iGTqOzvItSH97
A6bs8edLgnMyW4WzbrFCAvFaoraXBLlpXkV0RcgEFFgwiWkC4Q8PS4iC4OK1kX3QXhi4pMoBqwTX
1QdbU/sZAG2a+oFymlrfpJNi96sQN65+/bNHpZNx2lesLC8ZML3pH3zYS59dn5EgYLdI972/85UW
8BjWsmOP8WIepqF5lRflVp92vu/sRidYaP0caHtJ4xEMDRybC/QzxWgcZ3e0Khnfy5lCO39lEQSx
nfeT2hGEWC2bjDK/o7CwJAzYOTSGRYy5NkLPTfBH7U5IaFGb3TS7cXLRUAbmuSngGCFE4Io9kN1b
KMAavh1iLdqZb/vmiwkES9n5dje2qFWDZjZgLc8+It9RmqKUs1scfvC764tFF2YYHHU8aKQM7JNc
YLuy2VAYj+e1QU7N746fAvdk+OUzYjB4VSidSB+5UHqN6uOE5Feb/L/7cvcsF5AF+1wow5CskuF5
X+PxzCavvWVvKTHjhHc79f2G+qlLExc+0fHmHbYtmSLqEd1fp6JHbK0noKB2qeeEnm81yckk6Zq9
2WclgFQVmWvi3m9WIG9rbuMQQ7BfXYfqimFccOOfcRdLu/4KYGabij82nuSLPC9I1oLz6K+lTvId
UOkn+GPpYCnaIzEV9rJ6ph9SWyF3bkdCPXLD1aarVx41qlDy/howRpj6f6N+IjPPI9T4tc0e7mCo
rZf5E/HHmYa1q9HRGpD51WydVA+emB5WVrXG0qeoq4ACGOMvN1J1UnjCaIIKOLaFE5EXDiYR06rc
dwDWbpIDa0IFwDCi75RyrIFFukE5u6Pke6RnTEvB71SJznjn1Pyp1+KMrcXQ3uIiPCcn5xviVin7
ECy9bCDa0eDdDszYoDXg7Xbw/Y+qyB6aPB4IqOv8kRSqSopqbrYd4wfimIqSCSQxQDqBTR/CfxSH
rl15F6o57KLthrQkdweF1fl2o7UFtWiDWWG6Blzk6DVXuz7GxnEe62aDC3DWoQt1TviO10iUX6gz
EaO5b7VmkabxbW/FaKeWYhWSVeiLGxyTO95ykYIfVvpyQsQw6R3g07+860emQn12/rkAuN/C1enb
Pj571VAQ5c15ukHlkAujgLX2uWmA3EyDXB2B9C13J3+vnKKEBJJL8AOy7wpmqR9aV1VYXmrmHBJb
76CTGR12xg48/ytlPNDlN9B/TjbJqeRzajit5c83iHFXyZdnZRbnAbszfSerJdH0fwgh4p5dnmDf
0vu62Ny7U1iX94gofYCR5dH6mTgJT1toLzNwtgmbokcwfR4K6hnSAnQSiC5aieYwvsfeDoa9d1Tc
3JA7NfNGZiR5N5JD/uvfSYcIfLQR4f6C2KpSXzpe8xU773lqA8mSkB3uVRg76lIlgJqgtKSSKQgz
ufQ4zgZsLy4F2UHaXP62cFOUMV0JKsaXHHnnQiGnI/8l1vF9NXeSjeNXx2wEjuA+yxVWXvbimHMA
FWvIRu0nE0htKjM4ovDBWvk+3nnUb3xqqvQHBznkSbq46AYVr3/G+g0DBDiNvb34jkQFvde18OEn
0WEWc5PquTJQ0+Lw+Ql50efKwXOHyDLLErWFQGR0uZqdEk1tGzbeilHgeq9Q5gGrNGW7hg4zv+Ix
mp7e+evIE297R0aRIGiyw5yTBaoxTxDGvJJanBdlLtMDsmiR1W+qMsduDA7NFH0g5ZGGBRZEpYCX
u37jJdbg424lfpAYR4X9JgCr8ZYqdDXLo4s++8pnNhyYIjOv6aBZxZ8Bf2ftKTn40U8PgJrY3gJ1
Ev4X+aGoKxln/iqrumMBJiEQ3dg96kWvC0DGprOUPEesIU+Cu3ort7qbX2bSbvxmnC2Bbl48Qq8r
yVq1Vbb6az06vGgTGor84jx+uI7Qngn4RupqSeyoNlOiTZaamtBKncs5dD2eO0Yiui6KZqfqzcV6
xk2yAfQpRbl7DhOI/kdg892DJLUN069Tll1n0cr/I+jBhmNulx6Reys0xHS1wpZ4gksT8KoPPcQc
+P44mMGwXH+cF4zDLI6ycwT8AVCVNjQu9IFGHlx20ecMbbXZecqJAzL6T3AbEOLVwde7L3v7tC5E
pRyNKEz07zTWS02w0PqYMHzqPWQKqmvLjJTrSzUpCEY4e1+LrgCMq3uMKnWHQbjusrHxXdJBtSvJ
GPTSKyrdrGkswVyWrdX/i01SvYSxa9a+aQCIiDOpT/n4Kjkbld12dWhHRwEJnm0IUoQdFnbJcPf0
3P/rwTFTM6zT4o5OYSAWK4UBLTW+n3s7uNobAH8t2DXTHLxEcQE6T3mCq3aSaQ+tuBMcA8B6Ogt0
bQany7rMcJFOS6P58Mwa74/ZA4rkHFusIrQH1WV1hT30aQM0A5ei6vGGCs7WwNVwI0nDPR52EsF0
KjMrk5I/5cjd1hnmEOav0hY/3gvk8XVQlFNqyTCvERKpEN38fsROaYfIEOyJUE3Z9zm88vITmQrR
IxFG3a0ujwymayuemPOfqxPJVm6jcHh9dp9HBRq9rg1gmT+j715zvdtEWUllUiy/bLJQ9OMQq6pW
CFpCRsEn6YwbcSLoafBVhIsobYsEnyQurL+FUk6+6VKfhsJhV5Lkt6/7SL6/qAHC0z12d4aXhHFN
FRtOd+Tfux3Iu66eOEFLNF4M4MPXFltN0TbbYKnWp7sCi5Uo8/atjmVo6g/STpwuFQhlFuWgUOxf
/zoW+KcdSqWSfkO37yHcaHsN+VMCg10UchVpcaaAaE716QW7XtNzcUETFh2EuAqaZzjJdNO1PqLn
2YfD9P56tUQbvG3TKv5SAEsCK4ZcYDi9fWwlRKID16wiscPvckTQ43pHIbmVMKxHa4hueEo+wKzS
6/L6+BUQmTO0vFDJEm6u3uMgtIqLHtjIqcHH+BKsjyFLjIPQwgUdyc/QAAPNgMj9cEbB/4+dknTZ
+272zEpSoMFhj84Fxo6qeeuc3o/vA3A5YEeUel6rR7ry5CDHLDzQkkQwUHG6OPgQq7eAzc0irrh+
GLTHstxqVsdW4ZpolhFRvEzUOk5KUyebe6efPlb5lvjrBu4f50p/lsWF+2sQ+rO9w8tFdhsGMdZ0
oJw03ro72wSlcKWbJ48996nd3zAs6KUw4Xh2Iuwyl/cMtPvlmLwiPNhYhptlWiD6zgT3pTESzZz+
4VPBcYpmRl+Sqyv7fofc2P+lgOV3Wgpqt0+ip0pavi5IVz/Xrr3NLIQKtPNpgQttQzMwVE9HRauC
OgmsTjEZ/yu9bvetij9PlAm5uYvFomU8nQB0UatY3Wm4NIyzjoVX2vTiwr0sxVmwIHAqkQBO+oHH
olY+ZxxXF2Sf1nxPboAGD2/EZVCC04jvlJdzBO+kPB+vXBp+u/JTsiVHS6m+xT9qBDMW+11cxoAL
VKtrExIR5sDx2QatrqM3njtrHcAETNdy4z8EUpkUp+RgeksCRc9dGxQHdU+prXfAdvz9LwW8z4oc
VwwCY4cDrxBg71ZDkM3HdAXm4NcDjzq5y/BfsI5uZ2lXUlomR2mtb7YpogBuzBt/SY/r/nYfqWZo
wGKYOXCPY/o8BGyzF9CJlb1fqrEXK6qhslFAuy6jl5JC2CyB6kJcFksjHhZxA0jVbkABu5LYYned
KYPLYr18puZPvB1q7vxWLb+eM1WuPFGsJLyQtSUPgAyUScvUzCIHfqlo6pjN8f/yhiATpbEGhLDE
sLP9J9eFACwlZdRvgKOXg53cOtmC9vekRPk/ehAhqbx+iCOcdXBABKjnmumvGZNuX2r+QLqmFI63
DSns2TAY/mVEZBWaYSkHQAyqZdpspKTzStQHVs24YtgPLN9cPnwrmYojPMNcWlICfClkUeTa+v4K
4Z/mhlwfuC4F+is8FmR5g0SvAwQK7HUDcmgDddL/2IBYgQbPZAAKeeq0I1Wu7cI1Egmxi1k25WkO
eGobBvCc3J1G9c2bta0L0Eicr0QRqsrIp54d2abkz1JBFZ9f+opXVBK2M5Vb2JvXRC24ot2L++71
zYZ4lfcyUmv5S6ggxzn8xk8w0/6XvOorMT6MamGEY/LqfqorL9/Q88KLwa6KJAqbxDljdKWV50WK
GeYWIDdTLB6l25vxZuIlG0gYTujQYp2sfW9nXXprZpwGAe7eidG7Z9FFWriLXpxVq+JjWDlnQ3o8
r0twhRprbXyolH2BrcUUV2cwiGBGoPZVl2opj9JkkS8xETDxFOUATXBduB1211scHh26NNL4ObN1
2YsWiBYA8JOE/h49temgRgsEhiUpPObLJeptDHoFJFhTJ50XTR5dCgPVk9FtsA7o5sMYw3mUX3bY
YJPFKwiP8rAaSZ681yRugxNMENZcEMl4RvwuFkRuyPgMkrJeR8F9NsdX8njow1i8PUyst9gY1q6x
/+LLnf7CtqkKsPnW5DI/MU0AOBIkHjJNpPmJX66qqwGu2GuoI5lX1UJrqhvkFNMNHZJpSMp2cZLg
mxVsaS4qj3wCuAilJMdCLLNouaQ6wKXdHOEID7nc4CczkrVMkimUnzctMqpDHOOaYatbfYeeLTRc
PlgPrSVWWkGM+6c9GMo7f8MOt9Qe95ewaJ75JfluRsjI9nITvYwFJIRuMi0d49iTgz7SR+7+cepj
4vu0Qwuc+dO1QP3lFNfalx/9fehiqCTvQuyxL1QNgEsMwXwvQ4t29IXeIXluUc8tfb0rS55I5vGs
1IznXAMWFt7FFfF8LMI20WFNvqPbOwgFJBcWU6sSsDBsYo4bpA6a1qp2O9qIGjCoWz0GwdaQaoO6
MgOFOuAe/xovUEkFuyBWEEOKKYxlV4+LzsvRJb+6sqwTO3scoZ/mpwht/8dJnaaBUfk8lzDraJ6K
tE2TiB4ZObFdE84/jS7AjUQd25BSzyRJVm2lIBjP5cS8q17WxOZDWAlsQN0dhis8Ydt8LPgcgtq+
EqKojG+blB5S+TW2VMdiezJBvJaXCvTxMQEykUJNByLv7iEpOWGfVW3XEx1zU8cde+3TzoM7XNMq
Vx17RYLOP7kXxBAStx9for8LXsns+3ymXrU/FXid3VWw8Zx8pF5jHSo6L9gjj3KiJ+WOZflu3/J0
M0Hr3qh4CAqTsIdbx6EAkweZmUk1Ee3/oUxzhRB97ybh5cJILxdhi5Wo/tqi9bBbAjXEDgR5pS7Z
qLXWX9Uo8jKJLti7k7L8wa6q9+xxpkeYB8J2RNPJVhjBAAsfQbFfHyaqxDjRFw0i04/zUqoLE1aU
QbXII2+ivm2obunyTTDWuR66FSHD2D/R5JqWtw7S6vIdcRg7GsvSRY9pSKCaWn6RBL7z8aCUwS1e
EKOYtYAQc4Lew5jluxqr/M9zIrhtaNxJZP5Jk4Ubef03Hc4RBQvx+ZzbbXJ6wqJBBQHrBR51NCQl
RlUeRigSKvI520qu2zfKbFOezxbPtZIrNFGOxUhb/lR1K4rWOc30q+1qFByUssE1d0dDlUaOCjK1
/Y7Sgyl5giq8Hj3wHtHhKfFbM+MMuMnDLPPcdl+r4gRWU8EBR9zW2fGJQ2b+xjV54Qx/vBuyO7qa
nWGA63SNMi4gGWlK8CF6ogIJHQ0zxEcqxisPZdDtlepXaz8boTCxjXtu3K98NkorAw6QxJeT8w4Y
R0uHK2yDdV5hZ3KYw2NoW87AaY93299HFpu5YndLAQK27Savtsg6E8I3n1RJhDS/uFQRuV0PROVU
9FWRHEhJFlUENJoZMPIkV0OorSc1JeglFpF3zw3RExXHREEhDxta3zsDWjTQLN8owUiQL6pEoXzA
hb8Ex5dAaJjAKn7ypsUMqJdj1TPGWjGI04nd+qXfBtimapudY9QFp7ZTjmckG/edu/LAJhnDg504
D7bfV2XZpOsmY8uctZW/jDhpqqIkqNhgeGPR6TcRmxdNkU7CLOhFCt5ShjRuwalHhayQd/5NeouC
fKJAD2tFgo294xXmUHPao2P5RAi8txNZh51+8P39xW5Soxob+gTBa+i0Ox8wYwTgWWHJViloSJWs
uy7dV+SwhsnlGkvd3uZe0cnSl4ARDpTGl0jd5QYIEx4LYorkJPOY7uUAANrlvI7n5g/7BdHPQXcj
dTI8tPFb4YsIS5eGAKYTYrJWWSPkTDNftkVL3DrCa4NhcBG86swtw3b3qZ+DrU7GXF/gbcVDr6Iz
xW6rn4+UONw/16hLmxXMWRJ5oc3RkJpiScQig6/fGC38JkaGNLY7eUDcZ1fpD6EomDn4RxBvzv0/
VzqPu+/R9kX0CC12qPSxAWV/WdPNeZ7A4wC3AhX3TADFoTWeM4DsLtUzGUzLde8Q2fxlJQTvBXdk
wJLtgfw6Ts+Vs5Gm4+925d57kPUs2HOJxoJex2V5Q1Q/+gRHY1ryLzfUttVww0YgbBRZIYaLQIdY
rXlkf8WTANFWtU/h+z7hw1YpwyUcBkWevUwCyTz5xi5qMyk2o1UpBRUdUr5DPJcMYPFFOJwTcNqB
NUXOL10CALMn6Rqnd8AOv3cIsoQ/pV8DNMXUggzCDhCd+fmuGO6UuGvAe9VoYEeXiEtd6X706H7I
0VMxEVjb5yEENWI3TakNVm2iUDIP+p0+GdmXbQtvNimAgRxbE/hVWAP2mlVqZzKsqX/eVpD0/Nvd
5YxhtSBv9fPsAu/G0UFoTTOUkUqbfQUToac2mGEGmmmKozq3OJwvspSuZ5DvmfFicdaIKbHXywo4
iPILB/3VGuXIBrU4cpxvJgbWdL07VsgXrDSvN+SkNLHLRc5+Lwrji5bDjHpVFYhSJ6LfF63ogtya
ftnN4eDcHI+EZNEaJPgb3DhwPK7XeXBTBg6pBm3g53ttv/0vaeiG9AxKubXBT/rWEHWOe93y/XqS
+agQUFYRQolPOplzWQYLfe/Ygfwc4LcXzYjb3Dms+hDuyH4egjOYTDWnXTkrHqZXh9ualYZqt7q1
3KIca1qZTjtzXdPiyIBSsWZdu59XR9iwRB3V9c8cvlC43HTACiBeNKKEAtZzYLMIV913ahS+LFmH
xmZ/+Vvg8BnTFfGOPHX+H6VhxFczSimVtMUFbgouJlLNNMb1ex4j1U3zh7/Oc56l/bET5O/ywHLd
MKUeRRffz5mGohSDbPQKjcQgRMB/PoPD0o9q/ZJFHWSs7A0jR0eQfw+GV9jeltfyPDEUU32B29i4
wmaq6O4VXokqt4rrMJlNapCD1r1gm190Ysn5Lo3m+PcGFwDp+O678XHMEwnRGXBufwiSw+9Hbm9f
cpZyJYfI9fbbPh2ZPT3QsbhVV2KlIERI68hmMldyfpa/EMYvu36FwSbkkc+K2faXEdQVhWm9Y8S0
NjNYlg/O6NMCBW4oKfMty75NSosq/d3UC2Su3AaT7wTQFIDct3TxlULz7pZp/U8mfbAZXLkGsxHy
Z1zFGdUxzTuQz9SM09RrWH+j/tSdjxetJwq1QdYrRj7xq6BBQgG4Wk530RzKKMf+ehhCCwUZxIwD
w6/PyTjqRnNFChFoigSlz0wG0/+rCBJE2v4RbCj2cNoH0p6GBHEQwXfGMWnF8nL+lgmTxds5yr1G
J142BQgd/1BQq0NGXjatKLzsjoQ/iTJwIKE62hJXnVmG0Ces33Ab/RurHclQ6+3Fmb5aJpwe63c2
SBbyKBDWBsmpNxQCiqoNHdfStS8zwp7IwOvuL4pZhwbkg//GAgvIRM/Oro51K0zI5DEeFqlukalS
8ORl/apJuvT11/Pm4UGFfck6fnWCkQ6ixCnVPydzUdfHWUxe3LHejAZM5eB0Ae6k7PF2Ual0aca9
IxfEvg9Cl7M42F/4XiQhpe1BEzhWKsfu+IjGOKCDFe5DSoAD8LIQ1Yi7+uiIty3N5su/2sqXBxIa
7OAt+PWpUeZqY+5jlmDEW7R75EcT38ieRSJJvy44oSuurab5CBwYxkhBeS9Wlw61fpG67t4fty8h
nZhOpJWnCjFWFvzHdLKOadAUGa36SxIuARI3ZSZa26qy5dqVu7Uwdk8y6WxcqLKmzA64wx0TOsyP
rCg7gbOfXjHZYjf59qs2IJsZ2bqJ73eC7TuMhpdYA+kQOiWgyUsJKozrtlYoxCe0tJl1nyI8OjHc
yLo5OdgXSzFVTFvdPqDybyx4TUXFMTcuqdBpRnLXyum3v//xEjvsoPyUZZ8/xfbFxuo6H8OBT2hS
YHLVbY0Jz2t4sIg/XiiT+ieIJydVNAoZK29Qb9uN5cSAVPJKmMCYy3B0DgJqKb4/DgubEzXAtWk5
26Fe8Wfq1PxrI7mKP/YrTrRuGgQ9vZ1aId5DE4ynrcDlPVWqDmUijkVO1av4eu0thDMZaohY1r2g
YDOOH6kBFUsgai8zcx54NvYR2kuSmdOIM+ewKhpxFQDLkAyBGyZTmbOQhP9qtbDLTH+r4L9esUiq
14Y39MoFaTi537Aru27zFBuwydPBq2293a5nGaO/dNGD+dizE/biBZUCWvjPxpLBMhJkcSWfTl58
Tg7nVFfOpDPtBMw57MgFNrjnFgnEeuSLPNr0TRZqxh3fnMClpHrQNUr6igtqyp4UkbzZ3V5RJ95u
GCplfzwbvhBsM6jpMj51GZy+jWjCdIRnhNb1rg8x8G/+TkfiKqCmgTomviDuusLBh9+vBGnSSkaW
a1cbIsHoO1Z4IrMp6buXmYTCCgowm/+hNKlYo03LX2jBPOBYgKDQ2Js8NVc/tipOxGDhb0KPAULi
sWCxQ54bJkscSzxPCECyHocaKiZveEfUdGXs7Jm2rZyYBUzFlEQkGSOCd7M0790uRWzrXWV50gZx
2V/u8vP4o1DxSWtsTRG5dEV7V4y9vY3EOf33+STC5f7fQ01ULB11ODLUDrioQOi1/FTJM2j4XpVT
GEmOF+tPaN+gIHOY2Trv2KOfVYAcRndAKZ/On0B8nVrHbn2j+shbptWHmvidTmFcBbytF+7t5gSJ
nVaNScW/TSzLbz1b5uBV5LF+7qqOFMhsgI+FuDzMH5pSs3thfIMzosLsh0ERDgzHe8cz8hozfeta
DIdJNvkLeXu+tByH0KWu1vu+q2c9p0fI7p/PT//7HStr4T8L+gYLnmOSVR8N2lKeS0skd980oQ8u
/LdDwDJq/TKzpSRDgaFl7lugisi1xVkISyHza4Uago0PRXC7h6zgRYlozg0GKxVt5MpkpGbeETsT
uTl2Lh++orhELUUkLzgFkXkHApzMssT7HkgnKXGgWuMgvSD8zxuEEhdZEzZxsZqWTLuEY8uH7Sp+
r5VNpRfrDO4w9d/jYRnWE4d5hhK6fCLEFJ6Zp/8aeSpnaeLNTBaFpC19JJZ4Ex7j49IfeFgAPpVw
aLm65wvi0GPygpgxnJSj468NpEEyimnl7EcgU6tLLp/PVQqRfHGyQMlJpfKKVyXlLdSAdNaSG+tk
xIk5N75GpBY2zom14Mp+F/2pbexGCzoqjy2aUyNaoxBy0uP6J0kR5TyaOW7h2I9QPICjyh2Oqs+n
YWGifpV7mA322hhtmYNqgvgFodKcC4AfNFQ1Ce9WEH8f6fCxRo5Q/UhQ68BP7GVJHy40M2WmSvwm
LqVB5dP3l/pCtBI4hHrcTAa7UrsYaXIQTPqJl3LTD2cvsAnB34yWmqJG/3eHOMMNVUPYyOYFoXfj
NgFozz6+z1KA0ZYuozDlQJScvrmHa0/qfMISBd/+qmxcN6NBbf6lGv0Stn7tw4PSsKPqTas+Y5Zx
rYbtMqHLejdkQstr8NH3ZeRoJ2zft/kxbN1RA9+auV2I+FLVcKyKQJp8JafcF/X7Y5pf5WsNh4S5
RQ9W8/FYn90Y1sCSZ2/Jb3exoF1h2/TE1C84hfAYlTLjmnbMyxaj0DevhcHW7nhJmXUdoo/oZWsQ
YUhK/zAFINoLxujdCcl6ygjY5JAryDsqq2Xcct/WaZAbmoecoUVCAmm4dr/InYvoeORV0fEdgq/s
D79gfqE3bsdg5CtGLiS7U51Ej2c1pcRs03pDmqFm3oCuB9HNI+qtb2dIPjH0Dyp4e2nus2C0G7ea
26Fzry+d8UBXFLNLuzIZh486zjG+ObAwIUpavPMN75BCq3oY4/tmZhLaBySBlDrEF3BxTQDkeakO
PNuAOXkun/GJZb2Ft0TwQG9X+zJxZ6f9/1PZ0QqpFig3+q1gc0qaiX/CHnlb/jg2B89CF5eUSz9w
TKKLjH1cmTEigNJtdKMkT6GluPXfWEBvF1isuxsPW9e1aXb69jTvbN582zSPm7nWFPzkajufjrPT
pnFazDUentkGbXUAz5NuOiKOiJg49ls+nFdjvQ2erFs1LOmQY+P9Vk4epQ14WAwUUc+Sw2YZlAnY
OHE5FPZXe01z5hPhviL/texB0/HQAJWQCHLzGBsBhYS9537QEP1euXIYC43tUEjQQqCOhbiGaW8y
J4QE5gmNT9UW13jDKEm1MK+MREiBHsHJpmjpnLSnWAR5esDuqR7NCnb/9O3m+7td+okg7A7eCbik
+ML/50PqbmkdccfAUZWCIJ9TmS/1oKyEToG43U7zJDlTZXoB3Vp7oWvqmql5v63WaoThCMEz45tP
gzr6IvenK8EdoVqCHd6uwFYPuvw/hLnH/Wznlv9LHggs+ZaVUwFbc3yFC4VdjEIeOZVTBHhBM9sG
w7MV9A3ZvaYuGCrz+B/xePJQ9I06xLSpR70lYldfUZyIJia+f/zI+DAPH7IjvP1FLouM9ch8HLSv
Mah47b+OBy/1UwkXxFK5OYyugSX2W4LNfbhanTAAq/zjBmT/o5Qu+mkU3tmHNQsr/y6YCCD9kXHG
jjVHcpFe0wz+lSgVRTUgHp4dZk3h0Ogfi0YxwRiGkJB2hodE82rmDi2yXDGG42zwgS7YThNFSTl1
LKSC6ilZjd+RfmK5mwoXIvx2ckQxpol6sj5NHjHWxtzHHJqjiS00n/prQeM6PQko6pJKB1C+n8+Y
wYpeNcnZlnTSW/KNYBVjhWo2UsAxisb1fJCPDAxuzjlHF7BSe4b8C6xVcOK1abhm5pMdyHlo5Vcd
VpPZB5CgrMaMtuUs1/Ncbbyqh0hfLVZFkKKrgX7yorcjoQh1QUcR/LqnA4fLsZ7xoj7K6tt9MT08
UhZDj50I4k73ZEO6UfQ7M9gFe6IIjldVuxrQs/7Xq/UftR3wJSIgPQ+7/JkyNQA2CWKhmBWVo+NE
C0VDnkR+njSf0brPvl6oPNcr3r1PrHduE+JlDIO+pMB4Jtewa5ilFWM2XrcZ1ds0asHU6Tb0cerP
atqameJI+LF8EVDkMXtu6hxvwbmiWZeb3guXiZzCAziG6yw0+5nx+zRyhMDpGbc2J53nCRQdRoso
a+82kBkvBgcy/7vRGef7Xw/mQU/2sUueWJAPEdOdUuozNKt66PkUQ76QFp4z4kj7S7GvJO+i8qyG
WjjaoICmMXZbJQDCq28EdeaWDkxP0U9P2+p/7eMgCxvDORFCAxUG80LI14S902Oioe2ntMR16omV
4ULgKfne+3CmhTjsA4Oa2f5dFVGhgokqkhnSEOlymBdadQoesDjWj51PryCWteiecUDpAJSjPbi0
Nt0qh6QMFtgr0lIsrpvpZM2ez1dc8cl4s3J2FQTBL57o4bEeInVmr7z2kdbNLPUxMw6vwqbOC0pb
I0vM5KWbEUbn5JRsFYHmDD9TXTmQMIJeK4nxHSUxIxvdp4RTtH8CCwZgTooFhmzda1zCQkjsN6sU
EQ2UwuTTcOXB5qvkz7WjGASySY37QB6U7zuHKJt/do6smCX4YcvnfGJOlFv40eR0g4pVAU01FJu1
ajHcwr6CJQqqqUWNiUEsaUSADkwP312yM6bHfhQdWcZ9LBkL4enlpVMl+hUv8+I2DVDHZ/DuwJld
qittS416K7NrID1gU1Mp+c2fyPC/rEvLu41VcZpYZbj+bsewluVXkQRyIyUhNalvgO75h7NE7rFB
yGEsHQ4/OHW5gLUvAQ8NE5Ou22NSKpdqiwUENTyH9CuUj39cWJKirI+xyjnWrlSLyCz6nGU9V2Ts
s+xbdgQCGfkj7/DLZqjXWslG4Il5SiU+WBv0jwWp91Ls/yfh8HxSHHSdkM+QffDOgi6WNgJKinck
F6LDjfRMTUoRNiOq4vt4WJyPgwwfRugWA0LfGRnXBL9lyW/avXGL4ISygRgJj+ivj4AjMRN+MI4+
Qx+kIxdZoKJoDtGiCfYdiqaqvtGhEbiqd6FjTQQa6sTedRfL0F+5LVeXmqg9BOCcs+Wb39uMu5sD
FEWRROYsYUKQr3atLDK6GOx3scHmHEM3MdQQtS+aqy4nHYGTPjamwfB/Q4ACgV9XHVNmsH/y0Blg
eYOEH9esr7AhmXnl2rO8wQYvgzsQpGqZyDHXrfCJeQiQXAZt3Tq8FMh+A5Z0jGssnU+X7/AMbv03
jadOWGS0++kMGHasiMteRkcJs+2/y18j0lGNsOMxN8bx/oQachZoVPhY20zENONs1WDokEAK5C0n
cYg/Q80ZEoEe9GpDht+Lnr0JJSP4lCvjgJw0R7+SWZX+WqSCqHYt+20nriSalPD07bMQWYQ6gfPK
EFXYObRxt1/4qosUVHzFYGqDgCWgP7FY8hG5fHDyZG+8rFPfHNNVXQ5nTXpmn5E02tWtKzpDKbxl
mGVaU21tX9cbskN+yCkibj4C0vfB7f05FcfT/bRkIFT/I242mVlvEU74KTX5eaQreusKQMFszqfV
y69rjC+LyRhNNlLPLH4MNIL7DcE2XNpBGdjoos7MfsLF2KswVy3kfmjMQT1zYn9TwRsOEk16twbw
PDbyw5s3G0QD36tXNsCUq+NqugjDI77XX0xQdiNhtoXL5k4wRW+at4lNU2nkzcGAoVPA1agsA6Ai
sqk135msZx+rd7wc8NC5+Qh7CaWRtvwaNp5YBcIpZeuObw7MXhCn4dPeb9T64Qq651vJuQWpJsG+
lAtbAl9FdowFiaipOvixv0S0OXiM7i4FIRriSD96sVxshbK/JRsUHh/HYsrKnzIriy1cgvAVfJfc
GTWiJ2njl8oFg7TXXna6E4V2adxuqEd9wHN+cRicPQH9M9jmCXkDFUmL0lg9mH5cfXPeYUaLV6wg
bu8yJqZayQLBGZ8jr+oOz/CrVi6PKBcgPwHzjGlA9puaLL26aLMH531/Yisu0xM0mZ37rf+9WJuy
zvwBJoSQtVovk6ffRBPbR6Rljn8UzZ9W0Iv9wS+BWHdOeq8OzKpUI0bVLAWWekLZ+cwAFLuTcYRG
KqfiX252gQ+Wj+tcEp4Neutbb+8lJVgELI+yo+zAU9j18yZrZjnuZahcrVN58oQtk+jWJLqE3cv4
FEn1RZrcuY5DXmE8L8kwAWoUTI+dbTc86kMozLXvs5lLj/jcvPzdVSp+NX/uy3A2JFGsqpe170m8
A6AL2tPfXMShE6gMa9gfB3e/YHLXZ2/emGVBuqOV70jQrKMwv26w5b0GQolwaTG50FDiiFf/Blw1
6LZ5mlbyMLLLIz0S41w8F20/cTIUvnj13QnFgZ6U7XiOzh+dyeIbr/av3Hr+RFrSq8j5YdajcM0F
rs5cvRRVi1zq2ViUMgLEg49rQkpiqlcE5SPdMRhqgsAVgT9rFE7Nrdf2CTcskXzktpGrFW/fVe1l
nU0WrZFYItHRmcenY3yNL3EeUs0Y2V4CipexvTXZpHMTxFwjilxMh7cmDKicozVJLpJxvySu+Zs7
70Xf+CpXBKGVOsUfD5tLWG52iI5WBAmO7Ma9Ie0pV4k9mrTfTUUXylctwWqcJ8sJP140TIimoB44
p1t/1XDEbrcyseBjbQdWeWUg1NfnFU1D/YF5PJvxDeAWphrEgld5JGs7vlUKfpq12U+SGQcSXCyd
N9oc91AyeRGD5XlYR2lSEvbEqEvs9PJnLzwd7UuFw7HCkk0QF7KPeyIb5IRc0BYDCxhEAzM/3kLJ
xYQfdyUoaufTX8wcrm7b2PaUw7IRjJUfFKKGMGfFvsKTWsR3jsqipcv9rMU0fOJkR2MItIzX9H36
ilcCGt7mtVRpo6t8kaMKNYLrzey213jqOXuJ9kFQfsg6pjxfa+EqE+jjkXhJJc6DFtwgZwwSfVeg
rCDOFyHH0KQuVzcmRL3O+rjbcAJePdzmZUB2UIcC+0FQ3tUqiKsJgVpnaP6DyDc4c42QXuNHqhGp
2YtRCqpd6mQlNNJ4wZIJ49sJiTVlL8qKmLmtAt781BCMB2ME7/KG336kO6sU9Rrh8J7PuHRv54ux
FQwijf1TZG/1b3yqS19dvbd0pg7rXZSlvRL/bhhfY1wfCmEVEQsXs1jW/gdU0NFEd8R31tsuZyQE
W0CHrrtm/i5lLjWxbJujSRch2rgP69riK2JJvZ2Dw7R0/ccewkyRg95RjVHLKrh8e5Jw6JUzviQF
fY5yfTy8SrGZhcZzG3f48oo5FmHZ6GroxAsUqZJpDqIRFFY3SMID2RJHRAw2ZxKi92fdh/1N2Ral
3+6DPOxZB6Z0rN+8ks8HZa71dXpfnrKNGr6QY40QgINIHOmAgECtytBX0MkWEsGjii8Dvfajx7Nf
ftuE2QfjvotHW2PTgJZm2gIGKygeqQk2/JPLP/Atnjwjdtfo8qe02nfvpJ6GYTiVLi98ga9Ey3oa
Davrm2/1vZZboWxA3nlG4SF9MT0OIxzA8xqIZYOqAhirHZJiGl8thXYWVtuvBamsYkTGTjkmetiK
qf/x+eh+Ovi71JLnbsj4OiecWpZwsF6OIcdBFZu7V2n+ENsBTtgiQlJS7pdkXeu1etIdKtKfKIid
4/gYA4WNAXq0v4P9eTbkUlbS0XkZ8WcDYjZ9HoJXe4f/dO0NwyobE1kcccNC76n0R/G2PtQzKDcc
uBoM2i1WeEcXRQIpBsgfQP3BtZWGVXuUuysVIgCy0o4HBNBzIVoA34FeOdobP1VWp3kbtQ4/31d7
Db9fsNkX/Ic3U4ONcVukHCigXrCbdcTtvPHN5e6pUq8McRvENzXzfSa89pS0spfp+PEt6Gp9B89i
9Qkr5BtluySmWlG+HC59TwNm82i7lok9S2E8ErFpci9WCCVEMrky5f+CqB4zGhk6Bx0eYToKvbGP
/JJ2j6EjDlN62JO1HRghccb5nnXRTCMRtKqdejSmWC41fhjnbuaniYDjNvr4x0vZggrYxOicsJpz
kI0L1VSc4qTA8eH/tCiZHbd2c1MwABlPFdhSVqW6fzwhknXP8AwD2zBjXtzP3phtSiMNz9ZVXGZ9
uJWn72aUMt/Byk8H4U8WzoRwwjLvWVrRV0w61XnLXCkt6r8hIOFKniKPvPVB8WbiIkp8XMoZ7boY
BehdiNE+2/nmqlIqsB8/hb2QnaOkXZIr8aNgi2AThdVaGXGt9OpQxMrLYQWCfJp98P/Abggo0uc6
7oPrNLIPvFyqG7Kyf+XX7h2A2wZip78gpXTtN484ixZffkjc4nN2yHMIyTwtdGMkQONrg9ePaRGo
21F8K+WqE9vEiL62saXEWRq8cfPkXT4h/1+xLZ7ux/93hWOSJBAW3snLBKNFVTFr+ODNOuSueg87
tBiUZPup58cnRImm4Zv9uCUcw2SmLPywKC6YhjvTKlYYlgSgDq9kFbaJOQzI5iIiR1kq3lD6PnL5
CchpGtL+wwLHSXBf9Ucp+4bLUwqH5F1/o1uSgA3SAL46iQ5EfSuvbRc4yNgAlMwuNP4OXo2015DZ
Vv9cCD1hVZMy+HwRYqtRCo2uHwRUCv7ocIB9p2QGZldS97S6BxxDG6q7RAq51CDKBpM+B4dsiHtq
A6s8mR9TWsfk8q8eFsp8qqimvZb66rso6CSKN+bnzpZrsAm7o/cwZ/0XuEDIFtsVDaR5+5iAKpFL
tK1bJE3KDCbCuj8qK4Dwsy1ZYR0k9n0Ymf8ZlpqHIq7/kXerjvPVY6v5bvpMBqSnPh2i7bCwPjOe
pEydeEcRE1zMIgmsVCAgo4frwjTSpygcrlVB02Ua1PpCc+CFpSOcuawcJe71hwD7ZQ3S48c7Zpv+
hGUf0fDRXvJ/uojtA7qGWasU7k6ll2lyzTuHz2s6rCuu4BvvX5kuSAaA/aSx/+idfoOlZIC9NH5c
iABcnjb8G0fmuhXJiaHF3UgyJkgA2jFUfv+8VsqGdmnuY8xgWETICzMyBIE0GhsoRsm2vrCzEGfF
Sv6BKbAvBcV2bsDsSOYCln3YJqj3db4k9qjdm7aXKuyFncxhCjEVKgThCkghjlSiph1bKk/+40Ym
8ej86y+kxJz2b0x63APB1QGOgxG3y4g/ZiFaZXjNguRqErQrK3CP/PWgEGmJ2lF36NxcmAoAXESQ
sZxPMdSM9xxH5uMyAaIrM5EqY0DgRcDjwUFbOKBPNi7CLmgWQR8/L2efnM27nWpT11zB7cfiLI0f
sWKz2SSOOhqWSVYRQBSSQuiQR5xilAP7fQcjwiHaba5gv8SEWm7MRrTk9XlHYk3xIawdVnF3Bw77
IzCeASwcPNFFjX5dC3Yt/NLjGW9lUMPiUvufm9IKBNw+l8R3y1kbcHYL4yMVVz31raunT+XJW027
tWz/1DWpO/W9Jceh0MCOQeI0UoLbUMee6bZOxSNoamEMAq90+XorBUrnqF7/wasfy5dVy0WLl7hN
XOHvleMEBN9tJl/haJOdww174QXtB6WcCaxHd6tKO2SXFr8pbgH4NPMTyCBmMaJG7kRpfmIcFYzr
9Z0LJ19IM5iICdGL5xfzqWo/ELdu74lXc+fRUUwYQuzkZ67VjPzUqmsBdjfZDI3O4ROrCfbeWnIV
i/JhudtY1SooJ0Aa8xwMWVZUncnjOuzFVN77v96rYOAYJljy1HgPnHLDRNQhIFP6d0HNMGYt7DXh
ry7KT75g1uqTiyiWqNxT9eQJtG7KVjwlX0ziFCtY5rv03k68p2+y5OUjPVC6s5I4/VwvyomoPLmS
UZN6A+5BHEY8roZRocHpDBjH2F81krppWkVEr5eyKI/wCUsWAVRLgEoPj2KE5w6DSbsSDh7rOixC
zieEl/7TH6DfwXaClyCcR5Z5Kf/d1gky474YYh6i/iMn8/q5imYWh9Qb+eqbNJcqA+Oqx2OeFGnh
4gtByHBoj+4n3ZaG1e+OCPDie9XTMefwFEOA5+EKZ+feDWfuatyU8adsrPqErHQNDOm51zQ+L1ZP
3ROIJX9cEVOSXc0mE+cwQfD8ll3BtfXW6/UfpCRmFGka8/wNPzAYZSnYcrv4Le+kgh8D/+e3XK/T
MUUtvSyVSaWj2vh3OOXEo0KuEjvPj7WR15RfmQkys+Xeh5U1QMfOpN16QgHjUIzTVbqTJe9rN8lc
wiR68hwKvIsonJ6+pJMFeouQkvuuAUwaujMAA2jUDqrE99eR8LUd0a5Qk/cRjJZNLaHXC6DwVWkG
+UIHO164ZOXEUOhTD6fPbuuDSUqHZZNf0D7ZJkRyINr0pZ0iDUIg/KeWiUMfvkXhn2K4F0DfKvb5
zUClx7ba5/r7E4CakRp4ctTjJphyrUga5crB6oH4f28l40LfkEe7R7aR6lgQw9k1pVpDT7Y6dzhy
vJQ0iZkLK807L52mSUdYq7rYd+6odD/XNrDtVq4x3BDSa0PVSXi1qkUdTIMPS5XxSOoyfYyS9PP9
3VX8y0LcLodR81TbtjTie/HtLbi7Rm5jQLCIywKqaNo8QdLzVfpr9KJVRwcnKuVF5ZwKIj6drQQg
2E+Ww6sKMdlCp2o8mYr6q16WCFjZw4+8RtHrEVPwypSrfgX5/z/b/Z2sqS3XbKwyRUw2bmkO4Ilz
RWHSGJW2x+jaME3J4Bp3TgIL1d317/hmJc91RonBVaoplD3Kg2gcDH4aNQ8rJJxRvUSYRJtOVr+G
UJ+4PLFsYV7u65xK1RMlvQf7n8lRwJlp2ZenmU0cDYlUso0NfHLBQqmmWyj28Wncidf7jjf6V7C7
g/x6MOuPR25oIrlAqBTkB+hY7LmL5KzsVVuCPlmmcqG/ySR/FL7Xg5ql3lAKLlY7luOJScKmzlSp
tTJ7zvLOVaCpEVXl0rmmj44ZlBaNPOOzSSf21V4v+s8WzyjJ/mS/3ATFqBxFXXi4zFat9ATD8NbK
+ySCDxWD7TeBSQDgPx7aXxgksx9TrjYxESMDomkC1DZO5fo0xfRCLV7v1yh+s3DL1gfHQm/jnaz5
Ou6GOlQ4BdzSDQvMSULMZqApwMSi/U6ZU+JXbKkP7i2JJzRdP/BPeuAShWX8Ss4MU06uR4T98Ot3
Td+JpCEuVdi6uzu6v6KMF/ocIFFXZRp3o+MER+ZvlCIUrlK9fS3avKrmGduxeApUQD0thX86Ovna
Twc+UIruiiTB3+Rlowg07knDItJ6jqQd5EPqAD6bHTVObky+/32rNq26oebj29X42Qp5F5ya+tZf
obpvMy+BRqXI3yWXZBLs3sgfGlvrU30hDecW8VW4beN8y9UMooAQQRUARXCSUrA/+Vn4VLiPIWzL
ERtLyRaAE8pt7MRMI8Gapx8+Vsc9SuHrpkE1O++Ic+ql258GJKGxrzhr9H6IQbE+Ez8mzBMji4Q5
hD623JpgujkIyUwlRjN4Fjv+5HeSgBWSufyUOtoF5x98SogcSSUcTdY7cguZlS/dOQ+VcaVfg2wV
389nk18gD4zfp03tAa8adoyb4pMJJMqNqms4GApfsDZqFCC34Fs74PlSDrwcdV5yeV300rMrPqEL
c0yjYPx4Quk0RALu0vxamUkwBvGWH4VB8EE6CWylZ87LP7d0F3s5x/oKJTCE5bF+OLTOxkVNvJw3
YDAv2l2M+e2axdPOtDw3atBaTNfUmYm6i+xwx+dxaRrHEi5J1wneFYATiElHZ19krcGbVJwk9ybV
T5RXCLqj6ueAxRWe2O9DA3CwKRQlipDex6GO59ZEohYlp540DrVTwhs/D5znSWX5IXFKPBbamp3v
VgYRN15k253o6mkyK59o5VGpheQ1PXayVmO2ZsoU5pPyljsVifgcZFY6QZKcbYRq5M1ZN8+63qb+
ruoipAcmEgRzSOwaXnm09dzLFKf8Asl0vipRoj2PAvpsa2NzcRBdO/G98C3OC7CBiUxAfFeF+CD4
yzZCgfdL2+H9RoOjOY9fOXE4nPz70HkWWc9LsZ1ffMRvnRJ4RZu4+UOk6D1Aiqh3k00KdYRRQOFN
E0XfE6L9rlxuThQyKHXKcbZZ9f6dtm/kOnaHMupmTVzDWJzt5x46MyVx1jmxPisE68YFZaDIpKiE
ceUAA3D3FQc8FPXP0VCZI7jIXTXErF0bC3Eb0W334VAtf7xKPPKtbDmB/m/j1GmntAlCVhnFfD6g
K+dS7ydsNyn9bTRC7y/SFrsXk2F5Ba9W6j62WYYmHBle+HrKOuXcsS04jELXKUbDkGTsBRHxoB6/
ic8b1ntXlMx2qAIXz8CKYhodAluuchgGVk7yzi6TJqzHRLAUh0PqtXCZGG/D/riIkZu/YASd0iKY
85Qzdn9TAyPTezNqfI8s8YRNBknKOjYu8OK7dEair117L9Xt/oYifHHISqSyVy0JJ3IkeY9v3XN/
V7u/BIEHE+0Y6gUfwzImfosVu7TesR2S422l7hwv6eSkvfl5tdJxSHthFT0TbjNVQpq61xcnRLX7
kHrKpbEoI5f9Ee1R5bfLaPVeICtn5bPMC057eIiNkJQi3ncSvb7ehSN+eVTzN9QF9bkzLUmKjEhw
GtQ9Mjj1QTF3dqcSlx/pkbmQw0j5Rdhfu8f6Z/dM1A8r8DfJDtRWKcWDq1Ro+HdZam1YNUk4Rwqu
Z1SDdmc+7gJCmRl0bV76HIt46XR9+sBRAWDVt7o4boJQSYdve5UtO7/72iBrQzwlOdKSYJfahNFM
zzLiAaYMi/bdzoKVm/AlukyoGJOy3wWve53q1Sw+vAVX9MEe85QCJPn4hy7pVLoymXd1SNhRV2LE
YqiePBwr27WCVpp+BZ8PqJNTZx5tXSM9t/iqcLSFDWziR/nn4kVCAFsWYsKf+3MLrhQ5XheL0aaO
UgsAzXFwyeafLfOpjKJxAdm1P2yNhR+gBOKr0ZRztwYBH/l8hJHjW+OpZdu5uqXyWTCwLjTWWr3D
EuS73/d9xZDLTfrHVPjt4U4vb8PLyYUF+b1m/eO0ugxpGw/JucGEhO/sAfQ2fUJ2jmXLx8/Cu+R+
k+MHZpvh9xzO3X2ldxbbBBi9zyXFfUWvDsZEZbNInNGjzZ5zpIJhMU7xYjq3Si8I0jHwp/eIwPOx
iRYl0WisUF7aD2NBXJ0HuCCw+epXXXTmvCUcNvjTM2ebTqA3cYpb/c9X1uLSlcorb9BZFMrt7xOD
BiyRkQFdQc+UhRBesDJg4yJChU/GznlTuVV72AJlDNaz7jojh5ehGmz+hXnaUjD4K+OG6TL3Q7jp
9R+pXY/zQ8Z4mogPM0njoLEmYm2QXzBr98moaYEEc8RavwOoXYiRfS0KYH2GWMGLChHoFjAKLWf8
jO0zlpCyGZy+pNPgt6SF1havddi+Be0xGmC9eEs4j6AJOSBldhbUxvsxkZlU5yLHRjLzdcuaeeT3
euXg0td99jA1G1/KxTevV5P4fr9oxWb4Or4aTOFiSHxFUohOix/xrlHlI6W+9mfZMpSN7d515ngC
Hqq98P10qOdwA2Af/BM3o9urWjP6B4DM5u3n2MwPeAMLrU4GVK3kJasRfCDCdnyKo7eTiUrN7hI4
dSaAbGkaqvX69blPR88/Crdxbg6XWaUbT3ooqh/tAVJNknW2uLMiLG/ZYgIjOoodu4VTpQDzShHv
eV2iKGZDIbOMYg9H6eXOLtkSa4Q8f7DeoI8LuGG3oqyyCav0t24REJ1x52laLtrpjTDU1/zJ7xPN
mQuFmhynKCVpuaOpbgrGW2tAZ6WVjMcE7hIOub5bdZKsvhAIydbkzp5S4GUMZc0JHrR/x1b9jkff
lrkWTX5PK7mQrX90oRP3kMsBDecqwNqrLpeRpxoG4l+dfYMV/8LueqIO1/Ei7nVtSJLw3u6AiHug
mHLRYBVFJ4h8jY+uATEPrC7bullM2MU+2xvZuAt87UaHyngqInKPUXJ9ZcYgz4VeHMitLKrQPFKQ
8zaJXABVSNoo+yYd6rc2KvqjKQ5NMck/RzEJLh/ORZ40LdBy+CQfd9x4onScPSHvcEhyS7j4u8nn
GwvMbMSHojH4XD0NhSapYXKKrk2gjr+/G9RbSWQQ7zYSSxYpZfU2JiVc18MFmUjcCOdh/dAnamKO
D6HNhODGOag3alVGoNYYy12wF/9v5HrLnIdhtIJfk1GKpCTUbOygD8vkwSpfsFL8hC6nc+iQ0d3I
egEwIudFZ5h+gOREfQOYTgozQ3fNjGbO54701IZ2yBnLD9XF1cm+hc/4eMwtvD4195o8S297uROC
gMV3WeZB4Fv49BOI/c8m5OzzPntfvXV8S6WpZQBZG20ceDMhbylEastuCHRkz/U97U4/K8D6jxii
H5n4gMQhjiseUvkrVDLyyEzzKlGPTqWXbBRp4k6Xd7X4wbmB57R3R5aKbFZn/Ztla9/N6O6SBEPe
/f5E22dwyWT5JE0KZf89eOGhVAIlM3fNrkxmBhOrfPlkKBpZ9oyDxipDfkpQ1JkRzHNMv4EXrPAW
wB/uyObYVjaAPVAzp1WmBh6Nz3TElvZLauz5eR41x+RK9iS7ZNpNZcInL/PDkLMbXYSppwXEC1iX
64WJa3BI058fDxnqOvKSfn76XJkstnX6ynTQKTNndNiiOe1EdKojl+JLtl8KYLs7pgBWTSPNb2da
mYUmFiml5biib9h68C/c2tLCpNK3WJMZsUzxtxKSZK3sFWmLiwuPPhC6NMwEHKSNdBKr7VQH5Y2D
1qomqABH9QbbaQhfEmNK9okPZA6rEpgm81AbUJbJFvkVWUrxXonCaE3t8rvUZq9OyhqqgMl7t64r
YYE3gWZDA1CJeboVczu39jq2dXFBvu7LFQsFkDnsyF2dLchEbfhHHZKAo0I3MUE0SS1uhJDVmhQ+
YXrtECX9vWy/OxHbFlOW9RqVyhIY+oh5wGVr3G4XJz+1O/y6CAKTBEH/ZXHr2a7AB9MftEUzaPAT
w9zLX5JXDwRCPLvc0KD6y1cE3ajbZECc8oCuTT46HwEEe5N4CTZ/MAkJ9Iq0OkzO/dise/rCvs7f
AW3a+NIXXNSGtPOl+6WG0C7CT3E/8quT9sMX6Qbv1nE9xdfzaUOVlMKLifbkGkYnB5PCgIq5qcW/
j1ZGm7mDYVRnkGK0sjUwSWp2wmc6RRzDKcFvBQ+1jglmQjTrIjxhLKpGTt8Mt8XQ23GVNLw3/IqC
5pEfCskJBm/6khqJqDsBQ1REd9M2305JDpgexoIqb3UEEjgEHPmQpX0OxTFd2O+qEX2EWDIBAHYv
nxdh4kYH6aUevOOAs5FxetWxejFgp/klr1GcjMLONMKX3Xin97MUXi9DHo6QEHftWTmCsrOk426T
4DHBVQQnSnKki4baK7huf1ZtXH7lbrct11J+Njw2qymAxStb65hg0WOB3dxYkGd5vlgadqWEiynV
wMq5ajyziOb1a4PnCpTllMZ+Ap/zo1WA4YZx7dKnaVuphmezDB32Rstrm3I1M6z5T8O2Y4NEaUG7
ib+QAbK7tOzMK49+7LmqDse9xScY7dEY2Hz4P6pTVM/R7SEGHletgBiG2cB+xTfpGa63plUgo9XR
soojY/YlAfXLxyodE0URuhaPPGiK8rk9ra8Yl12XsXlzvtcEnpgoFP1ib7GLQdo2BKpSSR+5Z0iM
/NGKUKpJI0uAfuvkOqExxXFKxcERM/SgnACdXwVqsbdx+piJJQsdmERrLXAwzk7x9u1wFLIcHQ2A
Pjlu5l4l26IohdZ01Rkooz8oQ1SQT2LAI+cU32stanvZG+HveEYSp1nY1yxVaotitE2sXC/McOvF
l1WoHrx6O+TF26W68sgosDP0O7Z4/08YEaIJ9pYJmFVGm53kkx6gWWgrNciS0WPSicow+MSUZEHy
mKkZbSG8vJIDWwWGMNC6sch7GXowmyncEFiGHFoi16lG5ST2xGK6OMcKGOFUR3UsCzPa6MzwUtup
qfOdYEk2KOtaSp5BJMtyqUqc/oD2yfLoAAU5bW7qpPPU7E6JNvm6KrtQcY6vIDFrpQEvZR4LKhBW
K9ft8oet3a8rJfjtUFXwIHUgFzscrxqdiUgtQjWfGSl65b5Sm4NBthCQf5zEusTX1IgNRt+G3Zlq
x3qXTFQaIGdEXYVIct3iR7CRpgputHI3fVV8dwnxSImV0xIPIPcF2IhqYEEYj+gDJ5BBH3OVTgEn
zUQLZTKUyp5eNHUfc2wmXksz8CSDnPrHvXl0eH423Wfcvbwu3HlDEPzQBzKJ9BnraL1JeJIASdAy
aUFQXE2ehTHierKqZoqy+d6Io4XWFrR4c4N6NVqiDl34XThlwUgzpeb1lS8BBDkItMRTzP8IasZB
uFrtea49JaO7znvyul/TTM6scXbc2rJ7DNr3DEBIcCkKBsgFFgDbznrEWmYVr8xZXFoOEcZ2FjIL
yteIvOcIN6ZRu4dXqKhQmO6pRx8qTexqjCY7KypUOnzq0NHzYi8e7rdP0W8PBl71MF84BIcDj6ZS
pPGnwHxANk2hfmwnC4fB3CAKqMqyGOMhLSmzGy7bqJe576449xFtDeTjhIhZCX3eozSPwP/asyqk
nQUIDILqyt1F6sKnURh1rufztla6ys2jH1CIYP/uWG/T8otprX8IojJ3S0rVZIzA6LIs0OKTDwXm
GEpWvTs1C1EzdznGeEsyvoQW21D9eDoWlnSW+Buk/pNq/2pfUZzmnUARhl8QFR/rzoQYtjQrgsfi
5gtq7PftUQxoEA0r+XQfBXIGGvXlKDkI5RdoXXlhyrINsJCTq6RNSaYNnAhQX/7P0ytse+e3a4El
NeZWXqVq6e2G2VubfF/hhGiwncx3RGbbVQSN+P8cpznoIRbCJh7MbqPo+69WYlalMTCH0Ibz2P2k
kJzDviOSFdTa9X+JdO5GYs6SvDShOpsNEQhV1PE5hGUqKxq4NhA2bzVGzSv++itWlJRk8PY4r7tG
F3vFKeZGjh0YNu21M/4026C1iVRg0S8CN04OhnjjB2IiWUFfd3Fg3iODrhivEjbhAFQ3/IEyaTjP
K4fCewaBXZ9dufSOugDJ894YjajWzLUALj16KibQgnqQKAt6KIMW1f07EuT9LkXDFZMKs091R7zy
5RYE5g0aJ2qub00CkkhQxfRwYvGG/0PxSaHlL13E6MqFk4HbRE0DHyu6oHQi/KrgMNi+IcOzaKuz
Ti2FBoniBVNyPST9kROCNxMxoEk8cXjt71/caY6h8U17QXia2WBx7V0jqx8I2h6d5Mwr9uLDgX8G
TLEkKPJfkan6+KTuEwMRiqMEVqiyixi2Kk8nOWVZTeGwKFLB293XwyBWM6FpXcFtJWvIwPyPCSKM
/oV3aepVPM64SdJBpuJr1soXpzHz3TvDx36RXLsajED315mzs1rkrAHJRjYqyhSRQJB0lfXLf25s
7iSC8N8Q4hf8hwL5r1vy6X4vIuuCUpc63RESkHDuTfSATr8ugzKCkOuNyya+5qYaHXhgDl9Yz6Ch
HrabxSviVuqiDmWChzUlN0BeyZINAx2T3/T7sUL+wyS+5UkLzOVAPbUiODkuTa0TpJc443fa4ZbF
f+0lyRwqEWXAuNQ6NYyTxKqFxmL+egRFVrfAJgGDG4p+RFUM0iw7KIHzMZzSaJiwoapeRuJnRHk2
oHKyYjpGH+MlJYSQnDEI+FZ1bTCbexMNIRd8KGm79AuxqQUwEvarO3555wGW0v57x35S82qih1da
G2sILfPLA3MmExSOdv8MjgQ30gQlzqHUH+qxr8H1Y/eDsND7lH15UACv/LNtvRxnUeU4Zcrp3XZf
+jO73apgjcHsJgPodFfMImnN64DH1NIhVotll8lsmObb4+5gT9FbYFp/sR+Xf4131B6dJYzSbFRe
dcCBkpnfbcFmWTXyjiivAj36n/vxneoWoFcxYYgoZatJIKLiaQnPbB8C1cAi/8Bum0jE/MsmFfHf
IBEKfuw422WR6Es5aPvbxTeGfXYRNo3/o/fuDXZxMGyXeiCDRyf2XWbHOSwQJSHlq6X9Uial5WBh
2gTfQJDCsI7VGrGMgS405xNxBBdDgRRs/wJY8jwjan7relJEEYJd61BYumMRJ1NgenfzCubsCDXW
DICgtJItNaYb9JYniGg9fU1AkRVbKfnem1vb5KoueZQ3+duZZcMvPQ/rwVLevlv4rST659npn80W
sqZCwC7FtI/+yRL1PvTrTHeX84Lb2jbkgjaSyVimz/mkVOgbazGGwS76VRlafKCSNPss6q0QAbzm
Jlq+85mhCwe1XS38Fg2gqADSvtCwpduPkaqta08N8Y8MMGqrcWdb8bUShSipDhVjk5ai4NGwQo83
iFyCCk/jQIsC8bmZhkB6N/rcyVNuydDLSGi15rp12yMVpjRRQrOFj+DPix8SI25TfRGWOoNdyh4d
EDakYMFmRlm2ItwLNzDZvKvVsZ5/No0gojrqrBxFUfJ9cd3Kf1GBJwSBG9/QKXe8byh0a5eMOQlL
vr/RMbWREl8o9254s+gzVMdYsAyPPW4pY8MNuJ1SBIaEi04PL8eQkqlajyBZhe9MqZ0REv/d9vPL
44mdyY93NJWql4e0gBlsNyKDDUjJjBhtADZwJZuxjC5tnYZtSWBhSPrdh+7SubYeChlw4zkRT7FG
llJDafDeCza5kcUidq2iqzgbmTjq/5LI0hBJM5qNybFWnQT31ZaXFr53JfvZqadyTd7XfhPTI4iT
0D6q2ayWnWcwf/pYPcGSkjSm0IjjbtFvwvLjFeUj5LogYWd2hKmkIE75q7sIixjaspmpOxjkUAEF
PDxXq0y9IpH3g3DJfYp0XSJ9ohfy0x6blMz0pPJ+meqkQjG6EJlqACE/Tz9VP3koNGshXm0Bp8m6
5iIbXSWAAURWRQUBs91F7K7vmUWylWcCr6kJk8SAVifvkHcH3wBI7e2Ph+6cuJJeXDFo++Yi2ibf
gr2TlXcrGcWlujjlHjNKg+jbTJ5mlnlNurEjnK430ppIExf+HaYiakWWMoZ8ogYvVN89i9HNUp4n
vuY+AVleRKkh1Bz2grvgsKba9JeBe3HtdPRQm8CkyjQGs++Su9+NW9rO6IqA4nLlt0xhRZOkAcP2
kL1emHo1KNLFv7wJk6e0RL492673XipUfmFUjGEkt4GCBA5/eiejQ/7VlUth8sDlr6BHg9UGNFYJ
hNl+bAXaseGnltSTqqRo7QeEDTqnAUpMUg/DHXbgV+6Ljqo5BKh9V96GmYR4zk1gyelA1N9HO1kM
ngmnFTzhLzXT42//9bODLJBjX36cPtXoRq8B3hpOizmf43w5AOF/D27iV5oQ5WpUIYaZm6Vmg/LJ
7iVqv0DPXYeJ6faSoS0jgF0O29kgJ6SM9RGGvvvYn83366qTho9ad1+YEDv2fW7JM5o9fGg0dci/
mEx8yMGn20/wMhXe3dlwcJtqQX98D023W2HhhJqQ1KSQMhUzi9nxHybCh8gW3vnnKFaDDQhLqttc
dMdYVy52jd9ggHBSX2+GlX+cgVBe1r25HkskXN2NhkZ7X2w8cHcjtgKDdDNGZTi+iRpGX/OiPO3J
Sw4XaaQmt7jW7iylNHpLllZez3jM9q7mJOmmAgMCmFp54LDnkxjfIP/FH60NmaweWzkUUs1lrojR
LXI7M2qAmiNwkCuuVIq4v/MMt/aA8Zu4UUjF5vM8mkjMDD6F0we+Da6tH90CVsArqJG/eJH2wmQN
uip+3bq/0VMRFgAmIogXrtKQM1WoTwy8hwoVukLre8E1lJ63odntvJuRutxgK/b5k5tK4zBNeekw
eVmQlQji6ppr3DW83dHVl+CxzA5WKD/stYwF2dWKpD53UP7VNiMkutGSyH3ESXcG7eQv1g4a383X
/YIa6nDbF1feMvcwcsIzrncohoa4TbrE/adzGuUqYTGSXvEbqZXYzXtMbWtO5QpPQPV7ooydBVUo
D65feFgXhlOf7neWoVslUItiw9Ac2YPANxW7Euay18FqwmFXw8GpZZwdsKlSJL4ocXLBHf5L2Xix
yD2j7gJOKUjet49h1PRqkYb/BsyRHiffGe3sqWp1/B7bGEUprEO0+FlZi6b0rpwiuQ182f7Uv+g0
cg7gKRJ7bX25gVwExEaoD2Bc9LmyHM+Bpq1QNjWfEsLg8fbL5019a9GghbezXRu4qBFDWddGFi8D
RWkGH+lBcxyA9l7s+4qB+YM4lf0w1Wd/du9X4HYtDUj8BujuWDrBZ+rDj468xsQ9iPA0mx0UJm9X
Bltw98VShA6xqukMeGSMNYdSGOnodTsbhyhL5SONs/MPp6PaOgBUni/nrZAelnfJgaCIbJIXMXP8
eRT5+AEbVucTGnvTCfdZZHscrs6+9yAS5EegTi8SKzcTzlLsxu5RTAUig3scGxHomiwFOWkq1XOZ
d5g/ifXbLCPkQuQGKNqUMltEAsw33SDa7XG1Rc2m3LQjL3NXF8imczFCNmRGY6vbVwxsCKvUHwAV
Tpsl2tno21NJ7bSTjVnuw5xGFqq4Sgx+iRCNk8kTQwmfENkxs+36JlM9VY7uuePGxh7rAGs3x/DR
r/6qDHGoOxDnl1FojdrFm+rr95rLMOk4bWp6t1X9jFqHh+SooqrOwNHUPZjgCzobSoyfVNfjswnc
/8+cUcXNcbXjrvWXTxKIOVWcYRux5+PRPeN7LeFeTxf3fBWyPDbkPue/MvcOem2Ycho2zXsZwm9+
/cnKkSVFgPEooKAAAtmfhIYE4nzwUz2CWTGtp0CsxYoeeHkO/8tmsLd8v7ol/LRl8F2nx0UJzhYe
jddPi8qzF/IXm9HVZw6usWMMyc1ZOL+p+zRMY5R+Y5QN+OC/TL07aUO/BSkSFhnIP0kDAmFP3Mjl
61usWvfq7wK71irVMI+KLtG3rFYqyDGpCIjTG4WtZtgJ9sM1yYsfXXZnW277eO5nBn4oRfGJqu5u
L77DTQgu2p9Q2YhQzdwFaeSNGq52YrrExWR1ph6DgrxuJHgDbrWkMQCE6X0IWlWVeYI+kfEfOkt8
D19CP1i1LJNtewGjslim5w7e12mHPb3UQFEPExx7MIHp4JLkgUmOYvUPd0/F+KnNQ4+9h0BbC9G5
wdreX5AqnKSRZTEEkf/yoLp7X8jYnjNiy+DUEGt/mtQuFEhmWDeJeloZK0LNPCdJ8E/p1DLlFBpc
VXnXTavz21oSACitTpR/QNVt02tYnM9MxU/N0mmFIoBgGemUeZIxLQsZuMUaS7tzs2d5H67DvIal
SbXusFtaaUAfxe19Z6JSJM8fZjqBEGWQj1YrnxmfL6L1tvJbXDlraSgj4z44CUKpdsdc9oMZC16e
OD7Mzz8yJLl9lUDgPfAwGZ/K/l6slZQaOka4F6D7yNts8EidjgHE6ymXDTQr1VwBeVq5AicP+IUF
oN6cEzehj3bmkB9nyUEWQ71k7Wz3KNUFxPPGfPvWOnKG/4oYs4iuVVO8nzUkVbLHFL1ctCH/EiJG
IJkeoUTxbU5pwpeIL0GZhQInJ5I8zOInWHyiYt6g4IWVDpFoit3bhPgDJgvTlzk9RmIq6dJlQZJ6
7ZJP7OJcaoxJRYJC/e7aDTFMtN8atx/fSysGaaaVmOUqurAGHvtecr/Bs/9oTMBqWvAB08+oQDcy
QYvI/RXEZzqSzJLJNjZ8TsC5ng7otst2daMyi5w2ti0DSu/qE6yDdhv02rePE5rYRJqPLaKNp//O
geu2Xnj4KHK3QjLKxsFGi9HpbrC4aGLaCWHuQS2lp4Xl69OeBszTeYh+6wAC+D/cfg3EDhKiH4cS
peO0YnY4wbPeQ8bAGpo86nUUZj++g3vy8OXmdIR42SV/2UhnGJYpdrSUeWVnVEYQ1S9K34f3vKhf
LU4WrLe52fonHhGIZQJN79exoIKTtJsPzTm+9pblvkH6m9bCBF95eu2yEulk3K14Q+7WXXduvOwn
DfDtXMP3bwfGKr+H//6lyHhV1kYADCN3GdFCr74H1ed+2dzZNn4eyukhRCOUb7NvDHMW4jilypfD
ECOW7GlfIzFdc6vTIOz0mF8IOz+bt0Um5RNX0lUmlEm8ueljPYN2iT6/OgfYYMLP3aKHOtS3tInc
YavTve4JD4e/bmSkgMnqA4MsZ0brjlBsr5ikbloMZyBYf+UlUXv6aj8w08wKToytbZiyuocpZ6hX
MopSKoS/7kjoYnK6oNEZEBJfWmr5F2+Scq4AoMh7Dx/mH+FQCPgxP++9cBLjSbHs9zn2P0jmM2ea
9lJ3rMSbmsvBvmBffRVV0pcvQg0q7daJifWJMoiPzj1UlMHqNOxzfTw6BxfflOnvAlu579GLwnzp
dOUxCVPASye7MQgDW9aKx0DeV64Sf7fBSWGY2k31m9mDMAXpom23tddIagrM+6HNnlQyp7cuRx5c
2POgvuILs4AR3fQPjIH4QG4UhOOX2okMH8oz6TZzLqfJ7tL5fvHsm2ILUvh5n2wXQRAL+Cb0iPym
s+we0Avpth0gangeZ7qVDa7ztJ6KZ2d61XhnNYhTilqpG8H+QuUMNNka7S955vqPc89dH2C+OdXg
uPbCnQx24W/D68RVl2rE4DwglC1Zn51LY+FoMvjDyOtwslMT3K4HCcWALlaAvQMJuG7B0NeTN+jD
IU58JUeuTYFAm+HI2FQrsovw306xgR/v854OF052QF0Vnd9DrWJHcoyIJSIoi704/9lT8ieb8wY9
EkVrjJy6IZlUtfauYAFFna6WdlpwLV48G/YHj73prkfVt/LGCBEGFJ+797LOaHq9FRPJFrmoT+Xb
6hk0+Y2tXnC+FJMIsTlzBK3kecgXXwtYLdzMyRC92CR4Un5npSABaOysOYq9KlAq+/WoLRzWT0dl
Xugr40y1pdhG1TqkFu/1d6LgqwvRvyZ/I8tHfMj1fk9+1h0I5pTSWcPUVFdmKocqTOwYeTSf/faL
O4iZlVfseuzmd0SV50rsXYkrVTSheLAY7L7kM8hXPMuhTlWsNCHWRJjVh0wWA9XZXb/7wMINQUcP
eNloPUFl5snJWTFW8NOzPfjooFIwnkM3LbthcwPuiYxbngtQcPYpFdoc3CIK8lCffBlKN5oJtrN2
4+O+NlK1NZxImIpBmRfLvWRqk5g6UI1buXdRAx5CyRdkHLEQxwTdwfmcG4KK57EIaXyfVo9AhRx1
Qn1xPtFdH9sBcz1TZRRqT+g19sKwuisSX5NXytnWwa789pB4S5RGXwP9TC/Oy/EONvlFJdMUuJPD
Ui+ghVNt4q6NOVzPQOjXi2IAZdr5XfaAybb9LscBW2Ov5q0h0UeENoAkIgIaH2PkmdinArvvjhCo
p6dUunMEyhncmENjxMPyvzElZXI/BhczPNrtPoZx+dgggOh7p0brPLXON5PoelHBWwhf1OJMEmfb
OrVXFT9xWljIX2lsQwe6siqdv7Wo8VsblorKDxSxxzx56SVz1xp+rF8Mu7jRjESgovn0dp+Sv+Zu
Pe5eqs9mJB0vqmA4JHaMlLa7nY+Ik4KMyvvvmGx0WNOlgbthu35h9x5A83vGA87Fu6lXix8j4Aw6
l/TuOYRmmZZaDKoJdfZaPAafpAdBuiw9+8uLz1+XUFN0ZC1ct/KT2abdr22Jqea4Rh8vGKk+LRg/
dcsz0TtrNtIrXwa8kl8pmn63OGFBo2JoCvos8zGYx7eMjcILKjnocus8jZ4LxwiMG/VkQbtBT9n7
ikmwH9HYkDMeAehwvO0/VzyHtEL5tWgyaxEHF5rfz8W7xbGuR+rjy/s0Jwbycvh2oWcNM1Nxhej4
JuXgY0G9aO0QML+AV/Rv2SNTdHovXR3cDabuWvv+FM90NjKe9Cl1a8oek91OLKAaw5v9w4Z72OrY
ifao8c+gK+old1OxDWZlH8FAqe+WoxlDBDJR8WFsa5jk3RO21At5QH0SN2tzArTEzdun8tnpABqY
t1GPctVyzcNKpbet6LLnBig6IuHwJTlpQztT7JOtSUY9cL3Il3LguzKzyw9p+OtXCg+9kHZ+nE3A
XIGFssss/K1rsbW8R3/G/2ERj+3HL/fDDGqAKv/xQVwQbIim/5OwwKESexJLA7B3p8JZ7lOgz6rd
1B6y8B42ptpDk6SsY8JJrFgrSTztGLiBSipS4w55oLueS6/JXmpGVUPTtSIbtb/cdk6PxRu3Rfst
fAONVCllWInkfKjV0rlIYqIGZ7HEMZVVf+WT6Rra23cPEHBKf8Kxc8IMy7b2slX+NeEIZK9FTpdd
hRdOnw0a/8Oxbd1wLjXqBSBzqhgnHs30yzwLcf/HhNtExHL2BWjuuBadprap1dAnvCJhPx32ZrHE
8c7oPOPXoJmAZXpCzIR3xPMhMq32eh0PJvYLbb/bNF09o7XeccOtVclRp/ZzKY90J5xyE88Z8gaT
sjT+XURb8VPGUtG0toZ6XMk7BOnI25m67y8NY4Niil09XR3LYsm69ISIs+qAI/oyajiTrt/ee/oy
zXjBkFYlbXiOPstsS8C/zFx/T7fVwv4ZOrMMLEUEz0/GQBmvrIPis9P9gJyb17bc5FKo0ROnwYMM
Fu/eU+EiWwlsiJtJrWEq0v2+ofGjUCvFbKua9UpPwWn9/j7NqFAPLZku+urUH92kCpdnzy+lYs4y
/H7HxCc1QYN6rRpBka2LRjzCziNu3suqEy+BUh3SgytE62z606qnk+SRcajn+eHszJ+8HM2vrbJk
heCkr2FLUtgpTSeTmSfs7A0V1qOr/vEcOp7NYNRs8jTQm7JUS/Is0jgke3BkW2UQX3krQ38JTjfy
HEFCgFZglew6Hme5nvcHiQU4xRoH/pHa83JzlKoV4oPDfxsQPqGbfMHjjmlCwkSBVhrSk5+DL8+e
oIRpua1rZCbMCVweB25W2zItgaOBllF1hgmk6eVUyVBVma2LONiTa9pex8gVBALUS4+glibsu838
kVd/tAi7SkrzgIWX4JzNQTHbxK4/Bv7f3IX31bypxD/h4A87uWweliZTHOAOp8YB1nCyVqO1F0kR
mZueRLqjPqIdgYd3by2PVRieq8iPTPCPcTXN4W7aZrPj04Aq+X3pA3R4dwrfKXTJ2FoQHlgBDATl
V2+9hi+4797/sNhV9/Q7qQkraz2qUBl8s3tMApjJ5md1gW9JDVCfFjDXIVMd70AihsiihsM8A4w0
8fioI8fq/ZvLzvz6qHd73uIlUBbwza/5GEKIrLWVDTnk8WzjGMErgq8Xel/GOAC0DM0ONxdbHKRA
BtCrcACzg5fFki7e8LEZKyYuX0OfP+ZRDiPNkCKq2GfwooUufHNYoGUozPaXqi1ToIrTafbh2WST
OGRtEmU1W5/TfIGHLlpY9YLsDbz9dngtfSkOXmZuqNfl8sRxSXu3JBGTpQLPjpKLDNtCVeJdNvsB
dGohdJNnRz6hjDvFxIp88WqEgg2SV4zxQnmTRbMErUm3Uwki6Zfnz2teM13bRU/0DDd6VKDp/Adx
WzgfaIj1abPfmhgXuUYe3NQgN8s0H/0A5Lmo2lIyVajpE3hwN1fyzLTocUqTdKh811FOigEwzDjm
T64EK7ckkIdWr7uKvx64oK5P1Dtk8hV9fgzedX5ggLcLFJ61/5tpl6x/GGRa7JHYmEI+rSoXwTP7
yuGrJPNMfdEu0TuiznMcqOSvOjGUULbcsiT3m252Dao2tdUjblOAbMpve6KWGbRrw8rFwLOeE+9/
DqmHgGVyoonU+i56l0u252F6sIHGa1fMBAEjZSsz3rnwreg3U5S2OHLqSQ4qaDRQNZoWmQBz9J9p
7lTC8UqHHNfxa5Ag9VanTNUAE1apkLkDXe5vxDAPmqa+CSlf9CIQ88vzo+6eANkr591lFIX0Litc
e+nPb02xana16rZOWDD2YA/gqd0JrZA0DzVb9yYhAS19g+WaY+8lEnjsn/RLLy/w2NbBQY4a6Fof
SFZWW/fkNKrRNT3dp/0ulwuSZwCH5vv7liisPJDMsJBlzd2v3NiF7+cQt57zgwmS42U6Y7E8qt0F
4N33cYDnmgm6Y2ZqHPmohG+uhlbhEz6UFg2ijRn6/IrohquVTBDKlGoYYEpMBJoomjLJJ0HuVNN3
0JHG9H5OIYpwiEJXDxjGIvyVuqR2IeIHqNISdZWmkPh3ztHMqNQ895I7UN1tgospLVrDNAnToxUn
9E/EKG5IOiOPJK9MOjVJFEg5nuDeKO2Zc2XYQIML734bjKSAJVvEotYZRiq2zQ0ZrnVAZOoeDoAq
bXlZltXW9fDjX324C7FO5jpRYaQXaDDe9BZYUsodOoc20TXNe3qt3kZvsTrGNtegyhYKJ2l1ISAq
55ya4Z3q26sJzJzsMcHl1LzmV65RsD1LWQaTprEKfxYoIJiFFXb1vnsRhk4t4EECU9LvvPgZOh4w
xq3aAASEQS0Wkn1ifG1QyC/ISU5j55pRRXm+EqqUQfPWYHzpEAknYsVoRFXHPzbrAOkTBLoHCTTv
iDIBqd/T1fQM+RhioR9D5L69c3gSbj7NZkLhNWUchv/0wLE+u/+rfeeoT0DkBbQiTqTiQcBZ9GK4
PCXGLvuljU+o1dsW1JsetJ4OnlBQR9BiE7Gz7zg/8dimYBksoJgqPcKYlCT3B3hasrSSWxhUUUHD
yms3zlbNEy4vtUe0T2gO6wveoFvEB1MTeaujgQGD2eQbeTcnUPEJ2QTw1jEI6ElWmOIIeg8DbtcF
BHHin9EHfUynBC5tm1vM/4XM/wdVx0dOcocUO0eT1Z+Pjyx2dySCFHLiqy9QnAaoAdxDRa93+UUl
feNpJSavSLYZCJO90L0MjA8tFqplBV2nf4PH4ByeEjP3UR39FjQTY342k8QjJ8dVA/U+5bBiD7Kj
fyaVrkZQDdS+0apgwhPw8lggmzcJVqvr1mIgIVEK06zR4Ig5gNXFzpbc76CMYgMeW5GwG2O7IMqf
mW4z2NNtYheH2pZ33b06P37NV+K7f7Q2YM38aktuptk6WGxS8CpRwruZLt1pjAh7nmHzkCQa20YY
Aaev4hWty+6pxksve0cBDc1GWncnHI3mxWS2EOs5QGQ5sSnCFyhsDyE97O2DSPSDGGZnGMBidBwG
QYDm3H2Wb6UVtiIzGuFn81ckq3G/CHYSp6OAsNrQ1OyZJu/LqrHID4CMesUpi1qQqUUAH6+7kokw
YMkKctJbBUEYVX+b1m6RLN3s0j6d9VLiV9rUseM/SjARTvZ9pTvoR8QwNoS7ZIg3UkEADahrB/O5
zPskSBuBK93NhtCBROcklCN5o5I3uLRberc1tKjGh9bc/0CgY+i/kAFfjuEPp7P9MByidB4iTt1K
iUVBvfAbE/FN87ODbR6pWyoOwKTEagcDAZmjWEfIzrIF+hikijlTkiFQ3GIz/cVIVyPDOTKFqrqt
1+U5ELFDA2Ah2f+dbedLlk0Md/far6+GdCf9nwjDwwSoRVgQd11cr4uFFZAqFFSfB4TSMojWp2TT
5Qy/yPmk2rv+ukICWZk7Se2B0sP4BsS2O2MY8QO+NbUgpn1CfdPogPBDOOK2iMDUG7hwJU8DRq9J
SYhBEhIaOa7Onr6ya/Fpim5wQmCCWxeA28e41Il+z+se1zrodFxbp+NqOWRzGVM5oQoaJKtsuEgn
l+gS9Fa46ZnKTEZtAaxP9sLsTVsld8AAuJNcNl6UndxJS5kR1m26nzCoy/kKUp6fs3OM99woE0o+
ASHndsqX2Jf6U2UJ9Qua4Rq9sC7LnGNxiAJYNRA7si/x/nNjT7cFemLR0rE6horsKlOKFm+TOE9n
rdQsirKo9Z1xIY4W58u0w2TTeEGhcWyiNwInta506Z2+vR74sjpxcRUYymPeMqGzfL5fwsuWnyU9
FJ7Cma9Zl2zc11z3j/i5POUTyDlcu60aJUu1cx3b7G7ukphlD7pgWghMWH/L9YczVJTFtleBBywB
5GN0oqpH7ql9eaqbs7BhWP2scIfGAraa2sPgNLZzTKda9+ZtcqiBR5fRsF+/ojWXsup53oa37SJ4
i1i3j97NZ+QChazOXhGEhLne5g34EunTOIs/QjrD8Ch4P0TJAvGhJ/Vm4gzR9Vkr4QP/lN477rJC
J9jMHB4wKI69lh7/Zc2GLs3WthW4dsKU6PnvMwK8WnAjvsIvuN6j8CV8DZ3wLDHxZOR3hMg5Dzkm
NO4sW5OB7qQQFzqT3APRVMVjkSnCtN+KCI3hGvGF8pknrI06bh0nxqDD+c/PnWYsaRV74hj8y/6E
dPhTyMfc2pL5sIlYiaHOTJs552d9KQkGg6DZMtVOFRgPi7kF3OMLvXfStyurbe3f/UPnWfS/m5TU
Jvbe7qe5BKLPx+n46tZ0rSowPxW1IcMb/uboY1b3UWkoNkpRFw0+jYdUeo9nsOtJ6rSTfe7+DPiU
NsWr15SG+SQsV3QdK5jS8V/VqWXOsRe8yNGqcrjbFYlYmfLFx7i3MQ93O2iC/ig9ttP61P8eK7b5
8577QzjZ81g4TuvJBpKZOYLd45bNpVTF/1rOKgBqD0bfc3/0vY55QuAuaKCvGUpFJgt8B2rSfh3G
iOPAY+HSG54XsUzD1bM2zmKR/iFtqg0DzfmGETJk0yle/I7Ns4OviiQ7duhwoNHLJBqHvmfUFs5G
aBMlB6JF6C4V2rBSyY2KCyB58K0vOtYAYSNBAAzxHqyIhm5iwdx/GJZMSB51U+/gFFm3sfqeq9FQ
a43fpwxyG4RXm8wDLqIJMl1ZK8K5OgBk6HyWaObqwJAL3tQXEdcxb0BDYZlho8h70vHPZhJsWgG9
Rh5fH2MNFvooo5g5WP/nWDce0Fa+RWMlJMfejQQZCrV5sYUOyhXq1Ib4aXoq0OhfsO/r0HBdwS8s
IE57qGnBLOySBMqld+XMmKTwCOpua+RvMZlrE2+rrDi5xE5xBs4AsDQCtmz/eIgGS/ZtfXC/0ESc
JBhlIu/9l2keg+NZcuBsckhBc5aewFebsfl1Zm1+rtqaTsYu8ZzXPqajeIMrUuTNnU03j6b2d7Vo
IrH+IRU4tHKwtAGhAgfMY27EpuLsZddpFkrKw8ecBhAmelmYVpj3dfwxaNGLMiO/Vvmf7hA294ut
XbmfIKdJdPpKDSBVQVZRlj7crDTMVm1Wg8IVrHQXlnhCsd1WtMYPwBvv/gMCpGvGIx059Z4dM+0K
TERwaG8ydSVUawbd8ZEPbNMyQtzXL35iRJrf7TqXxYx5bhC0A2W/voPtUGnhgSY3L3a58lKkpgOM
dqzmgvAh/BUNhw3sG5cOLM/Pvw5ioSlbL+bnp3kgNwjmAjnRJ750YXNDv/9D9XJXZYy2ra6kYr/P
fgKnquAHn7rXaPPXX2S7q17H0CPufcC3l++1ohlRpKXibSm8JXz99Q1km3ayglXW+JgcfgUHLjlD
H7KFFqrxEvtdU0cdyeiFQJzdHErOKTbOMLiIhhOYZflFp/H8/k0mUwSdNTj+A1A9Y5i3f8GMspRN
G5+oKRgMjhHEiXCB2AEz8gJImGkfZwqqCN72TnFYdFqWWrFLx1nHTCyRm7ZKCe3pQ5YTyzuKDI4b
8NPSq1sOPDVcvAD79mrC99Q4rPtkKUszQR/C6G9cmjj2p69i8bhUq7lm4rdUW07hlLangu5IVYd8
5b3pxpDUrmaDMl+7yPrubA2zBm/vReTAVJOdO1d2gjpmr86aczXsyCRYwfGxL+uR2y1IFYIf3XWH
IAPfw/TncIaRMEVrfq63xibGDmx9+tsLhRg4MqgvIIDIfGu+9TgpZhOidDk/X8X1IRtkA58oL1AJ
LETgCCgyBz2j5KYo7sl9BVVG+f/zghXtm+l9S5xSWZMALJjCwZaXTrkz9J1OfJS3qeXSAlNkoo5G
mHRfLGA41v6XRVMgkiUspGE8tTtsgDV5EW9wmP/0QdWbsdHDFlktnahWfg6RBQ37WFCVXoX4pKOC
TZVmsDpQnU8KLJ7Tb5Nw0Leu/lDUlCH3R5wnK11DrNLVXHb+gN2XX3sRrSk2lTyepIAevDkdGX9U
ZPk7jW53Bd9WSzdXBw6JTHw2FmDXMbUiGH3iy1MVLflWkjg5clpJjazq/UYHzaREOiZQv0xnoryD
f6N4nmc9iOPCqqpUCv3aL6bujGrBBqRkiLcPH5V34qIwSjrcqVe3KqjfRPamQrtIE2y2IoFkOl6T
XMnOnXB6rv60iRfnUm0uWG4HtfIRVdZHXzSE3XF3zbzNylJuguu6gUbd3tfZs5dpfVc/c15r2x49
6KWBlr71P8CVA4siAdKM5A3pa0Z6k4pGys0rudcDDcave2L56/wOGcP0gm7KQBFoJV9qO5p8mqvj
9KKSjGE51U28BnnGi7vgNsNdMvat/syIeCXfOgQifcamhFn5cYyVwnxXYdrJsHXj685vLPw7jmRq
7WhUIxBc1FUiVfey+9ERLZcm9opuuUJVBmOOn6FG9lJbMM3KNL68V+VYOyEhzEvppS/SSHegNoed
MQM/ilCsi6oGOgM+AawvnjuIOajQ+v/rKIs04NKf4RFefXwF0BQd2PCdscvcET+cBSIZw8w3HKOL
0DYP4uZq5b+vXP6jXT8A+2njHzW8iBjBg6q85lnhKfKm1v5cOSsvHQSrRPSErw/vJc6JUVFYNtvL
Iu4P3GCWEPReeITE12159ejL63LlaP0HZXZ2L5HYEVdbnEhSbwjJffcEgUcu1hNYJJtH8PXUGvqk
ekrR0vzqWmKboggK5Rsw0pq+va/qgANUpc9jVIjedJX7k/CV3IDyz4U0APEGiB2kjMumMSwjQogn
4Z6M7mWKuXX4z+CSY8lNC7Z3jhs3P4ZUAv04cmR4VRBLB+v9UvsoUovvZdX76kmk0xozac7aQxYo
QyTVtjCDd8l3DfhsgkZd1Qqv9aOqM2OMlrvCg18jASgiNlUwD0kYOtXTcULz0EfqAoJYXXO7jcBl
90Db93TQS6KToHUavy/x9gTgdUx2JQLlOJvoMzd4Qp03Bk5Let7G7zMl9mCGmrHLUrCr6JMUWopW
xYLnoBwEm1R6tuwPbrBiRpfBa09UCgng+szsfxyHmWEIaqIVpZQm5uX8LIQLHRwBciw3dbFdWo3k
I4JD908OCe7tIy0jfuj26yv+lGNny/Sueun0jeMqPe8gZPGQ+LBdQofNTy3nw0GTsNfnQDOoNeul
KqkcVCin5TXWwRQhsapDG5dVEZxSC8vBmQMuVo2afxZ/gppUppMAoguC59bjsd/NvDcYLFtRBDYi
ZE4HDbLRhKuWkOxh0jkIMNRg3ToxAlPZTWPu11mOt/I+GsyJsrWKp0WaVoVFDfSpu3DZZ3vgxkWL
tTntsGKThPtrF6T4vy03ieXmBg6C/dr37BoACYQayTgdAXp5NhkGs+S/IRJqDr5PA8bBLrvdpEa8
EwZihonrcWAu9+ixVdyXGRzli2BX17iVECHbYWDl5ZRHiOyZycmnaJbxa6bnS4rD5pduSi/KvXoq
iGolyqnwbaczhUnAY7hTd9dLOxq63YbwghAtfUe1bRrXB8KVrgGYdr8DMxPbL9d23f7F78OZXQGK
lifQwl5odm0XEq61XKY3qsw2Z0wNV2mijWDvnsHHlcs6du24M43kKhja5E0n7jtx3oRMO9xF+TuJ
Kei8DLw0rmxQ5qu0hQCFn2FKSx9TJk321pS30+S0SGb3oG+ADvuJHT0wUE+0m7dMbnZv/HNiD0B6
VRkW2SpowqgEOwkWjMDq45XMWSl4M/rQICNpCsHABzfeMgg5+YNO/Vv65LTwstTcj2FbTqPRrGsn
eZhyyn9MooEB4ZLnTPlJL1l+Oh3FfZpFpU+ejt0NGjBG9mbj2fHNZt26uuZUOyNt6KW3fxbUHB6w
MfsGhcxc5tsy1/49BDUh6EjlATG02B0wpeqBfpycDPN3sqW/A1nfYJb/dmuT0EaQRVaZHj72s5FD
GpC2vRRtYB3SEGfqirnpZJ0XO6TtXezhro5VaJJUkHj8BXEmBkZqsXI6sl1Qde/mys2gHfRZJ/qn
NKO1HMq3sVSdMAMgVA7lm6xzEiEejNdgenUTt6V4wyxILchI5kEJe94nE9KilHrUl9Bi8Cvr+/Gr
S6kbS9wgPq6jnf1fx9RwN9U0Opexq5a8sP6sZ2rFCLaNcesBkcKdWxX5fvlPFZ21/zOFcM8wFmhf
ExeqvULIJFdAerIWnajNHGBjZnVQeRA2Q30VYxXaZf5MxU+dwyCvey5l1TPXWfkoUHS4m0toKxak
eZI6syEid6YJY0uUizNdYQdlewvRn2Vq6zKgT3I8inAsGyrQ+T3TNZ91U6TE9d6Q/S0vu29tuMra
N9V901etAqx5T4dMQIwL9ifhhEIN1uzqND1fs56xkf+FeStRZYRBG1E8Zj3iFP6pyIPMwEQPY9+1
d364cjlZKACa4rJAi3kZf+Uqohan3K90Eh6Kv5GQ2q0l9mai657YNzMgbTtyyBYIhNa1t88XfAU8
qpRDu8JRvCMESJEuLWBR23DrRe+mlYh9iooKzZOnhQQLRy597WUIoy+X54zeXJeYqxJz+li/M/ds
jBMJitV/ewfT17zMKFrXRCNCU91fG0OQSoYETu3KEw2mTImMuUxvnG0B8l0CkbfjKG1P2do+2Lr1
YkhWdYCWHFzSo2JvNykrqBP40cRs7twoF4KJJnLF71/xrVHjyYFNx707YiWsbW27PpGYXYrKySWe
At9aRQmFntVbSF4Wo8Z8yTGB/K1T5Ahnr+o3q4FQ1SzSZ41q3PcXShLgLX6oUDSlEtnj/UMP7iaa
Za8FX2x9YF9EJiHGmw3wWZ+7LgBMmVHeU4vOS3Q6IL0m5HcbZuMwvizW3SEfiPXWflTydPPK2crB
cLS3Qhq8IfnfoxHUqFNqanxl/L3Ms7rWUftpVH43QzbqT8EkgSrveyX4T1sMg67ejzKqkmK5C78t
2y3K94Anz7POkIv77JF+FKCWkqBa5j5fHIrViM8dNMatxAThjiWhwTRe2y1GN4qecSZGowEr4fkK
7kzoSMQNnqhYbec5eCTtcsDNBc67m5+1dpjuOzY6e47U3ttIX7vlC9GrYJUymqN2ZlSdJz/z+nRU
KjsqB1kMCHYXK5gZRSQBzHXaCh+sA6NTQscYyEc4dmQKIWh9R5broKKum+43/973fYogW81yMmqm
+1ZV1n16NCMrYMIIAsPRrbMsU4iNYCw2SnIhB69F8qJpG2QOvzEpRFr4d/NmYBFo1l34DALRzpfZ
qM+uoyTCeY7d3g7+KS6uvLdSqBFA1Y9dVDrNruxTUt/Sbu9Ov2P2uoS+cd7Zj8z5a2lz77WJ7QY7
igim5wH5+FJ6qOoO+PACTS7Vf9XtRJlPN4DoZ7cH2VPA3vkAgn2QMmqIsJGQSSyHTpgmT6ciH4VW
8MQqunTvuajVltLgjphRLMvUhn0amtrz2Usg8x2U7k0bLrfno7shTSuqbdxv3VT3aV241L7qbbXS
a/F6+OuYuLGKf8LTsNeBEnIb6kuwM+CszJOumRw3ueX+b/khU36vEXa5LASA/0goTCIdzNc1cQjm
vZH0SC2wvAE+huaI37kbThFjDQYRcsCiQDxhbMx8amdLi9gHR6s7SFmczyz+sTYKgEPkcsUd6rkT
BkQgAbzLznwtiReZ/0vfnSkGnsZdxr3SQAMHw3AtINwGI21StOncR/vW8uqFHRxNSuyZcDwANkSr
gEmdHDIwq7Q3tnaTD8e3aGH40EUhfdw+XD75TUYMAmEHqfldJOl8+yaRv635fHmF59123sccLtZv
HpuK7JuI5frkxLWD3HpKVtlg4OdWa7a8sdw8a42XpzCFGQf5Io5k8cTmxTiTSomslEuWaO3uHSIz
p/rbjQUSdjWf9aAt9BPuf0mJMt5ouuWEjLn6DcRqCPWIIT2z78fg3Xmaoox/QvhX0gpAPlGJHJed
4gJD093JHG4/3rsMOw3fy6zk+Pvrjbj5IYBjN+j7JLmKlYrLRdZbdychjZNeq+ynrzMMH2/D0Pzu
f7FZHql+WBQN0Bw7uf5VkhALJVLF7EmgjKyi6pYt9olit4qAeA4LXt3Sfvaq9yWHMcazd8zb4b4P
yVHJlKCod7ZeAx/vhJMLnXuYxL8x/N0zntFTSSB8p/bFXIhk3S2z/ymeuBqlGbaJHGjHRuhhV3ob
uYSY4PYQ3uhcE86Uf/I+MV4qCVavFNUxcSLch1M6CRBTWz18HYgETMtvhk9J+UXAnQKgVRJQovzJ
ZwFPzPyEXtJLgYChriBA+Q7HxVY4L3c8WyDq5vnblgfeI5Td4LHoIIOn5S48K2ReLkLAoJGLjPhm
khlduVY54LfkT9t30Wp5wzo2IDR+Il4G2zn/9K7kF+EgSAduiYx5Dq6dl0K+9XX6g2Q9hPHklhI/
s0E5ES8H7d6cdM9B7H1bPhqsB5K9LAryptYFf0P8BWdwX63u15ThHvn2otE/0IojrajlbztjQKpz
QlKNexYyBJQMkhp3yakiPirQSkW8OBW4yWovVRd5vTSML7qGyBD0/rdizBgAPQ2HC9tRWhgFso12
p8Ns+DH4LTp9FMq/DQayF8XHLEAlH81ihLnVZJ4hzZX7Kg4CSV6xyPvUJV1VYXKcBAKRC7SnkKzU
RGA+SA4CQ202ksTgXN12J2Hh5bRFWAw9DTJgco0gmXWRn7tmIMape0sjiwdjLfJDss2IpB4mcVSy
bSJM5E/aIfrrL2eRYR5Zz5sDRsDfrL3JV2T+jutQ4EOMpG2D5J8VAw125arjpLmyY5m5K5WM0DTy
3XN/R+3L8WHvbB8NsVHh+QAeVEFDsayskIg3zmmbV+pFEudBAONOwC94Pj0lLhuPl1Pjs3Hs6VtQ
g8vTUhVcqoTv9gtnY33fZdh+s2PRnP3bcke1EUAccb1aFOwLiaIRum6mF1+DH5a9ZY2mbpXRKhWC
pQTdRMINlls2txK8B6YzYRs80VSQ96jA1zd5sous4khZ3MZNoKgdGu5kfMzV2/rMarvNmnrzqLCe
aJ7j1AaK9YLKwjMKx0uSsnXarAZDYiKzcqUoCxoBwlBR0zlLDYtXYR4K0Kx9f/F+vlcMxdkZHqbm
2Vf9zUUCjfdh/x5MV6xfZSwCKmiY/hvgTagZDY0JLew1yCpuCYZirU7nyCFaa3M6dAo94mVg8Oe6
jtnz3HGDbXGv89R2WboITDz+nJkKULGaYpF+L+Lc0Me3Q1o13B/gdnvy/ZYsGIW8q2FkXStP0l8Z
DyxnPwAUFYz6OIONIVMfXJ8Jjt6GSLTthH5zUHvktIRcOUWOevTSskz3Li/FU8l8uhD6OrsTHwtc
XxM1fN36kY8o5JKVqlZy+q3o2JermiHU27T9h8sKGdBdlgwmDN6sEntcymlpbVC6yDUalQCYqwh1
BtEYhX5LVlVsG2X31KdMpga2c46yhXJs0bmiQMBiEoTbIJ2UMXj08oUqZzKATxKdXPGt/9l5rECm
YMtitNGLsfRbx3RWgg+fYmOQvfmjZAnbUFZqVCytN3UBLXBJlN71VSwLF+W/YBZFkVRMM83K1fsL
KWN2T1x/ERD+cYn4tTd3vGyTKumcpeG4I0DN0xuGvOqzVxdQAK4BB52B1bW2FnrhOYFiSVOiIZv0
3FqP8HG38XENWETg/fs+iedS4fjBr4wygpScYEdM1gYzGGOtw5nw+Kt8frtF/FqILlVsIFb9Z1Vg
GsfjPIrx+Q5OeneRVYIIvVXOKWTy3MEdY1+M6BZrIvZjKTrNupzbcaGahupKXAzQIvb8HUb+gPvd
MEBI7jr0c6DwA2lVxcuTjDu/E0/t8Cztfyi3yL6hCvM1g6X1ouSmPO+zqHqDhihetQALzS8TIOZh
2J6moO1R9H0D9ULO8WDEqHdUP7Z09EA+b8IDov+Ta3/JvcWaIa6L7xBpSxbB1yhU9GG3uFz3nMFu
1de9FjlKI1weIVylRcCHc6XNM1ixhMZtipDOLnT/caviyyv5BNl6R/eDGmPwOvGeJZ46dnCC5WEv
JDw5AiVOq1fRnOkh5eFvuhwPJmywdfg3TNaglZZ0EmkoSURCmnMRJDvYEXRmzMOCaf+A8mLQRunR
btL/8uFBvrEd1TPGAss51DTmy06PjXAI7rmlg/ezOBpcofFK0wIjQhTvzOSsRjhCDYrK7x95vtgK
EL6+5IlTqd/8+UY5L+DVDF+WBIIN0RsgboBRQJ1YN6zjgnWScbiV4RconPKpUfR5K4iNtmeVNjne
gn6T0JjiyF4MEwJlzeYSLewzwf5wm8iz7hme64nfLe76+2OB5R9Z/pork0P5IktXX65WDU8XNOVa
ERaUY+zz70hRgSZn2vkCY3MCBQ1z2v+CS0w8VALS7WOtBruqrYhb64uG0mOqnv03xzvU9oNHTEgn
ZJTQSLrHHrjOVAn2QKDdIHj2CoD1T+g6PFNm5vsOlXDMIGgqZ09M2LTx6evm4NY0FP96AFPm7Zyb
IC6OofP7At26IDTlkFw0jm+3NrqC1GnTmXeUpcUXIsUQqXrH8zfgLw4r2jifb5izilIgy5Pdfgna
YaOQDA+Xx8xbEvIuAfxMpVQx+Ce1zXmVIp05QMuva97H8nR6ZLruEfhYemLYSJ9Lb/Khsp4SfHhI
HQ7/Hmm1tVnf5ccdDu5wJLidSAvo6ldHGk9BstXm38YvG9wFFc5zXFPS8SfwAOqfqwgylPJJd+z8
p8A2vAiIq53k9eziqyc7kXFIfpJJf8NvnniGRxWNb/1h5vB7vU1MorJ2L59NH8wjuZ+w0GFLGT2g
aINM+tVzUaJYyzIiFWO+xIgUDfbOYEECalovdjtT+eyt3BbvDLUGM5Ec/dtr0dStib9w0YjXWczv
WnZFdWi93dOYeZEwM7obcqBAiJT8F1pL4bS0RUAIAG37xZMbBLENEaUDp4lvmGRfAC7TRtu54Bt1
M6T65NqSOXgc+Yr2uI/bhHS8kBDhA9ZCijd7QdjOmnLrvfyFbk9TXA6a+PzMiINE6cGBpuJtE+4O
80QE2hIbavebqHvNQ+jnxVzCNB3E8CiS8dLd/0urWHa9ijJP1m3rE1KUCdpE7kzClRmtceU1wjNb
wkqIUqFq97UWFe+dgiO9HUuSo047agKKilSaNTaVQ4BUiKxsb6V5SPHa6KzLFiZ8kbMBuFa/9aCX
9rBfwyV1aiJ2JKHdxokRUMFTfbsjV606KrZuoklyjVMJ//OUb+T4MtrwKN/3i13y7O5ybXqWH3Qj
YRmGlHgvE8W+cNHZ22BUjQ4VsszHfnm0qfun5cks/57cj79DQXFSCVjRmoptlphpwGxUb8qXjMJk
/+5JQAgHTPKkdqXfZT7ARhXwM91weM1OQwqhAz02V9SJ6bu2z+j6dR3kjf69ARn9NaQ3f6NiRfAV
/qM9ril888NyA+A5qGWCs+70LsZluTL7U/AdkFiJMK+dkgGRxRmxpkseyLhNlOYKqlvmZQSZ8B7Z
gAgHOlnEOW5QYcCiB7E3L9qBgOgIecv673ge7Vo7MdYrzrV5FKZ41yHobeT0D+5zHEm+3uEot8wt
X5JKnXCVvR+ZR2XbRJd2PYf2zboCjasuQdAVuXBINotpQ2GEsKcZlo1iepSZsuv0n0FUaP+pwg6C
ffaiQ4rg7XJqX7tNqzjiZ2Tqtg/uGgq4cHqx9CJrjsiFzvyTCrCzHOPxNpgtu0OsA5AN13ngWnQJ
+FhdeibX0SZG8oTEUlifS40z2MrYfXJ7PbFrCyKT0US4WlONhyXRl1qM/f7Jun49Kl+Zz1ehyl2D
glwTQZD2K1IXeBqJeYC3CZCPKw/QH1ftsP73AG4mJwT1ebOhdjEV4jSPK5uO2/GIIx006eYk+ip2
1+JgZjPRwU0zVs+vUeAuVA1HMcfm65dQmu1+yydYnUdg+Vtjhs6+jP+umwj5USwXpqJ95u0OYuz1
JuNa+YR2d4sj7jLF9kXBkR0he38dgbChWujzOADKjcNtxqGh/rGoHk78b8dpWRKtRTKoS04MGHIQ
Js48VliSuDke7SlHQxe26zlNbFPjUvXVyuforz6NVtS93Dc8zc/+tukkNFJZQwUkrZkYuLPSTeiF
5M5HQWOOnt4en6ykVY2SPrx9Xoyd/M5bYgjw4/2vm17SkQ451N0Fy9kHVpXbtMqiPn80FRmUtxcH
uT5O0Lv0d+dl5a9im59tB5FARdQ70/5yrGm2fzbRm0OKNvC1sDG1AkCX3Uz4/WuEcqGkjNy+YKYy
kauwkcKUGfgTcyKbZHMyR+Tc/pThsJqIk244gO+UngxFi++h1sbzXQLdymyZOthXwamrfVLa9f5I
f2/A+Zo3Cy31TVwZ7qctRe5IeqxLEPmeSNludFlLu4Ngz3WziAf3HYlTjeesqVegaj0DbdujRzq7
DsP5yATYoL72tD84ap5Z2P4TN9QM2CkjYO2EXaJrElDtcd/+VUZIJEoXV6yWTqA/2+gp0deibvaS
yTP8VdkIsISa+aN8jBT5L+pAl0NkrRGHuYTlQzmG77/5MoiKlN1NcjXL6UWV/N9ZkzP5YrOhRsxy
5IjbkOIN9iG4SOXdKbB0Sjk7MfvcTtKdtXYT3Wi4fcISqewETyqjwvA9KxhHRVOeRuLihRhE9yXs
LJzamkPrtvTRO/ZVbBq4IVwsO+29RCDSQogm4+Re6VZpIN0dzyMZHTJs0Fvfp0hOECsG+OcruBCL
qz4Ja0R/dk5wmlp4ECUBFg1I7/kXrg7kK1J0q585qtLTd6/GigDwBrtKPO3fEkIQPW74yj2yn+mO
wlkysn9KCduRmmEk6+n6jSReVoP4MalAxSTwVQEFsf/locAlxwrvkUSsPorziojnlu1gOQ6dRVr3
TpZt2snCu0e0WaPuQSJg+j/r1+VsfKH8Nx+ceKijkLx3OlMWR6UBww82GI9EEWQ9QV1NTXeQNaSk
u7/r0osXfJx/mdlfeVpCTzgHrn1sdkADCv5tFK1Q5yAkc+eJ5N25dp8rkBglIvL0aVCEG2O8YPRg
LgjpX39JrbZo1gU7B881MfTxoFshfs6nT9hdztVLqn3QbMrDFWxcStAolKfWvQE0UPghX82QZyv+
k6sGulCowjNTYbZdQ1bXU6+Pc7eP8dG3ujn2d4bvHrZEs5OMsLTX1uQadJY45FNasTI4AXp+c36F
EjfLdO55948cntAx81kDlUropG0W27EI8s7D+FaSMJafV9U8qglmTTjs3s1hfdnDEad5CDaUFjy4
z4RXBRwSymGAbCnMiLgCA1/7Zf8V2m2GUiKz3b7oHFb/CUeZYhpvZ3u8H3A9oNkX0Yf1HH4mlns6
ybxUpPvTyCidk2cmYtE8X21e8PUmY6PlH0tE1mowhTW8zO6XZGWEjOMS1GWYhJq3vMAuoONViZZy
xcKpgJRIp6Pr3W4aSwWxKXxeV6WunBdWdEL7THT9eG1O+hCO88mPgq3bGTfsU4ocWz3jaXG+g/94
Ir4qWqbgTW3JsUX8N7Vq9qNY1vOOrfNYFHv0C+yxp0U81IDW86VGkdQSTIGx02A25mjsd6iLngFc
8aHT4lMV9/FleCLQie8xDZmgzPohRJEy3G+vtinz3zHh4xnYuxHf1v4zQh4/770TpHoU9FLex35T
F0dtQYUlg2ME/e3nSS+stIsvU943QO0jJj+k/9uAqwb77kzJy4UHjBTg9b27ttJzrRi/SmBVDiey
uLbYaxLAU/hw3QRy9x4YIlvlPQfxr8Ol/Six7nUsTSRYB2xDu5UOYTMFJUAUbhTU2/LHV73e+E2Q
mhxzWtF24fcH/QfEI+iCOpySGa9jCpf4RrQ7OLrvrW5fD0IB4d0sBqcb4al3OvNO7nZ/W3ZK5qc3
5Lylseh8UWsaz3uqpL3aQomW0pc8DW2hD1i4cKT3loBXFIUBeatBv97YIq4grWUCaAWibpJTBSlp
8hjFCo7UQt5TELCCMJDBnZzxM9eF9534xM1gXl2kvaLkLrKK7eI5NvUPl7VNmnuyEpT6KoSuMaKY
mv0AtY3vI0FOwFrlkDRm7AtsYai28nEgtoFVD1dr/rEyKZ4YBsHSKArdAcexwwF3jyuGAp5zPHg0
fMAM8BCFsHoe6ygr16N8Vq6YIEHXjLmvPwmLQi5vT1s3LmMIGMuOiKKJT3SUos5KA3aAjYNlEO38
x6ef7RpBaJVsm1lPqUXBqXJuFUL+Oq0lxidYBaalJys+P62VIO2mXV/jrfTjhu0REX4ZJKkVIF6L
WHzy0O4SkbP6fK2YAqB/o1hFcmRwZUfEdX/cFS/qrGSOgR44fNj1UCQyxkBuQpW2CdZRSdiV62mY
MQ5UOLP3PPGsUj/qgpT2jf2eTGd4jFTdoYFzu1NkhlBMQ2nhBFPhZN8PDikcRnmZvsY6CbILg7K+
GAkVAAmc5zz7iJpSRC/YIgH6oEecMFUa7yNMFqzkzH9hPVIYMnkxf1uvxC0JlL3T3ey1obTFUHol
o0qONANDRJdThLTu760qecvVeaN7sNZdF5uRenCzMP3u5/jlf420l3BjkQKi9HXLvYsdl43EMRF3
Mvo1q8k3emOASbmMfLg8lTRZUqvrUoqTsPQn70JUJTPsjQ7EfDSXC5Ii+FUNV2CYtlMlaXUEX/dV
aN/+hagMfBIQc3k2Zq/VRV0D9mcQAjCXsGuZDqMXr7gDvJ3vV8skWVptpaYP4Yc1wGVnBDSLSYAj
GZlDLDmlFb1d86GOOE8PyYto4PHndSUB6W9o3KA9ysURFhZP/8Q3oMcp23/iKJkFTHwgSNwdFBjm
vxU1oc4mVIqwjpy0WngJVorNJMeDkKVZTApDoWyWGJqbcH/0yrK8OhhnK9utkskUXV1Z+0GYyFur
DR4yZnJqXHAp4o4FjQ5MgQb5oZt3yRDTC7YR+fwzRxdL0awXACPy8Kdwea9U9CAlorm3/aovOJee
JgSt+eJjw7O9XyZ53UjLDWJ+sfSUyaXmUvP5ZRQ9pSU/Ar+EResEWgBhSHLURv5ywUO+/sBTuJla
4daTiA7qFbpYJoWagHBRXuuasLxzrVGuEiDdmp9pS/XoPzv6XG+1jqE8nmzY3aceEujK6XoyznjV
BeBq3Ziq1+uRBud9GjK0XPVcfIV8onL3jzO4tvY5GvAGmV5uFoCuIWdVKY+YADtodlPjVI7+ZRzI
oH8TsOcdqVHbAKI+HegXYwL5YBc+JY1UhYS++AFDQub95Z7VasYDBJvPhkT3lgtyQAdjNohcg3zj
ZLqeYiXlaZ1EaAD+Us57uaUNZS1Evw5agWyYN+hWDn/szoeXXo9QJsAs1FZGFTgy21dr6Op7i5DM
LLiMRbjlL9Y82IcMVD2lu8rBpdX+hszFc0uBgDtfoN0mqaVt9jKxAKqkj6UTQe8RiujWBAkfu0Y+
1GlAiZtTmkZgX4XvbjxuKQNjEKgUSrdeTYh+QI/ou6bhA26ikl5R9aG8Yns8W7WWMi2B87NcXokN
QAO8m8I85V74oaHzoRCLit/lqw4o9NOGJzT7cJNOnaP2pZZxWxGdLRcnD8+fjSr0DdwrdI4biE+d
PN8Dx2+/D5isDO2UM4OHY4nALf601n8gnwMwa4WmIFh8OaGvKCeZRypvonkHOqFOw++Wypc+hfa8
RUHMFhNMBUoU1Cze/stECJ7m07tOuqhm+MKd6hwH0/LijItncj+2GGepZWH3Ayop3u7Bsr747fxi
10JX92yRPAa3FlpmuV26Q5xgkW50Cy95QrdsC4xUBmmM/a8KGbX3etP4FjY/LHEV3MUrv+WY4Q/y
Pgk67GzJhusH2mzm/AHgVDsv3YhqGn1buSpDFRbGQbJWcc6syaE8Z6NWEBIttr4B0mCBlejBNZ/v
HoSUDe1lRAly3dN2KCakpWSGXmIGz0l2ZuWRPFDsMwSLShK/juvg72SXfFJnr0Z2lXXoGGDrQRpD
RPOYPmae7yMzHxXPj6clxIn+Sb3JpN3PS0ZUtSffKC8dc5MTvYTSbGNqaTYjZrsq4ZvkZY+gP1bN
LWSbSP0vYWYXvSt0x4Ijm3J4NdAP+iRLVBQ8WuH9qQB2tYguzln0B+iclNtmuEZGnYULojCkdISU
sEEzMQbqzCpqTvAP/kwNRzHhL6sp0yoT8ObcBnzYvmQptD3GIraORj9Tj/pD/duKuYXQNF5HFzxR
oAm6WAXbg/ct2es8r8aUy/NYoqd2I7i+upigwBhJSQAss8Oc87W/Pw21os9wsxEeRoXsUssP5eZQ
tgwsfO9DK0Jdee6cUbtAbaVNtwKSAYqJLOwFl7pYpOfDpLqVpjHqYNFUyWhAmMKVuX2T4RWg4W4a
FVPIA+y/WJqltt+p/E5B/5Kqc9N8+3DwDEvQ5440EDq29VwssmgJkRx/zgBJfwK9/WeO6FDmpBLf
SzP/vw0VDjRjHt4QWLsPRz10/pzRemEXWgiKrVgvLoQamnKUKAjqIjH+UvYPa/b6LrqKxQD+N+FK
ztTvAqxWiIjCLgYWJqeOrN4mxRD8tZbNFb0pFLd9j10oLM7yHEBK+52InfPBeiHHRjFvIMS+BV9L
H2CcDstZVDtnjZBgL7qeJrCjoeJLXj33O8WVvaJ43TKxhOGbqga2nAGrb8U2DADBPWi1LUv4vRpE
d+4SDfOpGrdPcpVY3KPvoq2GnwDEZ68nIU1P3rjCjife+wPN0w2eJe2AhIwW1UhFii2+eiWBE3Wn
bLeK/CG+bt+iQ2wlYXZPaXY6IJxH+wAusW0xnrAR6pdbjXBZklYjK8se5FZzq4lThM3k1/5AgcZy
rSh2PNh67wyzOJwm9T5No1mVrOs0iP5AFBbjKJjDaNTm238pIlW03Tl6RUvJyJq5kqsrr3/QB9GC
V+JP5xVyd5XZMew/IMD6Y/5Be15tUJINMGHt2UjAXXBjh4AljRTTCbpZPD32fh28ouR8sZVZ7tao
ewsNxkgoZNaqlxe2yccCNUJzjOlaebkc2LFgTyoXTnvhxhVi5MQLDKZTVqB9W/3jPaa7cIrHNSml
1uBh30+YfNxMBa5DrUthR710yh/YaempSlPmowVXXdlpG0lpTjgmmQTQhBUaSdB4XixtUlqt2eme
YxSkowOoEiAQ6FqeFbjbSNYkeTikicoTiHVixELHkKkYJy62zVvJ3dUPNCE9PN59tZd3+38OvvbA
BsXVdZiQWAtD6KF/dyvck41q6ETMY6LvSPaKB55H/s5HXl6IIS9l95yI5+NKCzfN1tN9dEefWqqY
SVp+C9KIw69+mF/oCzoPBnVDIXKVjeyoKljTKlSTuJvoFM4U9VcTr1W149tbRVLolqlQes0eHQGo
Hvf5/u5oBCYBtVc84G4d+U5vQmWYGZ8BWvT1zvGzz+1xr8HzWyHUSwD6+3RFaH4gWZcUJIAZxFTU
KQerwBjqq54UOfOuN9aC64JFQotgm4JtSLQKnlveLcliKOgDm5IuLCRX5VTc0aLqY2AV/1ZZ9R9R
mUbC3BCsD1x0ZBJurqK4rpEB928CYK1Lb9UItrLuA/vV+6iHhN8Xq1SlcspapqlHPqpiwFT2dlQX
+5PapWEOrK40aL/uBLwMjnuOkqq8714BsUd5z6AeEJYQX764Z+cu7uFMXGtNECT0OsWxxDrzYEnF
4EdaQj5RawER4iH8x3TRevJTl2tfsjOcOfon97h/Np4KgZm1Gj5eX2xVmR40Vmg6NwlZn8iDMlmx
6+p2fxDDGzplMR0mA6OGvACBaHu0hD6Auk4qtrgDb2+/LcEnAYMrItlFF6/JdVeFjjyvG52eqaEo
1ZGW0Q0FFN/vE5sCAPPu6axUm2i4cgXzRtAFEvd8LN6j49IiQjNWJmy2k/ralaKDDVWnoLjofcLX
BpxPOmvv5H+GtzVwUQiE/8Y7SDPxG38SQsve5+gefv4y2P7czPF2wIYVf32YYSCjVgrwaOLTn+WV
KArEyikmdyJdC6Kl5CGZePYdyTUGAKhociZ7zhCfqolMJvqBIiDfJlfeX2Q5XTRL/J87c6AV+FpI
HZjiaJ/j5lENvXLzYYEROZzPlbWdjFBOq8zUDEgnUwJktr8X3tNicZUeYu66cBteyNA/okUjXRS3
pkYW31yCj6M1J/yJxEdQOHyU8JuuR173h33MUPKcOsMejv7DoA7LEeRABBX22pZDXIeVzQWi3Y3Z
E096I3JWZ/IgHHOaUuyYFa/GqOE68+Upwo0TYAUv8mvVab7KSG35S9BDxY9d4oluw8rzrEdVGHpm
JjJP8LiOkwkNBhVEMAWrKECoUaVNI3HhMMCPDvf79DD2h94l8R09+Ql3RJHlLeRmqxCQriGrnTWR
Y3KrGTkM6DINRD30/MxA6XvceKnFifODYGC/1GuOrsjiW5mLqC+Gl0Kn+w7nWn5nMkfJIJHpyzoG
u6vkQZWKoGegVAdj1d11ftvNfHgObHUlZGiiqo44bm3sVOTFg0Dtei3jDkOhIbNi2lVGrRz86+HL
gopUFxFe6CqLW1t0rcgyjbWeLc2Z+lyVlkHMqE+yIKJHaBqmd4AjkwciNSxLHBmyKxJAU8h1oLd0
d/PiqJQZ0IOt4cY5YOlJvmmvOA9WiVSV1eGvjYgwOvSz3QVooqS498c5UaF9DebFSxJnHQHFhvWs
oU5H5ClDn5fNrLQ3emhGhP2y0RjktRbc+ReZmQT9OFT5xLCTw58LsGu4QNRozfvNR0U/RIPrN0J5
OdhxjW2ARKVfWXZGIDhIjEk6C5Duqb8dM/E+A9EAk+kYt6t3xQQmoHChKzq9TGYzthHY64Zjfl/B
fqRE0Ll3A4uhMCGRShq0XHzauO4vvGjjGSs7thgzo9ytAaSebPtjW/Y1GUcJYc3ABY7VeCNy/0+g
KzkjoUM4HLdoWD8BjxkSn4nx490qQJ4Ggb4z69u2+jcz0Q+6cKGUQsz6rCFTnDE8NAvjuP6T355u
Br8UjJNGi3NkPLQ30vHnZHtH+6ghVjHC1/Hf8SabFE1tChky2Hhn1vWoUARSubbdtFmA/RBTM8lE
vDIz1yk+l9bm9S/XTQdFDp59bQ6mVKJ55E873Xy3m1+JjxguTPhWoTNCBsRPFYB5ZE5p2zOEtZO4
jI0umQo5+woZYXBWBK+7gXGc4RBolZT2QNfpdyDgt/uB5oOatepx67gnU0QAf+Qr+E//H3L72ln8
VAcSTEZLjNdM4wmWa+nKnao4/2SgYG7eHZtHTTZFswXE0aXYtDnwTj6juXtyU8SWbIsyWw1vuRB2
YkIP/XXGdGUJUegEdAPj1rzgzt/BhYzKgc6+yPElrKD97gXWjA1kNYcqMVrIgJrml33AZQ7fPZNf
n0ew41au8KkzVzth/AoczhJ51GzHpajVGFklsFH73PgglZmKDDy+q/r+Uotfmy0W9JhTXL0mJDRV
edZjtJRJtx/xFP0kaz6EH0b7PO6yF+qD5jRlW2kPDMKaup8Ba6VSi/9eDHmCWZebQhMcP42Lp3/I
hSqiOii2X3PPdHkVvD0NeWo8rcWwdL3ohsq43KMyflWTvxxre9gXlXMYU3CnkQcuakgVNKRTCYTK
nBSqduxNh57/j1pWzysvyvpBzPXnBfBBAuC7puhrGPqNKs5ZL3QScqQpx4Ki9mJVi9PXr1vvNvzN
z2emdaoGDJMBegq67Q6d0SyJ2a/ZlS135kbizegHLKdEVYo0utrWzly/D//L3e9IXi/mvtjIhATp
w7NuyCAbAKkLd/0rE3u5CYS0SyNBLtkhUTs6YwX3bhoNKRIB6JWQ0BEw4lEEwzpAPdHdpFgoPVsc
0GGa9GiKJ7PyC/J7kGIw6OaSJMFMesG6nrPNq0jMepvlMI9OV6+RGWD50YVYZOgXjXqi5TDCmLo9
tbB0omVjHP7+fLdBL6lL2aT530eQNTXraafmQ/Xi1g9qkK2tvOwixdBEcbf/+S2ZF1WRLEU9A48v
NmYe0iu5ULl+FkyavxoJlJ1eaNcFcAbCt4ly/vrQym/T4d2GGUibEO0zGkFHWtmk4zOMEoW2yMZR
GCVPhf+YL7HTdB5EOOWwcRgD6tRVyRSMb4RbyqhdfZca+Z2xdFD7LduoFjUjX5cVVZ9PJcBOeKPl
hmCQ5dzJH6V/WUiIvTgP5emMzqXGU3jRy4OAORjRyBsg92r3W+4slMi6P9zTTTU6WyhVYwrZ/WrM
qNl7qtylWkzXHmbH0IBkoITEp6g/3vXu/lmeaGlMeF5hVqJAQaLIOqmmJKhyjoM237nr1RXCczz6
LtHuzjymaAMEtc5rwO51cnH8nqDwsI4Sh1ux243rEChQiJp74hsjsckckUWKaPwAGVJlkI1bpJqs
jlIeIKMO0gZX3lxOyPeOdll2aufLe3GZg4UU7JXvgyygcmKx+C9dLF7ilHOnH+D2z36T7fPByvGW
wq2yp8GPgrEo6iCof6VvJIQGgHC8QZjzW5iIJL9TVWDtRQ4ys4720Q4ysHLs6UkhdAvXoD37F9/c
dS4ENGfz4vpu8A6ONb07TThGCvjYP6WhviV96i99qyZ4t8XYSNtZQcy+8KTasm+rY9vvEmef+6PP
R3m5jyopFVDhhVsb98rr24ioR4qb0iIpewK21WiKR/UmQpdjERqhcX1iCGAxin+DxcbPECxD7BPx
wQc9bCSqLPc/r7JgHbRueak+bzCW64JReUhMFTdwukl/BA7yn/6BIEAZoeNgdcZg1BvELV7DIkCU
1pildzohR7PakDH0motCUkFh8+uIJ+3hvoJBfgEOph2xstJJ76hCrHwNIpJABaCSkE9o78c1ayjL
ZwopYuM8XXQumKcnDCP23TRu2SznH3ZcJRIJDawlslh6fj61o+mcpXBy/CXzSjicAdzRrnNXXbOT
K/cdzNo3Dh7lOOKggVuEG1Iw72t9lGKcO8UIZmhq0mAlaaxHsco2+MEjRk7k8ubkKYnyzYSAQQ4S
A+A4YNWEmvIIBk/xc4Hqp934g9w8IliVjDqF9d+ElOAeWcxjfhB0ueTPCblxdE+nBjohAOzlX14g
4FafeV8cBXZR03o6XaOJ2oZ/Rty6oEihCO+n7MnDqfodtItu93Oo37bTOm/SEGFbK4yBcL9x440+
XPV1Smup6NhEtPapLZ305NCcZCS8i62UUfApTNfE/XsEfAFjGCEzT1c90JvX3Yh52dpSxkSEfFBX
ytHz7iZahh5TqANoaCB5X5kRdo2gV9NeEzptwitFiddp8eoETbMCUzVNw0VjJ46FUqf+U2N6jLHm
XEUAGnbFO3/F00duIVzrYM43LQI5rKASVtzF+pOWvTT8sqIIDnlETBZ0TDFhYSMQg49XoqNYKk0N
FnaCiZFHrbA5nNbmW6dX9rngTkL3g70zG6eo3vDmssVUNRDBTj3Ed6GhZ8m3F0Nk3a96nHfPHwXn
U0H6kkaYohh5V1qlvO2minbxYfut8FbnPeV1pPGn1JCe4RYzd964ZZRm0QtMlSf/ZKdVgiUKVBum
pUj5qOdDIkvpnBseUTnRXOzjeQnlCW6p7/7L7U9BHmWaMtXKu0bveXveg3TXFyE3TmBd+Oue+UDA
OoKDOVqomyl7llchMrczaFo3g79RKXtNX/59iYPInhTDMj2addGHhwJsG7ZMXxtplaMa7D4gnqxB
4aE3GThJsjtXBmPZ7neFqSLZR6bzVCOT25a+yzKyzKlLHujhYMPASMId8BJ8P/2TDLSmuO8XYr4a
2BuccckfQs7A55KJQYAkpUMsw5+5k/PkFlJ4jFWzELaCbuPZCTjZnBfR1su7xQTBVLuigilQ50JG
YAjo2cg06QaxHlyb8SkXQs+FxTrn7ekogW5ZoA6UxrneL44QyVC+I227a+wV99MIy3Q2PmFewxsd
dZ6B+r/FBMwgIAP4VaFKo8EBJJEhhjqAVpKBoswPJmk/Ud/qZVriOIHgjEB0y2bFJJcC76k7+IIU
bgAM42zel0VCYrZKli+m6PeK/Xz939YjuPZuoH1rMOrhqw+lV80zv17+K36CiXaNL6/4Vv/FDVIE
mYrr5mC1seC592IM+R9aGBffQUXEBg7iNe4+NioFPQMHveoYyQIDWTl5d24lHiIhcTr64Vh4NCyX
7/pSk1ljCRYII7J7wL2X8HoTIDaz/J4d5V7bW2Ofelgls1g9lGy+8w92XIcdC4TCFJZTHpwqBqLs
//jS7FWcHML1lw1sMhxGkUFdUbhsiI2HwQrcYpcpRGw6Nt2Q2+m95LBRRcy/bzh2+ly8v/eeJKh7
Ldy4eWeE++0HilZoBnYFiXRgKS3YiIXTTuUk9JpbUSjBhoZBiSTY3Fv+Po/HKIMbvXDPBWo6pD18
MGeG5zJJQCbMqf5UABETB5reMYJpLUyspfQf/NqSqeuPlPO1R0FTFGYmnJqzvNWpyzj9Tb1nqDRt
E2w/aL4486PXY6Kkcn59vbx+SGuFfKm9ZgXZhdjH+xq0GnsEiFpcrGKTng/ApZMKNbKGyS/Eqdrd
I8otsqcCsm9RfvT/brWuBjnI7tkHYa0HUSKvbJ9BU2BTCKiU5KMDCvnVpnM+Uv1lGlxFkVw8uRgp
CHqvA5HboJSIO+zWueQzvfZh3iyB46NOM9Hv7zS6LY8HLO46eFyCvwT/TV7pQfXC947R0vP9yLfr
tLJ2o6th3s1xe32/Mch99smYdlfQI7cYKYq0t249WNO2NeUtxMsmzaaPDct+zHQwK/GKUuytUAP9
7koutE0Yx86rafO+80bOhVmgQ+zfxmkS/FVqBvkd1XsKzD3dTIlprAEKpNvUdGsW4c2GPCrpbLAi
K5KWS71ZqVHYz+7YfbcPCXfSQrZnxjl8eU7K30ZQ3hiuGz0jYUVNRv2wk1idI+PHa0uUfcnnSGDl
unYRct801LthsRE+HgzkPwbdQAvAz69kJJqGyjlxQM3qEKm79PwqBnG3E6RUgSWfBN8dk8c/0gW4
PhVpGaQaF18/wTzlQtd6BukO7ri2jdiICnPJn4wImBEugp4xN0Fk/L09N+J279vWdUwqUk3mL/2J
fQhK1DrEShN22j1Lh1XB7qLm351ktdaIT5cF/km5swpBL+OnRXUnw7ODkIjhroKAsQwsq5KWcKkl
wA4d0IDHUt2U31zJxD0fIcGeD6/SctvzkZgXfQrLOsmIUhh6MPBnwrtP7cWOyMhFG0Tx4B3lXICP
U8d5+guL5Bb4/uuFMzeDxhuBXttc8BicCU42dwQjoLO7Z6+rBvfZl5Vr/hjfyBFgxRqKQx3SQkLd
LUFHyjKzq4c6tmEjZb1u0HJlI74Pvs6xcvD2yhPs8JxWsAdTnp7tRsXbD0tNX6TiSWYtPy9mBc/e
we0nfhd0UCDtTmitDevtdOP7VgrnYYoHqX2xfzLKO2oS6O3JiN+Ow8ieWf4nlETPy3KnrtVagKqs
hZxn33x4OYfK5p/JW5pNZmRjpWo0WKLs8S2Pw9y4dy1YpdkUXxqHVhhtxKv9DgS7W7hI5r/u987W
TZ40rY3ZjIwFzh8nKBYniPgml9YMCB/G6CgWtGZ6YYhjwWnn8yqplmL9WccSobf29pwqWFLnBvC0
lOhrh7lW5yBwvZmD6zRqqKsQSEgiqCaflF2m23DsCPsj0ont6j73SkabOnTfgYm/IVwsW4KLNtJo
z2cUfASLR4FcEoTo9mQa31x9nIdCLnkDjNd2rqwU7O/RRA2Cgu6xwexWHZzVghePXG1B7hbhK6q7
6iEpkPgOn02sCkNAl6Y4Z1pI+MFg62JQqKKqryZ2kg7Ql2j1dEptDa/rEAm2Vw7T1p5pPTFqOHKd
UjfkwpyDcP9rBPUSp+saVx2xANPfUai7Z72mWBR3C1IT4Z+FKgBnP4vIm/rs+z3XdbqE8leGUY4R
gB9tH5mTSrecOpiYXxzlM08WW9K+EBL0/k0xTFDalhbBOFCfHjlO2xRoezqcgEfQb+oc0jVHhQR+
bMWiTWV1mGpd0L9gOAy7G4xsSfJnlbMM7FNBUAKfVm7wbg77jutwWJweGBRWXl0+j7/D5Rmu3RrR
BTFXGdC+u9GF60heYk4y4XJhntDkRx0UAyQX8DevSfPU4MI4j0brIwpGx/RUVgtCShcScZYL/NUJ
2ynbt8dkjtRkIp31aI5mctVuaLWTLIhNnu4KlP7r3p+M+a1k4X4HPuMzEc/mrcHyAz4eDNQpaetS
8SFdYsbJVnRWqitOG3SoToKhMlRxQWKOO4ko3MEl+73gCtM8ntlkfxkePhxzTu290Io8VfDeQg/W
c4fHa5fC+iS0F9yZTAWHXwFaID9Is2BeYNYUWM+dhO8zTp0XKlnahOwxlEITBsXkXBmuo4wLIfDX
AZfPsIr3TeUBoTE0Zqm+2e/f3VXTgAPFIUOP4Qme/VRanWqXUximTbbgzIJnezQvb1EUhOxIGKTN
Vps3rzyXCOkqipp1/yJN+t4kk+T8iuOIQnJEF0pdiO/VUremP4FeL4HGHHDsuirNirDa2wKCNNjW
SG8z75rEFoOYcoVZAO6nsd8gBBs8T4U5EyuhEqUADn8NP+N8vaJWVny/jjSnGXbAlK0ehb0GoqrT
Efa29tZkWr/DJ1lHboxRkiB2sLSMwQEIFIr/ErN4P87puqaFjQM9Tn5GLw28uyuy7L4pRvEv2DTP
VHHnROUDCEk0umpyCcnytXF6ahZ16aEzFWCCw7Hay0Ydmp0yOt10/nJsr62QNu83ItHjhsDiUxVH
eTsf6jHUPvQynlU25fAat7ruK3O8HZRvX6ZuBvrdyNrmWmF7J55am8bxWm51o8YuoH0e0sgEJd8V
8l20xdq/S3Kh0dpQvxMYkD1ytd6evyzWPyNBiH3elOLl36/49eo3Bfe+TUm3xz3eJtenuHdpzhZB
JiedRIh399lGuflOX5wiOZBP4IMhM4taJkG6M78u7tzM2C4rAjvPejO57Nj8anJl2RLsrtUJWUrj
Ha2D1bsbgzGNQDbxvXcMROa/D8Yb1KT5HF46r5gN78zNQNOOZwmTQdIr1h7tdaqi+aSeLEQODsOq
dPCe+SbAZBxqqIdWt8mJ5Ny5iE6mmnp46oFQhg9z9nTR1JAfy25AuCKfSw/Ih0otHCI/gLVyRal7
yaJ0TDPDKJPffB9iqVLYn8/B0a6RgslJ4cPeiv0ezmnVI13QqLqTA8Owvz7lCl0yWMpfZx7FXN6U
fhXX90Z4PcNjFVeTTL4ibZi93FV2s9ZMUkTPjKuICMlOGUiRLGz7pqqlchHQEiwui0un9rv+qrWR
gDOOlscz2vWBVb3RXAxmWXvlxb0fBIUrx7Vh1ay5MlYRdD2Ij2D25QkeMHC3yQvGv0ncIYIc9860
Rx18YgXJn2UUoDSlJBKb0A9/mxVOSTKOeBe2W6luITJzPTc80/tJnFq6Wnqia4ox4kDPtrj0MUfW
OhBwP+rMx+hs893yWOv+T8j4gsEsUgrsb/o1QsiqN26kwIP6t9K3AZTA6DIlo0r68dhZWREC0FsS
ySwf6NAspC4n6PY+ps+3RVbyCA+gk7oiJ0yBZ6xbLcMAzxaEEmuiVK6LwSHSu8Zm1iDZXJlIWDIk
H7N3SZCYeIPEsOgJGkkIZ7JdnDWUksI8+GJMYzWClihPD6aZUJgD9ZzGtYooKEVoYoCYtA/j2HnJ
X9k6Kyy8X08kxYlFgWtTFsdONfSjS1PFmB6qefUbdvxTck/kRBeEI6ndoxo32eIy9bATF7RXFt/D
6UiFSyN+SsojqavXzEhRfbVB38MLGvsCBMwAjsKefxJ+GYj38Ot/6x5naeNHjkhlZhoRKlXukR7b
utMhuVyGufdMRklf8yuOrbytyQhPQ3gHun00MP599GTy8tXVfp9m+MTPYAKJenpc4Xmx9cqkU5Pn
33AG0H2SJ9wcSvFbWIrfOameXHqDRboYr+KBAdUB0tHyAPXTBpP/Kl1HcB3iVhTFleb6Z1bQkpEC
MBtlB+bp1Lv2OENnx9HmiugnmLVeinp+QgDoUVcfcCL61pATQu/jRjTm9Jha+PtttQC7GaOa70ug
tb6TyMJhar3NFSzC1rsVcyOE54EfttytRZbuxbg0f2V15zMOkCa0fRV6e6ByxwxdDv+E1Zw+b7CN
k7hq8g/A1lmILkyQwoSNvDfYli2CaxkoiJV2O9ZJG0FfL3fLWqVcLpyQSlStLN+GzRhq5GLbDlpt
UkvkCyiys/qo5SPa94ixSxZnnHvKGkZPJLmcgrIV0cAJpW7tiVrD6e+jjCAhcrd9KrScgMsmXQGZ
zqTyVkAcKxJTMI4NJrWE/iOtBpbzq/HmHnQ+IPEaiiV0mfQw+mJ6FK97KsP9c+PmLAgiR8hpVz2w
uKG3AmyQVHklaPgeIeBqx+Z51jdfPxu1PMTZ1/8Wuk4tu1GM7Gd/bk9TSFCOQntpoLSAMZre2Gae
NdS8/nKgxHtPqRcQ4Qy7p9OcGW0TXETmbL9G7WUIFuYH0ieRzdhLcH9NjCDTJ5RePEhipDWjiOzf
jADy6msIg9T4pN8uL/i5gFN0i6V0CFhtRPJwMVkeWdgPLZlE0cByPKEXz13t2L9GsVIZ+wGO0QyU
zoogfOA/HQo9oegnyYSIKLbTRlTPLJvQw9nH+ae/SW11bpHMeRyDdTenm+8rhBWLWLDYrzcgxUbK
DAtWNnI3BJx/1xwq+hnT92vrb03yo1TKtwl/XvfJJEWQKxA+gyniNZVVR7nJ+sWAhiGvRkrhdA8m
POPM9lPJ5me3R2M0O+ijSzZC6aqMbET8+YqtzXb3AJbMHIV3/eXMiRLs9n0Tt8ys5QpGwvQDaQ56
IVDXekSjDzrC/JBqiyc3OF9LUMOmv6E2FtmMX0Q58aUnatnNVLQzD5iLcMe+y8Mv5jpGix6eq7uv
JdeJbQhJMMg0Bap+PxCqeSspgw5npZpANUEO/hdLCBGHFc/JwFrlpy3cYJcLJam/oIeVrcVeET11
dIWmI+1V0TYM6GETyCSntrmfxA8g+vTtq6SiuxzudyaFBqw1ShiTe752CJ6PxIYJr65MuNlr5b3j
29ZTgoZyx5TkmZyelSGNQqBa5/TNQmahbiG5Vf0zFW/k/3FGEQ6m+6xkJvlSnRZfdriqXMF6RXgn
6tVQGFWhXpLXJXs8w0qKnYsyMPsNJPwXS1AMLY983zhT8UQaLUMLLktvWqAjzZE+A7ry7H40zXMT
ZaIkzzxHdp705m0eCoHK4sRdetNcGnRU52wiVNUvAj0CKgCgVG0HjbeV+0TWgIdir1soGs6Ysi90
9SR1HJRdY/4f5vbcFo9IKdxAeJvjip0bv/8QcOmdF0etcsSQ3ok/rQvSGisovvCCi1SXYJAlJXZi
qP8Oy8awQWg375R5DIeDmDaF+YVM05hMiaoYOcihMPbBm3G5YyOK4KvKVaT6td2o55zx1wQh/S6j
T2k1vjqB87E5R0i+b0uIcCsKfJYLuty98uRGF5+k379tCgVrDa+6TuZdjlftD8SOBO7PDIu2Wd1K
2q9WPfGH1GE+j4xF1G3X5d8BIDXO9M5QAD5pcWn2hC8JIiGb+6DlfNFzaLnQVg+s0cnq2jdsABSO
5K1OuE8+F0KzxmOLdY5+hSHcYkWVp2fxWG1TDHmhv1KhLOzsYB1170ilFxcpUyLK+bStAzPXfpO6
Iowbgsnez+jH6fmHtWNRx3BdT3y3TsurGPy09yJLvbwGJ270bopSmMYoTksu2F/uqIkwQ2gN2pnh
ZF4MYTbiQbdofC4Iq+enhkohloPErbxkrxk93m4M4yJYYw+Ua1Pm4F/oG4QPW4hJSCyoTLF/NEPA
Id+P6uTBDiFGd1lYtNS9gFi+ylc/g2Jv2GBcanKZJ3oXWtUnOFVtjLeo/LWIyjqe/umGN2DbnxNT
3y4FvCwPZK310zwTryxiJUBI8o2Wy5iLgxcOtV4JZSNVz/Swf0dmOhAy12reFfRq0dZDL57S20sj
rPNzQm/0OmI6b3K/7P39WOfmlXQocRtc5MKBQ1iAeYkzk0JJqPzHGrS9aHTt8TJ4BSh3lFgndUt+
Jk/4sq+hsHIKDqQloe6jsxde04sMORUQmj308ddcJa1t+1PiGiy+bfrAfSv2Yd9HRAjj3Zsrca3D
WIQtjXsVX2lrVTU+5+XAfRLzRdPJHX4NIbYJE0oHcSOb+khftuG9Tkb42kujzDy48Q+DL/a+VDhk
s5REnuguJbbhQfiJIxh3ir4gJ7O7RmtVkYXQVHQG9X2thZOspKgMDJ9k97YVL276pVfjGizaU57n
TBz/EtJCi4yQE+pNHoIBQYNs/NLKXOrtKeCaY3y8IocJla8CzWJlZMVWhZZN3g9Qdhhze+OppCPU
o+YliiET+HBwBPiC5tQb2gOgmV9PFFwJ1SkWkpzrL9zrZ86pOyjlXPEKmFMBxmNMax+JqQSEiRAI
tmIoqLhwO/O1KbQ3J/qDx0pB/n/vIe7BL5QLzMXDcomlw+Bie92bBn2L7+prXS4fk3mHu7D/aGU6
ig/j7fP0isCsSAO8FXBTIxA8+h8yuQGTxhuHq0X3Omqh/o30XFxxsKbgl08Io73TrT6NqOflO89c
0XbJ280YuFSuQDYtx9kOgc5d9wY9vsIZRRlgq0EBs0b+HYdKQip/NNb8e+6B17qGTw+RdCDePi1+
Dp6F467c7KyN2rYU3rGsF7KlH0tDitJP0zLjdGgNvlmwWWNI+neCXPJXr7XmheCxVzqifTi1gSMX
c62UXYMspKQADXA0mvxEtcy1Q6fe+y7FRmXFswWqKJeZ2I4ar9Pbw6+8hZZnQvP5n8yakT/T6bjP
rQaCH1/csNkK/yp8diq1hLUh2rYAp7b0R4EYBXrSK2Aze6Gz9aDd/ftOrmMlrmnoWagwNL2+w4zM
WnrOOSyRdAuMHcEPFVRPHn+7U/34cRLJ/4vNo5Fd5hZXFyJcHqVRlsz6NLN9YI3i6pYlBvGjFyha
kyW3AYmuVITX7cNqFszECPpxdNlZ5sdI4pfw6IF6aSmDH/ZYQGf8EkgfDKzFtUqKI44KTUnMGeo3
t75Ar9jovvzQZ602AATb7VUsnV0xQMHikYaV2QwPiNwQgoefJfzprPmVDcVOhp5UNY4tVDeRIW7q
H3cseJ4xgtbRjlqpdviqFXocEWjhOutSGsJCeK0n2L+YE3Am6bi1nHf7bnAf60xw2F2SbKiva7cM
u6id5OCJ+jNcJOUOufuQ1VTC11oCFaFkpTl0LsOcl6wDXggfPC4d+vxyoZ4Ze+3JUXOj6065Whuk
RIAF6152zIojyA4FE8cHB1njaIpMDAWqS7z522gaMrLsuzTMR1r+PAlD12/M5tkm5P2yGeVsuO7h
9jkajT0nIAHifX5yWMz4EhXHQ+mUdjrZaJWFvg9yKCIGQXFu6HpNc87J0Nvd4w52Htx7urrDG5Kg
GBgIcd5tl8j63OiVIQkcUtIENyCKASNH7k4CwHpSbkxhd2aWeq3N7IyzwWCK6muuLQ1OusQX2e7N
ME/u/EJ4xFoGgxJJYokGchJuQQlCOcr0PdG070MOJGBhmjNrQdVv81AShzk9/EQITdzIdh7Mo4Yo
PGK+2L6xW3Xme+G78gvEdAk6362vbjPm5IrUXjQf/kkZJLejU1Kchgjqh7qxp66FwFYOO815vhKg
TEWyW5IAVubHlaXPKvgnc6+JnXzKtue+h54Y8vMXxi3SqvXuod2E/zIKrkCmO1zXOjZDsYuMIkJS
tLH8TSa7bxkgKcgaxblfkpThcACjFS3SBYnllbtdlfmO8Wkg0u6WthVRgbtavFKHJeNi9l072aM/
bueV0zD0/pOo9rFmW9xrNvNYomOuP4oeIX3y4M0wJHZlnmD3VGHfO1CZbyugY+si7/ppaF975YnE
yyELIeEtBQS1wT9FKNV4C8KWulOR3xthFBwPKaiHSXM5KlS8W/fgDWN3L8hQpnRkPhQ3UCRPJLvJ
KKhRQdE6Jhrg7QkTjtB4FqslQP7nuAFij4OJ2smztYtR2K9vHHMMrBSLOj0hNAI7npgBKJzPYoVS
O76irPx3O5v7fKmD8moou+7taajHe+ubjCrnyW88OFDHhzfiuCoJ6C90YMxYPim6eafb2DWZRo1l
gfsE2BnmMCkAIvxM1QGwBLQZXzdt2mZsuhYGzdrAKqIQr8MEApSsPfIyHqBmdeiqJF+xlHc99/6A
fUC21xwELMtfZnH0bnQ47Sr8Xhvgk8HxbE9oqv8p10Hi6JBMxlB6rcx+S3xmH5MB7UATnuqgU7+S
fsh99XI5UT6k2b2noP+5F2X7VYqd3m6YfG3KjMWm+MiSlz3+D29U4+RB044cWpmLiJZkFzKzfyY/
wHQT5NZ02ZmGn4hRLfOlXEthZP7ihukYtuBuv90YnK8YsfoA3UJdamgiElPkD/I5fAbHVt9lIDj9
OhtU/kyy7WK2LYLAXOw1njOGjkU2R2xxmVplcfSBZCgo99H8Wp2lj4oKUBp3N1etxy1EmRACh0TA
BTquSkz6W71gYDGrWbi94GgqsT14aghDQK7Oi1jQC7voiBrsefSFCBD9pEnjUhbnOmsiMHpi2acM
tTKeEPqAYKXvOAKj5oPP4bl4M8c3qg2arkiH8afLhjjwO73xerFbFWHQBA9+W3mrHcYPicrdJKIM
QXyq+p7Gafa7CBwcHnu7U9Ss+ZjhV50PiuMMEqPRmbZzsYGx4/TJjn3SdQmk5HVxWNW0c42K+HGL
SyKsCPF/0ZKrLuW4KbQZCee97wpi67DOPGnKnkX2/EubQi9XS7uio9qTMjGIAjTaXaJjfwTV0eJV
b0TyhMt+rQH6IKgt5v3QY82KAzAjPjjMdzmRMbdqD/WNlgVxZt5y/tNMKwG7/xg7+ITE8VWqr1nU
oANuAqCPzCxdcZWIv5BNFzjL9YA59P7PY5T222d2/BNpkZKDkwY7HWOsiba9Vzu+pCU6RToqZeGZ
Fl58CKvaex9XWZY0XO0o8+T+eKMyCKP8iTXA8VMFBbS0wRBNudBi0MSPCDTCheroDnGFsHNklBrX
wgxcRULS6DGCXIU+b0y+vho5FFSZQsS5RI8vImNvtesa0QrBp3p5tmcyW3AUMezKMcbXiGyrXa6e
VjrLLH0kofJwOtpbX9V+lhqwb2EnTb95+7OgS/30SQ5u7tSjDQMXEnvT+MexmmoqJikA2SzocelN
QTGQ1ZxCjszqbSujjxAVHt68MmOIKT5XQboI/+Wm2CEC4BdRvA1NQLnQG7ZbI7cs8Pr7aEHRHvxj
qqxLKeWPgfPrNlv7+I+Z6auu7IJRA6+5zNFPJeOAUoiwFvbnCu/NxJHzBIWaxbqwlOH8BcMDPziS
5vZ343bIcOciqEwSPMZfOgL1yqHEqEMH+/nTkMHWCOzfuJT0NkistNOBRJDFV0kLzLPXm36/La6U
hyBG+lbqZluEer8F7xnNt2rPPM0F5XuOvqVbZTWkA6WR3sMr1lBFRzNoyuP3Ll7yIBrUtcK94XND
iUiPMoPLIuKXmMNKL20z3oys4aBEyQSiT7vC7xvSPDAjD/z2RN4rnUwq1DrlQAYxx/M7VmvFNWq/
K9gaB6Mcc75+A4ai7w2VwOOSsgNqBXMyc+cmZHZOSxwwm/LIuNHOYacBtVbZ6Ltl9pC+o6UDvAoT
8F0PKQM0X5OsoAhLvhGU85P80xr0IAre/GwkeqyhZnGXJWaZTS+GBF7YAVmgW2luJSthDQZn8Uj2
dVeynN27R9yz5I0jDGdEzAExo9K544M24LsyDGW0N9CTIizRADRAe0XTwVgzBB0stRu5xu9sP+4l
muaPJsoDk434DoxS/wcuIft2m+laLffhIKY2wEjcgJNZCJes7grO3FTUxZnPwhb4h82Adl4Drmgn
T+VEPByn0NLQqk0NpC8quMmqPcNR5J+trugdGZXHHTqOLRAJnRKKQ2CyzHldZ1+PUr+Ld3b2pmSV
2rHhuOx9BY36GVrDFWFc+nb58BQ699T2a2ccsp2s4vPBDTQmAi/enPQrbXKSGQVoUSntgUwa1w5J
LvEdqgyv5blezzMiGXw7lCB/ZWprxOcprit6yZ6yFZDZN8RSq8jEpWJn7mAUexv0YCamgBH6sY34
GVinP6nj2KmWuVWDWqPu03w6h9DEBKkm31WJ2D6X+pxgsfi53DIOpNJ55PQuEbJgs1EGytmhI41M
XDyyOEgwEYdpIM/J3YUCKWAS1KMCE51bKX6LS3PGCuk7A2LdiUVaLoml1y16TXgsACYPoTVHxp+A
8octHUkj9FZz61VgnKwMgdyM6erKuRKi21a1U8rDkMGNhwmjni2bq1I9c3fyVFZ6UjaxbLROLJs/
sikAEexsQQZmmq6UVOz5xB/Ya8DxpChhYLv72X+tEb1KtX7DKLroPsANy3XQCYuk9+n7E3enllWs
bLhuNl8BnAMAxGcqFkbQLQaLahEarcPLUX02WrEYOH9LGtkan5yuxt1AHdCQYqiMSbqKEJxBjb2i
MynmCVqu560K1QkAQzGFJFD5g/AMNYuwUnL71JCFoV5ZmqXyLCJJfsUUuL4yJFD3R81GtlTahzXw
T5RfWbFLOy61cINB+Ggh/s+Vjpa2R/J+4UhFzdF8673Ac+QnAeylCXvYDaMCeXKnoH1mu/JzKiQs
SGZDRnkOAlfOvdBaj+WWVp9CL5Rb2wgTw3AauLUJFdkQWErxl/4eob1Zs/Q2daD0xnZTax14sltd
IFMHgmFkizDS5/kjTV5fBnOaa35maQN07jnTkKZHXMhdSS0UOyZ56/BvL8zzS1qoXZlPsUCBkpqq
6g3iXCveum5wO/nBAURlzYPvVJGVgZxMHQfv48HaOPKoVOTRveNEU0sxvf0XMVpZGhcjrad1rMo+
YqoQWCozeg7sXaUK6XfLu435vvaI5Z7IMVzqTKGCVYyGsVlczRVkG71lPKqhvPJHVTroXPgzKxBy
G1/Rt09q2sD/hmcFDtnUIggTA3g0jfUNyswxHjDiWGJX6gIm+QeH2Bgto04gG8mE2oMXQqTaaHKR
Yx76yFs2HBkdxnNLD1a1kP2MpeD8S8y0RDD7Jbmi/bIFBsIkWu+yBwbRoxfCc5KWYJGuOODca/Ny
iqeTe0MWOz2WdK1T99HAwLOPWvXx3sZDeSF587R0KMKHkEq1Z8hAEj+wpRrGnL4HCXVg5R5BQPZf
1qBdtlbHrZYNTO0RnPw1lv6cV7yE0nZ6WedVskqCoEeUWxTcEL0GDwvc93RnceLI7zhp6MLbLgWX
PuTJBwXXndjwaELGz9GXwKRi9SIksV/rsyTs5qtHQNkLQeVG/6//rHHg9Ru3HsfuWkqxsZPASkTk
8vVLL8dLVRXQA+j65rdS6vrDIXEnWso0yxR7fyx3OyJkezPG0C+EE9YhZW/fnsasLf9+bD/Wmu1t
rqATebMcYkRdy2iEdOEVcQSItaFmE3WSVaP483EXZrhX85IeRJH8RI6XeQF0bZMSq2hIvf52C+N3
3cE7pl9FfeY4s6YMq2Y2I48wihyrCYi1pHajrBIvdvv2rbI/5vmzkMFas/a1Ze3n3JtvE2YlSmA2
FHbYAiYA6GIHoJqgZa0l1ELfiDzndn4twr9Q868/XVw+tlPWkvT6lvGKBrBHXW6ZSCcCyMbjUbZm
+bGAMNoyZHLrA6kYc+TGlK4YD1UjDMTWNrT/QdaFEBReMZp/Sri+mSZLTBUz1K+4eA9jxS0Utakk
FwB1+peZsLtxBxrI0W6WxH/6KhYHeyHPTe7XmQsog2MRWRZ8A3JO5DKtt74+zPSneedWypoF5wt/
GAvOVm0JrWGP7v+YoCfd/1jADtm5UnXHjP3MWrotC51+rRJryV4X42J/qtEML5bGTmSoMiqKRlIq
98QIMycUUMnqHdQqdEgmT3P0pptalCrXsQAgqFRy6+RPaRiIFC92WKiimWLVPGFer7dJCOTYg8v0
jaFuQxwmbRjmgqr/jRO9vDIldKLk5al4S9kGR/HPt6mX4pqQojUDNEfIuJei8vQet2zOxGhi5Cyf
zM7fmkh8J8a5COYiIoV1pz68x/JMPnmBA2ItwfHKRdrmPklC3zN2XgNg+6ZZ6UWnw6g/C01Z7NlP
5he8DWnAZEJFW61LGwVRYrM2b0X1p+5lSobQ0iymXoZ6LuNxp3mhMLbv76jjJgQ37IT8OVv6dp35
86XSzX+8dPjUte5hoAuXOhoRmNYNQk+mIX3kZZy4QAwyG4K8pJMU1AK0u8/b95fQjZIeM2WlUBEQ
n80Dgjf7j27uGHvUh3EJeb2o2v0/gR+PkFoQY0iB9tGVo1Jfe9Zys+7iOQQYAw7aX6iXfiPNI6Fr
Y+QDH/iAksPtLrev6UPZcgbzc32gwPTksHHGfDwjNKs+LjYnf/58ONl6mdk30NPvYl9nv0MWVEDA
xbABJFzMsxw5AgaOx13W33EeQwDtRp/NB8jGFt/d7qJ7rAzFs28rZBVO98vyS1V26+vPJ40vrogn
7i0L7lI4L80lnpyFMxsyDrM72bEi8pSPPDME5VtniouF/KWsfYS89j7BEvVMgZQo/NVBTSWg4jTq
y+HimhPtO5DmQzC7gwpIi8IMNeoXHoekREQ33P5rYqxC5Kt2BYn6r80PAkYCK9yvYSizMUtBzpGL
hM1jgtYJ7vmw+dq5Jk+F6etyw5aWRdRkfowHnLVhkng8zRJ7oMt5MVGRW4dXntED38tK+fUcsCwh
T/dWAwRM9JQjpV4YFhrPHb7mh0finj2cBdlhWVtOX2p+MDBB/zd2pRfpxQ5SQnWHWJczXMFPYQaR
q7Echdh1Fg5Sq7wIl5eIER9bS2kY3ciy0VIMZzClgyK+KByaeCQ7Ez7LWaCMhvgxRksoKg+k+CoV
3pjz3BbR55nv1GuxKOB6q/XrqpAfFFvqOfE6HCAQwnwNyKnApghfb7gkWXZZkdV71h1/KwY/u046
xA3poFJgU7+iDevjVe6hiGtn/eJtkHXpehp1vw6vp0iCQH3ky2wbTdkGPRxH45zKdc14ndpDz7qG
LeNJTEHtluE653PfkLMVugVWCEq2joovfpgEAgPkgm8OZiKBO+pFjeA5A/TUj10hSG8xFefzdUKJ
lVdypasl8QPaQBQNRQx7/IXCjOr3UWvc/1gjcOt4GfhYACjxmEVBKe8KNcAUojURMrSYsEKGhsxv
VfGBicKKpyHizDluelmbY6W9MsI3qmI8Tbnm8u1VDO7lXEk0HKKcY7ncSw/cB2v9zF94O7TuaG2Q
YGaMxDLVX72y11q4PjKPUGQ3LkK5ERoWsoGqFJ43a+1ZiTKRrKupnDH0rRfxFw0XxnDSdh1Psx21
kZO9pwxtbT++I4RCxUAk1mf3KAAIqRGpyUa6IjXx0L+UszpNocuYNA5hT8WulpJENEGJl7LZgq7g
zffuc4NuFpF3gdmUx3k6HgfxlMenXGrXYBYkZ3szxyNYi20uWir7thA+iDa73NIGq7cx38+k5hUz
CbH8kO0ZfXHhytdIYYSqBZZqZtLYAxh4yIhXb4+HR32nvRqW/Hn/xthnUGfw0Yrncj4EJrgPzWpD
tAqLNfx9uvW9SWRhLY6c2pHes9nkM5K9BxZVTtfuxDuiJaU4/A2rZDhku90K2DRznUhdIzk03lcu
jdLzUScE6rjqtY0l97Q9H2+hRjMRK3yuGMaRadI/Ix5VxD919kzwoY3Fn5WhwpllBw+a8X34/nLj
KqHhonv2b0M3z2QTrLJXT5ZZGOVBFJ/wuffddCyGd36v44WMSv326BC/AqxA6FzL8R4xEBhw8h3e
5bRpuZIi0ZJG/2FP6/yZTlDjFujSXmdjCKZDUXhkoLB6xJcnMzw8Ol1XfSAm5iVtVkjFTObfzvvt
pT879uNY4CKZxo2NQZ0zsNGxkAVoHViJbkLGKz8ezZIhVZ6KkK/JY4pUMSAY/wwQ23bV9vhhEBIO
rMePiQR1mupnE5jA447HqmLglWVcxTUqRW9kVFmu5YztWCrDVTw0MKTBE0B5mKcw0RrK9ltUJJLh
y4fav/un2wadLjWEGofL21eq+zuR9Bi8+Rs61TkKV0dtH9WXFJfWxv6eFBdXR4o+6EpJ/O/at3ND
lBkTrBp44cdU6IUHbciyhTuD4rU8mgQ5GgMnOwm0nXiayH5/c+j3Mo65JT/R4zvaD3E8+2xE++cf
DQ6uZscoAUfCu1Y++aOvox7yP9k6LjXi+OWOVbPpD13xzhVzXLuhdkqGMuLSlvwUyrOmTSyeo3U2
JhXYNUuUVZApTxvZuU1bl0xGQcp8FcpGZA8QKO9Fh4/6tc5HQb83F83zqQioo4Z614E1FtX9o0Qi
S6KADdQ20atpPfVoJgwa+ZUcFWkrXFKfCs9z79BFNFCMGo0VCJycE+S8G9+rH6f+E4eA/xCJKSCI
WQDXTQ6bJYH+qt/6OGSDUz6H2CNpQrIdwcj2Uq/5YoD5LH5+1W5LpUW7GNspCeEVJWqE9iDYIwBT
lNG0kTGbBRURPPDP1hmUFXeps+dRqwl12LACk3lm9BRv+N+veIaPosM5678RnTK/WBQGvD5q3FCI
T80Q2veQUdco4Yvn5mRsoCODy8L2KMHMfp/dR5obePAOijHdMRHH7V8hsXFiCF1M/+AKcgpEDg6K
gNrQtlRLOA9CVrAPGix2dHPv3gRo/bi3QgfyNerBjvWtlLqU9XBqrzjnFXyIEkd9mi0S5Ycc39+o
GlkODBGwmQbcb0Adp6w/MUWayHJoDIMmyu8S/lqs2lrE9ig5XoIDuqpkEdz2Stye2WUEInztGyOf
g4L+yvWEcuk3kPIidYoo2wgLOAXEPfQR9gmT1XjTAZrdoGwbUKQwOOOLqr7hankiuT2XsY8FPags
cf4GAQTMcJTuE/EaDV8XOYdNGfpnVeob1hKbFI+nrgazQmnW6lJ5V3XtBAkvwVMU9WnQGIqBinDm
BzY7/YdNhzzjop4wL6JYZRGVJecyCjHLrslXhzq0Fh35o07M/6eh3UfFJlq4Qak7x6Ype0w0mUV7
U0cyiOl3BYC3G8L6z1+WNSGPdM/qcf2JdTNeWFNTMU4kKPZchcDKwL+DcSu2rX8Z2esobyT9RO0C
o340+Ong9REu/4TeTsJiFczBPW13N/1TmWkO3eZP3ciS7/9jagsfPi3yoLAkBSMLgT1EoBVXwKxY
p0C6zkoSJz/laHBPgJJRN1wGHn3CqL64Ia1GWkAKyMMGhZnOGG5vVf33lIudVO3GA5AfRGx6jAIC
f+2eYcL0vT6uBpMobzIln4dCtrvQR4QI/Ts7cdKdOjEsg68TWkWVhH5TNTGMNjfSbhsILg215+KL
cUNxdDUhCFxvqlyJwVNn4TVXxdFD/6DeAJcT9bE4HLoHShm+Kejd/monzenTXD76rXQWS+TYwPoP
UMhVYZlNTHUADK0NHwVArim9gsIWmkthZxQfMwWiWSkeXGXOjhyFapcWFT0be8R/jA49hksU+8db
oOfMFFknjqFLmfvsOzaWHpSdCG8GaWkREs0zgWpaltRYZdmH9NPkZ7Sy21NGTFueaWjkDWrqnSoH
7ae02SxFnU6c/OiZaZLD5TeZko4T8jjivcKOvaDc319AnoJZbSdxExJbdW3HPHgzK1SBvqZVze77
Fgqim4f3Fix7LZP5uUA+znFC6ODR7mtIzFQwc4Q2WX5LYXx7Dt8LojZGMxHPzHj6RYk99E+ZFIql
bjMUPZxB7+zbnGiJG+bqXo288emG/AJj+n/a/7QT+R8VNJ9/Q20ZhaYa1dtkqwXdi5qq9K0hQ9w9
uVyqjjpcLlv2QBvvQk32xNZ56Wop1Rp6WNODF+AXP/qIm3lsNHGaxBi6V4/odLae5ESYyuKTB+g3
PyZUmfgwqo/vxXnOQMERuiYMuB6adanDvgkV9IUuFXsc3E4MMVUU5AZR7fx9IzFa+gwxvIaoi4/V
JcD6KJhM7ENnM7Up1R2AZkIRDMmZfTZ6fFpOVu5EFnAFtNMigujGoPUS2I/ZiUQ+VtmSkl+yt+zx
aRs6bPVXDQC1TLQ1FtIHYQCJUZHdIhSHtqezPhemWNXi/xuSka09YZIW3GhDK4GAFsGWBPhifGgJ
6dVByQXCsCcIoxmEemlx9QT6gNKCQMxn7Qb23v2Ome0FqxFXSRkVbrSdPjFe9E1tLOnJ9rDYFwlu
VNnlGRigKqErGQuCU/Z1PSaBsGYZmuxx4m8gJYoHXH+4repsKiYoe4LIbM6mfqqpXKrqLQ8Iy00W
G5dfghww3oSC8HqHVcqSqfwI0TUZ+pADN7nAnUS6bdU36+BMKTLX6XWwAD4o2UuGXVRUWAo0NAkX
wn1nz05IReBi/zuDu0hbJWPRf1ztQSieusDQUW48MsDGlONZQ9GShOCKGbhLZkNtz40FLklNTAZ+
W+UhtmMQwG2hrFG8wZD/jKuntlNt7lExN0UxLNs1HrYHZbxtnAjx1m3qIPy8ObN5B/5m9vtnGgR6
AfjukwB9pk8nhyhQDYRwlf8x8ZMXsC6FgAn0Pap5u7DN2woY50CRwcwfvcXHwGqiQsKTthiL//49
gAGp9pwNOfylKyqfpB8bQaRwmE6aXTmQEE6cG36NPufD7gNS3bL6PCwJVFh+yZoG14Xg0BK7ioYg
XKHG/FeeWX1lb6OMA9fjgw4cn0uzDQl0Ct8L7kNMnKQ4EzoVMBdA3EanIl+qf8EwqV5OF7lUjlLK
5oef1FJqSvK3WrHfkRUEhkXDSVMSpXrvl3gqbKevDrr9fk+dMq5O7vrGUSuAL90AM+dZnE0fmbTL
6hg4FWtIkWD2Mwi0zej3L1BwbNBNMLTsy9dtTnXHJ1DuI27cqiOMK9+cx5kMRcW0yvDa4AflYcTP
oKOI0r1/eInIBmkri2prTD9REp8F3g0bk8TeQaIrmJ2LII3sJth/PysHHKqI7sCqU3e0Iz+oeZ5R
rn748VnEtzaqqaLhh05F7I57dP0O5HQYVEpsNnHKiHYObd6x6s52WJXVa57eyK0tcVLwpzjwfOiz
6idyxJWcGIeFUbA0TIFrikAP/KsP51juBqaWKTXP4IysXqjlZ7V2ynR9T2KZMvr2j7+D1Xkw2M0R
GiQYaKHUCPhnzGWtYCVPx729267RUjuwJHMG2g49oYN+JZEfC89W01EAzv9sMUGrImaw5MFTI5RN
Iw/1MRTtRA+y0+5sMCqRvWlAbKxSimh5q0P6LUqz3voqcWkVAPBCoQMOsomHjBNCOPLRrEs04ptt
zF5fLPPqO00rPUMV15rTDRr/iRJMO1eFHYBuwrbcynrd44b5hMF/126H17dFyVYtkU6UMrgePTDS
2qQTf9JZ4iHPqAQsQEqrMqCFxY15dHLA5zj0/Cgdj8Pm2i7sh3JqyE78huovlL1SOFF7s6EBf2Oy
RGojA5Gzs1R+wGdN8ly5n1OZa7Q/nkaQZ4+Jnb92t7MkFllK25lpmrXd4yhJyzVP1LsNDhsTRfvW
opMtbwKTsY3tknX5co1P2NMrNecNL7tyX1SEY3Jo0He9rjMrrPHH2KfnDoSIKdiwMyfvZGdaWW2/
BqLGzEThqANCG2wfUelwKS2ELquX7yMtJIWTwcb9kHynz+tLHvBZFcYww72GkvmZoME92ECziYNt
SAWzi3yFZVU8ig/ZqjSpyiVx679DeJzf6PSc7J7cvlRGPOJjXSGm/KJoPBAil+aXljZROe4BbstV
aL1ANyUOXTha9Rtne35Dm8CH1MaAykZ3+qxTvIVhhPb0nb8GepaQY9CkereXJxn7CJpdNvPNCF/p
IWGCSYatpkvxe3fd3joD7aBOBUYsz2Q+BYJfCSsZMqzrXEiD2lB/++K1CR58aFJrftsslA64hesA
MUHriemb8cwT3sw9Gy/HNU6LMeuIBCd79zMnN9M9Jy5u8sgytBH+jH/M+GEgFljD/g735xD4n1RR
ndCVprbk46hZeN4yT2C3IWYuGQV5IZe0eBWRNALZ4HXJC3lK6NM6QGOSQaFLxGR6iQEYGgM/KnNS
B6136I8jeZTeCqK11RmoBOKiSfOA4PluXQyjBhj7z/q5l4sKgp1U0E5k7yz0BXLuIMnn9kEAyAHI
Qsazh8FMXqtbJomYoFItlvpimy/y0Cm1yW/eUxCBLrEPZl81icAzPjRyCVTg23URqPa5lE/xMxmD
OhmtKnSX2HQ91t/4RINxo0UUEpb5I0qwQ4kyOJu+A14gELrvYXksTug5W9AS8DmN+i4nt7hLkXso
TlNz2z6f9t4s8w4E04ncmjTboi3tbyiJ4XOXJwj9isZ4gdDg8V7BZO5o3jG1zcPGbrqdiN7tQ9VC
A86IEiTuujPe1BvbNEaJyjx0pEvpBuGfVALLeIb3P2k6ywz8DISul5CE2P0g5kI60Tz6BvddUriz
+fBDy8w/CdKpqTYCVBytoNEJhf9i1kDQ713lTC43JhRj4VasI0RjOMrRisSocHQYv0GhKsaaC8ll
D1m5wJQZ28cBBlH8S/d0DeSvqdJSrvqX0BVF5vpA7xUH46/Bh9ip3lWINQegA9B63uKLo3LMSihR
eVCzT+b65L1/zwCUCgEy8SkXlsQlnqsc0I0cquXik6VQTuTfcSMINetrWEaWwi3LEB4WEQ48O7EH
zeKdSD56yFoyKEb9KylZdFsObS/oGhJ9GuACN5b3PPfuze2Q0djsvi8b7Xeb+eFR4gs/3B73I7e0
hUZ0Lf9iDJKsiJ8rW3Zx5PIs8CBLV/1EncsFqLl/kGF1FjPl7BH8Ok1xTrrWvOOFHVhbQVXVdR7W
g3XZsBcw1ql4lqIqrPdjOIbVfYjnfE4o/VleCn2T/Bq/IB396ZuNBBjPSnRTmOLOgbjmLftKs8Ri
u/2i2CzN+FBH8Lk+WqD+9IwtcvT5iZyJ8DNAbjnJ6yhmlUKlPCgYIINUPBsuUjRqdHSids0rw3nw
YEtBfropUddD80uNZJzHwthV/XHZUFNJD33ZPr5fVGgTmc0DCufQwnaDCbQCXoQ35Nncls4XuSNR
73C3/A9MAENTxHtSDzqfd3SOImXuWbkC4eoUh36AkmfW8mWKAXi+meBQjTNxIFTEuQnXndknTQ0r
eSJZZElwpaLYzPgf5eUT90NiPCEBZq0Nw506ZWejX0Ibd9SvhvboIM4vilOtRLp2nLzbUrWsk7CN
PThZEWA7HD9S70tvPluW1YY1fR9boRd+CCHUkJ5lUlfcowpjvqMkmu7JhYdMLU81ZYe8n7TiJPZx
u8RuB54WcFI26uDVOzfjBY49VTJDnZOgEw0Blo7hewfMWdZw4niZpkO5uGVFVqCNyDV45CRoqroF
YM4fhTh/ADQQztAEa9iQ+aF84yPVQDjUQr9R048UPZmAscOCBisnfGH9eMu7ENp0h2SPZJlNZWO4
cCcsy3dpsaS5+W/OYN/5DUv4GQrxrdxwjJ6PiIg+mIVxE1Dc3BfSmxz+frxBiNcW0B6QEhJjqPcM
E1WCY34YYOxqwvqLt0mzcakY7nCVP2CbXdJQgqZH91YBk1HqvrDvJZOlxLO2+dXsj3qGB4TZsamn
K2iAtoYOMHD40kD5qAtygic7epqX88HD71Ufzl8ksJY5xJHYt/qnxiUojWbxmF+u3vzw25iht8Qd
oyD7JAtB2eILqv/5exINc6B9OHgojY+PrL14clQtmRHgypbOZmtZzfxZO9JjEVjOGzjS+8zqrWgS
fb57nVR3jPC+F1qPy8PuFLOpLZ1PBJx5vZKiTUNGFuRBcohIsuNNFMzUQB610FGcwhG89QJc1YfX
fkEEti7Us5nD3zDLLA14KcpqypPym8SPhZoccCOCjlpCdKgw4WH0p3YyoNQLAAcYin9qBmJmfViJ
7JYEKVUOfxxzUQpXqHFLRfticzdU9Ts7eDhWOOhn9rJKMzAsxSfCOWwD3Xwd2ffKXQH08V/0sstD
aoUWVzj8Z6rrOw6iC8RYnTtV6oXIJaJVOF9L6n0LYm7LHMVnStAjFhVJc2HB3oeaZtB7NUXG+txb
NtmCl2uesvzX0MmYrjbIl0iFxW3YP0OqT1j8kIZlaxocba1xTh/kPRD/4MkZeLFZUclXVUJKAm+N
v96zvti4WZ3Psi9chExAinxVIIkUmTJaq8lBuiw3X4/oaEuaaOhMqD26/u1vbttCQyPox3CYI0kf
Ez+Wof1Q2fVCVxSV0DDD80FEnR0GZdApbAB1+fRmDehum23obGB547SX2CJokVAlL08FIt1HJwua
pZKRrt+8gv6zcCYml7ouy0VakicgeE1THOcStBnZWuHvVMjaK76B35p1btPVwKlCr8KIy9mQDiAo
+HDODNENDtXWUiqR8AmGpa4dkmWVt3rAW6+95Pjnr6dsYSJyfPiPQ3gyaJfiZJ1mGPO9FKZiAU9Z
5o1lZGwVi1Rylmgyt5UnyeH0EajxGdASHWGsu86fgR6JJcYSVB4lzgasupZKFyQJJ5kMElKOrNIE
Z4DtmTpf8eXk/NHL1wUwHQA9MOYxAKtTHwVKB6OLlvJyBu4rI9dS2p6O58pYYMuwUJTS7WI/He7r
JdW0kSDZTHtFEVQ2RqG/XZgd2gA40XA7JVSzCR8gjYyrztLitv16uZgWqFMkIE89vs+IOlHkaBoz
wW0BWoaOTc7geXMgh/hJdV/pg5hiqaVn1dY53U8juscvJzEovmoCWHh4dMEeugJKC7Uk4whNLq2o
Dg3kCzC7zLhvgUCdVfOJM2G3JuoBLD+IF39IxR6uapR3VamqoTLeLTdceK0Gc4VuCDO0jZu7JrSE
oulxWwW7F3F5JBwBwR02OwI+fHS2xSaD9AgTOzHkXLxinADjz/tYcoOzH/52YEleifPe34JB0wsw
yM7a1q/uaqtvq6DZOxqloUJlZ8+L4pIYkPa5C5BcVkHzLhYr6FxNkYRpN4qoqV3tuQ4v3bzLZYnT
UApDIp1b96GcH0SJqbXRq0QhulfxrQIdNx9g/BRL0xcpgW8WbzsOUiOMLPMQL0spcnJGt7M8WrIJ
cCb+LTjNXL2PsJaY5qKlJpakpaBrRAWu4bXRroG2bEmJGsocpcLJU4XIV7DoWKHHtMCe2SUPo+u8
2YTNGh3oX5YlZodyuPXKhB7fe/Zk12RdBNA8UmkYPKMOs5rL4kR/bGNzpYM/ie0HJGCbiaSL5vtW
eaO/Svf7yLHyg7ANHRZTdBAvPkhNc++H29h/QnCeAmgJTctZ3MVeSE96kONCVw3KBMw30JKVGkgn
8yPp/VltZa9itxhXB/hllmEgZhAiKCnHG3Ro+Z9PrVEM2fuhr7VPjISbspi7dQw5xzFPUXpHFrd4
un3rh05sJiu9vXHW5NYRX5/CqYuKSGPjgQ/0hajj1lsFIXYApPqY1xyUs4hWSfKrbaBLEf18hQVl
vcviltPyvc6wQXqD8TgsrglljCdaOi031lIu4E7yf12KxbRXs5JOmnfh/loB4BMnwy5j4rdBg7o5
EtzLi7gWpF5fBxQ0rtw+S8U1fYu+BT6AdrJgRh8j5UhN9/mEEQIiRkbUNWnVZX+6P/lAnHfb33jq
/8MC6iEYz2aMYGNROu5moBuQhFt0XBQcadQBrQlvYVM+oQTRvAn7OQ7dPKoIgaGK4Je6Mf+UoArN
sQOBRw1LTFekVDBslKyGpccJrmqgjq9ahSj+4aCJH0yr7f+KRi3z0z/oQiTgvKWCDnLTnbZXPCSF
RNdrh6oMPjXmLyPXXRliGMnekHIKAT91QOEbntqrVQoU1piYz31jMlxeI7pVkKbouG2k8LWpdCsi
hNLNwx7uwCzPrj0gkQmzL4tyBIVJfR98G0a6GPrF7XUpM9HLKv3RiL7wF13giAlEBWmz5OgEgSJB
wj8gQy2PI854tH4MxJ3dRYMPGMwUf49GEsOAMSah0VjyAFSbeGRud7MKcTqldHWWquVnN2iz4b86
mx4TUxUaBen45RDGop/hYacCZhcoCTH4giWXku4CTsq9xopMEd2E3PegPDvSf4gxhQUcAOXrU1wH
sBWl7WSIGevuAK736YCRjWI7SoMraxK7NRVuLFJ+A7/ojKKJJCJhnDvwuMWSHLuc4kt5boXRIKIi
joIqXS6uZimzV5kGw0G+twxI6GK4hmEbynmF4/eRiXGk3DU7hrmmPtmC3EcVT42Bzg3c7fCg12iP
O2nNvnrJxuzxZs1m90EnEErAN1BvlSDBmt4jYablRRX66snRx5CTYDuQEGYctefV6wDqvjTmPw5L
5Lc4fCyljX9bEbk0tIKn0iaZDoMQbf7cr1RMameV1XFaVl2Fu4eGIAcwrAO0/XliCWyB33KpO+Pb
9wk7RvsRYf+GVSVVBz069zeuOh3+f35j5Po3muF0WZsfUSGrrZ9+SGV9UuthWkOU22Q0ZqNwSmuM
Qi9hq7DMCt7wJBqF/oMXOxAPPlXw6SpV19tuI3iAe9uxTbFGc6FMnhWUUo57M3nx+8BleoRwSG+H
b50VdBEoT8R028V7e1pkLdRD+T9zMbaMrjzWX3QDn91ZIGooqWimLlSgQApcCwCzBZxx3AIhlaq2
EDW7Y5T8FDU+PH0GJr/gNpb+gRM2EAQ0HIyYtq1mIwYoY1qBM+DoQ1nGqzN7mvnCXpiDw0ubUFce
ZBvsJv4LBbBphXTLBVbKpSbM4ZX7NxfpBGQW+YxQtj6C03vKjj87v5RUm2K72TqjuBlJUDAGioZa
bxYOWwOn/himJFpN3+twQQZD9TM6eH6IObauIwoLp4yXFnyzD4uRodpIxKTs1uhDZcMROzgvKc1K
0AwtzuBCGXDOwcv5CnujU5ugOog3q+1PGSXBNxMukbWLnZKS5yl8xT7Up/Ke+TvOnIzIXvrGjvnq
n3Jwet8j/+q7EzCSHZnzFFBZE/mvA6XwLX9HFxhPfvURiysmIpLzEZMundW5I/v2smHfXBliQkGv
0aJjcqYeoj2bW+fMx/g0Hw/LWPXIkdUHwVe0Izc8n7vjetqyjzyCak5mqpFiaCy3AD6MkXKiD+l8
5bTTAeRHuacbrMjDctSMzJh4OPlD4dhhCH/MmtKUiibpQODWb0D0rzQcNxSf8Ubu0Skv6/1uPccI
CI7KKdS4rv6/taN8Vb8Ovb3NEYcX4DhHrbuQSr5JtRmi90b0rqpkEl2LwYfGOcXbyEa6oiV4C6D7
Xak3JLZ2rbB7HL2XBkB75RBB2UHgnTfT0ce8lyEMjfe7TfiA+EopkV3yRoupi0uMQ/HzJwpWzdA2
0vxijR4KIVa7YSdAsjklMZan6PnjkhpPm3kBN9bqnl2evZmFJB8C1wPdZBepEtTIvm2Jb0K9cYZ/
kt6hKsdyHHudF10nA34dx2sRBn4+yvPcB8kDxP2z8urElsQGuCtwxPvy1ZNJNbMzC4wvevEdTNWK
sIIMHbgRaNwe2vuolmhNnwNUcKsHoV0dNob6yF1QbEIWBfgTlF/stQSlos0aYhjwOr+RtGcKukym
fpIXK7cDcqYtFn9mWYzIGz+rUonG2raO+M7mTCXrwnWneK2pO5Mafz85fZfmyjx6RoiICIdBD3ii
EllPPl5ilwa5p7c3N95uAUXZn6mD09IqX8A6N3yib+ISvof5ce726Y2yYunQ7JMcwEziUjRZ386K
Jw6xOC6oCxGI/acrMp3ADMqklswFv4YgY/dS1Ubgu5XjawTocal+Lz7RLsIC3VRyBdNmV1a9WvFP
fztWkhfhwVKQnM9Cn/8Vp7q4ukSl0+jsuNlAzYrG1XE6ECqitVVQAa8gmwj9Mo5raaiSr5CTcmrV
zAme094MZj6uSH/QAzWeJ9PkAov5webiufQp9ylO44vzxadGzXwBKHFzyCcAgCBlMgDCJOTudl06
LOsXr54kTuYyUJQogRgw4xt7ThWaBVp4jRg8O3YLQNPLfPp/rL4d7lD9liRBAGIwnFIWq/8D2iSm
Wt+F8Lnnxz4F8hV1EZirdQ7zzxtGlwc2ZWyXMVWR/PW0jkH1h0TebrWtoS0i86Mn9h6SO821LDey
C7kT6DDjvTQkpVr4Uv7jHJjvclmUqqeofKHWU1GzD/T03NkmnRLlrrHQgB62eQxqmNtgqdmHEXys
E7LS5Vd47iMRZq2GgM1F8jaHAhrhIJLyiE+6IO2jBvL/KieT9Tcv6WsLTulPNJLlqQU+S6Eyl8PJ
0mtTmg2yBrCd1K+db/H5nqiMWY+yMxilM8+/l0TeaAbw5/d4JOLGh26nZRl4+cORNWVWJgyQzEWo
3yfVqHW08R0xIm39BT4QnXYAoTSrwb42YhCoghpBeXWmccSJxFWWvSLgDH1kDS79+fQQBfOGISIp
iSnudNs74ekMfgdA9ZUkzXpCL43/Gfbjhy6VTjnQ/GdnfuHaLl6l5Qj731MPe4mUQJ4ne0SU42m+
5F6lq30T7LfIM2oSd8TYquKPXezWiAE39TBXEJjk7+hvJbjUlneWfe4HfYINozFQdajb+fU2+54Z
KreZ0pigarjmnI9PIEY4uG71s5cK5u5I30wL5EyDJ5Jwmlq9JCAASKQqofGwuz2eehP9bDjTod+s
IqgW1Hukr65Mh2EFQ1JnsNHiNhCRH6Yqm17L30FxO9ZgS7e0/1RNAT13yRFmAwFzVrcti3mfzxQA
Vux/urcIMSGjtToHHt8fAszniU4m/1EAeUuhQvjYWNBK4qqb93khC2/2c3rY22Oec40GxH/21jga
TXVRHMBzNru2e4HOz+xrJBnGcZlcMS26J8mdYSuaNU8dJlvr24DrxcrAgP772EdIbyOhG8drypxl
2OO5MwgMrw6XpPgXcwgmsPi82rtCs0R7NExdWiXWIN2U5X6wnhXf/xPTph6xFcXVkoagG8BB4oM8
mDFQjnAWDbx01+BATW9P3q0Eq41TNOq0zjUYbPX8cPypHbv07yKJeKdLE93GVBBRsln+M0mcIJw2
8rRBql2FvcSwCcvPhZiKFaxB9KFPp9YWsVWhaZc7qA05f1uYqxTnnd4TTnjai7QwllDskTz1+mVw
8TPvDpOb0b36LTdkvXyvmOvPe+PHoUN9JuBkJuQowWvelFz83utuhbgjzQ0Q898bbVgACECX/R7b
kAlATOKfgTkzyiQat8aiXwcE1qAidZIyeahIKxezehB6L+tK2L8+p8gWofcBjfKLMv3rnC/6slTR
Lib2Z+K6zLMQKPnfn+FNvmICxz/1uJq7N6uZx5qZXTcEMXINUjlytl5IDm8elMs6RIxk40Gl2B5+
+JlvE/De1f9x+wccOrSyg8aXkBdSx9GuGshd+/nu7Wj3hgVdfVMcfCpY0gclFhEW5Mi1zjar5R1E
c/H6nTwefRLgt+KbSZF/1IwxNKJVUMx2Z6YUMFsPD02Nqy06ABnifx8/ghT8zKyQMBw9cw2zBnhL
AZ4cPDE7FkqpD7B8aw+V2YDMlz6H05oaRjp7oCwB/CyEkIcFwtS9snqdD0H4Lh5nWDUcjXVMMsCJ
AruAzzPcWESroHWeyNaljO51OFc0ofbCMY5iHkR4DWPvgTGSrqn71wXPqvGRe0WMBZgd18kbeKMM
j961aUQuEqOyk8RSlYm6QgQR8gOfgxcOpmzlfUai6NhrdR8K5ZORRX//a2guBgYa0Azlt0wcb+Qk
thOgnwyfQsM31PuM7V19gobLYiQV4jxKMD2RXo0p44CSG0nmgI9qpOFBbj4P8cD/jzUYXHn0MaPu
eJRZ8VvNVdhNLNq6iP/NVh5YXPVgPLc0U+IOon8Rec492OwtiCsejrT/orkiQnMdVr2XcCMoN4tB
9/Y6ymwHF8Dxr9ANfuCcwjNqQsEYvxHUTTEh6BPOgAsHDz5qTt24UPrLsV9lD5hT6MAoUG9ow9Nt
FKoDC3BDet2HOZ4R4WboUo2rnyX0/e8IVswDTPWiZQwzUB3dWkumv2u6OstuYItLWt1w/SCfmPo4
gzoGXlen3ITv6L2/tiTjvUZnh6kWBuZLkllxccMeglNxiQSQC6DYHqaTjlCUYyE79/+vyL3LHqoc
LYLWXcuKgQsOizwPnA9dGbaZiINMdqh/htuiLPzlzu9dnQFMifJVitZaYhZW/e+lxI/oZGg/wx8w
9FJVpMedeibizKKsZJLo91gLcpkUzNfDArQ5q7FOht4EvwtWXUdyfLHb8Pvbju/5iuv2hf96eJLe
yM3gWlS86NMsIJN/Xa8UmOUgZmkro0pqF9yVqrdl/d3NzKETFpW1HFYd5erKt3vkx0BUhwJvqpj2
8SNiP9ZWx7vWouWd82zU84sph9mnNGEZfy+oBOj/xTcwuipoDsypGC8F47X49BopnuXZcn/EfsL+
km8y5AVfXxZZL98bH7k2zJeP9nIyb6TvnfCTAcbIVqz6z7u+raM3Nd6cG8VtHz7rV623eSrBQWWD
dGIC7J4Nc5PkzzvwGJPAxsdmH2tXGKcktMquRBTFxUAEg+wRBbWLncvtbBvQekTN8Kbrs9g++fba
rnXXTcsG30DYY7sscNMa9YcVFgATm2DedSb9csq+kZI2BhYgDVgLSkl43gm+xT9PBEM0xJPSPwa3
Ic8J6BqzFWEZZAu6OaGe6iKcNK+hJ+FJfgOlVdgeKZXXalpd4k6rGMi0ENF3cwtCfFxSGa+P3PSj
0jSOw3wptJSAjnQL7uL4FBl/68HZ7PmJyybke12zoptaUReHC6KyytqJ++Y9kdi8o4Seo7US3dJl
NRqyAhAb7GRens/OcCQCG6dgx4oAH/AemMgUGqZNPLWS1u6YKkqwSCKlycRmhWONQ+UygpvJa/8X
wQqKwN4YMULceLuRmRiXZV94OFLCP2+wU2mQpCIBU6MD/Jpx12PfWP5BpdTKk+RtT1RWx2KT1gh8
nCRa+O1V0RRyVagpHswMb6jBsGVJV0NPOPbkt2u16ZbPKJiekufcNB2LoIA1ApFtoR0wPFGIZvl3
6W51o8X434Dv+BARmFJrgS8Di655iqpmZuOqSRBp5NWv/LEHJgwQBQzcb/S5T2btjj8kqNSZUhsN
fPEmzdWfIEGONzRfJOPcNa6+UxZttxh1n1PuYiT6IgRZJ6rh9Jp7lpMH+tDfKvpiNjSB3UbtP+BA
S9lBpJx3MsAKLgJcrtdqUA73t5filyRhY9HvJIpyflvPz1AIRAi1aigF/sv3kh1pbBiB2H82adko
H28IK2jzJAJPAaCMlsVJA3QS6NtCb95Uq+mDbYcsJr9RlNgCfRwJGgovbYmm2Qe9OKXvR095btXA
UhduJg9ZtbCjAExrRXWoYagtiXjPTE3cyhxZoMZcpqhGZ8nFSnsAqXq9w3wlp/bPqrOfB/2XkeCM
Yvm7BzmeNiwDcTww4QMgV68akhVFyB/YlGYA19NhXwa0EqOK0i8NZVeX8erVDoLTeRzF0UrNIrL5
CCH8MidkTXMWvTvKKoN/h2aUxAO1/A+nRZ1JmSU6JsFd7cn5NHtla1GbA7uIYCQQ48BL/R9Z+B0F
Y+DxNpPG142Cur4XNVCEdxJF1pW2MTVH4X+wnSrQcAtwyET08U8Yl16nOc+9yakOvqmEghlPrWqb
rkjHIc668c76NLjHFeGO6u9lUmGae6Ectb24ejql6DqiScdlyzbVJMb+TwhXlH9Ta6rLMZ1GNUoS
ogO0JN1t6r1TdcPhAZvgbMyikuXsSwhvVabdbUL/SfUqWoKWTbX1Xk9u3mfZQp4xFR/gkk6lsp90
uQ2GChI2Zp8Rk3U7A/00u1m2OMxdvCJ2w6diWfJdUTDdA+6fLYFZTHQs1bE4uyWuwXinTjKZNnUP
CuP1OxpOMybOJnzP3pQmr4EJHRH/UjjYeeflQo6rfrUCxi17AKoggZhI2tytsJo5PhXlK5UovpVE
mjIrhWu1x9d5cXCz7T4qRT5ZF6vmUf475084EJlHRqpwVILzsLqmbQNz40ioBg9xe5FA44HuHlOv
GeT5BNdpFckg0wlrBm7pg6cUWy+UVxV5OJ660DDznZnQwb8xcWGOvnIwaUAXoqDYZCTQX3di3xUP
2ev7z2zHOqpqgPEiowfTGiAY3yrZJxyhq9bRo5JewEfY2QT1o8FgX37v7Rr1xfNW/JpEbhRGplU7
MZMzmvU4DDFLg6j+W3rHr6btusaYcKUeU/v5TxWYq9HREICy1fmTC19NNOW4TmkBiO0mNEO5Lja1
xN+Ro6O18CVxIv11nOdIsJPRqq13i2gvlKCwRh6MCvK4PrGm00sxwceS8WncXiXIJeVzxeimLBFV
Kdx3DuR1It5QpCa+fXtsRmdYuym2MYPoZb9OxsizwtbUtzlkR0QjvYOg5ISJB9XBLEyoQiBwrhPC
lMVXtxlTuO1GhC30IibUZYXjDsFFR6h/WEMrBhm4gUC8wHAW8riUS7AVWS8q/vp8q67AOfDLHuuT
3yGWtWOxuBj1KDN3arcvFAn1hBaOG6456A/0mjVcZNfNo+/PwuHhmZlrLEbAF65qJR4dXo22A04u
sytTL4OrFaGao/+8/CjS19GZlOi/cLx7Qu5Pgqguj4tYuP6xdAoxWfzVKdAeu+Vsc/tBQq9Mp2cO
yAh6FG54AzlPALMd/IEEfrO8qodQuF7wPg3/vDIhjQePwjHEu+f7YLKrzPj+ctYE0UuT8SWzXQuO
qN/aEbfo0usnmrvqnibG3k/IRb0lQ58Xr44VTJHU4KY7tp4Is4SQWaLeNa1K4GdaP4mCTmkgVrah
CLS97oH5Y81zpOvTHp8wZdDvLWwTka3x9/yQovDMC0qo0NXXt/RTVkq1wQURyO/SuGQCseGHWbcD
683HLMWxN6L2ytxM50xfJ7LMU+SIocKbr5FJFdddVKNbgIt+WGl79SXgcaB6D1K7esTTpRttiBGG
Bn74LYhNla9iD3TnhaQAUPNnXrt2Yb98mrzDG+F+oJvgHUjHIAy9vkMSZaIUbqxbqh/ANiNdoITW
/TYIJieqqfcEVmQKNPCxHUHqYmN0875UX+mkn3IaAd9lKp/GWSZGQJLS+285acJM/2zivqL7Ctxn
gHSCVa4So2I+LCzGncySgeTj/RVemfCCbeQ5GPOsyVK9vCo3yRXvAo4vFOJw0ri/bIyZp0sEbTFB
6rBY9SndfWF6g/63Euey9iMeBthZu3KOWmBsWpgu/J3asrpPSfgkgfbnGySb56MIgNmPP/K+gHb2
rSzivtAxiTrfPoCudCRYCk4dPOZHf0FNDQFCwYaWSyA0I0XTbLOLqVLMtphN3JABrQ5sa1ePMkLu
saHQBWEBTgjqZo7lpYTnJkCCVVNTyq8JVFPNJEULC2VWBCFba0CeTbbzD4R4iNvxDs5zqqi7p5o6
leQF6iUZPL7u60TXYa57AniKt3Fe3owaqmpkMe1+qoMWukKsI6qoIopmGLszZL3pmNzf0S4rCaH5
EkeSlinZkmI6C5zP083pe2lsansXVW7wyOlqOPbZE7HE3MWmgYncclRk79BDFGKK8NwdAtzzQuYK
qXac2FTJc3WFfCRR9rxCrS5yNPgTGRhVAXfuOKrweoEovQHp7lBDAaaojEEHzhYZz9YXbCqNZnM4
SRSvE1Oa2AYiiOYA57qyS4lhWSg9AFb5XxYk4XAenollyr4K7Dzgt0uoIh8gRfQdxnnpEubCPml4
rIaOzwqvEgHIbgmBjKT+ZEZlN33EYVdjeZTzFyGIFpdPI6KK/ssg75nu6OKESIdqM4cff21KNr50
KA2Q/W7dt1ymGowZnC464O9bG7EO++23jkgrlFZTWjoXQsPlk9v4msqZ1ZZfnKJe+yFbs6ghBzyy
gsNIC8Lmnu/0M/GJrIFwTW/NOegcihl+ZFVWFDAWtwYI/utg8DLgaoAVooEjIK8GTw3jS5rSWfzk
jpqRH3WWkd292dCwS3HIc/AR1g6cNHOtGUK70hhDQkVF+t1DAj3Il4wSJD1JuF+tamp/yf4e6zjF
423lyoJ0zeR/m+SVM6krNWEOhWvT6e+VqVcDUxkMxSWwtELgcpgiOltKDnwQ/ZfTDkVtmUJqlXzO
FIuQMSRBIppB5ezhxbQrZ7Z5JjdGG33z1p/7IOAQgpVy3IdcPiaurvGFl+vZFapTG8fnGBA1olU7
mGrh9vTcx/esY/rwgiG9UZRxizHMpOqam3kfykhg2XgS5s8BLmlToD0ltFIX0yuImAZ/NiaVxt19
UFtM6YqFcKklFG9+C2H2+68qVlRieBgLddqDvDvQ9mgEKdY2RmMrz8NMQ8+KFRkkFw0z+Q0AvL0S
20/MKt0ss9xA9V+gkWSDDx6aHRpFQjwCTjE+47U6InkR+G0rhubxmD+gB5MvFL5MTI4/UFZQr4lr
JI/bGGpi/IC218em3zMz4206SxhZjUyivp7DTD70mOyPNSQY/808Wn9jAj/nRzwdPXcY5E0R0J68
MYOteg8uDxzUpipLaxaWscnzBJcpcBNqI+4xvCBjnL5TONO2ZbOPUllJBBnW3m814I/8nsj/uNFQ
6jX+nvunkyBRd4PYpKU9faJLTueeXgloWQoKNV/yQSm7kD4H/hSRJjEpGPZlCoA52Zt6Y7WafcTc
Q2V4HmYuph4C9mxAOJ3/6qjDy7PjwIhfqAVsUbfPyFFWSpUJoL7QGvpEFtpMZkefRTNQRC8tQtvS
pF0fjm2didZuaoP/29I4b5Tfwr2z3CxxPUuQ/D3qse+5ghPS2lMEFSnUAbgryFAhZgzGcO5j4AJl
k26RWh6uj5ViPDCdyO4XILDuarZlHU3bkMSFYwsnUD1k5Dnu847MfRnXgsrqxMufece7EnVt5guG
49JN5bcVQcP/6R7vGuHXGhRXfoE6H4wOYuqbo1zlbWTreRj3ur2BERuFeADrXEb2s0wWb4N7j7/X
djnPJpVvCNNk36UWizJZ5IJgLxfliHkZSv5FtiNDBn8KjJ236oR6N8Ljwwru6zhgN2/Ye7lkQFIu
cs0ZRhZZdGHvXDIGTUlxlN8goV4/RNvLKp1NYXzXzXMB2PlYEg72UMqmBbI4XUeWznRkeBYNDlTx
eYeKcbazW0EQSdIQEjuu5EH1tIE+UNqXz2kIBwAgNoAuAGMUPCBT55uNMGdFTFP2Qs31f1fsCIng
utHrgkcPZQrrisQQL/Uyw8V/phzLLbM1kov75H9QfbLOBx4upP9xWJKXCbX+8IHDJI1kOKfCT/n7
dbQtfnSrAYRsjwGIfzjB0kvCEe6UjJmpd7LEcu9n2fSAyMD7AK+JdB4+7gE808mhHdCRh7y4fBZx
hhPHRHwu7/2N77MXkJ62Y2FBmvlZXgNiGqBfSgE4dseNFEql2s2d7Q5eO3IEiUxc0K2SVRIIFnzj
L72fDAClhLxolZ43Me2yQCJeedo+BEQS9yENnt9jt1E4uKtUh9KrQ/pZPMwo7BZMR9RNvXqXWZrh
JffJYe8TETIt8CKhpQG1cF6pD5GgJX1W5pRUZvHIY8ndlfO3ubGs7cE1JpgEin4fZHula3YCfQdk
M73J46k52V0Pwb63In7jPQp+5Y5uvmKDIFwIiU8viuiS9arrHEdiNRvwd4s7lpSN6yNCpa3ALtCo
iQblDoJ/w6s2vxaK/w2F3W0Jp+IfJErjb/PSq+gb4DtBKYcNlXx/KmRRobfBKZE0tW0IBUgTVS+w
vDoKQa7vivnMIE8HSzwMJFpI6xHAQexcANJfwTa2aAstGRJJfdnF66ukeIXLYZI3EQmivDQ05Aom
pbILY1MwAHNVMhftgAXw4oigfr96bdMJtJ0Fte8T/zNXOnImEM82qI3dzB7Q+UrhnYMhIgKZKluo
Zxecm7dD+6WCY6u+HbKjKGmqMn6kYYu+UKxmjVUqRapygJAdIfo7c94QsrTBEebinx+ECqx4bfvs
Vu7mPtHSUtdTEDK0woI38vk9JrYpr1RhJR9SZl5FA/yiMX10weOlv7obI1njRBNC6qsd3bycqe0+
pZTuJG7mFXAOG88DWySs7oBd0KMFlW7zff2F7Dgx+KJYmdzOgX6j7u7dsbyrqcRxxEk47Jwc4yiE
aPhOPBRIoXlS62omySbR0i6Xm2h2SyexTGRqdJMU3zWF3+itgFZIUrkpskKcUq1bIx6JgGzlfgLy
rJp7ntF+ZIKw232AlsDgqYuJWNNAE/Ed/pejY8YKy8AwtIN5j+2mfOkypx4bgLwOMPGjRARjbdtT
APTNl7egEOQeJnoDyGlNMbMyfzB5ymRlftHHXFQl7BuVRe0TKoOgN5PxLqHUriZtSMR2762wx9/v
h0NwYIcxSQksLE4x7qbaP52Nku48SzfDn369vJqerD88r7P/1OxqrSqP3tKTSCOCmUd59KBmfGNu
xx/DUVgAsjfkWwFt9QtAXVXM5Ik9gXxy/VcBSE5+afKYVcw2bODsHpnXf2MPv579Phhx1ZiEmy82
S6Uj0Fp+2ZE1i8EUxa2eV2qcjzczcFF0trMeAxdhvAw0zvVFDBKpSuiFTAXtllm1ByzbVbQU55U6
UQwPJterSjOEO0d40wQVTlEFFHZt+dJLe7reMM05khLOW97ZfTZRUqw675q/4xXfCPrYgMawyBWb
RgFxRPZC9rUFLwkl+vfwM+04+mvAX06P9KoJ79+CqxPgv+hCqyhCa3Brsm9Kk1ZnLkM+ql1x2gmU
jXLMrdYMyUnYVNMGBcwD0wkOw8HzjOI6kA582mxrQlQu5uCGv/rxvyWU2yMtb0UNiaBHsEp7aX0F
FBw4EWT8cBrhH78GHkXDSS4sOyhCl4XHFiYANyVXDiZkzFS5b8fTGuSTIj1hA6nEvaibengAy+vX
63YYcXfAdic9iR30TSJV5OlevEi0Bh62jChGoWNl1NOQJI60COFOfa6gmZIuUIALJgrOIh94yk7d
YCgtjT2XRlybx3qFle5vo8OWqw6vUFl9xYqGZEAkm3lXaKkB7JQkYC2jGXhf9iZUdzS4ADJebWxd
L/7rhYoKiHqjn5xqpxTNTrNVmx3ufG1hYqnGUCfAML3GAf8gL9IKCy5564vUpkBMxznmzeCfXHyg
3LSscQaOBKc8VBMkkpyBUlmE19R8JoQhbjkk3TBbNmWhmhpS3wY9BEclqLMelDUgwJtbZoeDk7Xm
MTvHVtk27da5kC0fqr3Mrve3/np1d+xwGVi3YNSfRV2TvFbkIPAM3y22Fpft5F34pOqkZMxulR/0
Dsz8bZ8K0dUThjxXUgwa4iANL23c057FrLLrNDGzJGi2U8T6zrA8IBLK5muNaVBu3fEb+Kbe8A6P
jTFGsiqh8nuqUBC4AduG7DqquZOfhHGgkp6CcjGpM8eEbZnupaPdpbCxT1zTabK/JNbo7omuhaxv
8haOQM4ZASm3qvJzhHHbernhqjCbQEeMb1TrC6Yctlm+/pM6h3nr7WYjfW5zX7rJ6GlxldM38a+p
ci78pfsDb2A1yUkHZ1JobJWiBAacPoZXJmd3By5zqvKGAIc6CZmFu8BTgwq1rszwjn5NU+96AWRe
emDHjRh7b668JD3WRCFg9WhXkLDRRKgeOL1fDMd8z1QuvgjVSd+3lsQOOPJDzAWG7mCx1Wbh0xS1
SR3XfRVHEj61+G6DhUjCVLyelV6/TweTyc2xXfNtGessD7nLGnQxv4RhpCjccUKYqgF6JacPCcXY
EWYQt6gECNrbJBzP3YCIo8vj5ZZvUTXDXy3W1WLLcG5xRB8r2D8riB9BuJJLS30pe45Be3fxpVTc
VuO7DwwE2b3EuKkvPo3rpp9vobZnCeqF9CknyGd7DQhqOXXlE/bJq5ZO5ODr4//IuExAd8vw162G
U2aeYGlgzKpOBc1Ub6mPiaKLSGYuoXOTVtd6P0oRtm8Gym3WwpPqCAB7/I32sKQK3LnJg1Uw6bB1
jkeH2X5kC8CAT94qpFGK5ISOAlc6lxBJesfS0Eb+dFxPYX51F07+SAIAlxp9/GSBww0j52pz8mdb
clrmrOFsUs6RhpCcFa0mgazuIouNpyGueJURCCRbqy0IsIsPKaN4FomYC7ozGE6CAVUeY/Cv8+Fl
F6D7blM0YzDY0Loj8Mqf5sjMZKCN3yvJhk3OZtj2rmSXz49E5zUVlDURFWIEiR9C0WWwaU7jXlGX
FyLtjeCjhv53zv0lfSs2J+fgjsBXFy1OrEaCxoipvEhquQzMD0wXpf1eSTTdKFayCkUPJPydRMFa
mactGBv75dGspVbueZABRm+M3tiMyDy7ffxAzM61b06YflcooUIecJflzZHTNefwgpHx/s938Ndm
7+o2rNfmHUNQ59tW7cuTMAUykna6tdJVpieAVjvE4+7xXa0s1e652VJiwwa86BnGy359Fcz5hG4i
GZh1knwH1NrOJBoo5qvXoIgg0wB/TZgABj247+w9NkqFAi5DZEAwlKZhtKozkCmLAZOR1niVmnWn
7GV6GhY9nB576l8bO03wWUgiP5rdV4Q5z6+6QvRVG/qMH427ZsMDKeuIydW4rZtH2qUzKOoWMuQQ
bRQWgmiP9166Zqh3K6M0HqsQyaQvcVYjCN9vwX+LtVOGiGsf+XHiMgbvKg+CSRt0PdmEMnrCb9oG
7NgiaQHNqMXQB/R1VytOjl72Wxo35ig/ejNSCHiSAnr+3mqQ883c6BNtAKRG6UauzvIQaAQ0unvs
AzeQX/arHOF289JFHUgrAl1MY1Qwh6/OHUkzeK+J0WhTv9E4wnv176NbiE/VZXPvTy4Bk6Zvo6VU
2UYzaLuHtEwEMN/pJ0lo92K7iqNbKIbVoxdiG40OSWoQX549LoCmCpKDQ87SapRDIzhLDFyy7axx
PN/9TBHkMXl+l+3iyKVLOBQJJBaABjSz0ViPvD/FtKaaIkTYTVDCWIGyZlpW6WCDm8ao4mLINp9W
6dLY35vAQX+Bn9l3nTdnIJQxWq/nkMBAm9Y1RD+u/vMuNFDA4xNWdOiO9X+f2suF9U6pvsqxMLow
BAfS/3VbDhW1CKKnmCoIvptU6kQDrJg+FuV0tsMVbRgXh/EymiT/Kac4BelX+3qANkkoc2SpjO4Z
VxG2uSy7R8tbq0KMiNxN3UxW05Qx61isiSqxwihLh6sFTVAy4die90u4FJ5urMvSvpC8yf/ewtUR
eX5mxbLmB5oCyjdKLEv9rMhie55OlUZvIowejxtZlsE4OaiIwOU8rL9e0oKe07LBS9YKgagg8IAl
r5GQ0LzX1V/GIuhuY+oC2cJJcpTCYt1dS2OaD2KLj99bVB0DEVHHAhMNj+QmNtGW5zl/DtPARTWM
g32MyYSX10YmGIbIS49/0BxU8YDMyndtrucUXfjsdpuO1oquNP2rX82FZgRXh6JJ3/oZdSZVeThP
EKVNiC19ZpN/DHfNgO3u8ZU0bEuf1X/sMrSYHdDiMllbB1YVlz9EhO6EhlwSonoW/mshJ74J64qH
LgO8IB0n2iKLrDSydgP6/8GH+PeAyip5TdFU9VJObZf9h1ua08WAYjmfqZd8tDPabG9qqhrZcaoL
AOnpTjuEJ00O0OfUWFdm9ok23WhlnBkMJYrPD3pgYVyYnmCpsBt0ztNAXUPtL1Taqxf2izzpDHh9
BftNp2Etb0ByisZZb3qreILy+s16V7jPytVuXiQ46DIweyHN2mjBt8q1ZWM1/dYI15KrJokTSHhe
RHMY0QITmTWTjBXaxPVTg2AfMCRmuUO+d8pkuhXIhPKM1LXSV5/9Nql0kmqOrIhylnRF6v+XSx0l
sl2HjlKjjmhro9eLG9kYI30AtmtEUHYmC4gTpPtZl8k5D4ZatidddjrTkT/P6KaSJf+umUStqnGA
KU8tgCMrC8c2RDVvvPnlE90oMvvJ+3VhSYDrh8Njl35dSpR9Ig081n+Y4GzdunMfkQaBQhCmO/4I
Erpn9kpugimQHeWHSTYMRZgzrKfXT0Qv1ypLCHHQosD/cXbb5+yi4S4b992Zag579+FJnyqTBSsp
SSGVZQDOH9hpYfwj8Fu5WQcqEVGgeJENj+C6apHU+iNmRT325ARMw96O3ASWN20GQHYwZq9jGAuZ
OrZFwAJOT49vJa2nE5iNPSmyYI+b/7Rau15lYV7lhRxeNmoFqfG9XKHnzABdUB9uGrAv6FhXMnZG
jsKy5wjoLKD+uEfBKngz4vAN1IVmjIcpkRwc+hkuTpIFPTC7CnH5DC278nxbLFhiacpuy/Kv9cop
kM0tB8r8Ea4mpXnfBbD37ax8fmt/79YT4w+c6nZN8eqYq1pajKK2jr16rkCMLL0M4TK0XS0tprWL
mldi+uvlUUOYy8tl3xMU1n+1ceu9o1MxKn+yhx35SaF+6Aq+jDCo4Ry8TfhTgpPQUF2VJRtjmuvk
RdDtrE0+Nj8sdtICwKfukK5PZ4rZozTxeQmfsk/et9tl5EmOTJbeHjy2AVIQ6FEbxaH8PBnBN4ag
t1ovv23j0wvYWgLHuqNWxghb2edfbMEZAMhpV964SM/+qOhDX3M8WnrEv/G/9x8cT3uF6p++SCqX
bSp2ZzorHz/YRT1iu8CkLk77PeXlFIHDmxq69y8+8DH1eDKDjfuDvzLThB/HWxgjgjdM8+ocq8Pd
GcY6a4eodoqmEUKGTy9XnNrDT28LSl2BbYfmEByQOQbqXjbBuuN/nfBvguu2WTSDIsB2cqwLu7Ka
5m3rGZ1G04/kkLk11DLlvNCRrLF4wnG1pdL11PDYaGhUYloAOuDWieIXAZVNXGFlqI+T0N3Jrqxw
oGNfhvMn902Wx0/yusgsk+hd1W7/PEXTuCyRIW1X1ZnFx9GKEZOfwp0L3VdHJ3pPVMSnWSkS68CY
Rul+HhzsacV2qP32N2zfmfuvC/nj+Gldd8jR+h4i4j6QPo7etoIIOx8x1ov8/kDncNX0Xmp2EHb8
Ooth8Jg0Ifj7i77s0rI4PH/ykrMW1dOuZpdrC5Bshocc5dEbehoyFXofmlP+6Z0vjLnQTjel8mwN
86NOienXIQ0GhpvgfJiJW3ElUJhP0txXtvYHex7XeAB6i1ov1njPeaheU202mNKyScgdIKwB5QdR
30qA3wLzMRg6CHf8CbjoysUGLg1edSvuBhLZxJkrAbi62a4ucwa5gNVUxV4D5TBZ1uGRWKOj6Wm2
7cZKRJl5qcagFHD6OGFl8jlvS07343X36J4+I0Fxpnys7tg+9asSeUQ1g0Rg+TaQ6j8oIQhXXeLX
6YUD+a0ZG/4WEw/+WaTA58hpO/IgzRUqiPJp2I25EKueprxqqi8VxGExjv9D//AZNxhPb2YFG2V8
qG5jOHgh3oW/Q4ziQnrEKx8drDGdX/PB90yIeOdqSg0CS9kNJVFqCQbobDG4or0586JhQ8mfqyjf
dlYHVM9HBVhAsUpfVhF+JOlQ2FYJwp57r6S0P+6QC6gLtfBiQCTv36shpIPspKaYxriH9dPYm8uH
+nRk0tyTgKeuFMOFIrUB+fqLK3TYolDVInalmq6+hYzNYzjP5zUo85GSvrhFrDVxfYv7XjrOidTJ
ML2U7uDM5NFst8yhgY5/+SEj1J9Yj47YCLVAKWHn7RzF22kgzl4CuLE25BkRlLgQ0ziCbT9Ahp3n
0nVmRtoc5eJ0QpXozPdAqBTpnjFs3YBmfengc3t51GGHrMv+KncLmRc5B9HE0B4DwWPObxbrJsxn
dkRViqXmF6rEYFRaKwF+chiPbeNkHeLqnYZEy1hSvC/PREgg6TAoKY4hHhpi1L+hEOaryPtNAcU0
HDo91rJKzQzb+PapyPyTnN3r6/h1W+VZTSOsZbwSUwYN7EZ9M4r26/lwQZuwD0yKTbDKG0JiG9P/
knlqcUz0ue9CWQEb5y0XCkuP7oX0phuW0tjUBU7dQNEiSQNU71qvSuZ6jdCpEZBTPksD4mw/EBH/
ZQbRuxltqBi/vD+z8RK9aaPipa7t3Wntlz5uXJ422Fh05SckG1U1z0wrJK3SQpFODUNvhQeZSuin
qzB75gDhxVIcn/04/safVmc91VWKTZrmsRv2lwK3pcS8mxaNEyouSl2lhE9t2cdkIqsOWExqhgbR
IjEruPCaw3jYNMn3p46PZt970o67M+QyHgsS4Gmqj5KF51jFe9K346TQuuxZCMs7e0ui+2vhA2hV
s/w6+U8Lri9GMRFLtdd2xM+PRrtjrYs+yJCoYQgcaa4vL9MFk/43pQVehSEx1Bvh6a5reYxvyh8X
l0qWfckjpO3mkj8xbvnuMIffsYDK3fbSq/BJhBwBKldqzhcxrMW8UFDIZX89DgXwYynKvfDwsN7Q
sGZBUTtnN/6pqNdP5zsCoBQe7XyWQDFssmDu/nApaADEGzKa0CreQ58+FuMjdC4h0ScSDPbZkhvc
3BHzYOOgUkfkogzZWzPKmhmcHro+cwV2yE13SFLEvT8dpDfwqvg8hK0yhn3ncYGB5JQbqQHL+t2p
OeG8d251No7d0LdxPRho2Ok3IyAlkE0CGNj/PyhwNYSBHkXCcgLn1tlubv973qElJohZav0yLt2K
xkn4kdRWRFBOc+9qtHz84e+P4Uka3y8TSyAiPVR/kmHaBtf05TKRdu20l6739hZM2SCDAndgzkVI
WDF2/Ifb0YmWBNDvUfPPR/06sBcb0cmD33UbLHfBjVsySaLZiLKwJVVvExL+ud+ysxLpCtmaq0GJ
htLio23ZFMNphPRwaNAyxRwX3H2DeaTRiUFGWJZcrnfbCJLx7bUHcM4PW4tid05og9hLLUNb0J0U
6jptQ3P2iTvfw9ORIGKWzirxYCDIA/LQf2RKoO/eEkLpbMQ/fgWpmnc2LINXqP9BfiSTfeW59//E
0E7F+bFbF1j15XbGim7xrH2+OGfUN/izBPQeebs+hyWH2DdSPBWZaqC59d/d0BkJO9KKEo7CxMWW
LxfwtVRzceMp/ZZNZlqA1emiuU7j2cAJj/SEMJX12wTN8Rsup0Bmvo/E4fSDs8J7UWksJftXZV2i
3HFXH0IA1IsbtO+a8ELq4L2vHh5u6cltocmeum3Ybil+Cofo36DpDTH9pJXzHV4Iqqd22mX5DeLI
fiI+Gyu+qdS4BUJCVSN3gBIO677O8pG0RX6eVgCoWRdqG8gDmscDuuHJmWXWOGY16aiTrdbwLS11
yWyMkYxELdaoM3yh2IaE+8/3ydXYtxxbyy1o//aiCUORIWXkbEbj2Aup9CLypQBVGX48GYyS27yc
odQ5DZuvyI6Ze5q0ul884gKQ/xSbQoc3/bcPxGHHvCOFV23EdwpknL4OspkkyoyT7I0tZpyqNJju
C5ST2QQGxYUOa3rAH03fu7hsr8EKHrAnPrsQFpVewUk/Yc1mxeTEVkXOMTYeko7upRCsZfxNQHoh
MpBOLo9uOg6p8KyJ1lEBre5utoc/CEVGaxrZjx0LbrckXL9//GCobl3lIoZv3lrY7zWRRntlSkTY
gZDpO3M6yyAPCOajG9rXF8Qv465TmMe7OX8hQcFnUaSsyLPFN+LMsEYy36dInMbX6D2+0S0wUsWr
TM3ZKEqUZyYlSiucPFo2YX0Ctj9zmIrGFLvyj2TgQ4GDdoBVj6hG+oPZhxpgHG333QeR1aXbpE3X
A2yGtPcFGIVcwZGZhN5imP5WUTeaNDhJ5McpZ5N2hZZdgxXpnQnKfbOh5sON5ANuwiN8eVtUfLOL
cdkDntVVNeDTECdtH0C36Tv68Wv2QBz9PjSTzjConj5rPmX5UEwQMRtM037urSM7aOwLaF9vxK37
QG81Nr8KfRleZTDg74j02+QSJSkGhN0pKgbK0TtkEakpWVKqu/zi6GCmn904S8fvpzZO6BDDrP3Y
mUlhOrtt8xBg+XPj+uGjZnxmr8B0MJh5xAiILM23nUDFfZL4Ob0mzpgwrVftvZIAwNt1Q4jO6Kx2
ZJqhLcM3l8H4Iz6REKbvwxNG5TA3DFb85PLyW/IaFQGbfTzBJszKinEWu+bsdbjcuW4aEFJx+zmi
Ff9v18ZKoeD1FzS9nkWB8bPKOGUDqqgJAqSPLiVIlDbBeBWNM1Im+EvN6/OuDCMz3ZjgpWfkuFxU
Etc1WhKdw9A7RIm9z9ntkL0QPf5dokaLWtRR1ELXXEV5SShYWySi3g5OKsWFOHlBnPBhhq/pk1TE
qOB35KXJ66vTH3uaLOed3dweg87RJp5kpc31v/fp0FUPDcy3SSBlCxIr0ZB4o+wGh+iDvU2cmFSu
QvOmVEIHCMUSBtfeCxVwIQybt+qPheE3AW+/KTUimBRq/D33DbDEZhzrdo4wlLe4f4XfN9kYrbJn
+TY0Tc2hxR3V+9Y1uxpGrxMgRamb9b09jUtIL88uUEZZA17ZGI2kfMTv9up04OALr9ae9SuXClzs
A7PnECBfVtIwpciwoW16R523C+0RSHRFIZAsGU3VPhm7hR0bw6MPTaBMaVkomYqXVgqK2FLt3DVK
YE50OnhHymbAWUXydDHXDd57eDPP4tOOm25fTBZ6ZHPL4MdjyoIglIWzvyDf4IN08Y4B76R5kXjE
DZtVplHtMbd/Eu+IThE22sR5p/uCPC4gDLuMuDZNwyjZSBfITU0BEioMfmfnExpZXlChiujtT8l0
fXSb18a4PzdfPMZntND5bakkBi8Pl20bWk4hCTzt3AxnGDqA3EkvJYgJ/NUlY7S3LWC739MZCmJj
5ID6bP5ygZYdthk4jWZorgfZpuS5G8ExNdITEAHt6D5YxEBBb54H4zjNj+fkY1cevDVMiP+ApjUz
WSlx1PDHJJ5r7zylzF8z3pmHYXlKeQin1uamfmiElZCXx4pbAf96H5XlFjawZsNi6CSG6hZRycUG
R7W1J5fUmEoQ+pFdeNMYoHdA/AqgSUWgNj3lAv9yBIKmicgY+VjX5ENE+ZjiQceUlZcpW1cq7X6T
Q5y35zKb77AZA5surNhImMDGCLIno5PZIdK9InGSygdxDTAEZEKBZ1zv38hLZ0ElaY9kewdSsNow
7Q4WqTHZuRTIF93D1pkBfyyTUlERJ9b+HT/rd7u+xdtnpku/YfkAJacikF/X0quQwsQU/IvMGtlm
JmBri+IH6eE0jzFOmYbvpAS5Godd2TMfLCww9+243DhjO86CVwFukJGWpMUfR9veKMwVtOGZxA2Q
Ru1ejXe4TRZ1O48yNTrEXiBe2jbpzS4VmCfIvmodFx948TlNpbL2OGi1S512nawzSZwSWjlQaHM2
CK8IMF4/+kdv9UGu9RRet7bFg+ef8Wa9Q4UafLlxWEAJA9/GtjLWtBw03DykJvl9bRmapP3LzZCR
72oK1i88M9Cbhc9BwTYmoNnQdnxj9+RW4fLPOOVZwGGt53oXy+8Th2vLqU1bi749bX5YncZj0T8b
MT71HXTwdGvbQyUioHFe0+p5N545e1OeGJ2lACkvE+N7zk+svDsfun5GtjwUUZlRbLGKr90eTrM1
l9velIsj06i50EBhW8hZSZYPYdIFS2V2SXNhUJ1NdzRJZnMw8C4B0eiPcmS7DmCFNVy9uVcSDFaY
NFoOAZ/PATwNcN4zhP6eo7837q3G/UWigcezaLCqQP6qqmVFWQhSCcMVqwPEVQz3GWDehKuLc6lL
D1JrRMmQ9kqJ53u+Q/Oe8tzHee25TDR9Q4x5xicTtNCnQrzwcVvOC5Nwcbjph07gdYn2DGDVxLKU
X0V0Ne8VB28abFwuF196Nplh6TK9zUrBygyJjzIjPQbZP7YMnK+DzoM8Rve1ebEOj3HotlP0bnqg
yVusqHZRqqRp0h2BxNcb9LgCnvWJunHu5AxW/9JU7MssS2SNxAOX1bNUkPv/MEBkw6fJu0ubVusm
IyCopFTz6VX8O/xuc3oSMfLAKoRCRItk6OyGOuHZHiRPZrTAOGuddk1Dl+hPacOkfqrMLROI2fW2
v25pjAGV+c+BfWavlAJtt//YxuJD8jSPdDWDU4R0pVejVnedH6k7XqJEACl3Okbvj3TPTcOgMWnJ
WelFgNl23dNsfXKxoE23XCHDPbd2vc6q0k0GPpSVus549GwaCGYHQNZWNCCV8D2WpK6rdrtrqL2Q
GuQJNemXLkbPFpFLXJIxVfl7lhlCsq1AFQKdtYEXRRCuxv66xSJvX3xXzDIvOwxbvMax38EI53pO
NHfGIGgADDyr8XgFDclep+Bv7grgv4+mqRa+8/Hp0mgj/9OFcnlVjIE9bjccci54H5sj04z4ZSa4
V92Oxfsbk+0Vx0dfFb11obW/QJbDd5aqfjP80wSfl2rd/UJWDrpecKLBbKotfsvjGNkLQW7sUwdS
gGJYxzQZxjNZhCVFtbl2hhYtnHNIfOU5ZdLRJWNNex5PnO7+8cBz1h+heW5oMYsOsZNGe67zZ0eT
MvJOoX5Cv/72NLiIxvjjYCtymFfCd3oPFglJLxAXFdwq6qLWxuBRKiljHcib21RVrh1827uJY5iT
TPcjlSOyRcAhUTMr7+Z3vHjpUqV7egtH75fbgWcYTB9/qdMiuqHOig0XGKWKPbcUHhKHhZh3y7xa
I9S47yUcJGApwpMrDAxoidI52h28wMSAkUoLvPyJSt9ZxCrY7SdGIyqia3kjxbHDmMdkvsNo7h45
buH5FgA+mfJQqG8eiK4ko1KNrDaG/4sRJB6RbAJHzE524KM7amdT/tPv/xsCemEY8pZlAsaJYH/V
4OFoE4VFPUKmTi5wjwfpSxNYBZCYfthoRITKs4U41fwgd6MI/5QhZmfXO5cvkWPY+SOifmmJzokR
Aw9jivrVL1wKYn84B/S631TINYUV/4hDQUuL6fKiiJC2KrTSDhtWHp5kMK3TVHiab0PTkB7KrRD/
IjwZcf1Ix3GDkMY7hwmpEb+hNyIMBjzwgcgEoq9lzSyDXbkpueDpA9UjC6au598e52jHkt7n/lcJ
Rf/gKpyw203vkm9bZoadT/WbbNR+F4d3KFZllrQx6Gem3ZhiLyl0vFpZSosANeDcYAz8dcP5Gx3X
mAJksNnRnpDPhiNnSawWN4Fcif2tBVNxSHCyZ2wOfTHasi0cpXlFfd1mNRP+hpc5x4bB9cVEin4/
FFV68B/TnX016YFiYl5npZ8U8ZxQ6InXaW5dKQF/gh6SRCGwMW9eRCxis9a4YHAGUkLNzn+rs3fJ
qXyp7c+1ALGkPjMYX9p4kGpML7vzpamEVws4q6IYj6Q4ZnwVYbeDK21TNcgJlio4LGWU/mZ/SjoV
/ycvthQVrNoEK79eMHKLA6GxeR3mbPkk//jYJEeYW3OfuoPug+IWffflkOKQ2y+1blcxsB6+pWng
xCah3Zm/wiGw/KjI3J4jpu3KIR+UQcyHwFEa68GMvDIbrW0QRHySoPjmOv253V25jpAetxK9VgeT
im6YbRSRc34w88AqtpQuUsylbfLELmfrSYWXUOJyCm5Heh4Sj0s5hIfyoeZKHDof4N81PyuxGf0h
SR4n1pMJRwcKyeM73vZ9a9as30IAg8x4fu4wNX0lNJNNJr8xoqjFMTpeLvQUKUoc6Htp9xpZVTdm
J2QLpAEaLT7JdbylPzlBMa0Q+hqNgutbOkGnW+AEkw1iiGimtTVPXyetIPA9j6gdlllQBEJ5qPCj
fqdiiR6m5FFycCkSadg/HmMEWhBWWq0CEhx/0IRaHPkRH9OHZF2J5uoGf7RDykMne5KyroyxEtQ4
66TB87A5zdE7pDSJzM1N4zDswEpRCKg02gP3j2ZEPoE+nMZL3idawACSelTrHsP6VBxvJpnk5yFb
VXPlXh757hsQ6vBaAOLsf5knL/sAhpNEs/Q83BpYADC+88J8d+tYDS332y+fUVV4d1YctSSHMaH3
fTmSHBid5SzG6GUcnnhRF9TSe+q4YNlXF2KUhGSb0ONIppiwZwII8npKVVyEJpsbq6/FAmt3MkYD
F8wyDjBgBIp11Smio0CtnE+ftVAyN9ZxqVNJDaqwcXYWg4sOLQQa9uKY0RMfi5I4/axPOtr6BEY0
4ejzpu/pYyivluegljF22ilVQPBQ8tah16P9LVr1KPA44pKuYBcRFAf+Tuf4Lr5Qz5Pbgscene/2
sEHSUj3jrwG4zC/kBUrbz3S8KqRb2IRepqnYjQqIAt49c+fruY4N+lRB/coZPSfnbhq3onrf3489
EEGS6X0zFDFM2PnzKcDky9y02K1yaa+9E3lqlT64HW3i3eXPcQ6YoZEGhBDkLR5dZeH20kjuIRIH
Sgk4BssIJyJXBrLfujiPIgcr2GKKSKR5qx6P/+gxYSRwQmx0G4p9X2EJCw0PpolspM4gjC2EXb8d
/7ftvuQjONGw6x0jHwRatJEzpqrrVjAzscNCCypj0MTReI08s4okZ7HO51f3lrRe/39oLtBedUQ8
6p8BNz9Ij9edDUVb20OcF0xPorL5sr0v46lRcdoedve3vq7qyqygGsliRxw9dGJITqadFmVO8n9G
JjlNqTxJZ5bXcRDmTur2ChFjY6guyMA1GZIZi8E9z3EdQlDmfzK9X4CFcA2EGKU2I0PQF59iT7VR
5h+wDFycOvs5T9RXZXP7P2lJsBAb5fROiYjmDLcSoUACUpzZzQZTyTHdbr2oNF31l0DRztVnwRUX
Vui4oVOIU68Fhaa4lZGBmgTCy5fem7SsSfowVCjSW6RXc/sTV/iWoDgV8cmxl84nfDuVItTW8c/W
lqYfdbIYS+Yn6J0VnkJxYIBQ//+uHd26ya8AuoWBFSI8O9bDm/yufIEdq/fLK7wLtilb0mu6w5nV
ZxgTZz7dSOFnhD1zOJP/byPeCwnu0RQBp+Jsq4p4hCzKngp+AvUp8trs0Yht6yFce4sFGlVRx36L
jMohRGTG+8r5uYMZZNPNlNt8ec+ymB2USjB5h2x+9S3e30sCV37YbJvZ3vpuMjSxZ0wDqUXmz3R6
bfQgO+ei8wM8tgHShVws9mFIyTChZVUabLsWkIJI/tXyN6ZL9xeAOsjBr2TQtKaC1k8Ui7xTbKUN
4jFTo+nwQZyYQN/7HGVAQH49vCb5lXuaLZ7KRpLaP8L+B+EnV+c5tXBGYKZMpcrK5n7llWU17lFM
CUyksT66Xw/tSwD31NVCCDMbz0KfiRFurIdD7agmEaBJAa1pBn8VBUT9T3VQfLuZ2nSRhpsXDhoF
Y9+5WF3KnGUmXsp6UqDw7iAQbCivWSUc+bGwbfldB7YcyGwQJa3yLy5ukXQ5vOZq6+IqbLnLsc20
6IUNPumOfsZHLPbCkYyjk55kkQkj4iFvkYMSxJSFLib56jd898kpCsubLx2723+8aqfybiTmxAPf
YHri6g/CNnqobqy/aD/1UMBJw9OnB4PucSeqi9OLsW6h7Z/RMkfkuYZVw1oU9rIZ+ra3uCkFt6S1
WU++1+3HjAJbyD+5SmvIi3w3QeI6mPFLbuK3bHNhWcUfA35YlHCeeQUiGEtLfkzE1nOQgl3xXjHr
/G+yr3pWdClzl/A6W1PW9k558mBBmwf7eooNDhMHmB/5XHuFBw++DFGMmHH5ScUnlZYp1Sx/3whu
kofbAu6cH7fN8fSeS5Ne2ROMNnZypmO+DPkAYJ3O/3mO7miD5Z1IV5XBXTRwrTQ+yNNRArgN1Nzy
QWvwOefFBMMb710+ZNnbfUXQFMqOXYqdNnaCU+u0ShMYBgutoCX3xf/7kgPzD/tOyVZhC7N5aQ4M
rLYp4aJjM661suQRv5qZlIeziGccKyaJMz7Qp3a+Cpm4UtK2Wn7obgk1sNDUZS3mxcUZFIJNovIC
OnGs3i1C+d8lDrAMoifa3oyfqsSkaRRwO1lnXMZM7OuitH+IuvQRygxvck1g8WERAJ3fhdJb2wUT
5AEx/n07msAYGXJ/q4oQ29ccSSMGc4l71v/El4ufjwuH7sgX4hz6ZRlpZW68vmPGJz7K/fn2z9pv
DreAIeEGW6iTtBacaFJ6Nqdq4gSX70bF9o25nNMMcO6DxHAl6tLyIJ83yHcS21l1ALJxi1SIiiYO
nmILxIydv4H7wbSJXDD/j01Frh3+PH8c6hXAUtaRHyaCCq/7NIZWDE1nwPX7gmWHO5LkCW1Sr7j4
PMzzIMDtcG8qcTCO7nywGOJTKgMDhYgTJdao1mRe0vtORZKNMEAProJLNMapQjHcrLXyU25AIEDP
7G0biWOG4XDsMqnstikezTWvEAMDQFAmsfPOpqofaWys3ozqSLS4rVp2UD+s/AVmBW3ElVdsH7gS
PcHsYGhyCacufhNegAv6wCq5ZZsWYbMNMz/QUbtThDR6Xz/ol2S4aKojMtyYj8JSe+wxRnpx14XA
R5cnZHlaxpsxW0OuobPT9l46UJc6LLaEM1mNtA3FLgO8iWlKWfPbXmb1PDATqYl+eKQQ1sWzdsbo
TeOlyW07B1MkjJ3xc+ZgtuG3eIG4XjPWfI2zf3vjnrAQswcNyspHGOc3Yt42lNjR6S4CpqFshMlr
NovbCI/lq12zmmzPbaxE0KJbF/kZ5PNglDTU0AG2ooX+FbChQUhoSRjv1BFmxYfggAChkLX8LYuq
JXUx5kVDPi/kGdX/yyd8WH8F/zyTZlJgw8hKGBKyLpsZ6+yVu5pQnu8JJwbOquJME5A7Qv6B328+
D3ciCCkN1K6jBgV4Jso6XC12i9/yO65TtG4MgH6yUD1s+Ujv+KwoK0p/9u8iZH1nDFpiLYlqPeYX
L83xhgrJCtd1+1St5PIXhkc/CGlX5zp064lGtIJyZqMhi3Wo2HyNsD7ef6IERv0xeLApRnm1UF73
gPT4VooRmk5Gr2pNmMzsyvp06Q4HLYMPrdTsK8F9mPeOh3m3pR9vrPhgFFsm2Huc1iVArgd7u/sk
g8e7Ht6PRmqf48U4WysVvI+Xbpi+ZtTy/KoFjhc324nHH3E298E+W9pK2YX51D8p9TcP+CzxbGmF
5ihk3bZS8AZhT+D0Gj1IFqGFMhQCyVlZenp0XzzqQCZZlaBgMccgv8MlTFDx15iz+A2zbfoupSiw
YAhsjZj1P916ilXPVSZasNz4T+9iSgwwAqxTy2sP762yJscyBpJ/68FXvnZ6m6P5YQq5eDT42NYT
JGxRKyBWrAaZQnABYt9odJRr91pkT5rYlSbfG3KZ/j9eg9yq6Jhv81JJu/o8SUkpH7pOcxha84rj
mN+ZTYvI679JgxCLH/DYviWJE6/PZt8GRpwKYD2QlWWHMy1f3FPkIxIii51uEG2p3/Do/2k1Lu8/
bUVkfsGTxweZodGwA1qEJvYvsBSxlrtXcykMfVCw6OczkyJcCzmDF5kmGnpnkNdXnnZypZ0hFwX7
kCWPbRG+LJGabTcQNBYULKburJg/WFmjNezxTUM2Jkcx3uS+01lWroxecc6SVbPUyoc7/LJcIBe/
iZKPvntWRrVd6gMMGhtjFdtUTvZH0NvwmjYZqVayXLffjWoRkguSO/wQ/V+/ey/f+Cs1j8eqfoBU
s+aMnbxLD/+ScbWHpWOvaK3Ft+Eb7hImOfPWFSU7i8zu50kG2ffSZaLyG2i97ezkwAzcf3n+Es9/
Y6zGxdADLnxWfC4BZRQzsWNYmD2CPpVtrLAjRR6ebGi58stb7eV5cHHu5f/yv5+7e8R9FQmc4fkh
n0Bo2KP/bDf+lTzlLBHVRY12UAi61sgDTlfDWve6e1XjPwYMFdeFdCT6J1VBBu8b2sbJ87Lpk0LA
vF6MMaIbdJYX66BPj+SuxeC9s4AhzQBjfz7aqcFaS1dc1DABcvsc0ehnON3BGNAbdhdIlEIxzz5h
nlTNtYS8eApMingoHeGJUaAYxM4rAfLHls3HCEp4IXhveIWKbXfr4x8adDssMYjauCZNbUW/A4ev
1w4BXRCcbIhSqnqlwdr2rYRseltovs6BnPXkG7tElzb2qBlnQqUl94Xck7iqSUoBCewhPISVnOPd
s/iWpEIv+/rQhebKsysrrYsDqnW4eAP/xJHSIsNQlF3IPRLq33ZfU7Vcc8EpbLHshY6rXTKFkwMg
EJEZ6SVE0GvPz9hokvY4ROFDlVbF1hzeG2EmAF3Y1PEi/3BVhhA+iaT+ReLqYkWCQoYhSvdp/UE1
7+wYLC6qVMBI4mzljdP3r7MLrRt0uYHoR12+AOv5nb0z5kUacW6t2NBtTImtE95zIkOtcH1S4lnE
9eMAzQMXKAXR0PdjtGH1huLiXxw1CX5aln5IO0h5U3BLR9qugkO8lSvAIlPhv/DbhL6XE+RJJhfw
lptc4qOId8QwzyGwWassEwMie7a1fQ7fky/Niqsj+APrk6CsVRRL410Erl5USTC/8HdO3kgtEmIU
6v6uTnXz4EEqOEUwah4ezuM343e8sAizrY4Aq+B1VLNXaQhTiq3fhEs9A1wZ+fNCUISISuczFyYG
M87qV6WWjTe1ALCASF+tq9cvW0C5L9+/XWdSOjn//9cVm1KSIM6HzycUS1OskXK55MtnrpOAV4VE
sxUltIgbvThq06I0LqbBBibdTxGJxdC8/Dqn2tVbsFfOkxW6iDhxkAgPH2Jb/CQ2ezpkQmfWxzI+
1JgrhAwCIFzKfIl3TVkavuCEaWvuiBEbRsKey0tdyut+HT+4sW+kQ9ZFDwNOXV4sERTR9Fbf9dXR
zmogjrEM+Drf8KYmSQOqY2sGk0C13CZ3EOrUMZImOOOtW0OQWXxUetbEJ87h/31x9yaVdAjEIkpu
WiaNwQOSeYIhcgFCqtxiKDM05RNZ4i1U2O9rVUgG4F8w84rjN3md/rGg/4H8SrsWSnOUGfnjSb+C
FUZf7IMz+briVxzJUg+T2oTKIe6438vf92ISOA9q0w6HZyv0tusdXaZuXcLbdiAOkYVt4smYc6+s
OY+S8leinzMz73yfr6XTHurr27w9tdSJKUm2xjDxo6tQXSuIf+WqiSBjlQwerxZwdMaFqeTmXll/
q2cjl1NwMH4Sz8wAKfrCun4vOOxF2AxMDBeDUqfxk5ENch9PYRabduXITtJ67y2XwLKDTokqu/Zi
d1OTp2uXLdLQxHdjZ8YuyEq9w4qmWz+XoccU8xkY6NL6U3DcQUgfOOce3CaakSBtVEe3fIVwUlx3
58SdnDXKCrFk5zYtXCOAxH6k5KOuDrkx+b2zPgx2yLqD+ixSsUEqAHP79b6SGiMgQ/ZZBzJMh7ML
/hHCsljYBk4pmLbkiGK9qnHeAUpV97lATHuMRXY0NREwHz3CY3Mc3X4dSSauB1/XlZo6uOX0kJ6G
rE6fZjfv+XUTxyPRPuzwU9yLhgxYtepGMpzOTiXx/H+PybHBXVN0QS6PBaG9AGk03MtPz43gwvPg
JgVzAbfn3E95sDV8F2Vo29g8FhXyEbotiRv1isMxmfS8P+DhH3QhvraPDREijIKzLMuHTGzx8fJ+
PmbkDGu8cS8FEzRc/0sAXw1SGjO5xObeQTgZxqeZkGXdd5kjYJc7w0j9YUT6/+IqXvuxwGu/EI94
UcQ2ECcOPENWYohUa/Fi48dfkhlnodNLM/xWPJj8POHlUyx9ggSbTlHn5MoPW1rCHsYqObuEy9qU
5Oj3OTH0zTGP3wn/23WMX45GpjcoTSl9s7d+WBy2JWyUJqxDXnM2TdBmzA91QTAbq0Jkr9LqEmcx
oov2G9CHZeLrT0UR8FDs0cgVkCSaFu1PkVOQ6nDXc+qCjqKkSdrmIn9GqjtCbXtyegQCKKXW1TCn
D5UH3RgbgSBJ6qKhrqFPuK7Vx27nsz13+p3dKgGpqgpF9cI3hLQHbqRFU1QGGZ+B0icvdjYcUTAC
cs4zhtirZpRmM7qRyxMJ4mGOmakm/ohjzjTxyJH4aje0T95JtN2FZ/NCfvJKH4ajKAZafYG+XCZc
BkRhtSW9BTJJxIhd/2j75C/XAFFYhaqvlAapx1TuqysVz/aqrVvuqTTMlRcWnDl3B9jnISSgJ4XL
yZrb3lX5w+vMC8jACEIcre0TSvMvMWSwFvNYbszGirQDc2YlrwPa7L+B8CU5A4B6+f+cItrsmlRg
EpR0F9kJ26BTftHG4eVYsV20rbGcKZg8ZvULVkNchLFKMEJ57UMkSgesCqIIatolkDzxl7lzG3gW
FLgl51Ptz+q13kd5uxg0DHguo0xNMDte60uKH3mHUUEJFUDQqnbuytp87Zgq0hVNbwDeEMkJ2kCd
P8fPAFvshkrPqiXoEnduUYeJOICJTM1m0r0sBkrAzAJboghFj1NoL+WhuzBJqizzx/yZwVLkXLox
X55uvRHfy5y1fX+DRgIKBJPJ34t6eIMiRdqFqcDfv3lNgEakBAwaOYhNlQ08McZdILLlPrZGxnzn
re3BByg8NgbLsgZXltkkLlG0KYtm5FMf50smWcPThNJvn8eRUzsRzqh2BFHmjnJEzBoePF4BCQir
QfZ8llc6oOIpPYOshH14rtxoxLwrfm6pCdlYyHc2nfT9DqMV3I0cefbDJgR/xAO5kLS/I5Y4IJwV
NlMBU7oyHsV/dmtFllItlofKgYFhgfm/qAEXrfoUjXFalA9XcksNZfjA+9/f8fIMY1UvfzjmDm2I
Wu1nSh6dMMK/FP6Kh7XqNWmIMjPkvxBewdtklyqJCfbusIgSIsd4www8kk1ikwjp6hQ0SRk6Ywof
tWUPpWFEnMXGL9XqDljrRnFVk8ShMMjiYsynvVoJmZKVMD9/Rvqn0qLEX+8XAlwJpY+jSm/Jwweu
H3+67WazE+ZqFNaxcYxpaS6CommVABObVhK3RxgBTiEozwRIsZ+0G7xy1bGUjOBNYIlmJOkRU06E
IkVcX+xSDE/R7YsEBf9cQ+RCNuIk1JJ8Bi2Hq8wQdj5/2+XQ4isTEOQ6wf4K0PVGzaXMXN1U3G31
e3KWl+TjSPeENg3FjwYNKWndwtUv93vM581JxCyJNRcOyK69cCjszsoFGmcNOMpHTOdA2o47/Xpf
DHdYoNA2cBTlRnc5xJ0qyfVDfvE0WcV6AXlhkyNu/YdGV8nJSM9qZ9aoa0O1iOMapS5Vw2jEu3k1
SPM6nniJXUoLZ8Nc04vuZya7V+yf4/4rm92wNjeUDb9T9DfY51qSpifuz5gg6JJH7Q38c1sOGUCS
PsVVdlOlGROGa6lxTmks/3VOh5wW2PzM5L/TBi2p4hZ6Q+FPAnTa8RXo0hpiIFQasDTGDTKM5qRK
I9hrGDn/z0bjl/1dp1p2SBy4xVk0CAD9sHwGTMRAFxwYUkKGH6RhhUEbWeiDRFCYXKnwzM9FK7/g
c2uLCKp919tVNIT78V05YUOEQIpNML1BfNbuCGR2tl9bxhl3W0IvEpQkGQacMUQpjhHFXnC/E8bl
wQMQyKqQQ+jqzIuHwkhEaaJT3vmAHpeVc/9e2Fs7rSlBTmElytjovxqE/gtF4+NOmL6zU+VwE9Fc
oRMM6id1NTweUrU/fP2ZbW/W9QY8txzAQdxcCM40sZnRDTmXgJCbfhgiZqkW5hFa+F3pcaR4j/RP
4+Luob+/wegmeMe0NwKlOkQAfXw3EjN8XpYRP70DgO+qvUJYstY4pHwTFxHluj1kKVjH21QlueMG
kBxswa3J+2rMu52iKaPHBVQ6LSAYvsUMujfQ3lkmgFIFiUkHktfwymlHMzu4RBJ4gqqUs8hHWgXF
Atm0+6+tSqhX05jDsSg/NAwL+JoW2TIvyDHm6wybuRSnXBGZk7XgELW7vqrQAl/71ZbQCIUHO9sq
AXW0hioZguLk3MRB6Yugl0TCL0eAnYUD50Nk8074Mi0z/TxqFHfceGYeXornRjperTGLWTzAN1gX
jFrIMw64epBBrfESXbysq+B/pPpzcARyx5pTWKUehY60YJOb3BjskZZ5qNDUXK3ATUAaDR5YoGLf
uQA8WYGzYZpG2m2W32E7BbT8jIH1BANtaCSG8eWNaJ6hoWMTunj+jVvPjfJYV45dRJeDK9fDlxm2
9NkkKvyojmV7mMCDAKeRAmSsu03HJAYSNHj3AU1VR7C/42Qrk22wOOGFFsaDkowUJzY1XP6ItcYQ
KJTbcQNbiFu+jVjjoBE8n4QzpD8OCu/omFGxhHUFyLxIJFCb/b9arjPLHBf6bwHemt6EuqQ6X/Mg
+Rym3f5yfU9hrtYriD31wZrJoOLspvXso75ZBB7kMUrMt3gwkeBNOu8zY5CTyLCsju+9n3C6byAu
Sn85QEDqc4xeJMu+KbrthTrIYQ7Zkdehy68li/evhOqwqOLqpj0b7boNj6BAMes+Y7KZx/QU/S/I
LfaaZdCwVdKdkiBnHPXUGSkVz6+Deu6FxqVUDkAQzf0VtkfU7RVtH8mqJcPaw1ooT55x5MFbfak8
YaUTSHkTpOiIEDtQMsu6E0ZI6kugqf/1zVshpVgde+jpV2ZwExsREQdXxFUjbp/9G3ufjoSPe8FJ
h5gYFnZhPIjQUl35SNpIJw4NpuCEx4Yo7x0L/UUH93OD3jhkj1DyflgjzmtGOEdMjRXpGY/UrsbL
8VESuWcTlub5pNQwPE/VgDxYrR/gFYf8cDvS9R4XTRNXGQrY7IZBOFwbGZk9fd+81FcKb8YDkFCy
RKfSfh2d8jNzFi+OF2ZHWNgzSAILzUl6J5Mvbtj3tRI52Qkqj9P16CN/J2H0/w9ibVnPKW1OydQP
svXAFUuawYspzaIvh5Rg3QdzQJzCqQOG+inLW66qBf58R+zMmr/LShXZLFzNsm72bB01tcXaokZZ
tVrccsIMqn5kIK6UbNqdPepZOQZvVjLC2sUUTAVFF8DGCgGXp/I+K81zAz1GzmT1rjSiNgRpUAHK
ARQSnjBE8ECM0YJ0qtGez8kPwld3dH4n8Jp1UMgN7TzlNKuGFqiC8krQOE6l+BN20bwI15jjW/CY
Nt3H2bGEY16fq666CoNQcBR3R1xZi4ViqKmk4Wc33CL1RXmW4PrJ9XqGuxXq8Phy4EvVdb50e2IG
jDcM35yvUgvivYBMonYeMhPl0vBHXch4d5JLWchKfz30x/Vuj8CcgG5mld8o6LFaKMVxkxSjVS+o
bV1PUmiIkB93LiFlZuCHXT1g26xhxYn44S77vsu2WCMxzI/p7vkWt+dELyFQDS6eGLNene39JGSX
G+IWKAooXP8ZpAlM9ETDiBwyZZ/5gZcQDAs/elP063zppUTQo9wPjRYiFZ4nf3gyEhYIUgJAvxAq
OwsmpWHCMnQ2+LvIAstxRSAQkPbIQrOh1MsBPe9d9bCBv/ihYIzNzy6SPIp75tdKxjxK2alinx6M
SUIf9YNeb6TkJfkWGC1CVGpAWrEQDBruOscabjK8SINhZF9WTD365U7l96Sndm9tq1eZGr5N0h/i
4j/aSSHG/X3r2TLmcMObeKpXk9FwFmuceA2UiiXBYzX5GTDtg7OyQAG7vk42uhfvvI3mettJp5s3
wUvfpXREE/3fcwUJPei7b8AipJxHm1jD+lBdKkElxzOWjVpiIdoTuKbLal3jb58Vo7euSSRWW1kc
XE+fcropIsq3rLcR/oZgOxiBaI7h7RI5olesePtWFCg6l27xCQyfQT2rAZwpTU600bbfzGm81e6o
yeopaOdkY6o5GbfMowK4vUAm9rzZYuKednQ8WId1m7FgdJzJYFHQjqmccjWaw0eBf3QROckFywqh
OyRKFg9gvKyjX9CEkk9J6bFBbbkyW/bSwyIZ+q6IG+iWWHSNqSbAARvpnaQ37X02fXEs9lyEr/qi
l/hS1rI6yvwmxlu95+z93xvQzvkksLwRe7ixf6iuo7d2uFyMQY70SwuIYcCVaVr83v/YNq3DThHc
BoMo/mhUO95wTXSCcAQEzidzzYrBFStW+Azp9VYRhpTWJxvpIpBIxrRau2HkiJLVmLDfR6IkWG92
2/fMTLurSKjg2tAqKdRrJgyWx1W3c7FNAHDyKvaQ5mHP1nynRlptan1P5ZJK+F5wavocYpr0YyRh
MgmsFlYppOrueKSfcGsWf1ENLm1C6Q9VJsYn45q8BDMdHzDGFWZ5wRUXjzaM6GJIPo9rxkyoKO3K
P38dzDoByBE2xh4BcXO5pTiz7oK+QOJBznL7Z8YQWYQ/1aSbTAy3/nzbSF//2rp0XF+xsQNlHBRv
8Is89k9RYbL4c2Pw2/qc+7zM58C83s/foZCt+cjcQzZOF7/rP3UClHEKLSJNCRtxOUZbHnNDeWCt
nAeremLTYtqtwv50vxvmc2QWayIG2wZewdgOh8aBMCK6BmGbtKwRHL5PiIE/JF6J1XZ5k8JopjmW
6SkZwqOBJNUcXYmN6pFBBqTLtZL1xerMPobt3BcnqUcZC54Pjn6njmduO+YiAGY5s5suqd2+wnRI
9f4OBK8j854FWcz96ZU+VMLomk9y399IjsmMxkiVAuu3Wd0cnCrv2uY7r8deRGawIVNAgoCe2fEE
BFUUeTwbgJVBHg4lHc1f4inH2USQTucONJ6Rkt8rv4AyWFU2SJaCq+eFZxMPlqDu4sb3pXjCu8yL
kcQT+nQHsbLFyNWWUD8rIalugdkf5BQSGH4TLT/35kjpkts2UFc0Xkfv5f2WDo+HqIaLF7eGYTlu
SceGlguXmcehJQbsXLvHtUYxCM4qy4Ji1D/J6+5Ozy0CEDzDd57z6BFXd+6czzGJoNyBq7HkcJyJ
1ycAu5D/9XaW63ieifXrnXQCBN+mtuJKMv0YpwxmSvc7JccQfy5WdsuGfCsuvJeNA23GrGjdqY53
FJESUdEkmNes+wqaQAamh0lJP9vFrDvnPkk75W01VjTFDpyydtGPiUJ/nKA53dpkEd4L4dqhZZg5
mvgK+lD8XKqo4hj3sSj7AxOo6XvBMNjwdrUqH8estRIJJDTEawwqc12hyRvd6yxz+kKDYGgalQnb
sYAc2w1qTI6Qg4DBCZjImyP7y1bx7DNB52nnUyz7+3OwC3Kj0JrAcigVtoPghR0+aKHx1Q7wXqa8
X4pQeyWPmuTTVBQE3xsalPHUbThVdAtCaQle378H9SOglSwdocNbPvcRwzg8waF5Pp724YFI2i8K
MgispEDa5jApoTy/dHU7Kd4XDlRyr9wcCWaROhrh+ytp+xJqUdqetLtrdDQ94RGQAtut5OLyeyhn
nhwF5FCaOU5xp79zpzNtVI5Y9E9B3c1Ly4YGTpXCJFHHFTqaTt9OC8+/Hru0+xbj6yEI6iIvrjJD
U8cV9MWZtkIyH2eBvH4H9doCFZEpA8zolBQC7wIE2HsJLA94n6QN2XBa7T+SgOvU0BxndfGCtUm/
CCTctpg8zm7Dhwnzg7URE52przpCS8yy5zoVWUsSzE88Rm2aJGOm1628k6MchNcrOtJ92YSWPe71
ev9+8PEHOjSV/wgPznpIyjxNQnVQIWdPgGlGVSSwtb9OAvxGzcuO67v5EXZ3P1V5XBeFtlbM/I+k
35s6Hu51Iv4oqIP6JVk8axXeVgB2vEIQu1lzAndJ7Rd3fcEWuCSK68bOr61HTebElgO4pUCxbNSD
KrxJVYK0IFcktriyILOUI8GPKT8qtvWxtyPw4fFlgA/ltFx3iTpHKDYN5cUjMFUa7Mfbz627T6fv
he1njiyEHPUN+0rvjd+A/luuqJBDf9RW9rt9iDnigLaIJ3nCmQTRHbjnOn2CzJhrFVB2dKMoZ9ls
yXDls4JJqVbFdMW8rk8po6sTaW5tEMCv9UR45Pq4M5LBf611+uLlk2aIaBbnRteTeu/w1pKvCNcd
3GlqkZDSvojA+BV0mTZiqz4VGiMX7BWu+NZ7IJxEE2S+hknbTDLn5abF8b7WfWUyHn78V4alApfp
B2yC85OMWbWY1fpaxst1Y8O/BEO5u4sYFXHLbAe/HoHR49NR/jrcDG6LhOpExFZEtnvRKh2mthpH
o/l2iYcAAUmZr9hFbvy7XtgO+MLZlQwLAUq2nK6+YM+xGp0bn/D22cp5Rp1+IwXAySH70X6a8U2W
3hRRkQeM+tDxqIwkunujiqEzMV/S8yymrepI7SwIgkDkvq00T+Fr36GJGJLmO4ges+G9Q2nZ3fLC
CzXLUn0lHN9PdXOdNVgxew5tXxpUwBR1uD0q288mTpnGYxSHljF+CpwjY5V339YXwep5Iuni3wPz
8hE/EPWogjOLbTcuUyyx7+2qaMe2XSssKy0im5wZwyg71liuZt5U9D5yzSY1GIHmaK2pV/6MwQu2
jNhsM21GVsBeuNZuQ/Jr3gK+PXa0cCCa19UoGj46Trhs3hjTkFp75ZmNcIIKg4aiRw2IGvzRvgIt
jW0fF388WLLugjUyMXSWh4ELkfA/+O516Fgo5ZuN+8VeSQRyH9nTQ3JhG7tLdWUnj/2t8bikJMra
325a5KDrTl7NvVYg0Z3tGz58nkI5T5VQNP3LvflUa1niF+q+Kt2deXU93Af9pbs5tSS/001bZ18Q
jBqwNhjZ08iho4SzY++iKgWISTPP5SnKQNgnjzc14f+4eneFQPnl3Ru0cXneQSJcFxbuRhJoQJpP
gJ3ckcjIcoUmHlOLAC+TeMwZ0zMFOrXHc9zyE0D/ZJzzCn64J9rkwauuscgNlcDTtOl0ZUBkHMe9
nku8LD3PH+ejEOmbaLXHWFwaekGThKGKa3m8KOyDletluVDY/7/UpQ98sXvei0w2Vs8bJjYTQZ7C
iZbpfKqrWneo1PsH43E6cWQ0pUF2NnrBYM+UuQ5PA98eJ2i52HTwgO2OTKen2peYp5qcojaswrN3
v1oWczL25Ht7qNqS+hw0F4rXLAPwt5R/aQ8jKI0v+gWq6y5o/qaRpNEjk2CxrbtDg5uCHuy11XCv
A/cGaLnALlP4wIB5aFh8Xm2uLlSQoZp2EWq2y82IIyUnGGcTPhvzAC1guBl2tH/I6vtaksSqPxnd
DTPhbbBe1JOaa0V+kWh1wf+uX7p1LsF20GRf8JMngvZRhiw7oqxqoyOjPLQK1cTmiNQpwUwgb+ds
K2JYC00RNyneokQGS8jDgs7SlXDJfhN6ENRzLWhELLby44dypVnEYIKxrc8TooVuMySgDhZeahtQ
L/NzAj8wh7BM0SDFub8t0aeBvSBAGjleZMBRnFdH2HPIZ7hmbqPrjOKeBXh5nlMOn7+569pKGDZu
wNcxepJ+jNoB5aGA88yV4DDsFKYpEg/BSO4pE4huTaWkjqSokDPhf/NLaXutNrO3PeCPsqyiQ+ng
G+BIm92RCxqt6UAXiGk70hIxB+xIuHf/V8BxUJy1/n2H/kZ3R7pPXCuJkIjGJ9Zszi8GH512kqdF
xwkKv464PBpNJGqGXBrbFo/88vWXOGyzEGoYNwDTNvckoAc/3nsKo9iNLoyvwX0OD9v5cqFMX32g
7n63mdf0Ha/o6eokZQY8tONdO8KkReC1JGONXKffqycNnCzPd9tEEWi+X1k4LJ2Tv8yPdu18mnCm
S4XgVu+ZIQdoiNIyPQTfWzP+h74yceeRWaqPz3NwPXm0C7YhvC/eA+p7EGddeT4nTEnv1htgchQt
p22ftavA2OZ0psXVuQ1R60+rtP3rLnvEE8RM2FN3IH7WNMEx2nBOF/X9M6HBe1CMiOfrbvyOd58F
YvkSNFfXTKl3TOfA4HdDe090GgzPbFI/600OLX0u2UUhF868OgDLbpW9tlQsRlo8MPUtMpMnXzfG
iesjTQJHFjXccH53rcn4LaYlmpYPzfPBMETxKFb5WwYbSIP7gGYvS6i2F6AUCUCHQvUxC39nespY
muZh/bV5FGrzopNQV+LDQN/nnIyzX+rqAvFQxfXasK+x/ZSWxDn1PfAsGl5+PflYKU0wHHE5BUCm
5fB2KGhp15psvW+lSTcHccAetAHTkATscRmKXstZDbQVLJw+HXuJFgTYQHYnbJf0XkrPzvTZgSCK
sdwjamru6Z/+2Vs0SR6cWtN+N3T1U3qFxH3DmFcorx6Uu+cscph2xmIgm1Xom3J3H6HXlzm07s9U
dOylTgjfUHjADxyZKpYYCRHaHXaCus5so8CGwJKCU/NZFqP5S+igQD2XPLrTslaw9d/5gxnL1X1X
x5reYX3cDrOikALuPybcYsPNk6kvYbfb1xjuqWKxOKl/Vdw/1sxXIINXUbI/g3qFW9dSkJpGOTOl
ugZCuYBth0sfx9uLtZ5MuFLhlvoA7XBFS37BLJQXu8VIAClf+HPgTs8iwLpjGlsXVtc4Ut45K1k2
ld6ULzO6ONORd28Mq+de6CaXYF/ocozkapY41gULQvs+6bz3piCS8GXl3eFIW0nXGfhyq1ttpWvG
26E/NO2dfXkg44eOnke092SeP8Vi16LkB8CVYOD9LRm54zciN+YYzPm8ap8RsivJwpl3DWRHdUEm
XVqxbBuxImpOQdN5mPTHzzBO7cspPBWfs7obDjtR2rmt5Hh/5z1Qhr4SBTrSnu/nOtqOWb0ydGI4
LBn0QDWuF35uAHngyyVRlbzy1LRmLyIPPCjuLAWzYYyl2cbnvd9xVMUeqNcMeksMz15VkcpSqtUg
Vzeftxy5AeqhT+YuIMudJYFcBxL1wb5f7mKAsR/9SLNYNSCUaCv8PG/7zRrhmxvJDqTtM87BnlBo
7s2Cv8sO/s6TMic/Ze7syojLQodHVeVs8eLjldg9KqgYqxpKNKiQryhbfP+3SMm8SZE5hcRvBOfa
EgfFZIMEXZCQzQNVrfIniUzkt5OmXvrrNaSAArJGMh+lxg4hzhiGhOi+6YO4mQY6+AqU/kD+TFsS
kfvlwqaFktg2bYRRzvAuSGsLg7bmRM/tGPaMwWM2mrL4TLOj1GGuoHN24Ji+w5Edk24W1XDEYB+2
juCSJTBX8/Ulmr12ldFHLdh1E9243VucDB5jJaSC05ScXV8E4blCv/+YgtkWKDzDR7LApkAs2gu7
05qFL0l9x94GeEFzVHbmKBAQGThv4+D3uoTkn4wCdUestrX5viMuLgj3DAjMZiRkFH7GdABs6Qhk
6f7eHdGGx2oLbAblLDCRF2gHovnSg9Do339nMMoRndAd/sX/aIg8lJgr0wkvH8DQifQbmJMxBVVg
8xUe8LZDjKCKvjUDsf3BgpWd8WEo8mVs5NQ6b+J/JXZy6+Nw7mU8PHLShBhdGu32lZVa4FxOCRxX
uigkSitgVqdQTT9c76Z8Ko5BoYe1Rj5zosIkD36v/HOGm3svcY5Z41DwrglKFLNlSK8DLmRxTnIX
LnqPyRaF+uft3gY0cZLA5xGkWO5OPbKJXgYEZrHvpMnQp9qtolQbtIQrJbaEBHjbVQFvueX6Cj2a
FTJbpM0ksA0RDcSltq0445V6q8+EvkIEWKn5bKDvELld8gEnvywcSFfjoRF8hMQFz48GgdmMYgWF
qro3XHhqXPMVXNAqvMEd3+682AOYNsd9wgAzPGBexBfdEffA/6uqhdqND3nRL3QgCorC0V+XqneJ
amOGkeGCHBUPv8gSgP04tWb3tqAdosiPxLD3HU3Qe3SBhcjtg/2UFprPOgAtP8asQnCHMsonLCfA
xYElpUJucMGy4qZLpqwJmFsRNDX7tACyGXBAmvALd4PMvApc0ZZifrfKqOD3HS6dhs1Upr+GkjrL
N2w33UnrXBmoA/YZBxM+yhn5dtubRVaDGq+sV13xPMiZc6lDkkBKmF2gGlrkjZvw6HvA2iZDDoIp
1wAEsRKZJce2CFUlWiwn/nNPs0moXZh0p7Fk9B2emvl0A+G2kiBEXToRC79Y6L0Q2/O5X3IDWTuP
lhYf6runY18UtIKEz3rL4nJ6vwL8BcQ+SqBLu3ast9iNsq7YLejVDpk5bJmGZF8QCVnX+f6GRXOL
sdfTYr6nh6HHHzxKE8p+f6sYDHRf6pyrndUDA4FVeijOS/ogHkLLwukw5juiSxMK/aIOwKIJiyv8
spYtw8RSIMCAAArhYGKjKhNWqVjBMJeE3Itc+zeWCgod56hWGnTfs15V/hWZeyZ0jcrql6XZtT/3
K7Xo0Gbj6dPV6r1gt1i5z7XrrfVAaoFVWHqf9t7B1ptdpfPQSKIjeB4VP0tozLT1nz8zlD9AAv16
EnE9bWoH8PWx2uIvgAApMh5BbSDDcyi3wnEKRguEs5FJou0pJGGyIz5pQHBIgAVF6gKl7dgMjo3M
Eukj0XIS17wK7r1G4i7AD/QNMfng+5WGbcdPDXJmTUcRX2QWPC+tO8fbM/ptPK80iU48gj5snV3h
8BUA/hqMb8fqM5BrqvhLPN740iTvei4ys8HM+w5oa9FMcWFOO3PNLngpEH8ogATJgyxu+zXDypV9
6aXVDiBVGCggpF3SvvxOaqh9tuFvOBx4t2USVxCvEBkKwNgLC98pWB3bnpvz8wsPnzssIwW8WU+P
MNyvugdHg6D6hqoJKw1nngNsOy6RNc22uqdRNqtiJTT1KE9YIKydCFsb1JaNmPT+RHwDB2dCgpWy
YoJeL2WOiKr+OuDJdXqdwEuWyw3g2uYliH9VjSzhmmaV0WlYg/uLMKfeKEj4XZpepKC/JhXR/d2T
FBlSKSA6uY0Nx1IkHCfxCHNL6y5NB8hWuA8A+NL8mHxeQ6DfKp58sLr0DVvFQw7zFp+agDqoOgkn
XumYhs9N6BsFvR72eIg30jRbsdx0fdrGpHJbXr7FB2boYfQXiHB3Qozcx8a+LGOmdJ0BzMmJGNhx
6fD6ikS6mLzvkdER5qqjeCxhHPW2OIdYvxVfBWeT4ZNyJ/pzTzxoY55z7Jxgvhn9AOK/RfduC0wD
2DRd6/gws517UOOpOjq/2vGefLOX/zWkUUt75jD7SA4mkwV52WZouL19Z38177P8aWXD2UuNp24s
0H5PspMl+6l/of8EjtrwCdAXQ8K3gr0OqRRFkZ1THU6snDGDn+S1pnPrzMFVupKU2vMiuni5PLqd
nCQfg4x3AL5R9DfwqOvNL82XG6DNA3MPediABt7sDv0JLvK4ZtAJQipAjXCetzg4VvkBxY15tYED
OHNryvnxgKnIgez4chAKSYPbpes8qCFGIDeOZ7mYwkJ6UuyW3V6jcO5LUxychEErfwzUdd+jNRFU
IBvO/A60j5WViPSpBEqUebAGk4RzQNx4VgUuKSJ5ztGHNQx1Koof1ntPYgL1Yteg0vN5ujQqX4uJ
ukbCFOj4kaUNdZ9fCL4YOSK4Pi0fZgMPpolDMdol0O9kKF0vq3ucTvnNiwFoSGXzr6Kr2BzqhMMJ
cWAB6u08B7WvbRgrlKmoAbvbQC4brf4HqhuOGfvpfankQ/nUaxBVbx0c5AVY89hHJ/Le2SvdP4xi
nnIkhkG3O4E3aKdNDE30esjgobJIEye1UL7O1WD+HKff28HuLOkOAF7ryNaJTm5d70ZPwSVp4mxH
KOuuIJHsAi+lniOspPB3ywsgeCgI5ukYjfuyc1MQ3QamOnlXAnrJoRAkbioUHFjOmfJH5iXwd98W
MhWb3Gnrf7YYczsjRgvWWZptjfXBGckqBULu/aT5guUdJmcAj7JSD2mkGfMJaxdBKpmjJbxXM6do
6lwU0XL8lajg5xqk0YBUYwHKePi8gbTDyr6lXwaga+lKdyyVNnESZOZ2X+jTjT/6OsGlWgvDBUyv
klq/QjSRUaVAAZu3AmZl/kA2F1oYPktF+ZFxzc17p5uBSNLpdyQa17qh/P7zGOOCRcfl7GCS8NGS
36Ax9sK6skx1H5rJNEanTPIYVGj4633OHCwAndF4/U8TahCjwKnn9MXJWTFBe1W0Qa/MUCG4LO9a
rSgqygqCcxU3VbK5wM/nZq/phC5D3Gd/4Z32XznqRiV7GFpMz8t5Dodl2eOPHZjLZ4RzGBUMQYbe
6xtKy7tCqDwwrYbBx014Sqg/njIl9bMPMoJH18G83obcgQrlgXEAXzq+y/bMAxwBg92JxkQlAWuX
7Isc1eltiWk+jsRCNm56qgHH1/RvI3Ej468qtwyuw/d4VJmNMsXfrzXWIFdHOX575mc7zcNYR7GF
ofNaJJzalkehTMoVMgIw1N11ZOS4fgGpBe0kqV1VtUo7Ah6gv3QwOWg7bz8jlmLi/B+ZLQdLeVp2
N0w4hmoxpgSYAOauYtP/6UtHC5EJGU2evF0zvge2Zc5PjgnzmD2+cJ4uO5A1uB8AWDChKo3OEb/C
LCs3YBU2D3PHjvGsfWl1Hgyp9tylOpkldygGtKVllwB9gU+mcWhozwJNln1b+76QditOW/q8UqJP
7dEd+2LQOe0mPxD2w5dxxkqExUKEXO9McCf77PXEZkMNMy5q/xZaCEsHbU9beAT1pOfr86jhk9vi
tRd7RaYot690kal+WbbpsQPUKLshwwBg/bwtpRWkDQRC9z/9MvzsTDFvmfSRjTH3TVq2PNl2irob
oG6lk/PWtXNHUvf2Rhxrje9qNSP4FJ8SDC5Wv18efu7d4D/QCIqd3r02XxFfaIXsSXJYZOjfgZq3
Ys4JvGHZkO7lLJf18FJ0ZBsMCxmnTR8ukP6VZWWNU2m7WrbDZPtxBP/XZ9CYhCrp8qU7cDymOc82
6iVqDDJjqaJnbA5H/QpQBGa55hl7k7xub7nfB+1UtQdNxJdLDBZS0G89/Llq1sGQ37kQ3W5C0MTl
igluG8xQnRVLX44TrpnyCtJ/n15YChyazbDrpzZDWsqilKCE3TL2j2V5TUDAU6DqqE1yNq2sFyr9
VsTw/HxqCqtxxiC6C2zwmkTXZBNkpNF15ELxBKBqsz5MSvUw5kuwCx9LY152XXWLequRD9GgodR1
SAXk+9OxrmMoSM+cYGs/AQYie+TNm9FOfRXEpEAC4OFCzIVj6m4kO+HI0+Cu2drUXOMlskeGxYt3
fWrwcNiU0/kgTwtjCXVcfW/5hLvGsO6oCWJcca206WOqysPUG7g3rH0qvNTuah1Yg27jFh3HnWkR
/yzIVqp+EPae+WTQ/eWO1ZfWbj9mpcTNdSzSeOpoT+LE7++Rv1WjUYCUjK3vfApET4xxN2/FISVB
8zVq1IlN3BAzvNNSCfy7tOdKHM07jjygKInSErdbfIOHw4q2YA824vfYnDWod2/vps4ThZ4Daho7
gxz/pfDQcrT57Ff36sUr96GLKlX/1XA4URGR4iUu0AwQU/eD2ldFBAQS5JWYHYcY0vnRi/oVuPR+
GJL/XF5nRi+qfDc8KZHyxyFT8t0DYNKGy7UUlGqYspMHfnAOQGxE9IXq5wrPPPOoHfJfksR0P5Lt
/yLiMvs+QK7aMIZdvD1ZIxTyveL8+vUbYu5Nvl6FifAH7TQkPjo6S7CidNrSBf35nIwLWMVe3npN
JwcMjjROp7WWTB/etrqmq+vIdzgphJmCNbkGJ9ecdjm06mixvSIph9KLkbjpksSQ+ct/NWor1d7h
T1+1fjlSLKn1CJfImrxm7hYeQ2Lg3ec2m5lVxygtYRkZd8xIhr6qTCogyeqAPYydms400lj8tC5o
3ok8rr7xXKbwT02s6N/BvxIEUi/bzHXA9WtL90x7yoJ4rjF/4GF29mYJXscRllu3CVX2pzWsqvkA
hpLPZ1y2CnCEOYdzjlvBHG6KaSe2+NqfaQhCaTooPsT7gIhzMNvR2gQM/AdYK+nk4DbJJ9HCbWb/
YcFgC0N1Z0pJfCr+vRc6h9T2UNG/y1dWXDNbEKuUyEzdFMeBKujWtrSUHhwuIX5lCRgHLzrb3syt
Qh96LvjjMQM3u5OLdm52sa1fuFiW7AwFsjfSsL5mlN+LsRcK5crQypNbcKNm/oiD23c/z+u7eyZS
MY7VkvPXcmi9/0Hs0QkROHsLNUOnp6kYUyw+BkUe9+j6LhE2h/mnSmY/4sxzbD8LKf8WfwqD6dUt
dGSlZM523p6mLqv4YD7w8q2opsEJTlmFTA8kTnYCNpMPrXl9ZmLRlt5y8mlsdyP6vMXP9HmML+jy
HPjky7YM1KWIaOC2psJvInusyUoPPkoWT5vSE7X0aYgYBLnPmZiko71S22oDUtoxKnkrrAV06ThW
oTCfaeoWNfa4iXa9s9IE6lnWtCjd4SM5/w//Pcvsk25CrPplWHb/wm0KGamgJsgsmo0M3m3DfVFK
fD8e2Zg+MiBU3fD8YpU/Lf+kMtSMyhy017heRDJ7Z+mRJp9gbO6ngQ8c0TOZQpAFVf3OCFKSvhDr
6Zkanl9JEqYB9Q3BT/g3TFTVRv22LzQwO2TNc1pMxlbH9KYB6XpExEY9uQ+Dkf0aFPIFOOeRZHV+
6tCTkVyOwutYfN4vCA19lZGPJY6Vv0KJKVJ5J4ofZGDBrTcC9LtjQFOQcIOsCK64ZJnXy/ur1eed
Zpk0IZjXOU0rKqA91lYqTHzThwczIQijY3g1ZRZYqXLfUx5SIyiogA0lyXXuh4AUlhgm9GqQ7lg0
6xXoom3QStbjjnJozCNhNQSbqxUrRlQ09dHC3Vt89R0YybnjPIZ+r96e83o8nE66OAddxRHfaLxl
i++1S6VbGrSKIjW1CSySRQU0E6uHVxFwm7cVGd8gTlgdQF+T1HxBfpcui2ID6RM+/qB6hCJjmp3u
GGCdkN3M8TmDTQK5NogE7YUJwK5pZzQAd9P0tBv0YmYc6ZI3KscGKWtb5S0h38bBlOGzhgYsKsrz
WRYitkfQVrU1lW5g7q8kGaFbLm3WNq9UyxAjMsivS+FCP5ih0xBRsV/mdWBlmF9TCWgZy2TXv8Xl
KPzNTbTEKflM1XcSLJGJjVcfIpSCLhK5avjgcSbgO2hbDd0ATpAvTDhG6KdeBuNtAoRiMgGiXioz
ojRnuG2qxw7dlpm+a7F3gksKc/RCKgcE/nMiISUPU4A9byZ+01Ddeo4UvXpjCVIUAwnZx8krrAu+
MbzV/L4F+ORdegGoRf476WhjHKycm5dzArOQFq2+Mbauj9Di/lKfmvgMHRQpaOrPgSw317wZBJZ5
BiItLxwrKoK4PIwkzdYiw9TBEU6vt7njaPGBDMse3BHgSpdbdkTjOaHTP2Nji0QhLvm5z7neeUw8
Vvcdz79jFnt02vO2wThQGe5E6Fzxj1sxDj1DIqzxhuTbGR1S9aYVSYjcOTgznxLKO8kajZ4peMtq
JvFjsWKSyWRFOfIjtJbWRzmx5ZtgyJ7ncigk8PxwozPOX4PqGsiRhcYtYoWxYXMHJvBDRk8ls4Qa
n6q0KE5EtEW3dDTqRDul8ctArLtxKChDn6M/YY/n6E/A9tuxJfZtsiZ6c81wOsptXWyheXs0T0JS
a6vZc6Bf4O5uzajyaOJMiqK54quV4hFQigR/lWiuNmmxLUqkEYhB4xJtVJQFQOdhXPK5rGht33XX
SW6a1MrXJ9Epd37ayWg8ze/W/fQTYkz5ZNHWfNeHAaUeG7tTvxNVgfWo/9L2gXkM0gmd+AtygTmp
QKxj7qBSdtt0JfSq4j00mkZMabc882121Gap+APHqIMllVJJSHuIhAPK6DedknTt3cFM01j+E7vE
bU/d7xlNIz52licsmcIsZa7BmUv+Yie7fWrOBlnKuH/9zvshXqHZ8n/hIG1CKYi6+VK7Rwu74XBn
EYclfe3psTPLBTgX8ZVai63O0gj5E5dfC4BL9p0tjrcQ6JQj7GxvaTaIShg7ailVkntQq8iahv3A
m7H+UjDE65Ev8fS+jVmLWtxETH6ylixY+UkY043ybhMvXt1pb01CksVf84RGOAhhwRseG66Vfq4E
ohEmvm7X36MF8c2KBqOThaYGf0mYIijlWuru4HgaoyRxlLvRCTbhG+Wey8AMeE9mr2jibHLkcbUe
QZAujNymvA81NBBOMgRaVh2f16InDNI/SlAkXx4yRezGz6ero2pKXRETkUFN20wG2uY8zfr4VbP9
+5k8d3DOIrEYHqpp+0LjuWN5rJnvxU1FFQBIV46sp9quDdhGRHnvGh+ZHmSLZ9zqksK5bObgotDr
L5ghrdznxAcIclJYCn2DSIaxa8RO7wOHOodijMuM2CPR+AnPOIF7gkOEmN3BVQZlRSu3nnwJa3UQ
2u41bC5ATWu2srmgum1SWdtguFlVrs4myqrOGX+IBvrmxY2IrF1gHbuyAYdG5i9r5+j9hLE6sEJS
c2rKbp4aypmPNI8nSY0JYx6HqLcRTxkfurXIAf0cCwZUMLY24W/yds9pdCh3o77GgHDRr1kFse+J
9y6TK+WCan4Si8njBQluU0w9iGKmogyajI0F1uZ9NQ7DvHZFc18I3GQMnVAk/tRqfMCL5XePtjfP
Nw8PeIiOlNZqlUnTZpAt1ArwglvANwVhwBfzABxK+PNePNFukof1PdOGebT0YduCLwIM4/B+hPCN
Q4+xcNkhXnRmUK6f6qxYpsdfyal4OeKdNwr05J15DvNzZ+3JVY508BMmcLYA3HgyIhR3YgTtasye
9i7A25H1AXZNlv4eTxPDf/wZIxRsR0Ij83Flp6NtgOOulhd1lIq+jp9llfS0FGPo/JnnyqjUQwet
DCkAUIohFwBrujlQhxUe4CsdbzhCiceVXAgHPZZkc2S4jp7XK8ZXgk6D+52602zYqHOmEcivMJIY
/1kykoTM+He9Q8qVEnvcItYoBe/mbzWCpR3iD6598qGd6usX1/tkzbEWhAY/pB4SAQXSTJxo5dXY
Ve/HozPoM+9B/mSsLoocV9u5zXerTqhY6U6vvTwD7KQ6RZ87xbAYPTOXyiPa50OHqCdsO1m4UMeJ
b5jGTl2P4xSUczq3FPGgfccxCLLaTBhnHdXVLeS5DsDkpMWZEryJFkitz/sn7L1/PPkGmGjQnwQq
yZcee6p0ErPvvKHUH3pnUpbW5aZlLuxnprHQ68eOFUZHCbHsWuN5d1AtYgzgk1sTEAnmmLMDp+3d
hsqrx1HzVhRVxmdQ/6BwjV7VdE6UtQgHXCsskNf9qYqy/nDcbnHyXwnm6x70V2I9aLAjXHrLfsva
3ZD0NRCE8UwQeIDL4X0mXIWC58FGYsciAwepDi4UcnrORddopl6ff6AzVt9s6KADftbnt+mxm1jo
DhSP+2+qgZ8r7njhOvqD681LcYNSsV/gXNJIkH+uDQGNIR38meYXYoZeyv+Dx2SuExq4YEnfRcgq
9l3VEPjGexuajPW2RHh9laBlXRB+8w456rHItTEEol/0ri/zVbVaollrCdoqApASeJePkwfwRpF6
8h2PIYvLY442/ar7yYGPEBMcNHbHe6mThdb2/jFfWGH3EFBH82cTDrrvb4JPsPqq1ApYFAVFznu/
9rw8S4/3dG0+W01vZ9unMj8MnGb/2srrpptR7wd8ajlcpHOUbKATMQ3fb9AhmjC96OG/3Uv3hpel
Dx9AAM43t5uH0j9NV2VToyq1isTquZdf+saIn9Kdac2XOH4P2a5vwvl/cLH0w4RMjSkmafLUECXG
E2LWqrm51PH/f80cQ8QuQEkF+hyjqzrPAbLz51zhXOCSqI4tX/A94LCEs1Efbj9st8ANe22Q3Q2M
UhrntMPXaxLnTpmlw6R1gzjCC6RpV4Qa2+RMDzEKIcjNHDJUm76WQGMofbbK++m21u1AtjGZrlMh
OetpC5jkmjOGDbScoJkA/wcYJJnRlw0rOOnzmG8zmwNksvUltKHmQEtyW5gZegrkLJIiqa3Ah9r7
EKfYFHHsbsIVC2cgQJfP1m+IkUmAOiEJkZuL5VZ1xJAHA9/i6V3KuZOHh7/yfJenGlpXYIKT+e0q
vEcEMLBRPWgpZfF9YBBIqsk3wL/0kf3i6ADrDnti3WDtl36/aTJEoTFmxCvUpke4mB7UDOOg4gds
JHY+/+ujU7dcLzQfg00QTirJ2LuFE6sBUqOZxe7/MgEr6b4J03Jbg3Uf3jGI4QXnO9fb94hXaL4Y
AmoTH/7op4fGzPzspSjow0FOpUeBVPhigP43pqraMsjWzTFtPtJAux0emPY2CTNdxq0Ju3JHX5NG
FI9OMncukhaPyt02r/DQgNd7t6U9JoqTdeswNlx+feDQWjAagc9e9aBbn8iZ+gd04vfpQKsW1SXn
S1aOqS2OCW679ZYE/PUYKY8o/GMDCVBenUE9hnV2bepY7c3kkuosGu3tsmSKvCfJBFLa8QkH+Iwp
QVYFah/WN1v4jE+963UraGogAyZ8l1nNCDWC+CDQqf6Pas2PP1ZydqDNe4Orrp6yhObTPXUOr+Tq
HGdrMAsc93TxgSD9iIHjNcR04GfvAx8PeaI/LvTYoUTI8MPmyVZ2ubxT3xfvi3Ogy+bG4ir8n2BH
SwNvhNLTNHIWpPRv5lYTh+sLm5HK0tOus/8fVayw952UFp9J8PKIZHYdmIQt9/9V5g/mnRE/22nq
PS1FZ+LbbczIzQfyOyaeEUb2nFIlgrIjedMkrrsua83v3UzUL7XXqvjJTsIIbBG7OI4Q66EWz4xm
7wPmEH8VcGStjoDqEyTW+S44Wza4zLzKBAuJzuXcT87eiRX3p6vnhEhDExVl4uu6J9wRS4474a+y
J2Uea/Y8rrXcBU1mUbfnOCCfIxoLZicRSi6py2xR4t1uLDiyTG0J/r8Nrb4YMhdOhnUUObmothYq
5Es6MeATqzHeyuC5x/AiA2nc4UMLI2XgaO2lJgr7W0W29ObJJx81pH+Q49hjzTnonjaqh0mNHN3Y
9Utyp7lm9t6zglrKacc5pXJLJWKaSSGZ6kQleqapgiFx8sD2zNKZNdZ4V5xZ4pOnuBOtNcNGwibY
P9veTj5Yxz0egPgjhaBu0jpCqKrscXgvpIUneAZxENmBM42zYMzCz993OKnLrLiob8PIntMCz4ZO
WsazZB+fL6zJUrmmIHI2lzp8X+5Sg1mzNnGvpdtUtD7BntAIKzrpg7mf+RVfg9ZdELX21BIAtq6O
iVw5+ibGrF4ZkNL3+yNtHMCrtLKy4qGFzt5BH2QAHdE2G7x97VWo/tffJTyo3JFU1CSfTKyL6L1q
h1YVLqpG/Rvwz15zyRZrBmzOSxsvsXYnOcDKhC12mKykIoSAqOQEf4bEykUKqCgHmDDVy4ZxILlV
LlbS+IOMKBkDa0+1O7Bj0cGitvr2CgVXelmrbcnnpOmy9vH4td3nMdFbBZrL5fAWWfDhcLyvrd33
lMyg0hzy4zpyuNWLhz/C5kspKDD30nQMEsGBdvkfobI1QE6maqd8T054poERWAe2l5CFFlKZ2DF4
iX9hvDbP8HjpDPM9yaK99MR9/dvETKJqahPTDzoc+W1tQst2yDzaBqDEB/1GdhmdlYlB2gDXWxdE
IKmjCyq/vdQdnZhJQ6KBc9hgsw2g5mnhUXPCLF4aY1w8QS2BAIcFrxf40Z03CW/5u92gKJ/yMw+R
pbFE3BavqSXbsffsnY2zI11hyZ6J2IKQQty34x5+htqRRHCztHfv0CRfvV5hUMaTonbNOEK0G709
UaIlkVgj7l3dkw8EEl15AQzTxlDH3T+JIq2dT7MPRSvnI7u0Icxj4dr32VWJuLXTp+qqAANyES2I
rxtQLylep5/dzNfaovcPgLN84swqPzDBwPKyEctXOai4bhZYHrjuDrrPcGjRltM/7Fwnl31kaHfr
y1F968ISUjVU6x4kyAohPXGjsvAxAf9GC8LW2miuauRYawIZUEe4emPP7mwilVCDYUz84WFnCtEo
/dyUD0x5fJI36wn4ZH0bJboc47ZfFz3pzsjG5jac0Ko7Z8vm/GwtkGgrlImp3h/K4vbYVx3JDzqF
FV2TWkUPWmhzuqACJfc5el1rWZ26gnnDe9CTeMEupX7OQAsU1tjTQzchpuZtFYJvDgu0v6LHlgqM
GMeGXwvYFbGqf6r3U3m980pHQuZnzhQbFB0oXqhGKnApnyZ9Bxk1kBJWsTmAzmKNRhdIXKTe+vbi
7cc92IKzRPzyo8q36lj0JmLRMg21AIqmWwtEaIWqAvWkYamx4OhDR8u/VteX5XT2++HiCJsYkLzC
xlsUedPPfElRLuVWOHs7cofogsTNFkxA1qgyaCDSHmOMmUpXjr1fRMFVBiSnCjsO93SD4HWhGpla
UnZJDmUh6wfe2ICIFP47AKrMkct4UgtrkBbDVKGHqxHXYA44Hu1alEmqXpHCt9aiq800XkjSLhEm
0KWLoRXderF8gWffmfft+BYYnUtrHgxb6F/pXHL8Nsax6TIWX5MwQ21ZKXaVgJeV38bMLgjLx780
jma0CTYRDTUPDcQ2rBgW+YZy6UUbDIg+VJerr3jnJHOOYcf++Rg6gZmlhdFHQYCNsURAx8LdZ67X
Ws4/GE3NLpyRQvZWjWMfzk737Yuub7BPtxeFu+BqzXbPyrTqdzVCVIgq2XTo7b//v4UnbtWZWMS1
pslBqpMpDxe/apwdXmuSDwjTIV+lP7H1vFGCDymj+gzgeYhYuceDXq4C8i1ICirZLk2onc3KQe7B
1QjG7vkhbInRyuUMyde0etRaFuBx6Fg+CqB2p4vcO8oum9LgEaHQKVDjVfpSDDLleVM9CM+Sq3Gu
jOnNh1D+Jqs/j1KoNSBmiEavTEVaYmyApC1o8YuqYUMaoRdFIpa8sNWgLVIxSkGrB/EKkAwpYpKV
PHGV5UDxx31MItKhvwoION9wZjA4i5kFtcq7FIhw05t851g7Q5dMsiQUokiuLPyHp9KGShWBVUL8
DOBC+3IUrngGwxQWAXLPnneEX+4xgbcdYJ0jQP49UTXjJVIEPRXJXv4FGXXun9PU6IA/5IHrfPmd
5zqXdYtCseKcFzGj3+zgXWoryUlr/Ij9dirUL6qB/zgq/hpSJJdJqogSvm7DfUA8M6DmIIKSTqGR
nH11VGHvrT1UR+HTtVr9sryGCYvhwS58Ns8AqaIByzMskZ//16fvWVbkMuwLRSrBK63zSRDpnyU3
FqT3UNSCau3HcrNDCgNLK8LIRN4OHEOsXwyl3VFrBrw0hAZu4TaUn6mjkcKz5LsaMW5Tware2UJE
g/29pR76zQknFKw8zrJAxAKfaMfsusb00RQD07NbHeZsZbiwFIpz9FU5nTkOFv6KOtkbO24SpUib
9UA9OOQAEepfGsg2zxsOwJ4V8nxABw9+s4RuDfb6ruwxBXiNz85MkvVEiOCEFGT7KG1LJmP4vphw
yixUdr6igGjvhaNEdKo90XeDKe/yJ+s8btlh8hfAZ36jNjfla9sMuHuc+fNSVylh/IVNICZRSO3A
U8/6zW28HMr0ELsKYhV9Ec78LIf1IRTHWRoucGh8ohDa6ul6U1KPddDJFfBlZkMRTCKMFW88DVcS
80CnTodimXaNn5ZlLfkYhZ6hOSlCSDjUfbstf+CroKXonFCmUXvzzku9UbPI8qFkHxGgtJJ5XtJa
JGiAQ7k8pyKhokRsqQP8jv5yGI6Hm2LXnByyE9R6MaXWoV7F7baVUPqIz4HWZjgLWTZHqhByefrI
NFN3G79JVSRx6EgEOf+b9xXTgfsvButo2B8jhc9SjpajBNpheFlduNhm+fLSxK5JUCg1dJh0Gjuz
ZEyqK6ODsAn9D0O+km6sBBnzZBjwU8pmCx5hXbRAK4vtwBkXMBhG8NoUZZUCCvaNblwByKBoDcX+
Qrj1HaPfdxu8H7aXRRCK9cNJHPYL6cXbdRBulH8CLMaTKGv0/qUFikcXyKvjuGTXaVL6U30mVbvk
1aX3IaZy5FT9zGMV63YtbzyUWRStcuZL66+tcNc8FLaUkTYf2WCgDk0QXRdf2SJarn4MVWYFnpk9
w7hslWUGfucG5iSffMiAQHW76IXVaC3TshLzU59D+NfxXOtSCHh34t5PufpMbyck5lV8THVU9rjj
uTNRXocKiVekZoxyUA8J3lUT5c+GWf1wYAmElaHq+cskc/74bF/QFOSPMZS9EpcSA5M0uPYiWQlg
mpf5IVHGQmXLvaoCNvFprdq+IKcj+fCHpyVzNvMGZFgbEn9FUkQUmQa8lVbb2Ss1kmodge9gQ7wl
QltAB/Kp44912Gl4x1jO704MMrchQ4Q6HDmKLtnBqHQfSyNSXH3zo0ExYtZIjxm4MXDdrMcJxSAJ
UdqJKlWjVgfSv7Vu2f799uM4RT0bR2rpOfGucX0Dn8UVctADmpvdOnJYaj2ZrVk8vyPPHrKuivyv
0d28vSccyRogwhwCF5FJjnSwcMJqlErroRGXuotBG5EhAK+n+cY5SA2U6Ho2aD4NuVUiBWrm4JB4
j1omYpDhRw1pEFtNHjVFSx86VLCkIkQp1zazHABY9bxWQIar1oOZ0xzt3Pqc+H72hxnZWA97QC2V
gZtP736ZIQLxr78mszRPaiX8H6RQt5wuMligMAikFsBHgME0KodbzdUiLAaAwct1c0btQalbcKZM
h8LLZj15QZtbYNqYiQ+c3lW30VWUcBkiqNf/WNA52c2Xx4BwejtLlvftRqvkgHA/NrVzxXC1PCQM
H7PvLo7GahjiQzjsxiQQLrDm0kIaSzhLJVDzjTmHGgxUVYqU9hYNCnzylMR1lsK5E6lBugsMI2+H
qt8v8Vbzs1PB3ZYvqbltvBSuTbrL5RmMt0VIZ+TcYq7F+SsS/H0cFzeN5cMCh88W3VvFVvufkyG6
1jKFtZYrltfuB/Bv+k7Hl0T9x8BbUgd3np4C/HaleR1vKiVWelbLIahXBme75QzYvEPrs/S7rYaa
ULOV8uBV2YM8cBtDyQAoWtUHmoAvBa2mKvNnikejMTijV5gelQ+zrH8pslRGNYQbTOvFoO/eXC0l
wf9v5DCOBdMA0r9UNPQHn2az7u4B+KHqnNdcn5PdMV215kdn/EA7ZNF5YwRia2kIOeawRoBuN7jF
QYskZV2ZBrg7qgFV+uauUJTYIFfvcS3cHowTlT+e6tDLh9jhjC2grHfHP6Lx3VG3U4O+qAuz5G/C
KfGEgNGV9B+1NP7YhpkGmz+zknCiAMjk9PeRHidLp8PjMotwAlW7y0RtyrklP/ayBRbQLwTkcsj7
uOzWPZTRL2ZBN8DSbq3tMa0MzeWhuC9TbEGi03bIMxzmNP01SQddC8mx3tEd0SAZTM9+fyDCSiSf
f1k6C1/I0wRfqc6+BtXH/t9IDt4FfDdLYVX0Xhd7991LBiYgWxhHAXk85JTT408Gp6PsAXKbpQgh
6J6BSvfCedrDyUjVwFnPQfHra9eNiq6+kL1d1iDwir/MUk+2Dy3wDswnYs56mPeV1k2MPP0mfJNn
2nWaumHG9TfY4CptK7I4F/lR2AdyqqxMYdHK8hsBf/bDuxAdWfw1/Zz7SsLplxeefp36K2PquMqb
ijXUicJuOf0U9qs6uOw5GL2eZVE1YkyT2gaumVdWFdZmyttt7+LncMyzD/213fG15t1/YAFQuLXy
7i6WmDEDf1+jDSKV5TSlRqwnTcBBc7p35S+Kw4rMArpaomYbxTQxnyDAgU93WSG8APJreaa/y8nP
Un5cFyw07ExB8YqzMQVGnWyoiOGg61+7YBIH/H7hS2q4O+i3IbuuhgBSw55hZ0hL38TSE6Od4QXu
w8KpxSslamOSotIMLFwPBWeQW7gJ1PXwzLY3LOxbKkUxlnmmjco7doGNH9/+Npa7iPhm1qQ/s8By
S8w0qYNIifPOFQHyk8avXkjO/xea1cwmT1L9NLWK5gB7KyQSfeBCeSDNesjH/MMRokjGkWsw4gnu
+Wu25kco1lc0nGCIFcYAkoKm6Im59uNoCa8GmeM5fcN3eNz3bQ/F3gf2H+UsHBqqtAhrPkoRMinH
V5ECo9TS54YgVYpu1y8h4cjaK/oLtGcUPF1DjEeb1ujZS0llX+jrHCvv7LCj/oxyogOW0/RiZcAT
eBEbqyI61MTFweXRY2kK7wVcLYtB3CReqbxyhoZTTjb2m7r+F0mP+FG+ND93Bexs9NY8aVjW9Nxo
8cThvQ449je6OF+I2NYkGdUTdR5rOCLRktv5vatiDshWJ0neuVIkeYdTeyg60bDOm79MKwZJn2bd
JYqgwPIl8YEpC/EKMZuOiUm5PJ9rc8cSHikTFLhMN9FgdToPTD6sTrOpfIG7RXA83hwEdgVy0qW9
eo0m24e3RiuUn9UwbdpHS+L94jV5vz+bgyB5IFsyLqS4oQv7dlnLsTCAeQczRb0AFFEoUtVMHS65
CEd+P8vCZBXVVQsOSJ9YAVoNKUKa5bG3q/niYa2GhYshIKkjEDE1kKsjo3z6n7qMfN3pfFk6XPO0
ZJiDw++WQQx9elDkgtvZLgjLy4WWhsvxYjMICqc7TSVVP+OzEpnl8Q0bNdAQXnS4T1+DStnbt5cu
4tHKwMaP8aJN2hDYBiJAml+LWIiZPnrdP0zWRVs/OppRi9x7ILhkK5kYb+fz6pwDQ/Lw+s1agFOr
j8/5ISOOYIZpvtQHiRbHzOadrbnezRvNHokvI9UTrHFSGq+7rF21UpCvsssUpv7SuZx8lQDFlItO
aFT4LQ91rPnL7byf5AVBvpeQNYWkV/dJr48klFYJvT67cO2M+tFld3U1Gg9+yo55ie2/xE/lcXdm
kxdG0WjCgTZsrMwUYFEKG2KuRjyi17517N0Ruc1AUgbhMi5tQpT8KT6+Fr97cqnOIYiHq+VQdnKf
7g+dACvvcjRsGPSnZ2JHaDGZ79andiSXYx6+w3wC1R7ahVPUrpqPFREaPBymmEl6U4pv2/IyEIRn
lqQxKgoj1VG+XNhi16HLL4wsPiKSyyHcUDYiwn7iQMYAH3Y8Caaa9A2bRCQPhIfq5aWV8ehT+DZY
o3rRNvOua0nMkdhBeifkH0ZUn5CHJ5YuyvBhAkM9tvvHhUNqGGuPa03tW1Of7bVktiQu3YE8GmdT
j5j8BV0P3bV37oJqZlrEFEtan673v6/zzfMPR17rawBkG807mE8ieIN4l1tEDLwOKLMHOcoq5JW1
dSsjEATirNWqGegpYagor1K7smnzNYhimydyDyfWjb31YK2G6xxTrovqulCGp7ZrgdxZOMyZ6KL8
J8DYpWC+6pwmhIUmLm/s160FOVK8f/VxcXN2LQXrZCHrCaQlspfBKFy51rxcCWbveR7EOgJ7eGVc
devDHCLlEdZwVp3yAgzNMo6VzRyXNEh76fK5fmKLQEWTp00sJWeVDGqHYwShnxvWaC4GFvIN/Klz
V/3G3HeB4bqIXYDxYEFPvl8MMP4G5exczZIKcNEfxG0e5CjLM0Kugzw683nriX9aIG7cxU3EQWYq
DWlcFAUnjC1R31PSjQcUpYuToEi/W/u0tU/KSFyBXPv7fYBz/xYcYptlBbe3ukon0XATj3WOSjlT
fz2QyarY4fpDjZZXHN8IzzTRPLLo91VENEJipcibxZbr+8yPjZvcTuc30VsPDfQcJ38cVwZc/5jr
vZ5aozgzSpXS2tSryYL/865nON9BPLU4P7/lPQpqha0w18N9fbRxDQoi3yzhtSkea3foMv5CMryJ
vOnpl3aQVWNuJOdzsPcOvTSDgNfwz+RrqRxKPtEgdmRoTrKz36Jb8Pn9dn0jTDvR/bFAKU3s7F/X
zxbbsy1EEoshR+A1CzsOysm7xvMEIF+xLQASpV8/et5RsdO4zQNgqCVOiKnLWmWworDRPOmeJZcC
YXZORux0L0UjGXMD7MQQVwgk9n9wM8vYvnPmZVk3Csw2edGClArgjosDZZt2GBBbr9mep862Z1jD
o5euh1biP1x0q8O1DF2/sLkYpxe60JEU1kj4j1hAaejB4WmlDtPWWb1P+I24TsQa5glFsqCSiBgl
LVIsBXmV0UdCKoUZ6QXvvUwrszeD2DtRioIsjGcJxS0U9zTjgHnBL6YhKr4HMplXG7vv2fMtMT1y
wnBipxpAVCajOjjw0qGsP8v6Khm8CfUU5hMugicfgu8EjzCqtkxvaVFNLwqZv4eF4henAZcPUM7j
IWGwch7jVodOr9g0sukWWHSx8x/zPB7t5fy4S5HsvpSKcqK0p6YDPxfNO8HG4/MexCYYD+Z/+sN5
miP6Fd75B7onQGgQYUUg4q/lWqcdK9SYErm229QIoh9SaCkjbQP6OyJxFQuShLMJnRXfmfgzqJdp
7dIMsUy64N7fbrth5g09LzTtbyXjBLp9hSaWcudqDgnSNO0a0e8SygUE1NPA9+1R8niB+3APFJLR
zaOAUp/Qgxg6WY4vxHByohw5gH+2KWuPiXP7L5wfyN94ZopQ3lJnMib6/rxCOtEQiLLueTc27oaH
WQXHFYUJxZSpyqh9cug8gR17m1uq75dJlj1UQp+LJqaTh0J1KXEmVDJX88HHgnY6U+NZCquod/t8
x5cgydCA09S3wM3nIGx6VaYn6JV2sw87N2e4YnOYxoHH8TudXQnmm3EkV6hoLmOjkwiKOKwrn7fy
D7hV/QOezaQ1SdwSfFnVmr1ZDFhST64TCZaiFvrCuFOmtWeRq6fZUb4qrVqjxMds4Lw+2RC9ipmX
6UpzDP614BbP8JmnHhyp/fL4q6LhxSX+H0FaCOgvL6jhvpEN2nkmv2aEnGTYPgQb88e1Dwqfgelp
z4hDCd+MUHorO6R4dey4XuiOWf4H1zM/f3rTtCfQH6C3mJKLhoJAF4PJR5qC6Nb24MmyzFIucnO4
jg0Uw/cpT1YtdCSjIiVJAojbMZPkVmeJcCSq/N1s8FI576Q68aBbWxIkttlEJ5xDQJB2SAAMuBAd
Lbr5oGk8jPCg8+w7zQoQE1fNw0OdXnJjm0XOTdl7iHm4j8v8Q+iLxmL59hl8EP4/4VLBhjVStcEN
Fj3YILRExQ0t0sOpAN6BIqEpXRLGcuInOjB4lgGB+ySo6M98hkjr4htPSQkh75gOlbpCVwPUHl/g
wVWja1FV8Th9CbSiMhbeArYXfJnkRPMMqlPnDawpxUI39jUIampBCIN0D81IEZs50kvHTsE2Miuk
2sGj7aEHo9f/ZidWYzvIww9iUQCYPmpOxO4pI3l3dpaixkf3Ds30hVY9kkGobHPSxJqAxXHlVslj
mGqmFi6526qNMy+q8mq7v0xLqugzdWhSLgg0KbXEGRgRK6uDyNWzvC3oe7+vbgvssSDXucp+5Hjq
tGd3kvhZ6wxQEn977IJ54kH8DsO4jMmMeZ71VTUfMBGKTbGuT9EY6dCKORhNEa2+mg7PRqN2EKrY
nonV1ubxJGCH1EN0O9/r9Ped9YMZUWLi+Tq+1spGeXZZcc3tw49WGmVnte1em8AZxRuQ9zO4Ua3j
zJ2KytExINLielNdFL8FiJmj37oQvjm6XIyeaa3z9Yz5OZ+DpSF03AqBB+irUDTeQr6OE2wE7zdK
UeUYC19qsYsmlMi0JVKWjmCA1wvPg8Yh21a11yRdDzFFayJ5Y1D/1m7LYNcJupKC4nfEolK18Fyh
6c7JOd/+oFzZb19kdBZr3cSGk2aIIePuND6b+kUR6F54xgIYGYUD8WGXpoksmHec4eQkP/U3PTeL
9uGHVz5ivmREEaFSmAaw3QcHbr90H+YdCzZPPmSq5qlLEcfFuX+2aYnNerYeP4+b//47253KlCOJ
iIliyvi2xtBBljnpqmsk3rkM6O9WxIwT2mzexoQ/tS87I/80Yb9j5blJjJlpEOhTxIRkYQXorMFz
5UzOatp1kr03sW8mehuZ414gRyCxTDeoNi8aMH8aw2twqC7Xn0Uxezz4tezZm3HqppER/3FG+1a+
CPu3N2ef/k/BbDS9NcIAL+iojXyoAkZv6xR1M6EZ53CpK2wg+d4Qa6drmPQxI7MD+FiuwVHMT77U
bpQw3r9fR6ePq4Xb4notHgflwFuNsgffSBTkRuVM31KbzoJ8jf7H8oyohjzoTp3A7q2DCM2RdxEP
IhmcQrJSkqYIlVSJcd2NKpOeoajR0XwR7AqThM9OJX6rYR2q52RXczg4Qg77CIsr8oJBGyUOfc/M
MVBanPj66trR4smbhSThQx6Uo0YliEC/4cXb6Oyg/xCaEvGtkQhw6ufGRP2HcYDTzEJstYU0obLU
QHC5zEsH72v0XmwtStT06qF18xfyk8bHZRJGgxPLRLWpj98wbsLB4tkdD1U73t82EUtF7dqzp1Cl
vo8pbU4v98fAA20snSbUISFsY/gJvngG7EWijRvXU9BrpXZd9Ex2/sfYhW/0QzLongyuM69Q/MiT
vINZ7AVxLONascKguVXuPF9t3+WUVbyehKQensFMh205F4DYxXe6CUebXBMce+ZJvA3iCLy8DvNG
jxZOJceSI95QfMh8S44863ydjkFmQR8QWpoX92ssD7GXkJjXBM2wm5zYKqtlYWoUTiTMsKqSL7ue
drenbywe6zkblVbqkV/7fvTq7g8Zt7x9q/05J9GuX9QBod+1N+LHKyRG19piMNtipUwFByRlu+UC
su7NFnvqD9jcxIt7UDKgJGVEdvRtUxuUvNCgxKEz8YPdl4jsex+pUxd1AjNZwNtHxF8Xm2GM9o4P
924SPj2ZntZFiQceC4AqtQP7nu8bX2aYdQJAX7v86ptd8mvLL0MBLyCMMev+tw1h+UtnqIRwgtIi
F+u8K4UJjZsv0jFAeoNa61+zNJJtv1jCCUIFYQBtdMf+Npo6CMD2lH+TWsSbkXNLIN7duZSCVMxe
tO7kqRwPcZxzL5MbdMqIT3tMHevbf4vAU2PMzit7vN4537Jdlpt8GV6rMIQrvvppYkAvb41j7U23
GvPLZEyLImcqO5yVlMV5A/usN4NowYHwcSL1qOYmTVVgysaq26ZJH8HaIZBxtdJwyFxdBu4YgrpW
9tJY5u367igf23dDAK0gNHvSA34UblicUcxQX9gL17BZxhwJbezP4PYQqqeSKqz9fnoCjUYbN+r9
CFeL3V1+HsWZ8VDaULcvgB94uPnTE7d6b9SV4Gh8Nr3/h3YSxd6OAVJOo0Wl9BHUpUTpKIIHMrLf
w8DwUyAwXJNYdR75yqcD9wnrU3FliXNEl9WGBx9AXzMJHX3V2ms0LjyjE82uQwhmtmLF4bVJVejq
nx/TKqdt1PriLOg0qNJX79ZO+u8i5JZTvP9x3awqKZc+apuoL4GrDIBXFG8qi15SVYWqGDCAdSo9
8uH/gLe8Dxs3PJGUBHm58wb1ore//W/8R8RTWxCnSlrg6eTKXnHyBkhlYrPUPDm1ND5GZi8LHjZD
fNYNQGXoDId2oSBzKXXZxp9xzL6jdcu554YMhjW6H2u0I5o2nM6PajvaFir3SUnkOqGE2XYJabZp
DkX2PM46lQ/yOboJwUUmaZ9mIBXAZhyirXkbg3+xuO0Gv8duRrliHTQwt8MtXepG4PnxKJYImGcH
JvKSTFI7efLXwDxOWhajtYhwLNZLbV7sLraquP+yiU2347xxcZLYw2Xcd58lNEye4flnWPHRLKD8
/GV6ubJm8cIQE/9E2h0NV5jZNmR4fpR83rWkEdXZTE6kJH8S8FkTm2BTXbSxPc1QbRZRQKfml891
z61Sww7QtYRhFfpp9L6/FZkODnGvY3sXVPTXpJjI9Fz7gto1YXS6OwhodhBR3qQDYoTc5lAmXkqu
ToMvvojz08ZxikfFtijo4wX0y96oyHDpfo3lzl5lAzmW8TSWmS8AcXwxrUmaKYq1+Ftfu1qGvRxN
OqxRpCRTtWxp2eLwqm99N90uUGWUfcfqH5aL2OWi4Ks/md7Jd6xk5a4bMzNHB8YaSL7uVF441NNZ
3lp5Ibd1y7Bj1UXwyO9K3EAVBagaLznwUBjGIlwZn/VGhdDR0judWN6vl43qO+7wWAyXkWXqBPZ7
yjnRlu9NDYBxgijgvM5F+bg/XJftAnXEqz8jRV9zpbora1RkXR331q9BagLhS217YpjCNqt/NPEx
6jl9KiXGgkZrmV3Ls5zCY9EjsOOl98sh0pdVLVA8yEng8EfhLoAqY/xY7jd4qaVCGrrLR00PE3wM
nXPRG802ML5G1Tc2+DfixpNbGqkGSEKqt86cR7+uizBtTKnvKewk5u3kgJrrCO0p5FfZN1YyMnHZ
NjGbDZ7RYR9Srd8L9jQ+uXysQ/hlTvB0SbQJPy7EzWpCBhcJA5lsxw1kSg/tjEGIt4nTLW/EP+y7
CiMGNGi1ZqW6ybCR6sJmucnuABkKoGOIGBc/JSIybZLXfg3wBHYc/NmL1Dnvb7cwEE4PtQxBxN1D
Tm+ZB/DBifX/EuUFvr204BAjnNpErysyl1n8hMJsbHcBgYXsDINcB6IYwWi2tgfAX5OE4tvkzWOM
msQ0PjONAA8BqJcO3x0ulynFb6kchVgTWwQ7mYFOSr/lCdWwmAPdlVEk5MaS/TZKkJtSQnu0YUHY
w0t/ly6sIY2gpQvHgPRSrUh02D1LFPHQpjR6vYnwolKh29JmSx+fvQ7Eq8pA116DEozBH8RSOlrm
5Ynl2TNXahkUT94hlh5T08GXVL1H+EH/CEv/cJJbQilKOHKh2fS8NehJRAWli1txniPyAvUTToW+
tgLtH28pPNJv9ouPBUnHHoOFPg5jj2sxwcZ0zqwVO+N14zD0N2Kd2TkUkxrJxMpjM9VxdoUnE7ZR
epYiMCHwGwgBu3dWbhHUQyhdyNRsAbZFKfiTP0RSZQKl7Kyy+eHeptCe3jlWQS7KyTFv7tjpyctF
+OBUFdXo3O1V/qseAOqLnCU9FdAL/Z5usifQT7v03yKa+gS9KqOoSz1mOfFI5ykvqIcWBnyMYCwi
Ovsx4rUHti5W3AO3ZdpMlwL/V0CP36Jcgu+6zrxO+9GSaVZGmFzgZeZ+r01NQXJGv6Ag3PxbRk5G
/40JM1jCCIPwbEKVxtI7XpGuIC6mhdA4jywmYmziRchxS9eX5VDA5O1woym8M1fY+zoB8wswHUtX
W13yeSftVyB5eK0ZpJjqEHIiLXoE1vkRUbxxI2+lkQb7v7CZI/hSxRl1Mni8rX7j3fkwMHqL9iAL
SIVgYXQ/lEAyXVtz/kQ4GI2DDKIX35e7we0QfH9R1Avo6eiGO1TM7byZKuX/p8gn+98olCQ6AKys
xL/TQ/duwIbTmx5wtgXYTcQPLpId6AIluBzac+MfME7CX4P3nanApt5/jFc1ffMWYD1ud+nYfYZX
2xjxEJNvFZA0iqYQKonDWokmDnwNQQcu0fXNdj+37gFgekG/7xi8shNiit0INveJAIq0Pc2DHxG8
p6N0g1HUibnUWae6BfI/IOlL0teNIGW1+BDXp7MrcRgHhs8jF1I6AtBHn+fRPeTEUxvoeli5hJ15
RKsey7rCRJc85VHS/HpmgEBxIJqLAPzn11vnby2P+uvctRmKU04tU1if8XmH7cZsDscjjXlReZc1
f7yUZFEdo6ONAqeeVDb1Py2UC6yq2Zc5yK0NKxoPUd2NbwRD2FzhPfOPqzfjhXV5GAAZKTACb2dp
wRa/d9nYP2GQpZ6+7ktfOB4iZ2zVxG06o2U8l9pcako7KSM/1VFdbFjukhtJXr5lZXJD+tDquBth
YOf5e+U1tomw+QEw1RP6gqnhR1u9VI+dja9WJkGB491ecpP3NmDFCGsq/JnW5eF2hLgBDNwOeQM9
oHQD3aEQZwUNpn/M5HySMgvSlZAMTs9Vt3Ewaqc97LoXJ6oaXhmjYeWwLC1Bjp1DCs1uu/Hprc8j
sEM+1/ePfeX8VgLc04HxG5QDsKxXPwfUVir5SG/qpIotsUcJCzl3andoR7rc9/g8jlgCqXorJuL1
IaC6Ja53Bt96cpS9a0LvQEjZ1VV3nQNMHMyqflvjGzMFpwhlg0Jv7EnD1ANY/Qzk0TlSL/iJj17M
7bWv0zyqZVc7disLl/XCVpsQAs/hVA0LhUmoJIU2IUKgQx5k1ijP4nzQuKC0ca1vf6EUHY14Ni/z
JNLooxEe2G8YpEfhf9rCUCNbwwv8AQJa6oSAen2WHMy09+va/KRxLzsAd7DdDv3+6WIWsowcGubg
32PxaBx7couUz+tvzDj1fjp48r8JYNWIf/oca4qZXwjbDHqFV9FgkvcfFy/0MA1eOVEJ+XURSmHc
akoz+gsuh0bxtpWUx7EDjrX4DqdUrjQtzMlOOQ0AWDryKlFHwWtEPFE9+7Ph3ZscxhaMY0A7v1sf
kX4ByZbnkoRzZx3tWLWEoWsXlqP7Y8pKrqsp+bnQEPxu8SQH7gKFKYxfv9zvz3Au5SDnGuE+yGVH
Z8rI5c6N/bf+PDpmgkgJtSy4HaM4YGil+Cz0aMenKQoUTXLjozU+1NXAQfOw14Kp98iNgpSmK52z
0Iajse9JBDZrSqLaGa37cS9sYEugxKdiP+SuYZkq54SmeYVknwR3QmKIau7Chb4i5CzsTPIfgZ9q
zS3btmwPIOAZmIJhZyQtVvbi5qu80+p3MLZGyfo56qKG2QCxZ+XYrFSraJ3DpE966wYRkEPyuRRS
0z+DiPmdNZPTdn4uEsjt4GKrAJlmrgx1ZBL+h9PaA1NI8wI8pozUoZQiA45poQ6HUD+2YKpADadX
0Bt7F/JK73r1cw4A5LUHyEUtvd9jCV2vdsysT1U3fTT1q8oPcz/+rs7eY74zKLNjiVOQ8mjJ4Pf6
d1l6rCAj5gx4rAbeW3fNoLFqbEVaPdzb1wwH/6T8w4FAmpoHxwaIGQQ1lxzJYlVzbXpzayWlm4W6
35m4oUm8jxqfobvs80T5BOS0U/rpycmW0lrPUDK+l+SmN4p2S7/g+7qqCx1oT43MIfohY7DVooeh
+gBK5YGHaX6kuhOmAVnq7IhLcZKeHjqnTlHF4Blw3igfGR0pJthfpsQpdIh3GI0l5HXogRxDEeIv
GAR9Juf/NKYvFjN4vxD/8mQiWGBbpLYQrvHPUrGupOB9jgp40Uuw3H42uDNa2xF23H7mBBJyhHj2
Sk8lTBmKSrOUpWg93NHvd7blHnxifl6Urpzh7ytwxTfWp7ViEzaTxO0cGOULA6+ZwhfPIwx/SBIg
GtzBMgn1moPXL9M2AwA6nl2aQDuZ7wUZnUaVOisRUOdYDX6RQ1ZdWsYDrMggDnNCTXWs95MYlm6S
y81ynXMkun5c79ETyesIyD04xOeK1Kf3k6Ik8wB68WDEaVLbJ6bZ/JHhO2Us3i2vzPucAVpuxEHk
IsyZlHyWkl0uyNze85gKWSSZAJANFH7acwJP8qGrzKI1jMZ40DXWQTgMZDM5wbjtkluw/eQut7xr
03d65ZeLu6rktPUgq/+ijE5BwpCrkmXjuAqvW+pe2ABcAsoIRXJL3FaoIMAGhYvZxZky2JhHBQJI
qX7cQP0xIHpECt6Y0FbaDcXKrBXo4qRwfuJFCAuvzUcCbJMB/mt4MBY3Ahvj8m2MJk8DWJcX9nV9
BC5Ykecub6mchkhuKnqJH4it3LHLy6FzAVbcLKg+1iB6vmPTo5z09yer52+NqsYeyafY87qLRZ7t
GIeuz9hQX0TkD8Oaej7zN7ZoxyLqGNXNke46Ew/4krior/5pqvvFigrA0+WL0K8+DuQgmLEQWVpH
r9eZjH3iMcSMA2YKTAsKSvRRL0wuEl8C8X3PnYCzuxvQluFNfFaDbp2nmJvWkhWEFTtPhGHc5ztG
+53iXz/Ng0fSA5lMzEN3JMFpU7olwJO+mj+6PjNJfi7za0ZVYralfYxkLPFGRQSIdnq9y5OgLip8
9SYEVbibrIQ9Bqn2ssbkEQS+86TcN8mEpGhnLkg8/yg7XFEukua290BWjRZhy3GM2VvcdHIJO774
dy90lpNkxhCrYxup+/CarIjxx+94iJ6tuMAH4B+1oaCO/RO+tsHtdLqTq0xG76+YYgCJ9zutvYUe
u2BTn32rVPebvHygv6F/l+MhWnIYdAGw95ZscFQKpCFwgGx0SUDC7Eqy0bA0GwGBi8q9yWiquiag
UZXeWpUGs76lGEeu2Me0zySOIufFcqQmEWTGyaUtCme3WvsjGAhoJz8w7bwZuMH8qUD3JPZeICf5
EhpFjTb+28l63OacTNBswcJWUKZEIQ8OA4LehVmvBJDN4sD6qUmmue7UyIzuAu7qGfHTmWIIq9+b
/xPJ/Q7eyUT4251wxZaqRu5bTG250Vhh609OjA+AuUZqXf5pMlnFMri48C055y/E6IsEFIaKM2Da
lYOy7/N3cTxrIhFSrNTvusnBOH5NAj4ZXzsRZqMDryosOtxzmz6IJjO98MrKLhrdcPLyUCGmRnh0
BY//227UEwORV8zDrvGeQ2JSNI+HmIM7tIDinABKDRLL5n0LYZerqEhjsUFJEOSL/qQ407jJJqqx
gwFn3QD8WwUaaJGa16RmEY8A4zaBrm8s/ETKMPA6OphoXjhV1DEnRmwOMVLl9lUz3WGevzxYHshB
1UgmOp4nTJzKiYRkX04Bn2g9SdpziWgQgXO8GFSsHNgdo/P6BBbxYvc+uF0eUTlEzw6svpu4lBI0
Px7rB5DqPBu7k4gygFyQHB75LtWgwEINouuIe4D0vzxKfpTyjel4bh1iT4TB2KDDyzDCWuAQ8AAW
RW7OEOZ0lWWnB2qYXJRNNHgb+da5A7AOSb1CWX2R/QrpU0mlYdXa9oVGT+NAU6ygxbKRVZkB3I1O
J5zi/5XbKpk8kESj5EzzVLswzZTJjfF36qj+FmMwUfn59OdjLGVnBbA6Y+J16PA++4FOuuVVbtKT
SGyQIG0GuxOzKFteNUi9y5dqrBrQlkQIKvvQKzUzdXfM+bJuIVHSww0dZv1vbe3vBYC5X5cElbtg
TbNmqyLZWlfvLUDB7416/hndyfV4eQl7B/AOz8flwmB3aC45eUDl/PHDmIXSYxD0+R9yr6n+2pWH
Naloylnqe4wmoCKH7BOWFmyjwzk3QbeVBoPUAY1ITS4I9ajqvis/88hHZ0rpLNBSQaGJUucrQC1p
ayTLaqujjqUOJylI+aVSSphtjXY17gsyS4zAW31sXSiIBqS//vUXVpBa8ctoj896/Y4Gdwy5ExS9
kVXBgADqlS0GcJyLagPxCECXb8u+X5Z+w/KO7l2i3+6+QU5H1NF4lXJQCO2kWXfdLlKq26cKG8mo
tvNST7MtgARU2GrAi04vl/1yyOasQANkcH3VGX/ubM1IwDTNbdDJ6htWysgG0wqeccDPpB/cdeUj
9Cvw1wsyREv/PQaW8dDrhjsgarLrGhH1HPBDV8aq9tC6FrlgETKkDI5aJPn1seCdwslpjigKfEtf
12TudmEO27JggakE1BEv/+9C9X1KLPgBOUV/808X32+sxXYC42IYkszUd2M6kFLEfm2AzlNTsUiB
O+7jJPeSlfVp/xYVnDwZSD2iHHL+Qa5PwFGclgGsugJzHSEwjHjOzbgxvT2KvURZCoQU2nw1GbwN
2yyNVv8VVXpBhpj7jdkr2OH9TEbPLfXNtjl2I+/hH+LaYyWsHUNS/UaMnDFhLTdZDwTn0bNutNUZ
SpKt9XHA9OGr0DOMRmbLvJt57peBqlCDZ3I2aJGdwKyv7EE8AroZRl6XpGSlySGKwzU5IesaGpyX
4sv3LpIwF8DcOcR/vyYGkr1IjYzmw+TixHPZhhP7s6AO46u2CUWEFfrpMDUCB3PGOssPOriJ0NKE
IFRyfdB8wrW2y9Fn9CNNUEjhm3K08CZKIzyVhov9BQpeMXlbu99Xoogw/m24vO8on1sD5Yhe+7Ht
ITDYYYWaEqtENLJgByYRLzOsysK/Kr6V0LUevXxIGlXpilkwUVWBCB+qvo7pAByvzvWyqFRnaAaq
5uWExDvdFLEX+kFD9WQGEj1AC5nr42Owpg5dnlGNdOLSMwve5CHIPlCWAWGThYAJYuW1JoeJYiO9
vXkDeJ1tuG79jO3SuWjVfSKNJrwtBcost1irXGK8kGoxmCcLVEXLh3BrpZkm5wp9Fc9SoAOH0rgI
8ciCjKfS5UPtgKtQtEyxMQMs/60jjYfY/B3yQ2q2U9Fmf9E6IrSAjUjVRQgOa0fsH+wbq/xQgA/C
bqvbxwnYIHOYVf/M8rQc60+ATWfMAXoPEy+fpmRKDV0Ub+Xq1GpbBTzem6Q5ZoYiP19SjSOfhaxp
pyxUbSMcl+QCMKFoA77pjnp7At4V+Oe+RDvG0zWB/Y2FnOrN7CEkzazyBb7zVkLEQ2gQ4o0C/KAA
EVl0Aibg4N9cMoQ3IUkD0W+xbNYTtRowRmB/uoSELDAqbValOH2LxA8JsyRNUeTgPTYF5s7lvme5
Of2xuE0fO32gzyGNJCKAIiHrQ5S+TAqPsw54DvRDQSBJTR0EMNyY8KvxbyHZWS3qdBghT5GBAuhi
e/NVUjI0S532UZal18nKn1jPJn9rPcIVNIUFMJyhcNfbIYa+FuXJ9+0Pgq2IgtcfM8Pmd4nVXLrI
jsRZ3aC4tev6LrRx4GpFJdL2JHyC+16+de2RsQr2BjfFYEdlxiAuj8r2DHazSgjCRN9Ve0zcxR/r
avSFHGfmpVLddbToadudsH2JsWgWX/5GBiDd4l2bIbJC9trEBs6I5ZRE6Xpwg2mQoCGu2C1HzAkQ
XH6vd8aotACob+udXOfGO8ryoFLZGH6QlrBCxVr4gySqQ4Pd8Z7HQ3WPZozomF6w9+flXFYsB3VS
4ZzdCGFrwpSnqNf0kV2X8zcRM1UbXL8SxuUDWBIX2i9OaKYIClCnb+MkPIRpC9eszx8dzHFozVHV
GhI1j8Km4OoDg2q/FeovhgbkcaSqdwutAH/irnjFkJ77BKzJ1k9VmRYyEbpI4zbs5F9W2UkAEmI5
IeSANX570A0fTra4hpeLkvwkiSRREa6AwOoZkOuvBDL8cHbOrHIjVXxMQ/1yiX8ifAERl3VZveiv
/glYzbMPwpfc0t8GSbLwzMWQ5xMndfnAlC+Oe0DmznOgUpfxQO0/2Y6qR2n0JpYm7CeZ2BFFLOj0
arA0HSerK4/qUfteKKog3lYYv8O3OCjz7MDL4njqXoq4Wcl1mtPhxVRm0OGHk8EFC5Jpoq32gugs
FeRchY4Lz6FB7BG+A0yG5jDfH0h9jgj6U1cVR0nBgKzzgyOCOnrsjpPpncHa3XdoNwWvv25fYfku
QZ4/0KgF2BMVNXQmW2qJVt8as44Zv3lDA79Hzx0A8tEjxynbLxuO5y3bju/DvNRiIOKwfX07E+VJ
1s7oyIj//IdNu4cLvmJ5TuZSXMjfxPhkDHP3gr2kNDTWuaufDTJyWYFnWSjUny7+dOKfMiZoZ9lC
KQOXKCp4QptvoriuCyD6c2hfPP25ZgLu91v2ojotZjnUoHxSjtTRnhwtHjiydVYbMI6uurDp5YbX
ukidf9XFZYN3RiKiECRvO8ZKRsL047jy7KjJUQO/k4qazK/h3Dxjn1dnIectAtnKkDmDIB0YaL9/
9yU6NEP5DWEUEn91/DqRX2Y9/lfnRjrsBDUcCXNui5xSGziP3WHFCLCOq5vRMRRF3tptdW0dmLQ4
bI4yweCWZZXddjqTuope5uP9DKhhoKYNKrsLIhrkNmE8eP5Xe/LsmAt2aE4VKckwEKCCWmKDeWjx
t7q6lwN94ZU0v/rWaIajg7VKd4rJlsVR6F1/pd4UWwGVg0qnwzsUkbWOk1zZyn5Rg2MwyRgtPWBD
LXWdNH1QsOAopSpMwC5PebZBv7SSX7wDmGzkc1zOcggTsX2784TWEvXVmXBGvgary/cMrwi/lTW0
jGHfTKAj333S0NhNQmemqhtq99wlJtOiVPl+05HR61Vosf3xGTaWteXu0YwdcDec4e6rJ0BLex5v
rrfP68Ky6RiEJRk4dxKajaau1d4F+mUEgCSgeEtLDLHt40oeVggA/ND+YNmlGURyBSeVw7OzT4eC
U71A9iYg6bmpeUedwoFVq1Ar/eqrUJy7ZTQajVqNWchciLzGFz26k31nqhzc6k8wxwEO2ecAGR7Q
dt3X+ZP4p8aMoYuFActPa3oLBxsAiY0+RGDSAlhRIfIglZfkdF/tr9/G/j2gNUNXjKe3/6AynM3L
JlQ7hMyy/iE+tNa7DAaL98fCkVdCuLVknBFdXIVEBwTIPgtda5b/phqdhABDE9juViK4wCaT1pN9
90PWNeHTRUc4B2Sl/UlNwxNewIbM1CBwasbNStoTAxSlNNziAZzEecVZB6RiBFbbJhnlGRcX3USm
0QxFPM6/5+Oz/p7e+q+KAsFP33earn4rMNKe2/3e6OUOYk7c1SL/vDY3X7wz+T7lV1NTxhNNqi+N
ATyIXfd6Pbse9tnQ1PMQ2YguDv4ePd1rtunJWyoCYVslp5QzNUN8tAjuQeu8oxuHQQCia85xpJee
NFfwh85+gFuDCPS76uWKr1a3AEzVs2MhFW2+opq5WSEUsf0sTOgBeYB7goxH6ea0r2CXcyjXf51m
TiaUBjkz3+RVBT+wY+IIlLB0N8tyi25OIONe9oZdx3PmqPOSgKNeUviGc2J3PlJCGbiBbV9RWuo5
DXGBXeXZzeNi0MPmoviEBQgQfZqVR/kKjudJKsd4r1jbTA==
`protect end_protected


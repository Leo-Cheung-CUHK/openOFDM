

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
p7OtZBpltt/h9CD5IsJBmAQ+bQJxazkQVbRBjNJ7LWO+cgudo/XA7alKhPL+qAE8nYmt8n/nhFV7
1FHJnU9EmQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o0V8lbvMs2u7Pr48iEK+soyjigqgrrzx5HsGK4k7Ph8gI81XWNRtIljFPpaeGwucYu/H+gPVGgh4
LxNZUBJhgeC8kZr5P0UJ497gR4WHGLQSo0hvtVYHYDlrxnVk2S/+il/2gMAwvI5YF/lKiRUCJMb0
2mL6cpx+2git922rE9I=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hIqrLT0Q92Qul/GeORaSvJHHAIqLk6EmPwtSD3Sw8K7TFMN/pzvjFhA6g78oxGwtYju17YRUOAPP
BxWjMZac0YPGSx1A1AySaj/jWf8/sND51mJS4hxixMPKgd+iJln4gROFDpToYNAZ0eBhqGsKoRPf
Exo4YtwLGOksTW6jkb5XyScrMy9eg1uc2W3HXgQfQg9hr9gpWWe4xqhKUCFXFb9eiIDe3eaUQ22t
Qgz9S0YooH+uhgkKhXgOsKoG8s8RO9q+oyyLd0ANkoAdDySOy1H2+qKDhuJHoo8oHgkWp+t8x1nO
sbVK5ZibMfLbKeRbGwFkFsj+EKfWfOy4ck2AmA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
O+omGGx7WVLIBeJijOGvFCJZ1IO2vxCm1x3fAW3H6+gw883MkRTmRZO0ddVzk3pvzQaBPeJUDRsY
1XbF7OM1C/khYSkVv9TjyhihrgNNT2rgkTkWtfQNoOMnsmtYkK2fHBBMyNXzHPZRBh+2VgTZHxjv
olfJ+wvlLAdf8BqZKWo1gutmRCut9sBqwVpKtMbEKFGRBnt2pETIJcWkewW45hEmUxoPlXpgWrRg
sESpeoKuutTTWJor2paEV2RoktNIWs/+x82raY47L1AIZ3uy3vEVemolA7/fyBhQXHdXuWEXntN5
bzesBXIrWmoZpCMSf+IISz8dywoKgC/dpdCKGQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pc9IPtPXrLLm2VmqSrmdhsB2/sqloTepqxhS9rXzXINDRuCWOADiBYd/5aw6fJ/PtHP6hvfQmgPM
pe5Rbb9vXhfZlTdZe6IYAV6ajOneMnpE0SRKlyLpgkbpQbwWF8Ta9x699vjybNfWF62AYBS3D7DQ
b0t7dD7uNK3C2oBkpBFbB3y/rTrUlQxN4AZtlp8BUDmTdKIOwvLfH64R9omltAgRoa9eT5fKR+NB
hJulrR0XnMdnz4MTDv9F/TNStcRrNIf5MM0b3o9Lm2heOPvkpoBOr22fj5c2jTQHuYFT3gyiU8GP
rFykj34Hi9/EcnhfJs9E3mtp1Tszf4e89AyXHw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Rp2qWT1ngiwszVInFfAgNDsqirvFBRH0fhGMVLdTcJjuZF6cagj0r5deSp/lHSGQXbQ6hn2NE/pT
sVS4xwCY2B03TkdpZqI4G+dZXB8686b5iwRUQ7S4WwcHb3WXRb4Df1OHJ6dgH8h0dIOxvwXXNlqh
PKzd3cQ77q4ZzFc8bvI=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JmHrUUSZT8PLNYfmwBtqUH6qJ1p97BdaA2q40RVMw79ZG2/5JMAd6P3xNNzdIISzZU+jzu0NYPxL
Z/zfPbolJrCwAck6UGljZ/OOpPHLUDGkBAu8BIP536kFNfmsl2/w8PHTByudSnwDI/YKiNqfsxGP
M6Sq3+TkXml3dJEoLhHWDNi1mL1f4wADZ5vEh09j4ryxXNWZ0T1vCwLDq6JQfC0fF5S+fWguWeoy
y4GDwuB3WNo6v4nkxnIBm5jk34GhklMVorbQQ90znGRfAejdTRlBiH1jH/CASbqnXiNzj4+1wJ6K
83Kv1+Hi6TU2vQtu3O5wYTXjTMpJrASuG6iNvA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
SgTZSMlAkWPOykrjOiKAR9fECqWB0LS0Zq0qDF61+KDzjiMnBdEKU89hBrLr3tHtHhArBsJBrZGB
IcV8UMuapF9SCyeBwJLWrb49f8kQlXTlWEiO/FDXW+Onxvxj1KjOCqs/plm5KfGAfvbZnw6UIFYu
ICgWhZ5ZCTRi8xDn146NzCijlWfNHQ3qhdrdx1DTq7goj3jYEcsMDhrGtvD2MeeWppI9W4yoY0UP
P1BVcjRktKRQu2W5Aodo4cE69FtmW25sBw27VQI3tV46eXz0r/lCVroDOLtv0ydGFpvzFGCL1k/w
HXuHnHEcQLiM4eGFx0ND+qLVdiEunTl+v9CHNWDsd0SrrVp0LeUZ0DYo4k0kvcVlHU4BRIEpbKjM
+z+Ado4hnM/JCiYpjlruLDW1tfDKxxDrDSVrCL9DNTrQjdR/7ft3hn7J+wC34FZZk5gV2ixW3VV5
HFp/Ng6bbxdDTm/Kokez2mu90WY87szwcBI3qrpOF+W0I4uBcQW6ny7zNGOtgEJ++2DYVIzMiwAw
ospI6bFotJSRpi8VC1MlPhnY6aH6pwzastJhvbirRMtd8HkeIB7rxtN6j+pTxSUE2IjrmgjmOP8u
2zmfJBkW0SxpPr53KrW0ICgOj6xz+yc1t6dNotp/TZX/zUd4APC2Y4aOA6TmpcebyTMgIbw6Esnz
HFL14WrRksaUF31inFfAq2oTnwxH/sSXTeIZRg3i0BMoMo5V+u07cXOhr+8OrSzHiUN/jEHtvgfb
dvPCbMMKWk3pni7RvkkfRtIFENBqDHg4WpDqPsxOWEdXr9rutfd75GRZ2qGwHUqPszV9pPCoRrVO
A4/t/HzyoHmgESSUgaoxLdnrM5XGrzN9bPY2N3Lr1RFDoJhF0x0j6ArQKHWS6H0n4+oC4Vq9gxuE
FGIv3+lY7X0dV9+IuTyQnabyLFTbQnw2Dnu7q2cqeR70+Z/kY7YEmeNWurxXO5hyJ4B+OerLg8tS
xyG2MpY80b0rFh0a7o9GZs6lqo3dY0/aPg2NVysIdNofFKAy+BybWbklMM6EY2JEckJJT3fYy4jl
Cl3+Y1SWAf5gSWGLrRwSk+cJG75YEEuJvcpBNsMgl/mTIcxkWtobGiySix8zKuECIKOaxR+v5BxG
5fhgHubz7vegXsAEudrhTK12Sh5RP0TIFAiTyXzxJu67zvBOPNPOXHD+genpzW3IAj5FwYRysgdi
wEb0xNbvkijFnJ976GpCciANNPZRHn6LHH/RtUbO3NE0w/H+c7mb4sOwe4sMI9rweRb44jGy50Ya
I0A/mTLHayJO/p/MZn0KzYL0WS9mCq9DIIthweCeTwig76WkZVa3Z6IrugcWCx1Cz+/RoVs7rlxd
wTRjnFq4eA9qTgwgX67Xdc6FDPyLx2LOK+cWeJ47JM3UJH+XTBKhllm4isqQ1OVFqHYw0931Myzy
isxZTQxqSgMHdr3J1fq0YXtDm6JJ0SvPwdGhVMjeIl4xqImqiiKYLX52QuhUgccobcxhSeErdB/C
tYLhXlxobIoqmvM6yDHlHaqlAU7/UfZwbsi/J0r1MSW1Lj6Pxcpo9xGIku0PYVWYD50k+5dgDNN1
pckiMEzlqDqEJ6ns6DOPwOT1zdw7QcoZt/xRRe+kIWl4fUzz6S8J5R6m8g6zQhdSh7WKRj7+135a
ZMdsJy1ZQXjT0hFfyvKGblRAZ7Gzs58t9HRdnafIuZNDxSaEoJPHUkqf+fwVbin0c1/CjhTPCTwH
gU6Q/1qp1s5YNnOvB4slInnflKgFL+X76Awt6b9Imkm2bYY0q9Ei5ihv2QJrIClgOoKjfQsPTruS
qulZ+0LUlcMtmBmPLdQjMNNLckCtU/zwgaA6Ejevi95M3g7QCtfoVYWx4JQWFpoNwoY0Uf+DhS+2
7XABes912lhdgCFiOwunRIuubJZklaJQCPLY74212Wai8JnOPXeVY2r+pDtnN9jemeurHw7M+Cmd
VdeEEaSleatD4waiVw06Ft6CW/nDcYKYA2kV4v2BDXFI9Oq42athFtAxl6sdVuR440Svpqua2gY3
ZpNBqYWO17AhTXlqzZFGnmZ6T+ZTuE3llleyXessc204hpOQ7gH+gZ+hecfIST0sptg/sVBuSR26
dTyNj/XgFACsFyk9DMDHaWkubIESWw9sc40EPYWe2Y08DN8xfztmCoSUHIvyjwcwZoEdYWTFWlCo
9JXYMaG7JzvTQLo0+Gm83cocSQ8V8yVwV9H7QuUpPkpnsABdcN+ooWL2qtWk2cYEOqR1P3I0IeJ3
ZYTmHFDXvZodFcJ//N8pyHy2gt5yKU2K+IrpIKelvxLcs5k/LquTYBTlzThmqCFBvnVnJQnoRG9S
gHKvUf8JQi5LkK0wMS+G0pYjd/Y/ri+6ocUTojZzPvB3dtwpL/ct10Xz1zAJUjT1tf6zuuAdbAPo
nDlK0AyWsHlsnEGVbhXOj8Qcpg5T1mOjPmiwYQ90Sq+Ux51qLd8wuyfPiTA7+X5c+d49oLIuNwCm
gSNp/98JTlCftDUV7Oci/NsFVuwttft9xwlCt5M6Dn692Tv7XMJYFSz6KFns7aS+P5fphqdWaUi2
c3aW5hKsPcxiQd6nt2yO2HP6OIBOCZqt/ndug+GWMKLWgbnqmcR0j/9scI11yaJCZ4R3o0MLWBN9
Tw5pyYbIRTlYHXDr76R25MTU8vT+I/UfnFdJ1oLlM6ARrSBgxjvM+XTxCgUjXujJ3Jk4U7zEh4CD
6VjgI8OvFe+XaZLoQPAEUdKT9iBrxjiz6eV+XXLEYmp0HU2sI0LncqU0VkH46/vVfEgFIb8/IbfV
EajUsXuy6Y7hS0peViauCo8Bofanz6CDSJcN7RvLJkfjEm8zvzRemYFzKATajz3XmEw4KSf0xBp6
1h7TsULjArElwF5OL1fL+p0SGwr9Py2VHGd3g0rYhiEKFBXcjLd/bBM/hgIphY145E+6USAX/I2Z
VIIowvjN7FBWPdz42efqDMIPBXfeCV0HMMyaUHn5XHSwX9cJqoyCw8dho6ahf0i6ayvPWRVFqK7l
LsBQKloA171py48wyGjD0ruYd2c7nLuN6RBVxgZ/7c3RE252E5mxBKDzjNwaFElqjTLapmWoGTcX
TDluOgnHgevNV3ebZY8X3Vkazki0tpC/G1Aj+l4pVEEaFvCcDih5W0I9LJfKwzDi4mMLNjTi9kPf
ANLz99ldcJP7FROwjuRxjG7xKOPYcFPe8zryZ47bDjBJ9n642aEYbixPliOyYCrcWg6MHaD9IZSK
mFhBPnNZCwdqVRiA+1LjgCUUldYqgl+qufkP50NbG4BYCnShgDHAudF7GCD4NUKuIvsluGhxupWK
TGPMmzOvNQhVfBUu3XP1QofqsYXl5iPT5cfxxOpvhNMY4ZgU/j9a/6dqVhQLpJT9285vOB0J/HFY
wBBcwuc+60XZ/J1mgQVblQkAtr0+xR1/aLjWGEryAu+1eSFRYZgWDDqtWiIcdlyuIXioDZI7pzrh
NLvs+llZuGDZMW2/G/vmkLEcI+tKCpuMC04+vrZUo/9e4gKMccG3eCTuflvNxWIkiWnMnrZe+PZ/
rvrI/ysw4vemi+bDi8tft/1pFIi8YKPRjmS8GUIWl2gh73R0dHu6w4BVIjsq3DsdnvO1GXe+igu+
blpwVot7fEvJ0aydPFl1+eNckRPXiq1DrJdpDgizLR2Ld1Tarw7HxpohGS04NnzLSyGaIVl5O4L4
74orJLM/VtKqFm3xwfNvn6iBcmy7GP2Vs2sei1QXCTYPd0Aga1SeOtofCUtlABEW+QEpwCRgegeP
GNZJJ8zDt3QaYrvODRdNRSZDuk3/FeWznDiZ15Yq+1kw7vkNssI53APZlI12JdLhfPZ+EB7R7cC4
Fpy+SLuYReA9oX2WdSN7CQOGlZ5vqO5LZ7OTFAvgo9sMHpM/QZY3uiNO1k+Zp4kCmuCYo4m6gtlG
3PUDKmJKhESksvO0+HohdydFkg3bD/H0T7bNLMJ9nABe4VR6t+DGB4xgh8kn1Ntm2rw/Zs1zNVJ3
SZGFBjMJBDzpP8pnvoJhs5LiOj2hqB92UXbhqLnDRgAu25V50gLtQezZ/hvsnuefjW6LpsN9TC25
r4qF1+4QDjTdnDUv5B5/PytGV/zuY/zWaoEy/WyNCb6zKIXC0KCogkLq9eE0nmP698mfXmTD5O7d
oOKt5yWyXmMM2CqwI5nZY0eIgtaVSaPVm994s9DWXXe/JQHTFx3bKIthS1Nh4xFT3N/n6dOdSOQj
hSdULsYxNrN72wmwu+yWuEHKpnkKgXIMSdu+3+9OOzzYrBbAyC2OpnmAW8a/WtTyPSmsEJIHe5dE
Ruk/6qwWHUMSgfJRaXGYhhZg9hHh3jIpYoqrLjQeBbzYFDdd0FnlY07xLrA7PflawgtfeknQLTAF
yz5ri67v0IQ396Hrc4EKHEhJN2hp0ln4T+V2b45A6X2vh/FKVLK8+rICoimFFa345vm72x7auq3e
djqmSMs3hcVTqKC5Rnq1DPLHim/Ph48kgHi97F+/y7YejqiYf0sj1uAn1qfQ2mjhs4qOnq8gqNgi
df8yI6yuVf6G/JA8k25XCd8kp1blxsCU1mesXkTheN3bbyKhqk7BFFdRs6aY+vHt+iRU5emSDozz
C4dcZUaETnD3bW0BSJCylPp7tli0EmB0r9lNGjTQLTPY3AQWm11zSYWMqZQg9YNZVrwqvdpP1+hd
bPmwHOZTQk1LuXh5eS0ttQHhAB9Xn3We5efydyPGTmNg86kRp4NtZ4gmHHYgmNCmFNL9+bPG25pH
48DfDygenNFtigLAmDAJHb8XnSvDnOKUjZyWJjTSQW1w+NIo8QINTbclL8wLOnIS3uTXsplPt3IV
hv27pUpLg3oJHs1KfbPZR6jfOxQi2HFUlLALxZj7mN+49Idc+igK9/xyofZMo/51g67GbCN2lzRQ
iq7qA2EYtcx4FQli/FzLpoxa/SqK6+FwN9iVm8dX9hFqvqxntTNyyi0V8jB3qAl6Ljw/4JUU3EBq
btezrseOS+R89iey7O/uSAelDCZYpOWqsoHpIdMTdGeiGyWbc5DwgyrUYfjwQUNT7JVynTZA7ZCx
5UdHufd7xtspJa56wim9GYXVJ5vgSnQN3xj8v8NgjdJSudPrH7ZJmLACUzrq00fTYetEwiOgRM3k
nURpWA+YgRErynkPyesvTISJivCDeu8yHwxi5LIKFKTytKjgmOZS7mQZuse50QL5hOtUOPo4039B
FP6WZ33seowBys2hGf6vz2aCovSg7zt8rSaqVioTBFygekE6NogtdcIXHijInlC6waRqbVVBvDz2
HJ8T7C6UeDxEp+ZWPqHJxniIiUuee6cS8Dzxwl6FQIWPQbaJZqM/DmjlGO2fZ7UWSDhfcJCxSnQH
EA6zytAJUcwsmHBKZ+lXhNdk8JodIdEoZkCPRmJAT726eWOY/yUKBw1msX35zZq0JaTz5YNaPxA4
ztBW7xSKZVbaw3bo4Et1Vgwaz60izxW4EDQ/ClziP7e79uZHFFmyo7VTi+pueMv8O6UeMNo/dafQ
KxoA8d4t9nuuc2vp1GY3IRDmSLidA0DEmmCRlBPpgRROhY2XtFDPDr4L4gj8Pl30F6eTo27bpznR
EyD3qAYkrmjEa5R4ioPwArpo7pudJzJVLIPgIppAOVFgZhFfXp62uoNq21/6Kc5orWBGniSHUBS+
FhRykdznuQOmJKhGPrQMQjGXZqeP65F0ozzCMiAfQ7EnYdL4vwareRUy10nEaiqh+Y4x+aoVYfd8
LLuTpUa/5DePk7/Wr19/sg9wgajuzfBHiKqetOhFfTuDs+OFzsFtdJsGtR2FBtA7YynuRE04IbBk
tGaPFTRCG2tYMGsI4OfdIN5mxwD4/QCIPd2huteVzdzHcXs9z+mIK0ivAvsIFUaybafItNusproQ
sZxMfn5/RE6uTQkpNBvdaRol7HWKgA89UJ6So+KMQ9ZaUTRopI1bV3u+jiqMgOA6JfNiiGYxKdOm
ll6I/xNNQDKNLsCRgJg7CU28SYIcp8VPPA79WkOhA/MvrepQhnOS3MULs1CO2ejiT4OFoaMK1bz/
fLNxiMJbOLZwLSoeF8k82TEwYFnK9dtuA9dhgnpsDS8JgSQ8eo4O+ka+nuMCt2h0W842uqP/418c
F9q17StTorC7nIfx4dqlNMJk81gW0nfuHbce4Mq7p7CIVmJLzsbuNDY167kHqafhGtnHnjpW5dw5
ZSdErT7DpFm/fVKUnOp8SRTotlEkTPyT3pPY872B5GzR3PhXGwzkQmarytl4rduZK6pN+FNl7Ags
ErVOOj1qmOHnrXxPJNZtQfVSsgT6j/1l91aXy2KPN0wICk97l+Mm8CwZ/jWf2m3zufoF/FOm7/tE
WxKEfi435JIVKijDt3r/ITYsaDINcBFi+IjOsG6epN6c01yMm5ZmjhKl6IX/g9lQwRdGDLO0KCl9
xFF3SM+AuWvRe+msYoKY8UROdOhDlmkWgWiozQG0LgD6P0FDYBqv7FrwJJ1SEfJqFxK9pQ0fuTHY
rohrP2+8y5r3JT4yjRvV2RlpayZP434LQojJzC9sD1n4D2GIYrkBXAKnSmdxyQ8CNoRN5jR8ema/
22P8azUGpclMB538g2v9Q9QU2Tg5G1lkg3x5SZat/SetXPlUe2KKkyqc7NPcxORGbC1r6vdoCuCE
9I4AkQ1/zJtGSvOoTW1o+bwtEqwoXhASY6WRTKiNVUB2sB+yfAP3m3/SDa8pG86YADX7qyHlvsZ2
qYoCZCEpyZ1fCY650StKmvxOW9dFzZPgZ6HqYJ5wEoH/mhW95WJvlXJuf3BVZaJX/P3dtpHDL+Ew
gYAKXLj1+zYCVKUR2H8unQsLkfVZKAI9d72GBXWSAgCJ544FNHcAAGPTlFwNr2AgO+ze9CQszQFu
vTj03wKQyyqnWb8e/sW8wgsjXGWr899gksv4pnByRTgXYe5CWb+zrPjwd1z/ls0IDBqWxi4SA5SI
QOvMdNzIlfgek7MKJ5kgZkI7zigaxEsKRNYHuT3Jm9LT6yg5jZi4Ceiu3Ic3xjTqbQ3kRRB+XaX6
0pwMX3eqRIURA0kWwBGHEdhzwz08rS4gklPsyaL6848xAKDqBkNjO80nNsdwOE+3iTvQvbQOtnJ8
n5AXlC4yNMS8VK3EvgQ7MCz2fQ2sPeqCjOK1aw0+VhNd5OmqED8bgRSYu8830Z2a7IIE0mC7CGs5
t4z9jpvrCEZ5sDn1KHOGgOzMJax/KoYOUczFX4b5ae9utZuhMBsv3VOUUxUajqrh3ZN88KzNC8t3
Xi/w9an6j8A5u6L5xvni73XQDONp8jJZjCANTEeR2GvCfttFUcfViX6hI7GC1jHJgzEKwZXcbq7+
HdI/5gZOetQDB16aJbfpeIHBmuc1SfiTrNKj2SI8wrpgvSZxYsl2ittE7mv7oYZPLWehIFmFlnOa
e+Zi2plo+ScdJ12BCGcx6l6HnREc2npk0g3VQEPzcc1pGCDQE1Au3aeLaxdrVeto3YjHXg3J93+C
DJMNfs3Ihr/uB0z0q6De2XIgFrlNRnxUNVamF4Vv8yzqPeseiGD5WWQ1SabVx+L1PeOeMOo13nSP
FvjJjSpAydv0uiS9xHD7ChEMd5CD+q9m5Fr2caYcD9RjjDgIW0bOINcNAQFZh51c46oOLVhQ57DM
aNjIVwW/aUw3qBNqYFah0wDtQPTsOOXGHD5PKB1bpJPZrLI6d8Aiqn3d+VUtFcm+PtDIy+F3/dh8
zrNtk/bcCbdpOS+/4IkFazIz9FRt9ohLDkpT0+VIipLwdUMYd1phfWk1XcGgxjUdpDe2jfdVPNeb
hpdWKXPDTgqT2naKqztOqecIEj1I9v6gFsvKP1w4xfiJx0QzF+ABTVbwuBZGwqaPLt6Ew/PDr96t
l8RxhmUMSk9gyr3ctjQEBgqP9KjjHI6c3WSLPqdCLNEMmqCil7/CchPm1GRqNuNJtJm8vN+RVCPX
f52WvVB7CBmVNuW6x1iAQQdSke4DQPtvFOaQUDKoVXmANIH4cVlK1x9wWCP4eCGSuHpoeX5tNONo
ucpgbpRfCyya9WW+b9cij8EGvrg+CKQABaHfALa27hPr94BUiwBlO1dUn29P5WWEZyNRh2COQOk7
Go663QkTSLNgsxSJbvylBqkgex54Ut9tCUo5YaFaPzCCJtQs+EJ8ZBBkKM+CtWxrS7IVpSnMxo3U
ya7Jkw9z4MSucJyqdW5agDgkU/V9HZn5bx3D8Znj3Ys2eAfGFFmqyaPP6pF+FvLedJuZLxl6rAS8
N7WhwTFBZzuk83Gvqxi1ZwsN5+CCoIrzwOe0CAbduAHWYprkDRPwI7OvolctY9ffafUoDydndHzG
2ZwNFhRynyKJCd6p3ob1uB+Y1DJUp3dtCEMCVEVg6m6F0eivutYw4MP7WldzWIT7PNgWZXzbWV16
qxMh1Ypr4+2olDxjlK1KEnqvYpvnwvcbE4DmzbN1efeSEHsbmMNWoy5IgrhDodfgRZ1Ub5sAvZb/
fMtejj5dqbFjjq4MieK0kNwEwyDWOndBYOxSRXzp73hbqpcjzBuIvxw4PSaJHzrDVfMzPnZaLBXA
N3iSK8iJE+/BBPzMUQ70b/ojvScjxli7X0FLoJ7/OGIU24Uk8N9sN4a4VgEjFO5KgC0pEAWB1FFo
44rq0Cc/VQr/3/NNXIIX1fLzx+rS+QvNqyaVL9GjgivZ4GUEoyPgyXMeK5svzKjJ8RrttazCHZ2K
Ai1Q51YA+HY1ewnAQ+Btlx+oNNOtQPShS7mwpx3VePAsuB5PkB4NAbksY1WjLmT1tF5pRC2vJkIu
JLkn2yFgsXiiTg+gjNO6iViFnnwJ/zxvkOo/omjKBrt2oR9eU5v98HRWZE5XbclOMgY55OyocgzN
B7FQU1IoxRp9v71KkWZ4d3eGh5kcN8WfPltlLWHej3LoNGEJdEhCQ8P926fHTs2ZJeistB3as+l7
XMPX2uQVyCYc+pPm64SPI0iv8iV0cfw9w6wLXYDATGKsgNVqtNh5CmEnv2M5BqO3JRFhNG7tLOLz
taGFAx+jJ4dm11OWBd/6z81HwhGHBTAuqF0p7VU8YkKE64ZkEO3I+YlLl4Z2+tarZyrYBHg5MMwz
ARoBaSXI+OkyGHgWQbyb9teDcGyiNEVL5eBeAxdPIZfvOmCsgAVd52HdAqzPLwt0bj4S1lz7Vuc/
frPzbCrQ1Cfu6Kv7il3/VHU4hcDV+nrI3LP4xjRcmwQatVkIeU3vbQPp9NxXBeGgW0tLmH9kK92W
9M5tyHNpaW+Eqtrei4k7x6BecG8nEPU31QS2aGZ/tFRhSlyZc2JJ5o7Z2F1bON/aEbnsXl1Tdadb
BDWg0uqeHRI5wVyLE0I8ryO3RM7M6pVSlI2ll/WWEC9wvX7TIeecx6nzZL/lN+weGb/91NQB5Kzr
8BTnn3o74EA6IXkHKEnCC8KSqLGtcNNLOuMswTKhgU+bwbZlXXdG+iPkBsl2Jdx4jPn2Xjd9I6JL
JGOOdoc9dL6XDjh349r7pucCxRGMmMeK6FTdK32Ah6vFCohp9uG84nmgyTxARtOnc1WJDHpjCMJo
U1xLpRnpHkzeKGvFQHh0iiVjvL/YLTxHdmDtLfVal2EHsKST9CVlEGI5GZX7NxSz7QCzoc9ACBt2
axsEbByeI/Yh9e/SPc7x10nUz35s0uU/5MV0juJKGfNKmg6kCiFLP45kXf0Rshh1gMxGajv2XdiH
Xs8mRkzkDF/4GSiQmodyOhaAhZESF2aMrFDIvq6AXAMzXogwncvmopt5bE3HeE+a3uVOzCYsBa4H
/GacFGacbygU1gWSLFaWA8PTs4sQi0iVGajCGhDIts3sQShfIaPli+0YCKX9wQfP9+peQsyCeXzy
u4aG3o38NrDxZHRkjuKCEq1OqrvB147bev0J3iPi0P8I1cJbsanyvKTQ/C3phm+utxVp5kQGRAIN
TdxFkErlcbswPan5afFeF41F/Pr+hPXzrjM17F+mQjQLUWZuBjPB40NDI+V5mBI5lbZDb4aq8Tg/
Vm5YQty79NcfreJWGw5OOUCsjMyIWeycHtC9rr7ScUvdOnP+gmOtTlfB+3MAb8/mR61H6eBMsoJT
1IoBUskQ9nTpnWFGCjekcgv73AkgpuNpF0gWw2R8rnR6tlLX+iMJnBhoThxN+iThSEaA7Qws1b2W
ixws6yJw7h7poFuwMSYz4OWJmXIU6i7Bu72yknapa+Mmgkt+MWX2D3rcKksGqW7cxrLUyBzSRQdg
Pe/wLkUku+FLyEEfwmelSYBKzDJ38Cl/KFm2H3o/0qua9QJcqkB4tH1IOEEtQAwVxG7moh/ZTqjl
uqDVyBIhWealVri3DyQS5Ca5wL19CEG8PjLh+aq2rJanyTmdYygG8mn6l/PH6deshaNiBQlkAanE
AAXH9AG8EXJk71wNHjaOHKNJsHa6hHEKFXkOhCHT+YlEp+gKQu2V4tvLgJRmEGs4mtBpbEP/Xswq
vd5OMi+XSEzNklMkAMS6oYs6qmDHR9zDCqs2VAtxSxHOTIOxUhVHwXm1QM2e5+vl4irmRohb1poD
EG7HJibVD8dbZKrkaJiFAbf7fJtxGqrbSUIxXEK5iK79JtRYkGi/p31mhHDyCspVENYonr2h0dgH
5qBawznC+fx3icdNu2uxEGQ1ltNMLVzSbk1cxPxgv+0G49y3Yqh3Q1Dmi3Smxi/xhVxotP9njDZp
a9m6fgbs3c5YrgBp/LRNrBP4UYQcLPHnZn+m/inzuL7XFKXEBFyaqYvyDA2yP7aJ5gzbLyaO/W6m
7/PiwkeLwK8etad1khDSG3Nhgxnoc8RGx8dvMCr4I2gNeAqxLevmIH+X8JbHEEE5a2MGlXGYw0bg
LNQhl41uOKwVs9e0f6UYM2EqbUFLr0kx/9FAYDEkybPnw5bXyOlWMpR67k//zv+7CbvKP2EkotWo
Q3tDYzEk/GLadYP+wwvO96AGviS8+3wKwOtm3SF5P/FcyFO9ztMVB5muIPyvTC/BrqUu7joVIkEi
7nX5mJ5gQdBKToR23icE/xvBmQ4T6q0xZBgqxmH7R6NrDobZI+4+82TO3f5Y3LJrdUpxyBLs2Act
m7QZ5HwQH3oqfQ4/I8rMf4k6mCnAN/mz/J4G0l3IIbiWpgJ/NQ82SpWSBOOKb43qMECRK17AjpJ9
NgQyvk2P5anuSCjVJB1uEeQ8btEV+r9p08QupjJB6kp5qbHFnAKgzq5+z12nCTxXrfzH+lmpZXW9
rXKe2d1IqxGP4c0aIt3E4Va/eiCY65y5l3Ogf4TiRUoK1gg96sezcrwiy4j3o5MgSSHYzF6hDtes
IGWj3ES0js4CaZm4Nqa4P9v3TVhIXZ3UvJcFT5jIKSx9D7FKhbMbDMFFwgDPk66EGMUdM/t9TtKR
DCsLfEiOcSetff6wcwRPTzmdJoQ0VmP7p/mCIECIcWn8H4mUJzkKcAQqLngeDXbE4E2/gSsPSm4E
8qZrGjckIHmpZHFE+TQy+P02GHZ0I+/5atCHZMtGYj/I8+ohexOx3jq/rSp11V3/chMylRFXxuaK
t1WBsksQ1mt3DOz/X/ZYN/b3dWvt1+PPRaaWWfM4/JUnmvxV/Rb5fRTX4875jCqx7wybOSiV29zF
7ZZKFzCq2kiEBDmzqdGyVa3y7QDEVtJcxe+RggceCE4QyBr409Yk1N141J8atouVeu4f2qKoJHdA
oWmKVPAtXKbVYmje65qdZGRvCMxfB/sEbb08XBx7BIQSY4KC/gnLm0TXghsV41CUHKylNGZFuE0H
djOglilndPTwl42LEKuNoDiR2E8YaXrohsvB1ZNPWQkh+tH8/hVq64OvG/rHwxPOoRAhZOPYEcwX
gNBF3dZ/TvthBPJ7YEh1bDijZG1AeXFutIu4C9G/qIn5pNTCIauCBsH+PKnqocJC5OyTicGpcB1c
+BIhiq3oQCOZdNPzJPCwe1TAEnhTuULOK0ErRT9g6LTlHVORhuZbdnM8w08BCQDvZ4Ccfey97Vf/
kls62X8QcvGEv7eTvFZykNwwfMgwBVCLRWeWf4290xvKreTXeDJ5bHXIgGDqUrRheow7vuHruL6C
1RR9YdJtwF+H1iN26XlpQDOW7JMPk4qb4Zp6Llql88AZ173Bl9lFLj5hvULKzPy95BbgJQq3sJz2
qIWL63YBWILR3a0hju8GXReWTZvpHpDQG11zTwT46SRa6FdZuFUF4r8YwAEWi0vt3eAkgZi2wf3y
QU51/KRwzoEtNXJuuP2yWmqDxwmP/yFzmwW0LFi5U8vJSrMDfXn4G//GXuHq2BqqTi3e4WQSxKZ9
gtfTZX9SIOi1AD1yOVpAezGloDhEg2KgeAl6wI11CS4NxXeBc+/WzOghvexOHSdp15xVpOnUG/SG
Yrg6OTFW4nC5wK14p/Xt5jrZtfyI+LshaVjbk4lYLN4MUXHl4f2+qGUxVxC9tRco/ah1ItaOgqQd
hdQ5TrCh2O1qr4sjVn8GVvkcAtKyQmgYqY+gHssj1LLECPGtzZKDhOpAJbFLFfsJllJc2ncomeGL
FYu7nKaZq9UvUazuvHuUd6h5oBLU+/XX59wWvtF5CxZM/4PR/8kgFA2HhIAnVZ+PgyeuOtotpk3c
55ebML8v+W9mj1YS78hLZcFT+DJBcLPyvDTb75DhYVofSAlDf4mDItZ8OoD/52bWTeh2ZzcjvQiT
MfJ95kFe/JaBZ8Bs5sQVxYD/UhqI2w2QPcazbrMYEQqn3Vdu/VUH/sVLw4W5o3qPwAy86LEfKZtL
ObgAqLTyV+ZhgDOWux+wZz1nQwhV4WtVs24CUKh9Akq/QpvDt+v83j26MszCaxwQp/f2VmVV4CE6
OLb0xCqNfH5m427ipQfJ/3A5qLrG3MlDL1bKnltLYUoWdus0pX5xibp2gPGT2w6eBqGpZSjnegDO
9OHIU4BeRG01VPKY0RAOIGaDXZZOZklWUkbaZBLM1hAWlnq8HUWCTVHhT5C/SNyaKBjZSiZch7vE
L1FHLOg/q04sSDXkWeMvlBJ+I1fV1Ez1GngUvohpRkrWEpBQ6Yt3FE3bV81YJgfjzN0x/bM+iw8x
Bse79QP0pcrpnE/Vwvh6LJOvxrTVYjZCigPsHTOj8yg3ZobBjRJsVQAFOCqX0CaXXQl+ikH+XxvR
LrvuxgsvG6tcTyfAd1SmxPQiehSpemXss0cyWdEAlUA5ycA6ZyDxoybFEHltbWb9hfHIRdAHiJG1
uWT5uhBBB1BUaNb62OpYGQu+A9GC9BnBs5/SanovqcOM2vH/URUgfsOR+fbOxGWwPjQcL9xl2XEs
F/N3F11N0xjo92fFNctCdRsNWm2p7xrvju39dxbRtxkPxa4eB8NWisrB7xacsgocfj3Zz0DFLyMQ
PA80Gs3B2OCdzmPdRcAF7MO+5G8bpGdn5p1FMWBoXu7irbwGmMmfdLE2dH4PU2qnivsKRKMAEvEJ
8bJvF+9g9UzOt92ymQ0A2nZxoMA68DYBbtSN9+3S581Z5ze5798TYKHDkZXqWw64G4dCj6IuLacF
C/y1dU2hMxFGV+Pn2xcLhlyBmbCDBBSVsYkZB9q8DGF9GjtVTUkETuoGIO78rgg61Vso/jzNcqFL
ZT0IdwUfFAgAraNtgDxygxZAIaKB9raaMVGEDb6EhjHS0FM3FiRwzCTe84/bDu3er1PyknPkcOjW
nJPZbPpV9R8wVeEo2YZHV/r9pdpIHyBk48iPWZU13iom6qw4vFU/TYuC1kMRSZvfcnp624DxdMUL
+wzVZdhvMuegCWSOieEYWtd5ceamFtw/fHMtmSCZK33zMfz8XleC8+Y0CWHoZ8i87TZOrC2UAWoc
bRI3DdXTCshU6wo3kR6twLQjGR8mnlh+nBJDuW11QNFBiaEPbH8Js20WeTPD1nx6UZ+7FF8y5Fk8
OuJ/CjplEXRF24k2fDITDxqZgRgxoiPX4SC+nFR9MSUbzXS3Mw9sqLf91Eq/m48MahRgYVFUnjAq
Mk6HUTj8Es5ZF61C7k4WGjrjXU4LEolaMB6hRB1qX0TUW6Jf9GCw8R1n2OpW9Oz1PRkArMLCETGP
3o3gogX6JlnAvGj0WD1jtSte0XLnwzQaSodfNCOsaknaI3dLj2sJsWuYCBs5sUkYKo68Y1933K0n
pi3T+eL/Ubof686p8m/M/OH56e73sS8ttGqTKePLG5r+QyZ+JMDVenlv/FMEEKFPKzh9gtfOTWIe
fX9tmJ4UtzfFS9lMbvyWKApe9N3x+MSv4hURS+ffIJ+I7St3auW+LdP7mrYviVu/zcM6YGOmt3Up
qKm0PxCo1E0AX6hxS8IBEgrZGVUOMLI/H6JgmgGRDGAba+GIE5+LLMHMEN8zXckL3AQy8jTfcKcd
QNX+0u+MZgkrCw1c78SBD0LqAQEi2JtlFB8TJucUmbRyQn+HNZOx75BL0/ir9CXliil/83/XTs0r
Tk+oHjiAMIU5cbXr1sPwLuuCH8Qvt11hRHjia/rleOLh53ZH+aAz26Xb61fTrxFnKJOVjOFKwOKh
/A1mGskBgH5L5jamdTy1X3ElV9w2ZrSkjfV/NSsnh6t6mIbWaSkK/hPYmqeOoHWRARKOZCKgmB7S
29LHzEMK7gGlhZbNwljTcnBDLAY0ePsrT73X04UsqRzRXQmXJB8IubjE+7uDoHUnVQQooU1UYdEy
bemQhNdrBxBAwzae3xOmv3P78HqzuzZ3OSg6HT4ZhNEELoaS+xpZMeMz48abyZEeJKFFET6RyrJ9
OBuvDx1h0NWV2f5QU+7vzSKSksO9SFuZpnaxEA1CsUORTXj7TRb7688CgMCU5HH0HCt+a7SNoXrJ
9Ix8BMTF9q3UaLsqrk4DAxAdCPa5PLjzFMSJXys8On0Zo9WI6h8PxU3HSq6byT1JVUTyq/aEKt1y
M1QIU2/rmY9ectIxPc8Pfi4blNvmlT95Kick9A4CFY8LwQXKe8D3tpCKwEaQ7W8bPeNp0zNo3nFg
l9nQOvjQ6+3HbtP6f6zatTNlkqviC9O++5sWmADSD9BkcYfjxDoovfmO39/x5MelhXcat7uDu1vI
31nynVh40whc6VJqp1qcv0N/27Jdo40zZmEJE82iTYLzXm9tRyB0f5icn3ThCcy3SZNyzY09mAgc
vu31VJKI7l3DhE0YexqQzzc80Kp8v1nNTfvJKQTuLJ940CG3RX799M1qaA7RxbXAIGp3eAdFJvgj
zUWAgzS4peR7ZiiFBuHhHjIrUBjP7k12MIy+sdv0jHm+zh3uczbaIYpcN4VnIfu/2/+Xd66s9a5g
BboKynuCdXZncKOcW6JjnvTTcteHzzwdYsjWYpP6mGRyQYdK6bipt/hrfP18Ah0NqYzA1r+9OgkT
V0ohcRGZrYcMXNrbaMubTJDPTPrEDck5ffuE03gmt/YIlHqKNadHlbHTF4jkHrgUWu96N96tz3D4
v3mQpTBsTJ7pk+WAa1ZintowC8YK7pLhOuCUfUIIUWTAcg8w/PRQocBYr2Rn8b1a/k8g90rBQQw1
rJ/9str4IOfDSSCQDADPwQNHMMcj1k5i+qYj4HB2jz3+Dn1rVjzmc8jioCcP+wg3ljeVG1DM1Kz2
nhdabFx3wBc8saL7mkFHEc41/YtgyRygNKN9hQOSP24lkqjh/yzDT7MkW8QXuwUFP8dFO1Jq7POC
xBUskmaP1L0rdRP7V7Ck6SXBVQka6+I3rsIMYnxWEnp95xHi8LgCv7eZP4hv0UPD9o8WfTGAKYez
jT+e1Hu8NcL3F0h+lIp2aGxClynjfY2LelOpAadMBGDsQGSgZlHkAWsM3g+XOxrP6rI6RpAzyGg5
njcTvCak5ZijGpaS2TYjET9VYmcpoxud9evCZMJW0wt687pnVt4WiGEwxBDTnKgx1EcVG/mL4QfU
4I0DN8lw63r/AQ8KgCdY65YN8pApv+I02Wq5gB7J74Vd0qPdoScU/U5RDd+puelqL4F6KNc2DudD
S38Q5gygZlzvnmZDirxR6jhY8AEjV0/2OOqyDAtba9cq19Z9iW7Rb7enDQblw4IZYvRIV8zAx3YF
spxcBgz4Z020lXQ9zo7s5cM6RkivSDWAu8VFusrxFQ/1pCluKr6kuUU3nuooEzLPgcAXhhT8byih
beCS2lYEWIujC7HHvC1lNj6wuKvdbqAfQWNy7EqTwha8/4igd0sP70LJkktp9lqsczoPIoPKKa/W
dvMRgI0HFfR31kxt1o57AJWZcFHdLy7q+wXJ2voKAVoNR3JGxglbpZlDN1EBSGXXqgmnFZavwfnp
6gIV+kIOjzOxWahMtmsgMEOid/HlkXPJfEIfF7KONEPO9HTKrjh47XPcXFNoHvr1cO9kbpv7F6m2
doRXSBDXn7qoePcYyt4I41EWGJr972M6ZC9uYcciHMzcPV2AbwJuWkMS70NcygUx5eJHuqChf9Bn
RcDsW28jhepfBAVbpCaoxweG4392zLntSF7fctNOCFAiIvLxtBiprf1IUcTpErfzKEcrUQmMKrGD
H74nmrUBoOXPPCa6TrljPZb5d7Ra/KPIz60L1R+pzYZwYkC4c9ilv+Vi8hM7WumE+gtMOx8CY8gR
MuoB5T6Y/ySB6xNd61MsTBSVuZ9SU7XKBQngxSJ/4RipA1NUcNONiT4wAZBwS6v+89Vurqh0J4yP
E9cag95MGoRF5XjGveYta6NX8zI5VV4IYfdgTbUyv2fo5nfHRgkcpz1BMU22QKtflv7DiF5V+3R1
U1+f10frCzqdiAa1cAvOTEIrBcnGe4yVBEBxhATm7oOzltEitW6tePRb+XjE7fbsW/lWgg0gOXkx
7f2qX8QIkicY5KRWcjs0plGRf+0OYH1kLcevCSZraFN750Nw/OY1ey7CCidRo23bPcAntgbK1X92
RtsLfxD6vm3EWJts4KLgLOQ8uoJENQlahNgAips3AoX2Y9BCYjSX0htC5nCZy71UYrjyMMfv5h6n
xDpgTm6dBV/l482D1uM13+A93JaD6iihmp71H9yK+XzEcw1uZaR+WbBo9FZzk/ZOA5Ym80fYuSGz
1iTVsv3dKSGdp4pFkobGIDQQNyfQQbKgT4EMzB/izkDbJhhr+KenJ1OtXzUCdpFA24Rzt4ZR93PC
CRzu83P5LrwQhi/ZvW3i0Mnx2S8bfuJna/RhRA2kB9BJGmrYamiKHsfLaNhoMpB9HBtvIG4t1XwL
L93oyRzvMNxcK5F89kSuitSHH60GrbLKI81QG9zIgqg8XB7xi+CmPaWsgt81I/pDAjaGp+K4NnE2
Uv9gxoew14cvT4u6vE5JljcpHm7kp196J9RIzl6vAi+E/3bYhy/G0Z5frgkrXz7ed2CXvPcZ5eYp
LAoRj0DNlwNjcfFkt9GlG45KtAuUdHJ2jPJnE8+rhvi6lTP19vYznSEVW9zgKKVa52hj3Yyxt+Bp
IIQXpuwRVhXwuRvqPInz+D1FQP/woFiPzCfcDGXO0ibkT97jePbC7Ac9SmXtuWcwtUalNibdmlUU
EiuKMromkcL0X2GOWMThX7N4RXDqW/L0+Nv04o0705foZuYpLpgarQ8gNjVozSlLsYz70GYY9MJW
A1cYqqHXCVtfnk1A/71Iu4aizuRp5IrlkzEYjDbXBTTdE6LLQetWsdwE30wd4PgYLc5VgA0BSbF4
1GxUYKarIDfee+AwoDeuZNmY7JFBVHU10XdihYi4n8BL66PhCEjtfSG60dUuAEKuk70s7y3472/p
q1pk49eHB+tWOd/Udamja98CA4lpnJ9yB4LfsRIJXT3uzHzEVmAw3lucHJByCtHZsS28ypAyiJme
Ki1thaZrJUWI1zzmrAc7RcBYCpATZly2Wieg1/7oFUENAAupkbRpu24x2Qkchr1GXV3R6ffcjJ6d
9skXj7cvlcy59PSVeV30XXIGjMO+LLYNAVB3kCwKKTQnJyvrOxYboF5pWGUWWa1+YnvP5PghOtk5
enNw9SQ6d8hFBGV0WVY0j2IM0mg0QrEpSFgLqe0IYI8hzuWaXkPOzbjLH0LZ8yQP/0J5HSAGJVYV
l6azbpacGBhJU3HRPT9U1gyn3cELntlFYj/jtO/NMhpyygaUODw7raKaLaI1lCAYwbQa+2qFNJhY
EDMqYdMa92lpqcsfaTkWQ4PfLQK3SxPjD1bmohZDbDdby95YmjXYlqGzOulipQIvJepLdjW6CnAN
4QRk1WlUkxdEPMJbfHajUW/FoRUGkKZTDhx7W4T4AbyLXyQb5jwSO2LQlT1xhmIx96qpIMysxIxh
BPshw6i9epaB6HdCqT2aHlk0wi6jVV2BoozX2EyIO5Y5xyXhWMat8YEpYqcSElsQJHBe7zSLEeZK
Rp9mhsZY9FecHDJ3sMrFbcEBnx04EodNEVFYOwGt0MFPhUbBU2Q8YTic+vw6mVP6xE1cuYA2QLX+
R1LwKneLl0K2BigE0bitHlzX4psFL2S9nlXf+7vw1Cw6gUe20tDmxZmIRHKCFZHRvMPcoHMLQzvI
YJexNbcz0LUfm7ugZJcjPXElkt2beM3kaYGNzkq29jMQESz5v0VvgipxkF3oIMo56cgQZXzUrTsb
IXqxbpAxJrARig9ne/YUEYeZa50bb2dwT8wNNhdKGh8aFJq/upr/IEiUtrUyXtNoXFdIXl05wmyv
Vz84frGiw3piNcXPSvhqir8dPsdOeFfInS56x/lDbHFsxip+eyEk7Z0/J/5qEuUkYzB0mNBGXTEo
9oXlAhPloxQIF/VHInc3uFrw+HuHb1EN6k1Ufjp4qWs3ychkSk5p5qMbWh1xppZJpc/TMEw167qu
ynnTIvQ56nQzwWfKDFc3Jbg3PL6Xp02PsdKMKGUL7uxKgVGhzoZJeONZcvOkIdJkavAmyqb0gfUX
1w33LWwaaaAaTBrLOvlkPnHvmbTi0HLNMRdLDNextKn2NBcd5RbYQInsNGagQX8S55ACCgLMvQ4h
06qDrEgNwZxPYEZteGn8z9dCVrntqIKBEEhovro5+pXIh/jnnsliXXg8SNOv7qodnUGJqh+N7Lzl
d7wepyIyLqHqstG+uAI1MW/YGWLmGkywcA1ce+EbjYXvB+vQUBWvtj5/D69+YGPf8ZnckCsHr49D
ESDVJvf3XJi6skobqul0ANyjQTGCXI5aumOIYHvmI5MyB0lmYLc+BhD+phwwHDCsfJW07pZrFOH3
RKXwz0OLTvnibQN95UzdXuVserlWP/wrgswXwSTJQ1lRJYGEdYXj9aDuamm2BPKxNaPM+t9WxIhb
8ftbFDoAzX9yhIWxiMt/BTkAvw4tnU2DvPCb43hk0nTvM6ouS2PK96VimGChJZpjmmqnenOiMzuh
PJnC53YvWdW+fUcSOt4eNWJU/cgEFCJ5enHzD7ADkuMmXUefbux2SscxIeKVrk4boaSEUfEbO62c
4EI+YsvSv2vDX07jV2JS+4SkgeEduELyBANGUR4bTbv4adeJOmlh85hXcMLr1CZv+709NveI/+1E
EzxUS5j/UXvfunUrUpMrbl+bLhj/XfI4RXR5iwvZDY2+UNRdmpdUHstxekj810yaPZClk9MMcVGn
cxsmyIMaBfQlc07aUhREn5uUM/ELxiK3TjtW1Pk7eVvuSTz2faNJ91fkCcwuZMf3u3r+BhUW6PVX
GUctXQ12J69A5Pw40yZXehn+4xt8+77/9GBfT1yKlhdm3AlscL89Indq7Tfqachci4gUb0CbXx13
8rcgHugI1S8V68z8VWp3XgJvIia1fLgTuWovL67VRbx4wseG0I7OiDaEqggwPyMC/Z4dYt1DFqUa
C9fLiTpnLIvsReeZoAd0sjz37NDQCReo2f3F6qI54u0bNixkVcOulTxd5P6QR1QxzjxSoPNtTthI
IYQdyl4baZYTLCaMfPoBIGoQ9pPRxCYzCj6H1TAzkOSVEJhRN2zt9UnS6g0G1ALvFZwkf4tNew3Z
aVDdXeHeslxK+Rb9TsWSCoDD06LukmjhBlc7V1wPnGNBoRQq2NhqLYxuztI8sLix51HyT3qFEjrB
LiFYpSqqmY+zJaCTr3MfiO+FanBWa/bZFv8ieHAfVBIFOsrJIcZvIbM/Skx4M5qx2wVKTbpstcme
eamGXBMzWBOrO8/qHN2Q/dql0KDUcspb+L9NuG3ChoSqW6nGnhEEFpkwrr9xAiOLsPgf+k4fMAI3
CtpRHuMgnQNMiJIWrRYyvs1CdeqKf3/XIu69MWynZ9UKPFteAFu1fD7l5Oi0PM1XpdRp4TBZsxu2
EqBo3I2ayifizWqNZKxreGivDd6F265LesA6v+A61Q84H7VdSZC0jClodcZII3lP1yTRvYwqwN7Y
Jyp12zJGjMnOKBCsB6tf50JWPWGn0OdL4jtBT04O4Ws8E3iQFEiTwB9AL+wv3G23zVO1OV4z4L7o
ucIql+FdD8zD9COqtp39I6LVNX06cQ/Z2F0mCePNJKmHdGJsoGn4xSJzKq2DpQfq/8j4c2YNgrAx
oxIkLcFbeG5gKdLa3mjXdu8Dm9euGbdcHGPLOwcX3VGKkuUiC3jR3lpHbRV92z8c9ZO2Ok9zrGLg
DRTFjNzMZKqq2YU+hjq2MbwfX6yvyF/G6HGV0wqzRJE0UWVJo0dyL/Wu56hqUAxDmdrjfRRCx9cw
vJPhW3xg5/YG9J69+LgmJ4VmScawqaCgh2QYjHvTDCP1XJVv5fjrFZSuJUNt3lsdnH57hGHJjHwW
FHXs4k/SsAY+tgEdKtKCqbRZQk9kl2MsjtmqRnOfJCZqFygFidE9WeWDgGGDaQTWBnmwFaMdau9m
OgHZlourB0674vib9c3y0dhuS3fFKp+neKZ2dyB4eAYJ9Il9JxpGgjIU55ppCsGZVhXVP3BlRtKW
9huuWg3d8VIMLIgbL3F3uLSq/u1AINfhLRe95HvFB6YupyoBY4U1AcLycYQXxKz8uDlYvkk3Ym6D
1OOxLL7miav8si8Lszux8vb26aB7TR/8fdBuZXrb0S9oe2oNpsyFrBy2AmZbGj/9Jz5qEaWsqmND
cOw20Nov+t9x3GATZwwJ4gsL1fYGPWOTa3PDUyq9Pn1yAJ83cFtlWdqcHrs2YyZSls/cZNSLVlIa
8E1bUoTkh0Pzi9M/SZkmVyfbhcTgK9IkyS0trHriwc/E4jFwwBBbxc+UyR7aJa68wPG788bq7ZOx
VFDVrKwavNCLlQgSB73CMlvVNgEi0nno6Z4ogP9oMuUnAZUyWVNgprRWghvZ82i21r6tAmPtzLHW
+IgrrIZ333Qo2szOFcauphP2A7l2yJh7kLYOEtRb3wFKmut7KNDvEPczrh+Kum8kEZFWf096u2bN
sDv23sDphPLtZilbqrzHWn+fOsmSj+ahillYvayt9sOIfIPc/dFaGiirDR1Y2wwmrJghUv0itgMZ
WkhA3brQJCsUj5OuNlNmzi9XayLFuV+QOhIgj5tn41i9HXJSigPrH0ockn/j3WSwMsVrNCepsb3S
1wBb/+OGPNJb/hfnUwgkwhQERkqIizUtOstkdC8cDo3b15kWrWvYIZA+tlQkVN14ZtNhlNn2sd9n
32VHdvkRRggDU9wfTHE8bNiN/J5u6lTRAkMznyhm4IedXpqtc+MeH7GCPm73TL0AR6wTgr+9URnY
LZvDLuWE39odP56CflKyQfxQGIqdEycyO8rcXO4568hFI1wQfbK6z/QwfvwDqbwdN50h+LL8j3I7
qwpbcUjvIixj9cb/HAEyF2k8IFonUdBLhWhaW3RCQFWmoiL5YhXXg7XtNJjMifnxSJbC4S/KnwNf
Jkh5rZafJqkF2PV0XtGgZ6JgG2h7qWiKxd/Hm7vcmvMPtKUge0PDCnqHeifM8ojoT8cnRUL/6Tjr
YKm20tYrJoq0NkfRjnlkL/UouI5WFP7V/Jiv7AZyD3HSUqM1Rt2YfA2IYenGqDICVV7cbCO3fsLh
ZYVSF/OTmssetm0dzLLQ8uaDtOvL7Nk3EEMw97snHKklT9DaVhZXHVVwQ2rc1SvQnW57H1SX56pI
00wzG4HgWrxXKqb68tLSkUyX++1yTZGzT8/3fpkVBh5ESM9koY8x+DbJOgONPkwQMTVorTKbcilx
1xfG5tujrd1w79Kg6BSjGpgrOwLgeKfDQN/sZ4vl6rRJt/h7QUMndoAF7vE0wrDxd13xyxo/uzvr
Zjh+Goz1oKRfE5rEMYjL8YURxdIK2BWdSXs9g83syqJVkrcGzfaicBVwwHDDdKptMl10by28V4It
u5FdeAcPV9Po9rY1yIGM8o7G9CMu4Lsrkb31W7LTc+UcLCvH6B1GHct1gCwwtAiaRvk1ex1l+A2h
F8ZUHbZZBSNeISYkTrGqnqwlCs3yCjBuAt9y55xrHeuivV8oS6f4qfjr0apXf2DBgbOLbNo8AXrg
qhZmFVfXvocvKKRDnbHgDISZKpaEmy5o030Oe1n5Q0o69gylULwS3Ol/au36sVWHxZeJdDfZ3Lpf
o8sVwXy5BsGFTdTA6A0xFAf18hWIU320lwt4onqK7qwufJcXcxNbedUdE/bV5eIm9z8k6utVnh3/
umGx6oaX/IL/6CVjqxXALCCKZPJwTi1A/V7kgAhciCZi9zHobjhNieLyYfaF2appr1I2RJEwslss
l1tsPFx7/ynUhhsrkLcIdVn3rtq7bht3OX2tOPnN+9zy17JIlLdVyBQ/tTCcmc3mN3w6Z3oX/A1p
HoXESZk/ZkH2PmwFEABNQVFBo8RhRns2MinUS+KUloxReos2nWrcopzQ7Sbd8EyE1X88iK4euBDB
i5u3xntBNZX49OkhoHV7SxfT0LxVdpmhCavqKVtnS+Qy3qiUyb8pztEuMjBNl0sNlYAR3gK/I5Q4
kMkUobzle8Sa8AXCxIOjrRkCJHFO7x0hYoq9kYm3vRKYGSc3H4xJOsj8wrwYZ3KFS1bl341d+kqW
wOBzkr6fvRuezGodOBsxnLzWs/7p6u1maDYKICx/QIUv01RcSTeRANV9XZ1ppK6X3YZiHbWJ0+yM
AohZJG7k5nIHLg7YVEHcvSmRyZP7miYqwMLfqV9RLsvpfYB0dzgmSlSRMoxFaEZmYgJUI/YlzCVS
MTiIm5GNktYFOU7BysXvplshLlVcrxzxJbK5ILK4exlDeNx6k8fX9v9k24rJ6/EYcnMuUmfREwNY
i+wzjsoUaqwRVT3NpyDopbjOyCjnkMEwDunSGWz+4t5T3CgNqPQtAFrcLyZn37ekdYrw0vy8meX6
aIjbZ+NhfTCuhjELS3wg8/5vgx15PKeP7MEMzTI6LBBHwsIjRlRcExU1jWQu658/g870zfLuaeNS
nPwz90mwW7vhNa94z8MbQt1XvCGJwoGsqmDW/aPScU6IHeTURzLHWo6MunUxFvVXD2ecJ2XBbrrp
UAhJyqk3vSY8gMo4Q67ZNlf9KeBRBhk2jpE4sAFNo/DNDroMqqduZwXJpRHqSDJ7o9sA/pMi+o/f
lEK0HOGPzJO8wn5rdgv9IIv0p1r6S8e/T+B5+zZU98LFLf2V2ij4ug8eONT/tAvNcwgttgtJ8+T6
xBRj0noM4hMJ1T3oVh5VddqvnUh7+O0VBmZ3K+zQX/oUqAcuhetHhDu9DROpE74pNWeP3sjyM+NA
FaDap+H7JyCS/Imny8mgRrlyAGGM0Yltatwf5m0unTu8Vi7epnQnLeQaJf97TIXBqQ6VwBqHoorH
1HclSTsN5fnwYBzcKxdxAzDLPtXAgsZLzceblCyTGh+FHEXQbdQAnM65ytJj8Rf6UYrQutwAwAJz
6Qb+z8bIwNpe4AS3Q78VyDvKzx70YiykbpE2RfWkryIgDh0fBr0swdR8g9anVJ2HSYy+V/JSZH5j
fwgOyHdX1BvwOjC5WVeTwgmuF+j6H7X2kekqvNHKgyY5s/Wz/ZJRCpJt1NrV6gGRH6/wTq0FvtI5
Oyd7yZuAzkcY2u3bamwLNzISGZfk1o0AZsXkDO1Xf6oZGAZE904j4FlYoS+p6rqUgtjZ6q58LV+B
4653niAr1r6OFV/znvtSAi6scNSXhu1uFyOTzofuQFNPvetmVeyposTQwHIaPFEGoZxC1NqWavfz
31tEovB3SDXIo+0NGsH6V9H8PZauYD9KufqOk4iQBU4oLi8c7stNmua+SfZqLpR+QDncIZeLmPct
4zuHkP/WdmeJ6q1cNSzKZcojIl/Fm85nvqbIwBuyc4o4Nn2qIRwhjbK+ffkFLdSzbNT50UMdAlSP
rgeL/Uh5XBg8rMuOu4cGf8YvPoCubxjEJWKdyHja8Ka9H1H1KdL/SHlUZ9AwGIZj81PgWLpasbd2
u4uDmUdZak7Dzyk4JYcNMDhRhSm9oGxvkEqMyQdp5Du4tUVGs8VjJvH67vR4q2vteyMFEOogbeCo
4He1QbnGx9NgCruaZCkVngUomDfPeddKDc8WoAgI/+HKeTMV/RX6Muub0kt+ed2pyy0ftSkHjwh2
8LRaLmEpfyLT/TqO/PCZbp1APjBEvx6fSxQFnNWvRlF66GkIOT4Zd80xo/5GoPUoKzxtDLEEanmb
ie3pmMxzf4wcn259r5+Hn6fB+pfr+ADcc+lxG5nyBiAR+LA+t6cFNihix5y+scJUKjZoymIJLOYm
CVX2lIMeTwnBQQLSbtEAjdoqG5pVR+sOlrHqu/Kr7Ngg8Gjn1sYbXRgLlPPJGIHNdsLPCsKW0C1m
znYR8iTFR2saLOloyUsXIqPl1th+0OOJ3Gr+DCnIwd1jI/Qxo6+II1RrLxfsia8y70pUWvs0RLsS
U57CssqpesSeB90DZ05HWE4NMCAXv3089+0Expc+OQgrKIULK1HyoEhxvshKVszY7Z1pThg8CFJ5
a9hv8F0gNSNq1JHRONHbCfUtQaF2g+DoyqNKaMj1NULEMWFoC1xthLX5LdcLKrKNnVV3Kt4gPfdg
6fS7ZdfT76q9Jk6P1QCZe5nx4TFeMh53FYSRWsOiLm/qD3aOMKT20HaU2fjcL91NanHy+WGAh/ux
PoftTf4qjLzIhLjuYJf18usHIsKKhM6Xq1z+RNvVeZlNTu0CmpjygwGsIQM0W8WkqkCPMpWWJXrM
GMsNVnirj7JWhUmIXF5bGjSPRe7OK4kQ4Z0slHX3s4GXq5NMg8waeCPC/D1BexLC8k7nDkx/MudZ
5Yk3iFzfk37CMLrt3v17PgYZzd31rKESq0cJrbX5MxYWQm+l6umCLLv5Xh8yCEz6LAxVptlGqh9m
7HhAktHgLcxsDluF1DHUm6rQW6yrrJmu1Oy3Pr1tYEgzFyxe8gqzETVEMlPh/R9Abq23nZJUDp1k
Pi7TMttXnFVh3YB7HTcSngxDl4nOGVsC2zQybbjcUNwXZHrhwvvRcuAurtqUlvOcx/1jvIRPA0kT
Yn3R8CjbSWGRt+ZtuaQgleiuzPgKSCFKSW6vj/G2isBg2rGL63RklWRAj7PqttXJ4CDMLDTKr6zV
6xUxFfWfivcH+rqv/5/Cep/aqGLnSIFN/efqBcaXiB2V5732t3qX6QSaH2SNaAiAwoNb8z+q9K2C
sPs8eCQ/pM96u0vlt9kZAnQWB347O3itpB5J42EOeOoapid0D2B1FR2tGr2s8dCiwZCtWp8wlgDp
T180OO1oXurfo1xDnpCGV9N3+H8PpSPA50FRjDw8XYnCxFoIK9IdZdTSkIoDvdlHaprK+bYqFpIW
fYzwTRkzpuoHrfE60DBikqzIJHY2Dxa8z1FUiUslswIqaiAJ1F7o7K1z36UjapksMMtLF2fHIS3z
CYQv649QoW6+qZFdw1LpVHmK1E3pAkqTxngKKjv+265gn2CKMBRWpZWIb+QMfHR8ssPk9TjI+oHQ
IusYr+WN0C5NM/1w2spnQLkj52gpbMYismz8YbUC6DX3VVnVGnJ3tKFpW2k9AWNMuv91PeZPIp8W
QPrFWu6+jKe3HPsPYMKCqfizeVkJEDXNolg+YXdsXSH9H2qsdWdrUvliiS84NRNb9dgZ2iIqGsMj
yxYqGXODQnIkzX8vJ2K/KoKdttvu05+3OHPvEKQU4Qr3h9jVEi426L58rf7txVUDW09bTPAwia8S
lDW+jetOcH47pk5Im81d5OmooOh35tFOzmlWLv5pR2WRT+arrVaVXlei4WRcKzWELKkHe7q4dhrk
eDkxMgwIh1v3LXDC+Ilzg5IfjkINjlokOhrEb4X4GaK5UvR05gwhFTbGfcpaqmZFSOd0M0c2NB80
K19coBHhUs7/hEJ5VLK+hGK2wDuwZfvGzBsE4ZiskNWMizQgmmP1qjb+zsdd3yj7ZCKs5WcKnwjc
ixgEK575LSaMNN0dvbfsFbwot4+2g9ejYn1CrkgexUMYRnPEJkHQvIQZ2TX2wCYT7TBjb/2wnpOG
utkLP1T4uz0s/6EiR2AAFS3OxZ03BCQbON/XnFdiqIm39EO6WqEi+QDHdMNmvPuziT1qnonR0FRK
S37gF71QImiXgA1XaPfGxsGrhV+S9BhlgCnfNaL3XFvSwOU5qseWr55gs3teQeWM8M1lkugoLQeX
s2hRBBmPjaweS2Bfy6HoHrTc227ULKR4cD+ectEbCoI48LIKfMsOtoMeTE8pWGeox13cQovA6tBC
toMD5J3UWLnjFb+o5khYVRwoyajRuR1s1bXQ5v0+iiNKlyzgbRqlSoNkUSZDX4VrE+SVqSHnRHj5
1vz0gk8SpaJ1omc7g24PUaZ87qVLUlQtidvUpwAxFtKsAfHO+7UiwRnGGxyyC6LeyFtMaIdbIfZL
wRwQW09tZbQDOWonV4LRxfmSbDJXlAQCdiALgaIHAbs4ae8zqej9OE4SxwvJekqxeVsf06cWZPFU
w7YvjuIYU0YXRnqNfioSokrMsZ5rGeh3knRu0XhNJcaCIWYpgkDb1UNYnHyQ5FYD5R223jeuROiJ
kzBiQ2IOnA==
`protect end_protected




`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PkyhyBb59EPgq8kANKUgNUvJSxwVgcYTKLlfXroHeM6zPnPHm+ATuJPY2OmCojZnDY2A6SHiMUmx
ylnsx6jVAA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XgKClVpS+h3z22aTgNZepCZW5Yffl4m6nNLRjY88G0b6Og6dF7wA3of30X3Vr2BKX5GVSe+jeu6a
q3D7Qa0T3sEnO1qnWdbom/P31G6nS7/pQCPaLh+suxznQX2imRfhfTkmY1B9wExxZtZBbss2GPfs
EFGX8a+efiUiZLAKaSE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LYMHL9qwz9VPPAbHAyLFK1YM6t0YBJUbhdak6y3IQta7KscLfLakFo9QXv7rXKj3R5WEjx6Vg+9K
QUgoa/uCYy+n2t004DDpVeDamNuGIrJU3WXV9mo6tEi21Rm+kIG+CFgVuqLY9JSjwI3dhmEqYYtS
wC2GIO6hKaV0keq1ldvsRFBu71kLY+jczboTe6EddpUktWp3UM/RqnrSfHPMlZWhHp1k3YC0SDq9
gvcPn9DB3vIjXgn+xRbyzZOt/j+s8RfjF446i2RalkF5p/den9o/OMG5jmv4rZKHj9S1V3Z2UuL1
c2fxe26sNIvZ7tpz8RHVWRMloPfcPVakam2zhg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BACIRg239ZSAZHpsLobWk7IZyWSAM1rsaZq5LesIgnba07iijhvT5s8WIOIIgHZs1XEDKelSnU1J
+5cyEbU9WgPZsja6FQEw6J0GuN3L/1QyrvmNIJKsNXINx7R+xaY/n0uby2eFsFE9luplvdOyrCEw
eK82BghXwPdasTT1ZUgKiycyGYtNsp5ZaPIWXI9ezN9oHowcWp7Mn6v2jrdDl4lzJuoHgqRtkZvG
7GqevJFheGfXkRPuQGkNK2Pk6XN9woSB1a9C+FUsQBM5MlIE7zrBQAjONIQj/nd82Hlp1H4PRxBW
1mmFP7PskMeNR2hH5xwkvg4Q3IfYBlw8gdzneg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vUWbACu3JL9XeVH21XChN1bLnACIM0U/dLRQNf2LGaDFNW9CL0o3SY9pOtV226o71+9Eal6i7P4l
ht62RU2AHTweJsgWkXtQBI0/jHIw4/gxbBebNbqZM6m3qjEE5blPsuzJ1njoX2JWCJElO3p9FfRu
uHpC+4hYoccdFayGku3vk1gwz9lLJ4FcYG9mi1vLIY+tzs0o83THQ8dLrg50Rr/r2n0Xf4hxWe4U
tJ6iUOYBQUYjeOwNQOOxfjv5PKfLIgGA2WC8sJb2GFe9MkTDoMAo40nBLK0Y8+klDIJTyx079Bx0
wdRg2JxUF3+TGlXW98+2/iWy94H1CPEVRm18FQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VX8rVAT0l4oniSvb1X0sblwaqcWh2XE0oCAZbC0SVv8fCy8dLmmtqBzFq3w2V/7nyMmJzWKNP/yV
0GW7ICEfrGaBejU3VpwaHA69xE56Y/8NSHGlZOhr390/5/UqELcFOknZEPJXMLpeKjUn2ijACn/u
O0myDIvGFiUyRGWWYKM=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dlKAt52rb1rebbUvCxUw/pmWR03F+be3vApC1VuekYTvk7BFt7xopdHrqsvoU8rgaCBc2wuCudx5
nUcu7bKEyHKFc6bcbp6J84c2uG0ZckyqBn/OHRMbmq4Vbar8C3ERI2YmcbL0Q0fBLzMosVarF9eM
+c6VfE9hA5lx9qpwFJhgk5v/yx6kjgu+kEnG+xsdWrpKrj8LIxxh6gkrPOn+jQtKQSX3o7q35Rcv
W3vWLRYdH+pHsfJqCdT0wL4oBTLa7ozdsufX9l6UDgT4ECxLf7R1TtNj7XA1jaaefThL0F1AUCjF
5WuhMqBOotpDZUmvB91yVtbXLMm0r85tK9b/iA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26688)
`protect data_block
Hz9Izy02qGjc7xDBUcEs3w6cIUd/miMerfLZhYcvwamMPKWmO+WMWxcW9u0i20jBgJs/dLFAvPFX
lbwah3OGjYAt/pIjonB89bb6YxVjrzqOXi+rdnKbuLROYO9HcLfsNzqdpYvzxRugk8rqIS7xIVCJ
JFINcz4aHjA1ybChZgHlkB8Dk8Gl4py0Xx2W4urxS0+PKO3odMo5O/fDlbEvQaf//TCHJ4sxrJeS
jl5N4FV/jIFPnatG82duIppymDFoTIE8irrh8PbzQG7v49vytaftlxc9Q5sSO97poRaC/GKarVak
8l/8kXsWKYkVp80dlZLCMNlBbVLMzUtfDBhRvSaOPFmMd527A2xTng8OJassNOullBNkkar6o5mr
jkWwIUFCcyiE4xK899zUG52Eu/lg+V4iMkWroRNMWJmAXy6T2KWlkx2kl9JIQZMcR8rBYkkFMVWN
2lLtJMvv6YPRzMK43ydUBPKuf6DiKswnhfc5vC+/tpmMcuAPaWZzYjMya9/17GzI4RiC7RHqMTLd
WsyjPe1Lgpm7zQsNe59Efjn8sEUqG6fa6cDu3FxXkhsdbx6cYoAw6i6//PGPX3MAKWBzR111qA3/
aMwGVSaQj7vBETPYkBMaVbVkBXd3dtS0DgmOWPRMtTKdFlLvRLbblXluG6/lKW9Nh/S8YyrJIGF9
QeevNbxf5xRHT9/PCuUITropV5P/9muekbMaymHh6byDkUwoxe/MdkPCAFGb/qWWEOpHmTIwtwrM
7l2usxUzif+Uxrz0kq2V5nS8Q1/rxMlFZOs43Ct3/Opmh8gXLCfvjlBia4USwdknKE1gqBu/b8xE
1mmQJNQJSDRU+dVRj+SpDwd+qqaHvQ6SD1Q+pfguH7y3yFo6a8+L9d3j94y9fERaxZDCTJQcyb17
xne5tP0d1n7aWFaVmsVnBGGNicJOOVrN195rmcdnv5zqcV4SJa4ZsQxIQYt4NW8qM4XYO6We3vqg
VpQTlqbFGwqZf1hlTzJst2VJ/ub+i0eAbj9f44BglWg42Ls914isGvuxfvqeiadePtxLQMAt1DfS
GVOfmac2R6V9bxHSLsJ+68/AJRl+SeblioCmi2CGVNFEXVOGtrgtFxJxytwaZhdwRzVCwmJLKuVK
zxXD2diAllSfY4HRvgTBZzLTA2a2SUOYQUKSDR7BB4b4QEtxLJJZyPnwVJ7iZnK5od2y0uJSQSzR
YAWRFRCWF3zMfPlN9Ev368KFBT6R6bELzoPw2A179CCj8a43f8R8oYsO5bCBh1hiOkAxocdLFFk0
93ddUSrNbmlhSak4YH3PmI7wHj9Ccx9J/DbeqSP4Jg2BW5NgjSd1nNjesbtpcVS0TnJKP4Dh7YEw
n7j+UAA1P/yYOA5hCDKj494PuyUk2L+zGXWzgyAPPPkdULIUMCUBjVl32hxYhc/L/JiVhGmcgLxY
74P/EIG0yhZfxyXddrUzvM4Ejtiih4dldbqCawoALhiUuj7JyaQX4mWUATv367w1faVt5ARDIR8v
HPFzoKreLceaty3Y/hOXaDuvGWjFwjsxfUsPwLsW1cTY86PxXNA6ZtEEBIrqVHSAZ0Z6/O0uHTrc
CDJZB+ZfJZFLYyYRzwEum775EdIicB7kRR8dkKTsgSLZaMiXg0BGl3iXkrl/vexgXaLTHbaJN1dG
iVCm3iz/CdJLr7C3dt8JenVc5ZSaTNyJ5vuP3ndQtCtDQ06wCftu/8yhS6eUYDQZ1cOv2YiaaJuA
2aEIy3TFxxgAtRCZ0JO74JmPnuazsxGZGVOs8I/GA24ORtzqjjorIfEtKgVwaJDTKdWGaUSq/Mm7
MpSapcuHc1B5RWGbbwm9bZ+UHFlnOAZjjULGx6osNg0fxJObvgVqzPFPRjSiHcMwX19MRMotk1tE
uy8Xx8+FGwaXZ64hGOVyCqMySzMdmDuA6pWuD/T0Op/XqmoE3CauocsuJuphs+ceR5e7/ju8Vgk5
FAQH+Lr+8Yf1TgQ4E4Lydo2boAUELzDIxzrFRTPJhTS2BT7pul1cKynQy1A/+z8Ap+MmSpIacgGi
KVCewi9Db8ZVED2XWe8PajFXE6opWAZmqKobDqs4CVFC7xEi0tH/I7oyjLiQ4YlASYOT5LiPkCej
0v0Lts/JijP3fXyhHvCbusJu8TY9iqGqTl0LRPkxRZaM7XBBziE3nLm5XtBTrMghcRxfDL+9cGBC
C0ghg2li91NymUfYBA43KmS2PWfXcVI1LALUENpCCT7nyvZxFqdR4i4nVDmADj0P+PdghgoyGQuR
H5mq8ujIQzyGnKo9T/HyybzqWjukfYLVe4XBcHF8jsf9eBci77wJwzZKV/vcdxl8a0UZUU8DrZ0n
7aIQGmvQks7nD7NhkLF4MQvbRgxjfjNti5qRkptQlUE5g+A7887ScMEkXPIshPg9m1qfcfD4XrRY
hm/aIbipQcW7DCHnxMvQ/ztf8OhIGapVD9M9azxAY0GV7uM7doUtR6R6TEBaHh1R9Ijd479hICN9
KQQ13272jOzBLZ3eXG1gmlycAWSNo2FayXNLAfaHQM/F9N8yVHoWUaxt+gCXo6zwOqJt1BLYp43L
V1lFFNHRPkxGCrUA5ic0PQtIOD1JJwI9Xzgu1bByfh/YHp7gczSzeW8yjoeRpyjUaIBA34uqzue2
kvQY0FzJPpn9Mmy6c924Zeu1/FmencgQZ701ZwmFSw+NaWKymju0LTxcMgbv2s6L0Qs9akyREM0d
MNWEhVIK7tuvU6y6n4hYf202YQCrqsn6OhWxY7tw/2iFpzkjFAj9Eu2aCpgKLarmAhDbtq8zZnb8
HTzQANF7bkNfZL1m3OMgh20lixWw2rSgHFiDq9R7gTZvKTEpQFROKDcvhgA7c97CZ50WJWmyWD2o
A9nJjWe8wMZGKVYgcg7mcmgh6hJWtD3lsFhCBDoKLyb41Gyv0xNCW+u9QvaErU7ZPtouEuPCHcSW
EU32u8IIhWH3HXJugbERSBP/gIr8kMDpAZKM9Gl3lMKPFc6oQgVfz/Fq3gMG6xcDpJ2jRfB6sFcu
r1v97giNMW95VRYWwGifCDgIZKgatdpkBa7z4iNCoNW7QTa08ogZHUrXbHkOGSahkb5ZnhaCvLI9
B8mcsqUGc3XimVoPqKCseasCSoaprVWrm3kQLh92JdOPVGfI2y5FdR0wLhh/LtqhS1j+QjpPRXYs
1F2td+s4BvyGJdS6G3PiTmfQeghVExCjJDgV1ifS1iWrtSZmUjJ2AD+X41HJw8GgNTocEDq8RaGb
VMOOFkHbe0QtDpjMghb+UfECOi8/eCoqnnIm1oTc6LPopZNe3xxpCNHIF44s12a9HMSm6bpVwdDV
jyzRyqRVYEuQ7E9MakDG1lIXDYc2E0PbBAavWmO8ilVvzEmHlJjCutNZuSMUglEgM5FNvZXstSPt
qRrJpFrNmwqYtL+GN1CWeW+pvPaSg/wPK228frsocHH0bii0oN9sKgdWNJ81Z+pimO6ODOf2K4cz
8BGKSLqmwjRARhCpxKm48vdZnojcgOVPrF3Dp6kMtbFli/zLgsbimMI9Dvz+WYS4OQtctLMFhrWX
saxBiJ4L8B3BpA/dIX/KCtsV+XbMMs3udaOas6D7/vg+IV/OOGs1u8ZKNiq3c0a821Yaui1eKSsV
cEXdQEPzJWOiVEgxjePaKN/P5Nr/ugR3Ck3uJpMBMUN26HttJz5hMFP5xB3nKfeIQLtIXrE7jHvX
Sg0Ujkb95EXbcHukMCjhqaFnMhJQdQsupcA1f+lqI86FUv8BDORzfCRtDwulNdpRvXxvfwf0BLzc
E2oSIV/PP3BRa9+He7QGj06FnSuBuRL1xy0dFnvg9gUcfGcCMj7wQPDJsRtS4r9o7NlU/WV4FFKo
IesKIFzu+wCk7o5svCn1zCyGw5vQG/7ToSqq3R5tifXX+flDjxjExoUoC/p7Ew5Azie1JaXZ73oH
mfVnRpmWzBzyJmtZxI2RT4iRzGP7zhVlmaXamWLDZ8b7pQH6c4gbcRaxXl92qrtKzeWU06qrPsnM
K26CRHCnmUSYsS6SPja5bOQHycEg10vZPHRnhYZGyUpoXteMBHfGOatyyU7xFlyVCAyu91oamsVS
dAEspNUoh0Z4+72yRGSqT8yxuKk4+kzmzDl2wvgIRKk0E4D8kc3UD2pYyHnQveyQ9xpGMh1O64aF
WojdEoC10625C++WQhE0y6zVEqRroQ9bEY8MwTTzpCzSePniaC5xgUUHk/xWrPJwIl5nrH0AqyiN
zOfUHmw5brK7NJsdskvn3UgY1JOOTUAt4uu6SHuyqR3iJGnT4ZCB0KAs0agfQPwOUnmDzQNc3TO7
YcEAlu62Qaib+ojSH7cZ6b/qY6Loowy8q1+G/x31gYKEAQaGC+xUKCxlvBi8MZ7X/NYnIPWjqjQK
/NT/p6LyOGRGc+V1MqKclnNeStEHDO5CvH1n+9vLwGeauTfvcaYDW40cmIL481odNYGHYrCc1xRt
mXiYWbm+F+BYTN15Gh5M3zeFDpbwN5Tsljq+HIMT7Xx7fxflcbPJ2KXOx4APT1TcMcpiVXdk2Lt5
oH9NhX2avEj3KXcuriO2AA7gJ2iEjniaJaKkYdHkE7o4704xDCxFC5i7DXrsBbJk21xKvRKwEP4a
C6uq6EndqfxXsZZUqTY6Vpq2l1CwfroznK0mq2ZimdId4G0wOy2HATpNHiWbTjHYYdeza7V1deXR
Ue79/Cgp/YJ3idOZLybGJpBiNoUvgRcMjsXWGX5Uy+grcLA9iWUtSZktTykamsGuNEBexPEIYzI5
S3bRnWXFhRmXzai88dTZPXehByPYmwGqq+ttWirIbP/CGhJB0n9+AEpdICYk5me0C/FM4TyiYaEm
ZVgyeXlsxPilnMMiBFLtMyQ3IF0n6lugciT3iKyokgDYIcZghN+pbt1/GkuQTELaqH4tXPbzkc9i
7bWSAbqlAQCe5iIxX8Mk30yDR5d5cTwtPB20cUPT8T0sEAQiVdK4bvduKJMd4+ZOOmEJY3MmvLNf
ngIhL+GfEvGQptepziyyHNekX7dYzTYbYhkgK18myihzXCU82GFr3uOwYxsM4WsaNO98LVfb2oah
AqrzTjR44SzinvUt62qkHgeYCwBlvJRvN9lYF+VkzhU2nF7eau1th96Bk4DTfxBOTGDZVAEh1mSz
eIracFthYHqhCSBkK5nf2b+5bU3WBnbIw9bNNmNdcf5o7vdWURWrOEj1DQ5JuHqm5vs4NB9On7Am
bgGSIKH0eq7E14O55GRnjA+JgPDw1A2rZPodJQpO+ax0nBrXEibp4k3fYiFBVAbOVaDAytfZHCE4
6A+QcbUui2cu6kLF69WLuRZdrw9QwNj/7iJTmQY3T9lsvPyD5RhqT6g4GHXhg2FmFZb7QbK2GkOL
pz4yL1n5BzCC3fYN2JdOu4p7eAMvLUdiOuwb0W6vzP5AdGDor08ehBwSY2Pu7ijj/JuphFwqpS3m
6GFSroKVvB7Y6ZN/cOlDBKm4WXXj1mlyJKbrXMR3rjKS32jwwAn8lMJySD+KHf2taX4Ycg0X7xg1
9sg5F83qqkTbtKanuvBVmQLO3Liz211kyAGzmrBkqjLFhidY5R0oQjGvC3GlczK71K2s9J/9eNYd
vs1VrNqhWuwMWC7jHyikGTyq726axBSKLMjTFF/GtGezr7IgZH2cKsd5pFI2N9TnehhNxOcCnXJb
d+Kaclibf8ghBdFcdFAUiK8DG5VmJow/P3W2WVNdfxxtoNO7VjCw7VEOZIluW/im6i45KLnTQi8C
hMc9wT/52ivD8XYu/Txx/3A5IbKrR9bR3I0W3octYsnVTNVblHYcmUeoJpoztdlAxhwsY7wR5psc
qljpzn4Ic5nliTnFQlLXXNtK5/NQWOz0OBhn9fSkzxfV+vSIrgY+C5MX4YarZPanoBnUMPRkJrJf
qhxmT+X93zKXOCBq11+AAzIAJZSWzntA/ACLxEuOUaD0yy0jhZbpOGQYNC8hIvc6mOYsxCaOyQdu
dywbU+JUG3nmPtSb9WPVj2WJ/cw4VhTHbIFl6KLr1f2VTb+mKH2tAkfqEr7qeaMPLcqYhzi7lemN
cOtzkAvFyurUNf8wq7JiT4dlpF3twxlxREtQHVeBUKI2/byi3x2wOv1F5RQy1PRyghiXKLoxWVAY
7jcv1U3RORmVcH8psTOnnUm1a24ls6rRCvJpxY2ljSrTOV2qX8vaDwpEUPBBrcHqFhW8XQ2ZjObN
m5RkcV0QFNnj+UcxOYg52i7/MqlNaVWxner+qti4MthqKjCTbKaauViIBPxGY2xQv6BnR9Fv6bz7
XTTrlMSBh4BSXFU40NE0X2pFda+TnXkXesQvRMcaxhayh5GXVRIH3C0H4fqHQWLJsX+0ln5nJQpW
F1xR6qHH0O7I4vj1OeffBfRYtvWDmWjI75nm231t3zXLjfJuHGEEwZAzjpVS2l2C+UAniGM8Naqv
fa1bgzCRdsHsNmztj8K6dTz7JqedGdwCMDxrUnsfcPaMsvhXnzDwddZHSOmZoFdfIK5LW5mnh6ai
H5JLBaYWTc2bh3dgy1JvqA0OaoDkjE4DpP5HQebx7n/6p2HB95YdgazhZ7GMGWu/M/LKWYk4X2Qi
VZz/hMy7FVAY0YoPQmT6bBWUI5pAgt2kr7oBKCYyUSknPYM86HTbVaZPcLsbmx/s/MxOWMH4mZ2f
olYQl1p9W3IKfiTGJy/9P5KFC3Nc6UdFiXOhYFeTgBJGnSGdgfc4LqEsQtjy0JgjT/Njd99Hn8gZ
JvxaIZOSqah1mC/9KMqB5hsybLoH6zWiRQV6V+Y+oXZnYnyxyf1RhBs+dvEuB99RzrZSCpt0pnwO
+DED5ZOAXw0hFWXci2ItZn52UfGeDC39kJSyTYMeRv2XzBO0Tc7cfYHRbRHhA6d4mn4vZE7g1Jd8
BAqG+X+CoPJPll81PJlHVtt49xPFu3ZZ8F+0nsvIojfw60orWgqVv83YdNS4x+5i/uzAUNkXcZKL
Puu63oM441pJBCLapw9cYCgc2f/TodKnSaLbHmF2O6FadPawhL739vpFvDmqBhQUXHIB5MDmBVsg
Xw5rAisMp2PCD7yy2dsnIto7D/yg8XY14XubZKHL0fbSt8U6N8/+K0w5kDVxnrsQuJAgu2Vm6dPS
H0HPyDQgp7hdusJd74dYuNyFgBFwBeTwxgmRRK+KpcTxXUf4T0+gHqx42e4WnLWqSiekl6saR4Ld
KYvjY56iUmNQGm7ZFqYfg5AIAz7fZf1H5Otaa2x7EiD3+9y/gJKmPAvyvHzhxw+FOw4HFvjfmBnv
GR/Wp86EbZDilG7MEYdij/ec5e/X3CuH4HscuXCIlML/D+wrkir/bga2EjbPqbMvz2quRAAu+JhH
io+KeoRbSzmGTF4ZYWGDtwRBko/5fQ/yQTUIB0yPhcX7Se2cAtERE3c+BKXwmGi+b6yu7UUqsFNe
o3HxFuJESfHXuKG6Ig8MZp2oQOqy6WhigCfRzVGFgMh1c3hotp/8KqUK6iZlontt2Z4sPhqN2Fmn
5sHXhsF6jmwrjsbzEfsWoZn5wWsch+Nbi7gT19NLH9PEXpmqUKfF5cnmlIj0/2eiue+5GIAKc8AN
KVKsZ5o+1JzwognwWU0Q6kHSXGlpjDwy2edIHUzNPmfg7zwLhUCXlUVpBhqXTwwrFfsLiRrlpaPZ
z6OJRDjenH7uM36b8BEv6uxmwQb/BLtkxPD9vfoPxpKBOOmjd9NCyORwk725DaM994LXF3LgY+c2
xerSLfLJZ1pcOSNihHIIx1jTgc+Ztn0au9DDFJVQTzOLB2jD31P8PsLPRyUCKbJOOFCd6mjVQgdl
RqzXiqNB9bZV/J5dF6c125tSxbS4svH+Pr3a7cjbsukOfuTLBaM+9QlzxOixaqOL6SzxUL2cz+Ag
ESiclC770fh/YQG5PBMsj+jOao3vcCdkIUebsFKlUIB/8hRQnDmrI96xtARIeisyrNmZQJ+YBj3U
anLSsefoC8a2cBD5CLeRCUE+8aQG7gxRoNaoPdqRqLsOBwFhIjwDxNuhlH2IOKvONWyRdIjqZ1iC
GFJH2WsiSb2F3bif2Sux+dpqDxFiqJRbk8/M2SW8HX3kiUAMiu7L2xTGrSTMqCdEIwdupIWQf3xZ
AOi5YtuzsDN8RMzi87rI2W/uSa0ZCCVzIOG1vjC8ay7Q3c4HLwnVlG2JYLly9NxEzxM17JJQaJ3m
pIE0S7iWsxTaeojEtNpDnO1H2UuQeXWxeKAe/pLZ1gl+c4e2ic0HajQB4GGHekD+CCRfl5rB13Ra
KyQXJqjRwFrW7a8N/c1192s+uto6XRH+T8NOUFGL0fJsS/MRqNeFeHeTErqGp3S2oQHPBS5/rz4Z
tYSsflbsO3VMUn2kuv6el/x5nM876Efvg7U+z9d357/VTVhmwI7agRdaLYptcNsb3b5rvrctSOC4
8ARg8f2YPGbrNNMKcUspO6k+7kBKaZO2qmYlE4reZxTlKR8s1wVMJ+hscDlCHpCFK2MmIUXtc5kw
vOurWQPw8VP2OnNCLmakCVSghCntOR5+hkZI77Yw80ignrDzAJr/WVfPH1FK1GTi//qphM3nbCxF
xu5NWknhc+Vr83agCo9311U+PVHYTdNf064EX8D7NFvCOaKNisHMDU807/r+OY7bhPnSsJrZZhFB
ceh2kS/4VCcjhujoF2XPPFaxv7VbN/wVhATV0bUW6km5es+ZaSsnlPoJigD3dph1ORcrfKaCWGA4
EpcP3BjMwcTDxjAufxsNok+3dQU/GCgDAn6yEdAxHWYYqDfOYPImDeuw1B/IiulgEXzvyeW7SScw
8U320P/DCJ1xCSd4xNKNCIKO2f4jdclxyGHsx6ByIlexguOxCVrQ3Y8A5x40QQbhjm1pqWgMnXAy
WfaxlaHjMVJi3oUv9PSy6GVr6bKGptsq9ank4KrB6MuY/yKq5G/AloYheGfEZsRsryBz8gjnzuVI
nO2WmsRJpAxKtBZlQcp9wk79ZhCEfNalnMbBWG9dAIz7/tymMr7LZ3gSLMpA2vlLQyuZK/n91eb9
IXZdy8gJ2IAcsR2kDhI7qAjChPmolP9SnSNwDhPbA3pkLjCn/QBqK2M/F4uRDaR0KZwvoOf5qdf8
1yRtmcrHf4VbHMPzxAmECC3/I6kpu609Sz0ZktHPSChjCfFi3ziRPvZcLaJCyOZHQ8ZjRkY+bKqc
YIVFvQGCna5EfDxzj7hOFZ+r5Hq1oHGUjuIoZA8RpAWGW5hmOTRLHyvHfkvTcf7RZ0BJ67E7XywB
EzLjb5PFsqIicE5KNwa12pnmph99PVdI5odsdKWj82SVR4p/ww4jBHIfOTBQW0gKB/4Glll7iCfB
D8w7F++SrxCEjZG+ZPspoTz0BfkYurnuX80SWxatOz5ESuRop1tXqTcPT6TUv7owqJ402IYcXUGm
lOX/z/8EGsrmaoOglPUUcTqkLvKFc3zTOhbTfhRAZJazKQvx225NxIEmNjA7yi8a4trzBm6HFQG1
6yOd0tk0gkIbYnFTyI2ZpPEwI8/O7ADMqjK0qrGLvpIaMLbLetEbVQu0ezVN1jo99CvFQ3vlR9QA
C0/aJYQXSwRDE8dpt1Uu4CmezkvWbFmoOxrkYCL0l7rY9JyiKRrvkrnZBnOcflV4ro5RYQtGZkkJ
+IppilBJ1ueF6tdq4RmRZGi5aLB9/WHoLYGKVLr6t1/fNOQ62AAgVngJr/xhhM+dVLqC+bPHNd5c
4QE0ZhAtENPcWiAbtFOva9OcEqWpDYW3rn4iw/4V43ZKJrqjNOySUyZZshWvW5N+uS5tX9vpnAH7
kZhYCA3F1A5b7RSbabjzwuPgMIVEvAr44r/fqfoDmRDGDz9RUQjm0kD5l6UFfxxQEU7qAMwD5XY5
E+R0owuYNTfi5gP0FHdnZ9sEIizFiX+4JF5m71h9Z95DCy9wZt6xZJ5UNGS6Ku7Hy59QEsINRk7h
DsVnaL3A5aIQtvze9WQDoWvxtP3sm50NrT7270SXYmjTjIin2v9jZibDMJSQuh/zAdqYtrXCZRNZ
rhVUDeStEnlIi1fq2kU6KqYluy7qdklmVxhnnGHW56yFTOg1Kvsrlmk4GhfeHk3JFch2sOoDNCCW
X2tMNUdf2j/W+y9+Fq86Qo9rZCZHRxnj2Sa++okRrf+bX/N06qX3vT899jUehytNGY7YLCc2XoBG
QPq1nc6ADYsEyJB2xYLdTNajhvfCs5YQq9uwQYnYTiCXTHDdZsBdPrAHJ7nCDKLLbSVx6rRG460M
uOeZLKYuLXi32oEkHy28xmo3e5C7mmd0wlSHvXa5bZZJzhjl9gv3bxy0qwOJhldeVBOJaKU4G1nV
l4XxxGal8P5K2Sj4nfqMLqBOK10UOHb4y+awwsOsykPKJmLXh0JgM1jrESN1+DTHldlmFvVjP8yj
t81KzK+4xPEdyAF7BWsRHnvfUlfYnPAPGiKg8GW+vsEfaWeUD+w/jn5arxk6DBevYmpZywJ7OKXJ
cFSoMp/wX9M5IAKYwoCTuzE24jDl6+F6dsYmY0x5Dg1e0UIEpDvxnfjc/Xyb+ttAw48XJ+nzaVa4
68ytxewjkQaDogLPDWYiIsqzclz/dCfuUjCyIKdtGzMVhvKL/R5vPEA0vCSv+cxgEY++6f1L1Leh
9mYR/qLa5VjV69gY9HfSOEejy9u2ye4TAI9j7g8rBgw5/lNu/whvHt34etI7pb1VEQt5Pq8SsNxc
WpdFJNk/K09PrhJHCnyxYXx9I3D2Ud/xSaaHI+IVpeDn40H+d/GLPKZnIt03Zmhxk8hWwcNnHhoX
2r1KHeUjYFPnilbLTXJ2pTZxj90OC8LzMSWgxzEbmIp7TJylF6G3a1qX/zxDXgWJiwRgEVkUx2rp
DQA4Kgx8YmPE66fXC72V9Q1ZXwYFn4TGOo4rSYNfUbZmHFh0adjKibm6Q7x+jUT1XQznZrICPU3A
WLLvKqefIz9ijzqxuPuZ5TwbanbwkULLM31lv/rpj13IAMTSQN4il5GnFEg52xik3EF14hhPcNiB
7xuX3cDTCWJyEtPInckS5H+JCajpC2XIaAO6p4dp+7nAMsxjfYI4gWbO/cjrDqphmpylYAW+QaWB
YiXvLQafcvBoG2LTVpfJRbWEVWaNLfZ++pmsnfWEV4sx4/6Q97APhdcLJV2yFPZGN5dlprhwHyZG
bcmX7A1Fd6wgo83XtriHxCgXyZu5U+fXQR3xFg8QEQ75oK0lJgvD7xmucjhwZKJkYOVDgJyJH83K
dJ+odUGpvIdhNIIgLeHk0IWehDT/FepWlCvM3cJuaynuBa7Pj5LbGSOhiWLkw8X4cTTFAo/BMiuO
fs1c1gC6NfNHKOfJtTsHn/dWw2wyC97S67JZ8WcwgjW2Yjvc7yclW4Vh22iWa42iCmwhdTUt2qua
LrdN22x/syqxdAUhw2CaF8HuBQInDZbQCmV2Q2Fl85fpcO9bJRyxmMF1pqV1VCeQsZBdSjeTX56s
pdkAJtzgD3VL6Da4VOXPgwmae1LdZLTsYolnMsa0tjbbVSvZPZ6FYFGT+YSXMUPvOQvKnksFJNBX
YzhGmQLN3OFHbEHTAGG7EMpl0OL48z0G5XesdodDHw2pi4hvGEuCatST68+aqsoh3ZvBD/CyPXCt
NOTY7Fx0nntxWeM5SK0pgPBagf0Gv2yfv9h8QRmp5IjeMnULaPq2wEOlxUBpytib5kBzUw4TgIwu
YoyCTro50T0t1UFg/ixiheVREzLnwaCvXobytXAmAUthsBZoVed/OQzCuY7id4r2cAr+5a5Vmbsj
A6P25HPUJRAyVv7H3xPvDuCuuorjVShlYu9EknoxnGrtXYpdWUbFvlbcU/9Bm569RnRz/KwgJUHG
UJDsMYP+eWx/TRWDnbTlMi8MYolrhcQCwQr04G+FWYPIEUYsNdjMCh/oiFxK08QTD6uN7dxGNDIb
U/fCKVkl+5URZR6ZteuU2pXdOvuLNxyPUude7jyi0GjitZ9sXKOY65XgSgUBvMiSB4QOoTIxFGOQ
kKng/Vk/SZ8h0U5LO7SwHAEZJqdSkJT1h3tyNzBos0dQaNAJDitEI8SRlwfEy1rGkJ4Ljc5LkYqX
G5ivInQT9fFpeJiiKwQumbuPCrmOc174ciaSLZToxMrgGBVDquPhAgj7emwnTtbUzjH3ybpOfMYE
SVB9cFFESRLJOiJw7qWx4HJ5Hf8s8jGnWCvL/Hp03Zc04N9PE2WeIsoVFk3vhm4YOfQ2nqsqNxfo
VVba4ORVctQ8X+crkuzEJkI+Zq7YJ1ZWqf5oqNDyK4kDGKmPMtug2eVAXrOg4Qhnt0iwXGBeXKCu
cz0L1epeVLiAWjh5nfiRxUJ2fCv+BPkjUaJk3C4m21Yy/7d534wt+vmDbdFEwlu+weBYJNRpDN+3
CAnd3pCjYI7Hg/T+ezaGfiLq5teeZO5aN2yoa9jkYZSEojYy33gMGdIPCjGf4v+7vNWAl9RfPqjs
2cH/o6scLVSCA91UFdh0+1WqA/PR33h9t+NFjrCnUwI33/nJH/XzItU6IRw5cVofPrQSsgKc4+/v
/WnNezxHue52sOt7T8jnz74o4kHBXw8mrovkw9R++rW9HMQPkuxiAbysXml8ilPfh/J0pDElO0zW
pHYoSH7Fm5VrvR0Svz02dUnjlVLkg2juYW88puBZV6PjEw5hG48bStGpW4uM+ff30yO29v/XLwOr
Y3sMEy1IoKKrsQLI17Zy5Iqx87qRhBgmv6/RrLBMt9eTgd33bf0wW3rfwVM1GK31N1bI5ClOF1Q0
lvv//fMm2jXiRC/XCUvJv+DmLCut+AZnoh9OkIyvQA8LsJAO+YcZ1rSODRYzVxxfGSrSyvIPIWcZ
hdZut8ykrLhT4BJL6x3EjpPJqvyKlGMO38TX9pqcDGYcoDnTEzCVoLsBaUbC+XICuPSQNDEj+uYs
cX8G5C08L7lROF0M4kk1i8IMg12IPMGJLaAUm2pr/FE0AqP0pTDJRPdVXU15uII5wqaTY2Fxksko
wwH7gMYLsb0BRLIAldFueDlJDwK9wy52bezanxiXMVKcKT12P15uKphjxwJ+RF2Q6b6WGp7cHIcL
9Xnsnu1+8ZRorrXbn/Phcy8eZDWIZC4auQJx2H2sCLUcsumzRv6SsP15cF7BIBp3VB1IhWuD4D7+
K83Omegs8y17+WdAs8oLNvNLhnmGb5yupoklwKPB5kBoJmAkL3iToh1QiywfHkv/5rP48oINNsGb
i2L+ghg+HYlOPHVGJ1+m7LCbb+wrdSndgOnc03/yZRER4KA3aibiOov9HolW1NWWaicO6fpS24Kh
ysMiAckKBiwPbY31crYuuuDyJqxTadCx1qjrjNDq7YvggBMRwjRxhhNcWhNePHKXxkMU9VOobp8x
aTUep39+ggC536/doFsdQ/WmVPaO8fRmI7ZN45EOD+fCZFM95cwKcvJpU+R3Y0f1j5alQrkHYGTN
onheGDOoIdWzbGs7rfq14G49ioITxNtJU9QWDF1CvbGUFqwfRR0dt/QqO+bzKE4EmsuPmzV+ldcN
LZigffiCzVqqy9BenB5yw+GFZU4jqUTq/RhDeQGJivhlN2QIl+/hUu9PxvEH6etDs+gRGJwBnCyX
yk1ZqeSnjZ8W+aMtz2keyWtkxR5Jo4Fu8hBoZR+U7Jhmngvo6dDwvxdSoUk1NYez+fUpXb0vaQe7
0X2K25D8K3ZzlsjWlrKkqhUf+3WZjMZ/8EraTWd5Y+GJMv+kB2b88MJEL3YXfx4fWP4n51W/JIBI
shLO9E5FZsuMHdSI+AdOfAJWiHI7ez0taqeEYWHrqY8vdL98xkBzdupvXK8ve2+MiCLBplIGD9GV
7IUH62vy3EWl76T7diDeJmDgPxv9GY/0ROs9+SQG20xSSB1wmuplSc35SHxMmAZHKI2VBazBjLaV
V1oe+wsncu/ILiJFTWXr6awRfLUdI5UFryUNZSToXr1/D+vo+MuNqk18v9q1RH87kK5xqYdPqsgK
g5v9qTQ8vPvRiGzmsVBj2G/cUxDFOGxC7njZi8ikVSPC/x12VBPv+BJIlUsMHbAmnjqloy+FBbcb
/9PB4UEGNnQV6RUU10XWKKzZAi2oIkMUpr5X+ZOk19fh8vrcvGZXK7BswrO0cKE6JF3xUUEPm56U
bRKViKnFiS+e/BpCjWMi5yA9X8qkP1PEWnmZKlrvPPOG9dvklFsKU0P1mlAJfNVhawL9F799BVX/
ftqgI30RyDgWc67dXzwCLOscV+sA00Mlpx2LQJOwxsXsYvySx+CIuivrU5a0Zpx56HsZxUyhuVt/
z8KYebbzTDzv4uh6OkpZ83N2ui/sjL0Atc/pNAaLPrw0ViLXfM8P9YLeUmhhAZNKwU1MBLkPtzbK
i7sgIHjKSYo091lv7Pnql7NpXSIBZ+1c5POGLZJb1df7YeoIdssmd/8IXhE+k4fV1DofbR7CY+/w
57yObSfUQitzGyaImxCrO7Pw9ieQtw3XqSToRKQIzxt9L6TohALc+paSaexAAw5gQZq69Dp2fjZW
TLsbzW7B/wDcjhnHJoNdYVY9IzoPmHQC4tzMHJjG6A7FSyVV60YOcHbQY2D2iULRLECvnTg9I1Ba
5DFoa98QtSxq1eKUFJjTNYNMZBlP2ivKmMKobOQZMVmEXRsXEruq9mVcMMcoziEZkPFrNQpX7D0t
1iYuQYRZ2aWGjvfMXo8b+5HvVfxzZz7n0pvq/F0Qiy5NNxjQFjZ597jAHNtD2XiMlTOWkLT6iHKI
E131VQpNPMpaJ/VNU5wpTY9pyBnANxKlg+pce/rJVW5Hn56yhbpQDMcJb+QiQMeMiwmSlJBGCv3Y
wv7rGzraSWg+BsbZz/V8AVwayfcPCS5blzZfZj1dTdfEI+SiiaQP8pAKJLq6tFtP8yxq41F0aalX
A9rgMb11fkwnizI7TUnJBb1aT/Mn3ffvOoe14/2F8iDXqdBNEuRUvPfm6pGUdM4SAM8ob1phiGUu
bYVYamnkh6igi5ePRTSPeqJ/U6m8LLiPJzLYVA4d7cMxch6cerwXwkXdSrNa10hMUtpnG/6vn8JD
dWXd8A5JqVvPVRT20bu07RW033Fo5ILB4aQZ8MXEEkaWcukbdVNl3EoRdcGRFJoddQPX2zoORuUh
dXOm/JxMEX6vJhLu8GXsDxW4+zZWFCQibN5xeW+2MoQ0cSeO4muvWo8UDd5teLaFmfOBU/msYJG9
DrUJsbFXVz8STpLPJ/5zl0b/zDvav3aRSu8mSAI0j/WeEAOFEtRvTO5bs3MSQV76qGbf4RlLZ7TO
KmQe6FM7khvMddNoBACCwf3eB8dHkYmKdheWuq+Z28FSKksgVWMtAkSUzYsGbCa4PVRVvTBi1R+h
1/cyr+ZHyOGiYx6C/o3AW1EvD1AIFnToazyrQnmi9yq4ejzkPp7w14u0urx0/h+3HciHYLaH5sRY
knAVrJHQCOQymKu2fLhlXwxA3If4TCWm0YqGQHyoDAdIG9qmiTPH5XLNmPmk2ZOSutLWzlzia4dO
XTReeMaMq3vtkmNuttlOQN1z1t8SK+etELpa0j5FcrxACnbOq7kDQy9K+Ra2sTM0dnzhhQ3axD9Z
VAtG8dx6p5Y5IhH5Wma3696cWw6Z1zVhj2Iojt2HJxvxQ8UVJkIvOQQ7ho407UgzwbP4fVKN8O+w
hn5VaPkNOkd1T6UpRLxLBZd5W6F0R9qqv7KlL7djfCzm4WRPx274iFkFMLAi9HAXt4tgQ22AtOet
VBtgZmMcV7GHsrNJ4URaT3RjDGKa0TfewO3sDNy1nH31YZlsJEgeCgIicrKmZpdM1LtYq2GPLDkV
JX+x/4UXAPsS4R3DUsnCC6tDhDtNAEmvS57CikZ0s4J07dEqWPzzTmhR1p/zWMTem8lAcCvMwf9g
EnPViT73D5amZaGTAzqsDEpTayGBzE0Ff5jLXWgLHQxFEsvS27fD8SUb1g6RwbNJYNtRIS77WWv9
iK6GdJkZ1buSuZAlfd73GdKled4f5UVEH1mknN/junHC3NkYZwzTVQtZH76gxrKF3jYaLuwyNwT/
0HwhlLMFYWyADajhP5Lg51fzrubaZ3v7ILjYiSRt+P3zVsdvSiaQKF/mGfnP8H+ngZSX6DDUOXM1
ZCPZAHakA+NSDcv5IPS1ido/HKsWu/GyQAu67T4/BIXXXMU1CamGa/1enOsfOsSYE0ZeQ29S3H23
/C7nr2gghBH7MXBiGkQT0Y+ESRppfEe5BoZWQNRyBhYg2Do3dd+CqelFQ7OWt1xu12foJgWlHLTw
4KcMbp2O4Mbhjdp71BdVIqNA4qpxtiZHW+nxy1x1gZc6eoitEDFCFd0y3KRjsKcD3tRsEVtdC8MP
Sx3ukyZI8LCSgde/O8YiR/BNQ0iYkknIhbFrehnAnmknpisybAVubnSn15N28bntj9ByC3LcHy3P
4iwPhAEDVgZkTvJ+tbnJpzdc4DYxcmyCnzCVnOoEagBBhwIec2G3LNbBS/gFw6JIXeXs6aT45+b5
WeeaFrr/vIkmjGL7VJNuR8n3lc5nnM6jEDKpgOR4Z/nG/mBq3pj2D6IC/r/dXC1V75eCsPTVlwTa
QVzc8GL9e0M2ZkohiR0HL4WUzWR+Pq7HTQpE5Rds7bUzymYxls/rRTz6QriEFPHjRa8LJHJt44ua
ETSB6YLJ6afItIYYRo1W+nOJSC+/Ao0dUJEBUNFycpTUsH1QXwgeVi085Pip3NnhibqXnSwU4iMT
3HiOs06mlh5mKwR4tg0kS3BAkezBlxkBPce55o2lToNCHRvmXEsQ9l15E290iykH/AO7PLvlUVSc
GPXzxdCFyunwAMXJMBa0LaQXKds9cYGQtJo1gf/73iH6bhrzOo0aSN+0g2t8+SGR8Es/XwKrYeD7
pDL1lX5wJBu6RuSgfQPc8YnPpb2AfgiWr3b+/TLI6980ladYjalUCW2NAD0RuGEZfzOGwuOFn090
RutLuOBWLNJRmw0ZpgN5+SpHDF2BZXoodtOkt3uqMU9HAE9QMbUELBr25V3uLANZFJG1eUJtGWms
jNyjB2syBX0BqiTRZSc7A9Y6sryCC10ehLq6Fmq+aD7pYFW+xpXDavgva7n6qSviECNqcO8gbSh4
fnqyOX1niDnVXu5raeiD4UUJBdgdB13BuMKatiGveEAfMjXQ8F83Q1/1HKoe+FOtgO8HD3U4fhuD
RXAtqUcWoyYnidhLlML5//AmdKpvopNIUvoBQySjmDR92TiaTUY9atYPqHheU2y4szWNGZIPszhV
Aw6faJ1oPL/kHVd/0AY5NL0FcvX4OpzS4x53YEaorK55VswRC6dBsECMt3H1bZnjKz41G6tZ4yqy
tq8Fi0Fs7zlMVfCKJK9dIwejXBbnDKey/fd5Z+e4j1bGKU0rV8aZ1ff4PMYkxzVyQ5CgQrIBphmx
ZjXVaUXTZnMWR7FxdRZwAL03UGFQifMxfV4NeGHO9V6bFuM1pQiQm53ohs+Lr0XTAJjnnNxeIujn
ZchE24w6o4BO37PfG2L2q6d0ujIOP/1Z1/aTimiHQo9ZZXfn8V83BqPbZk9hHT5HXhlANHlbHWBw
0RHPbZWz6BAxE+Wg/rCmda9Gb000MF+3SE/VJQfBBn8I/BJ4L1t2cTNx4KvbGaA6Urr1fQKpBFl7
JgxmlBdYqE8Pz+pkyZXW7fYDoN1NNXxIDR6rI+sM+ZaEjBedmB/Gc2Gr1mtaDiGW8ArTzAsPX6/k
MfdkThHT8W2ys2cStuL0DnKmpV+AT6pqNaIAIHD7ylB08SK+M+rF/Ankhs5hFwq0vNspzNVf90Jp
4KssmqUCkCHMRvK1ZZklg2MlPizM44CNNNodzbiWN7bDUlYIjukPDrfloZm8dgK2yC1LPT76d6Ui
hp58DNr0d/WEZGVH5y0hxmdOOxHYLxUgsQeOmGvMJ5AhMaf6Ztlu6uPtVjsCpzwEb+u1NtIa3WJy
n2gxnn+pt53CsBsOXRSmOvr+jjHMPuTH56GC6sFtV5ZUvh5FLPnJeUoWQZrQspXPJRQ1xmpm3VXS
lb3SI5JWYJRem3YGTPLKZyjcr7JyOAa2gbeCbeKARDZYn3wDQOK8QYw+sE07O7MMCD5s2jrVLS2S
VybAmXDF0QmxitLq0op4dKlIamRwn8YnWXov3WlN87CyNCrgOfG5H2tFPr2oEworH8is/17ZETw4
nRiky0doDQ25ww6w6+rhSKsK6E3pgNWKLkzXImkxuvNJxtw20p8T2vlkemqemxkqR6Sns96W+AoY
PikSE9NS97Z6IsNPKVQ6iwbCkrbVfp6IvaHDk5kaDcVbtWkZHLLSeJnKTDA8DnGPwXB8KQoUZLMo
ofWY8tlVKCA+QKxmBdrL8tRuRWLthibpZDaZfbmkEf8Moxdbqr2tfOHpCqhSfcHhNY97y/KOntEQ
yvnI0SDHf8QCxg7sxps1wZsxNzwT71EivNlC4P+dHRcWoEc5pFAd/MfHu3RBvV0Zq+K1vPHMzhVw
WLsyFYC/wgKaZdjWWpOpl9hvRi2yPekDK+k9bXmbIatZnfW5b47V240UtiHsTIQz1uv1WjWp6xkk
xKhkQ3qwEAZxrJuSd+uYbYFLKBdmS5MN6xchH4WXMthmJRuX6AEb5MgHcF6iDJm8z7VrkW8qaoyo
u/HQtH5LstKqE1nD5OoqTokJqUJjyUmuJk3qqeQ5n3iDx6RwHYvQQ+aQ1S3o0IF8HWhbYojhtxEJ
wFjxq7m65or54hlyAFtdBctU1mr8spjJKg/FCqMwnyrZhMvBJlU/MGaI2JYJ65g3Kjas9vtAKui2
Rz5MARMpV8DE14QJjsTN2OeVDdF3dLbLBhO0g6TwK9aioeBPT9LOl2bgHLjLykPjJ8ymPyx0nEjx
FVkP/ZCr8xiQaWQQkBO3cMXya6CQsKZNkG9AJ9rwxRItpzPzblIIEAL/FXnqml+SohMJrtXzveXY
hbKtTaNx4AligI7PkUyapyPl7FCJnFkC2/NdGYi9GnkUxR0m6FEqPoswxwOChJrRp8lTGZ3Qrns6
It16WzlE0pzh+530zw2xWuFWqo3De9XZYo2lx22xRFxqFx/s6IrND7GJZgviG7paypR+MNKZ4/Iu
tqcxGrq2P85ArlWdPZVvsfjc5lFRm6DdGUyotqyGvqofbnhlocTii5qjbOn0tUeH2JuPhd71SICr
14DkCxDh6l2PUI9KqG1lV5e7E+ma41QOecU89zSAgNL34CvG2z88vP7wGDtLn2+1kUBZzCxkaW3h
pDUL1YMlTP+mPOYKwNCNY9PTPzVj6AojhQQ0Ro/wnRvdWS25aRfzZcZ0ASay0e2x1pHM05ulXhZt
69C1MaMuET/cBk+fJ/FCBXt8KC6dfK1TWr5ivBSbgFdASdzcPG9HLIAD3HOl6GxcKI4LfVPNl2f1
TNLAEoU82wGmL4W5jBuxmozsap9QFciZkOjGgqPoxzmHAoYQ6SpjgEhQnPEV9+w2LWSgBmzvTjw1
KEoxIL25Wn3qZjGXt4qjIA72m4OIKFXMK07QUP1vVsINSVCMNzoKVDM8A6pZyPRUkqk23HtRSMRs
Q98pJUEjhErUV8Yz3OhQv62YGxCsP/UlI99kTUadsJJBcSaYeltJuNK/w1PYsS+wuK/EOyV4C5x/
jNiO8mQee92On19f/D4U+qb7ejw/itT0ZWfYr3evdnkQvcvD6eJHlodnj9/07nM1L4zwRQ9ObEE9
bVHvfT572ot9YDi7IpQ4m2JqNfsPrKxf2oa/N59ieaOsBOHTIFGGq6UCe2lEyF+mMcj00xqIXSmg
pOiH+ZA9uW60UFXS6HugDGt+xROX2nYiCaZJlhYUrcp8bbXUzaMR+ozvmY02FZetmyKf2PQqrL3M
HmJADPAPwbVeSxNvy1/oSOhUZVCwflLH0hn5Y/3nPuNl9oFo2RMVJ1aoG3IIo2OhvtYRLlcz7bKu
zycL/DdJseOHQKyOHVeeUhQHZcitFl5P1eifN95GdDye597TK46LJfqZN1My8mGrJ1y14nRpAtYI
8VPFP1KiuVD7ou02O22SOQwqj5VqGffpVgJa2Ej44wCDRJwFxh0d4SVWOHOSG3ca6AlpS75ALir9
Z9yqdKKAAUMVaxKwjEBSnE8UsTSaA4mcFYl8QW246VpS+OGwnkIprEy9SlZ4EcEqV1FjHECD1P1B
VV8gUchSxjJawvikkX2CCSa77H8wXOd2aPwYbVOF2vn0rWsUc3vjYiJYmPS02hnUtRuEJGfV03lN
B/+qONYHsa9OGAAueEJxYoetN/lYbHdzrq4AB+yYDUTKUJCKVNnnt4q0V3KfCAIKeHna6CfaiAOE
f+GCA5zFmpyqmKwCapjnkfpD70ldHcPNhKz1LRzpTg0AvoHMqF3E5S2AnS2EkeuCSDt/EoRdCZ9z
Re1G6GiHh9GswJSWzKy/lP7HUgR7OW9PPomWaePtVQDqIJDCPcvWYhP19kGUWQ81frwFry5zrri1
7pSwzsXq3CY7qNsLGsaLkkDQSIoB6vwf7Z+FXuegH8BF4fqVvRYlVVo4DMhh3ByO7jyMqXcPVF06
azkz8tAZ3cwi4tKi8yaTHLnluIVwIQ54TChSjb7oMEs04ARZB0LP/yDofo5Bs0ROCI/EdUx9mP+U
0kb5OqAEPBjqZEV1z2ddqfJHMQFfFKQzat8KiG/70CblJ5igSwMIg1kmnCbGlHrgTroEQdB82CZ1
96R6y3gZ+eQpuMZYzLK1qCoTsX2jsl3v/0kwpyXefLRu3gg7qX1If9FZfhsah73ZkFnYh3SV2SGl
mJToNu7fCO6cobmnTIVM6Giy+GelJS/qIX5p2r7R8Z71+6RYeJf7VBKO2e8g5OJqb2J9Cm9Pd8lD
JMgVKndpwmpg6cfVWF5d+XyQyem4Vix5ty0BA9cCM8dXtaXrdM07ZM/fISsAnjfDxMV6TWyGyfr3
JhWocavvKN0dLRPB6w9UY2cXUPc8huhfiLKSUUI0BeUSgXZB2nnczA7yBzQV3cB3JtYGjrirAEIf
6y+n4yFvf4nwLmjWl3g9/3Qqy1g5yjj2XwHQsoDG66kowfXgaDb8WvOSqnoN5hGnh3mrPzKjTyLn
a2QQEiFSZbf+k2/5JqrMJ8UyAAwkOb+r8t7f/sigBK0VXCje3XM6h+pYvrHyH7Xd05OJ9b6tTXoV
DGJeUvBZw5zHOh03L80lze6euVswygbFi8JFsrKF5uHIexJ5h1eJGL5CjxG4PHH7qYB/R9xjsByX
DPqoC6W4f+2e+8+YqmArbHh3EFaL5A8nz4hULcT9AJ3zHGKCQUgepnYhojygYyMsbuKWx60YVlgB
bIZ4ghrQzZ9yOEjzlAoY8TAS6IvSN43v+rcORmvA4O/vefO+IwUiBhYpng95p094MzQq4ug6BDrP
QQXQ2xLX0QNZvaDDA3kVgAVfyBh9EEZMnvtXDjjMtiyiF79W3LCDaJuDuBkMI/h1PS4M/EBIHL1I
H4qfNltc5jdMCx82lFkEySZi/dHPgURd08w8Z4X6KsIBP7xv5FK47WewrM3XBAGmhVHeYxuiuX9Q
kruqEoWZdjp10VzPqkSUVal6jNPYmNgRs9LI+Qei07xNLotCdhyY7OPUkXiAUA+KsZq0gO/DRk+2
BKuO+DDtggOYu9EPCPZSp4TYfdTl96SuFRfCKJ3PRe/23RdRRxE45nB4P4FqVGa/fzwopwy4ECzx
YkF5gmTDxw9WRYADvNZKlnkuksZ02uIV2tp6yQMBYytGcuS40tM+EZUaz8XgejKcDiYzTE7W+9f5
19ueri3T2DyOOj3KOC0WZAvdJ/yIjqJV7WvuZnRWCGlFjtzIvAa1TO7zGh4J7bqJqv/PvCuYMmye
9WHOFGyzLIFGPFw2JM9eS/DB8uRX98Syvd13/XIB9S0DVkNQkqyiQztRvxIaGSKbhFM9x5W07Nk7
806M8KHUNpZwk4o4yTdRAVH3ieAOxYZMvVbBOwFYpRjqxiVMS6N3xKN538ervDyULHGce8EqVkOX
wt6dj9aI3Tz6P/k8UH9iHNG7QgWLrj8wAmf4airAP4F5VrPUp3VKNz/eMI1kLCIj6trebcZPcejg
r7DtiLAtjher8u4quZCr77RRgwfE/2EUwXtwaiV4xn6X1VHrNuQRw6iqPvK99tQsfPzQHUi8dNQr
hKMBjv8xtjxRDvCcQp0h0RtByXTZNwynb6Wn9bz1gfcDQbaDwc08J2B/4EVMAl4vdhtghtP9+pWk
KGO18RSSexbwKZiJXuEsA1Z9nWbsNeRfx3rIpjUB5kN1f4SOtySELghD7pMeBqxzQUReK5CFmIIz
7ei3f6RpA5tee57iDnbPX4luBe4CAEg1782U9bmbOW3TnAK62bS4XXLgQKQ/QMfjwTs8lM9zVF4y
ceoQ7WPY64Td4ntw1kIY+BxBcxj7SiTxGGl7JBWhTZaQrHC/oSSVlgiXMR3r7aMaw0VnC96p8evq
5Qsw6d/xK/Ymc8whFx/hu3WLUdCvERrsXuiq6jK4yJKpn9NznDTqR+d0TzQtl7hSMwvBZIBTNTLp
VJnKmGjQyxc4hHAVnM+JR0RD4zGorHgncg5q44StHsnP8K0+5N1/ZZ2zXq+NOlXi+uvS2moEaeFl
wJUO5LGH46T0aRQkNrCEe15a8ijGKkThY6t853s6wr48LTnROIx5R4tX8j3WD3iSsQCt6AeLEcvJ
NVT3eVXaU6CSoj3k8ZEMGtlB1rSE3va0WUQ37QQA1/UdLRmMvsaIEISFXZyDXebGd9Y3Kha2G8BV
9Ue6EHMP5hrw4+2aXW8RQWVr/NmLo/PLwRg+y6oLYKStSxPRIFxhBmIb6Vopw1O2N7vH2XiJdsCe
JuxYy0y0dR3aksrcMOb8U29C9AAMDXz6Cr9UKysdgpe8+y1hZOTgBC4Lbe0EZy6IaoWgQ08PGyne
XenKO3Y/12Urv4sOyvp1KrWPJlUUAsUZ3RNvGuMxv8k7vdYSebQJi9Y5wQ04HoUgeE+XhqWrOlFP
fYyctwqIdLH8P2iTALo7zOxjp/IISQ/9XwPAOMNraa0UcPyGCGeZMkVzNg0mXH/OUabasyyF/Mo6
eTgY6Nt7zQyqpLbNvB5F9Y6cBcPx6kl9QxM19qFV7vBJXmjNo6Jx1gsRET5KCKymjpS0753EIlO5
IP+eM8ZFYhS2L1NbthwmRsgthFIgOv2Tr8ZrWiYomex52LDsOLxKk0LwKp6eVKsubbHVoLdiFUWM
hPJ5rTw+0T1Ob4cwj331L2a5DCaVnhccopeT4UQDcqY2wryMVTYohi9yX/enkIjr7CPuWA38CnAa
e73+hIjf22Tdfn1t3HlCjhkPoFi/PxMkBmgfYL9+0VRFxsuB/TpqsdzUl8RQ4U4eaZzYgBMI0Tim
BEJFUxJoZXAJ+6LwD1nuHrneNfZSxA8yw8sWyfsc+8lCLKVFvmnDNxtbpUis35h5sh0YlCdKcOxl
IS4I78TIh1ly9UFRBI6lfPzBmf4UyEzrlaU6RNnfCs149MdpzZrWwhjWLTrLQ1KI0h9frVrc55cm
dswCgmZF57PAQPlxcy63R2gy+/wacdr61kyMV9HhN1oqy0RPEAbpwGeGpRkqEyApkMaG697WElkd
qDZZ41HKTJThVSylHBredZtMCqXWzztqpKoy0eGumlHygj9dDTCJzT7Sa03c1GofmYPExxHcaPnr
B/48uWOc4BQvMx0UyWoU/A8YDTpzomGK7dk5EAFe+JBscF/EHlG2LUWV8Z8+oe2nBWSNQKPrCnTc
3POfPeCMdxs2RKamiYh8o9LRi3mrsZPX4A73PeUOWhxx9UeQSYsVrK7f0GVd5pGZZeOZdnVtuok9
hXpZPZ6JTKL+x5oYfLQgZeKK4XEaCtE5zZITqGhd25WQzfOoU4hD/ML65CZDqjeFPNA35EekJ+Tm
pHa2h4GOUcnI8pqKh/7hoa+8eD7IjUlh+5qmDVnPwjFK2XYxOFuJ/raKXn5rfg8GvZRvLOdb+Kby
WF36VFr8eAw+L1Awc/J3WyMkz2VCXN744HPfrM7VZVJtew7RGTVJDr4pul3P/ONqCRBtJfrA80CE
/UMXy49XCNzjV97+F7/jIpu1V/09iz5txrmVqG4KKXMvb99xwrG2hpjvNRoNReJh+3qHAlWseTbB
+pS7BuigSoSsBrKFvS04rCp3V38SzK++x5jtqWPmQiRH5jg5tp0yaF06LXSGp6qnjOXeQOeZEAw8
3wKQDl7By8ovtGmz81iz3QZI1fvXstDyNRbY+CraaHgH+UzK26oJ4j7+wEChXVRnue5R3SqBOxz4
+mOPc/T65sGooJDEfBga8WQLgY0PLr8Sy8m2cWwCEW9V6XmMdIXb4YpBqg0GuQN7H+04C1ZYjqHL
bO3niULoo5tocLkRPBbfrwuUri7UR0uC9E5pH3ofv3nOtdlZl2Te2PdY4qAB0Ve/mMdQZ5diR7tA
na2/HGSbTpJGqVENo+yYwSTVoRepthb8IckmD2kiCF6Hqxhp63guiDVr/1gwb1xguxFZQxvouRY9
S+z0Tcv1md8SDkBc/o8yp/f9O/IlQ91bsOL4dsztEI0ktNF3C4G1ziOjEdodpd6N8+lRfSP7jIbk
EbByi5lV1xZq6PSUHDb4o3lCGdC6XSnG+Qd/anBxVGJgYKIhhoEFe/4Xlc92FJxF1AbGkZNX24Qc
MnU0Q6cQQqWM7slO+HjNuOQplZb5bJHN3l6yFHCOQ7hF8BjqcPgpZL/04BjI91RgJV1rLXLohnHZ
SpFSM++s/WGXInpjiimC9Z62JWY6OfV2ueLsjdNaETGt6hYucoz0Lpj21zOesJJqCGne1a9z8zTb
XK7IhQe5V1eu96dn1f8BXpFYpR+DWYOR2bTH2jWcwfOCWTy8H6bNtr25Q7iiSQuXE1ESiom0vMel
fvxvNVtC3vW8FKLWQftNKuN8PBTlEGI25R0C+wAlrt2pLczeFxESWQ45FzZqGX1H+HeWj9ZkIWpd
4M8HUwCFB6cBG0lOQcn/DhZM4K2Y4mPNZTgP1Zmc/FDE+x6QJqZU7RudEwcBYtYW6fsvHHFQgYfY
DQcbY/1NJAwRd5gsGQ2nYt1U7ceDN/g9fEZuOLlfsaEMmI6BNzWT3ClTnDyNbkK6EZuciq1uo838
MiWh+IF/+ih5FNgKL0zFkRhHaq8QC4tmrTTnllh6KDvcWqoXABj/8HfQAKWyqnoQ88p3V2JT14zR
XPRjDCANwr2hcfLgmmHa2zZey0utNbmSXG4gRIjLZlCjzUVHuLVQHp3x9n1DWH/pGx69xZS4mf8T
wVWScn/8frkVFxsTzx2sQsnfiMiMd4JUArx/xcV5M7eYihTcKcAcEd8w7uHJcscGB7Ly/XJWoAFm
uzcSJM8ulEG1UZ3tCrlng9AZsCBG2zBLZUmSi4JHIOBRRhPHWBpAhK3Apy5+P4OFgD6QS2hcZ3vx
Pgly4Xt7g2WoRfzwBsAa9OU/5ScQbDtKa3GcBUT52W7l5xljDGL4CJBXnu7q4B5n12czpHPa5ucB
/HuaMkPVbTt5CAsplLllqaJlHq9iztsHDB4fb/J5v0U+VHeFpM0om++czzpefGFIGULpLBhkeVC8
Xss057KpJRIOZgK/ifbkdP1F2Q+GGvTVrqcFgCxHw1IS2900cRg1BWBZBQxUoA0XyIwhQynwZNCj
N1kYqKxA3f1wGeyw+NcPRPsmWtqcxhRJRryAeF7UldK5f64sIsyEt5WwHMj9TwKQJqC7UsWY30C0
Qbcjn36DOpvDfMrPWJuY5BV4XuK4kuknzdfC1Hm527XXDRNCL8j2QbnxecqLw0g5SO6Qo/X90SJ0
G/8Lj9brJl23r/Z6fqWr0Uz4egb1EPR3qqy0KXbbRUpgC87NptfMhI4U1Wq+j69vHacYtsXdnKgd
o8gryBfhUX3c83cTZxOxpbZB2HjF3lUnoexZcxo4y05QNptvnPYa0XHCbYMlMpgl0CFzj4tkwgbH
b+k1dmMEpZCqZJBivu6PS7DKgd5LZY6MgTBI5E0+wA56AGz5NE9GIuwpRsH6m0qA6rLTNy0AREvw
YufgbkOOV5UH2sytI5SOyNdo1UG7u530FESDasz392Rz94mol2cS5174s8vJWQh6tuXKndmHjEP5
1WKQPx8C6PmbgftK2tnokK9mAuuh5xVuOksdRf1o/HOwBEvS+NZHJHPqOpN8eg/WadbVuCsMpGqf
iVe7EX6BekNrs0/iCD62X472J/LfU3KxwUlna4b3MGDxN4mfkSH78A0KqC6KACMfRBO7JWvuVEpa
CMhN0JhNh5TwAJ0VHo85dAaaaaqzTrmfZQxs3WKXEi1DjduMpqzdd/1UxQXEvlmj8MRBG34L/nDt
VzYEZFI3UjixJw7n2tzi+C9L8Qad0ArW+JiIwa+ugtUI8if1QScKTy40CXlGFX6J8LEacpw8mTeA
lQaQ26GGmoEu8rmYucEaP5KVBRD3JodmoxQNKQ7UaO8S8QMF+U0BDa/nfW54TKOE3G97JKRQM5Rt
4Vytr+O4GcEi7gaKu6GnoQn8rUy4BnT3sWQ9wCO9H2PYA1a71zRVnzBspoCjUhzydPGXABD/tBB/
EOekgKHX97LMaMy5MdEVSJIgPh6NEVb5fonfBdzOXy98+5ew+KMQBQYoOsO8RjQLKj2IHkDmFrfr
+oRqU7WPO7rb3D/AOxDPOIX/dv+LXHYIVc/9PgzH0Cc2cNs2a3MXkedW2R3FSwbkdaZJx/xChf9p
+MLLP4LJkqKWPAj0na6zAfONsQMqfVIFlAD/0g4hvHI5rnsRqDL40qtUXuxGmFg35q3oZpRoDbHm
4nUlBdhxf8WiQz0WzTAz2jDsycMAMTYLn/Q5CxVQ0tC1L7UELQYgWJzJZcyR0cqmmjutQSAg/Rly
QfCHciZo1/s+kTkJEdHH7WWHtkHT9+7SICaJTHJCPrzL3/ZPgoqegTsk8GtjZhap6nxG8Vv9eCdp
oXJQE4+YiRcur+u68q2EWuQki0hlcG/5kq/adm9LSABtMaXgEkcbZRwYbtsrj2V8C8kbp+KO2AvH
l6QMi+wdXKsWCteIR8TejO1A3s+/6NjGb8tqXRY520yJLe1L/kcLRYiDVMPqjJMNXgAEgqE/CnfQ
mrqPms3M5qfVlrf2/rmUc6Nu2MXqvYFv1KePHJmwVB9LRRnt+PWD2/CHU7rrJzTc8z15s+ro7LpP
7gV3VJZf0ygrlaycW7rMIQQLJ52dqAUB6wmjGAdCN7ULiAXDIvy5KVsR7sshXM2yTuDTCUF2zERf
DZaTfTAM++Z12PgL8QJlDQ2zZjv9RyLHy1E7NjugeayF1C3xtEcrxO5oRbhEorD/9hLnvhjVcBmb
XjWR/jwd3yapSieQt+ROAVI0wKlr9H3dXEeMvhvUTu0Hsgc9VQbz/OCzURSa/ZzxAfi9MBsn2Iob
Bfu6QGBqjekVIX4got1LL4UdbgRh0rGmDNWRo9gOyESfRw/5T05zmIC5k1ncmxbxMeSKhtmKCNzi
ZMAcxk6uiK3HmA+4QYdtmxejxMivyeCyQJ6x3J4vNJqOSh4jDr9cYS5O0D0VFybOpqNmS4XWv7E4
Hu1pLc/ndJSjbUIaLN+13Ck0X7EAocKnwQFWocU2dJ/ntbPzHqUSAYjjK2LFKaf6mCRGP6uVuDsE
FpYEVS8ivhcSUzPWJ//SLJ6CXDPspI+D1PiCRFYw21H+Ufn6VI3Q3Q64oeUywhNccXvGgtfC3Vj1
wGoohneDQJy30JLaRr3OJv0ESSKvEHfCCcRL31S8kO2c6txa8aVXt0ivnq+l4p8KlXXFn+PmYv3K
r27MV4Ia2t3MRqRFU0OAu6S8OQNw4SJWnb6mZnBcebPlUpn4VZCfRc6jBQ3NmwIp0Z2nxy+3FLc6
+OQDLykTc9HmyMb3sqMpVNtbFFpnm0R/Iqz2P+pESlnp8sJN+M31muqvrOb3rRLFiQaiC8mTl8TE
2LTLZplBd/kFOd7lRJRZGDqvensf1z6hbOh+mqFgrI86U9je8/tVQ8Zwu9o5sPeLosjkcCm09YaC
h5CGwTCVCNmb/eELYTNxrxGQMgMBYNOnYhiVP9yd+6s+CtRODmjFXFdcirYHBonwMWraUNppktQb
m5tW8UIfAR+TnGbjZHlasBniR7SBgq3BAA+v3at/A049aZkkMzrV0rMcIVLDZ3uVwf5Vm/05431c
y+4iiToDFkAIArxuViBTauMLnwxoOWmJXbqHXerysx+lmOWm+Pg0Q7seboHRf7eQd42lL1S23Q+u
6uYSoX2eCA7gGq+l/s94lRqPaCCpje7AZb2ra28GZSvNjCCttLnm/Sli1b5OOGkNU3KdwWMZ9G2D
NtJwbpekMB1V+PAuehRv3m9c/DKQXgwPUmeIO+7jUmMsXMT6G1NAdzirfk4GnKcD9/v6otK3G7aK
U6RwBbTLKKiL3NWSmdbmGMfe9eWOuOB2VPIeR0NbOxmJaFM/YFAOnL0u+limCeTigGuCpjIms7+u
UwCDc5anjBmftkfcxoVJcsp6UBnScDOAk1uk3k9IgPSzakThuoZ7XNLW8mslKvSk4r6juNwCH/CO
m0P3nZr1yFW1EsXetM3tfq0Bla3zTkfQbXnjhQZfb7SW5WsjHP0MhMQiWwb1t/zevuV9letSalmn
XoFuDOJTORF+wNI/96Yml17carfGAH+N/ckC0K4TL3krQ19RNfiXMy22Cz458YQXodpCOHcHkYIV
LqqvhOwLsTq22ofWFerVWqipIaO3BKudCT4gsOy+jG2ozEKqRx9FxSwpB8hYTnVYnV7OEh0YOGrQ
29a+fcPUCKRod5bt+/v+ZLgBbZKZSCjuELcdAYbCnrr/lONozO23kXB00b1utQyhG7T0ieuf4wj3
DRRs7M7sc55DDhJF4KnyAW2vECbQX7nF+yyooOY7Qx9l484FElt/IEOxhlbIYw84zxahAPWtKEez
Ash6cVvK2gqS25NFYcbFYkN3/DtDyxq+MJEU9ErHqIlKvafqYtfODJA+wtHrv6YZGgnM5lQoqzXR
Ho2HPIhsSm4GPCaHQ9xQTaZa8/WUHXwMb4ELtwjoO5qFO2KXV9vVZVtZykQJTNxfIsvhAG8a+StZ
Tn0ntTTq5U49fcb+rMMIUbDiHiIWqEh1q6JM9ch/myTVoiErRik3f57Oy5TvFC2BfspUQRor7QkK
4WrE4IKGZ/BUl7gwb5glTRC08lD69tFt+zeKYW2WX8wIeWZjI1STewbOrAV44zG5YQTt6FiouvSD
y6YKfhECykPTCVLCsQ3ozLguBeqtGyHxWU/0hUUbznKkcoNyYnkJUnG3ioedmR9eu2lcIJkEDQkD
w6nDHGOKE32HfDrrH3TAdU0EIbRXMxtBAZII3nX45nhkl4oV91doLFdelb6QP1C5ED2vCYhNXanW
GuCuJEBCxYrDgTsBvG4C5F9mNrt3vNj4F6OiF+WPvPjbMYASiv2fH65RSAm5a45pz3i4rdAMG/o3
pXH9v88EkbnzuIr/EPNusBpdv88XXKDFHkkP7r3CXKgJQkU78CPONCRZTvzIovqEL/2DB8szf7eV
xc0zzebQhqKELgMPeDezci6hsBd5FEBxoL75hz8P+5KtBqYnzoLlcB+jjS5J+Q4Lvo8utMrCe0ir
J6mmW+yO/DJmsuCuMQEnGaZfn0teSC2mD+UgkKQ7F914O3f6MokDQ5xAisRYfP3lLZk0cFQ+xDTN
FQLA5BWkORwDJOMo5u/NHMCL+cPtf+JghJ+dKGAUD9TMP0EyU1+oG3KUIJiY9InzIz8ImhiBlKdu
6+/OTvhInbnks/AafKcUBm7SjmlwJlZjiEAtxY6rI0XIszJnt0qlj0oV+82zYUSYcIzWCTdZdR30
/BChAqs+FAHlYg7IzW08XglE5EvKZAZZRqmpcTa6qIgD4d52Wprg7pKC6JYy5XWercNeY37Q1NYt
GumxbvwjPmlCydNj5OS18LKNWiqTZbSd4mRNzc7ueaZo3nzTYj8XzCT6NiLhDmyFgwt7T0ptxQ0r
jBaeL58XMMKkzLJ92p4GQOgHZAGYe5gDHKY+7sTuomdwOfrP+SUWWmQS3fRqo5orsWook4+hoYhZ
XBEtUVAmCnLTv2JXKiSGDTtuU9gImkKB9PruFlcsUldPRKcbHKrixv7G3Ol+JBi05u8pCdlmLQlL
lboI0eUequMi72Zo6FlUHgrpwJM8jj6LyR2/TFkvjXgJQT+BEWylNADx9gNlwpxdScYI8HC10pIU
J/PD4HgPtrEOnA0kOjjpBjmmH8H+ONIcGbNprn5HgDi4KPIgfrbo6rVUOqSqHx39+IM5kgvienvo
agyZc0fQv1YFJhIaXLPuKaH0CdEhlKPYrzsziGnkRi3G+LuUwGEymZ89bfEtzfcCs9VfSyDVvFbI
pSHUWh/w+PfZYHZHlwbRLgtSvIP9i6NmnMTsuUG1drMZeBujJHuBZ7YHdUgvkd/0pIjf2oYo/S19
XxlM6wrdIHXyqIZpK0GApkDwbZYjDi7GF+uQwkq8FNkntYe2goX74M8usPm5e45hIgzz8yGJ21tT
LCAwWWtHJ+JDny585NREWjp19GRSc0v/VDcFW57Itetl6IfEQhBnHKsY7HomWJhy0uN4NJ/WvQE1
/jOS77ditFxu7DM6LiJR8Z5GELwk54Gl2Q9p33VnU+hPSeqBo2wBwZM3UCG+KopMUX1AS/fldSZb
Vnj31z+4F7EYjLJPnA6lV4NSjDHsAyLo8eHglhxW5UzO0/vV9mwS1P4hWlnVMmNEiEKnWStnNquJ
e3AEHQZEipKVWv9sSD5Q+AV1n1SX02EY6RDv3eSxIdEpNEU/0KdSfw9O7dZyjK6zo3/fA9JHQhKC
rheCf1R5xN/E/IaQbB9xdOSBEr+choBukmlEK3E98XMnh28eeU5AjRJK+6aoMdyTBo2PY9uX3Dum
MscCOwg60G1Neo834+c8scoltZd69GTXeKH5HfLX28TPxXkkg+6iwdZht77bj5pJB2FFKpRt0FM6
n3bITEnHXxesoMVaSvwX5/BxWdAUMqEh5+CqJenHGDH6IgDYhGS5p2GsH3io+a2Qix69vh0l9CcY
IuyVesfgMhjJvhqsrd4Tf2ek67wTT+e5cOxa5KFbMo8wlBvHtnDMPBxmNi8xR2shg8VyWXf1rsAa
+RbUyVH61TwTeJ2kBJ+m3MxBF+OV2mXr8TbvgkpDnUVxr/WpkZmkaWj5Gibr/w6IUiMDjJFWWfQl
4cuSG2f++8Rr4cWu0OA3BeA9fBE9rX+1r+c2FP1JomjaSP2pbt+xnwhN2z3tb7bRBan7nHhotXzu
JBxVliktu61rDMzGmOVRJC0DjPyWl2wqpgExZZ6THNOIxA4ZJtb5qVuAKvB8ML6IOhswao8fY7XY
W/nom8I5cPCIDhC0f7GqUToo3pK/y1lJ3Df0g/kgVvrFJ/wcS2O+1B25JzHncTPb10d7DbYIx7Dd
SRkvgLvHB63nGwmQIYt/8MSCfMzLlcXD9o3Cxwbpr78KhNCT3E2BUBIfkIJ9HprAVmhu5WnITLYb
4mEQB7bKSm5Z+VyJzEpj6XNYu2sn9koWTRuClAW/WeUCYP98Zn2Ly1iS5EQIUL7IxbZt9x26Y/pr
okkinNE+bR3S6v3iZH4eSXVscepdPwj7Sv9s1Ra1drtHA9YVPHTBTMKkXUo4+VCEhlgw4Ev8qJ6f
mSUZILOsRz5pBI8R9L3vg487h7FXifeyB9uNvL0IvKYSXXOYT9w3feswxj817KvPW/B7QGtfnBJi
p44GCCD4+TDiwGMDjmG4YitVJt3HkxNRoibZDEX37Vh0Rh8rOa4UpXS6trmIMFnZJIpStHVozsMB
rwz0wZBFzCzBFfAUrA6qsvyIVErFfbZSPich4Y08E/y67lZ5G+ZlVpbx0KvSIonjQo1xLePpEV5A
WEbbjfYgjirTAr07Vfug0VgmK7mSgONfepPq4U+GfiFyYzC+TD9GD1stebpR2ZL1VNShVqHHa3hm
IIDTZtWsrSD4HC+IttEsJkF0W9k0ecptGf8KX6/ZvU9LG99dqK33ZqT3rkz3HhekVjeGvqJ7ktWm
nUFiaEHxixo+lz1ru10plDARnuIQEOjqEauBxL1YY2jat6ZOTB9fEgxEwFBZVSdChDuKCFbSs0md
iqb96jjcyl+pV57+wzrIbQ1SNcnUigtQ1mgpm8GbJm0qfOeCXwuxSnkIs1G1T+6Om5SR/n+P5+Xy
p64J18dNrUdrQJ+D4GqibdE1ODrZX0TMgjsZBjh8sg4Q+eAVW7QhwOI1sVICKTjmaQnGYLIYmM3o
LngXrT6tzJOsZLhBSiaoDKSL1kZ2XOaCcZVYUunJ8sAfhCT5/pO1j/m/aV4nyjF07xBUAuq3ouZu
eILYQUn7Y700b5cCBGVOBS8nCW+3jz0LF9lxxitITx2YHHHLcNu4eGos+iJAAldCDOLREmLq27AX
mqy2cKtY+CqmiF9k4+fZtqRKIGN+dmtAUB0Cu5QBqdku04qx0P0U9M8Eh9eNYYOmCFdWsxuEz4wa
3RePx0CPC5MxWMoUH1AYJbC4dqqS8gikQasmeokY7LfL+CiBVl3d/+tDiPx3rVTr0/b6y2ckNB9k
y3Kvq5wlJkgKacV03p0uW0Z/ijKmEkWo2wzPT7YEfywLM/oMTt5S7ToS0OrX02ofAm6DF4bohU3U
ilplKBiq/l9dGEPwNgp443y5oa/VQNPSe2JQd+WFi7jZFLmKNN5xwqIiLcm3WVCoOWkOUAe6YkSE
7bQlZJ4is6A+6C5ggAAoBsmAeaJB9h/y+41RJN1DzJGPfYlj3Otpah0jf/CpEPC1wvT1g7+HKJvH
5QlYoWngD1qNMmDQAHLN7xtQ2xh9oPk4A7dGBbRVVjiNOHuiq/TJ3OyqGWqtELYkHtsQV2x2qVkO
mypvX1ZjCGucaKuJkxD88WDMusHMI++ceIrx6O89Mzh9Gpffy5yTDYVaJGo9J7iDELOWzJL5uRCT
daBx2sEAURj1kK/HcdX65AJXQ31FSAbKuw9F5aBHMPeD1rmCmXHv5ukObsPJMV2tndQSMBghwTX5
sGH5X3r9OGHRbqrCCk7DA0z13HiwAuJrUjUnL22OFB52ji7hCWqoF26oXKFWn3qe91BaxF2FC+ww
8RotJtVRFzNiCp21OlI+7R3kpvPQ7xnlHn36ql4hZCNlYNByYJzXxnsGufnD7RABJAvFZfrhfaGK
1hvX677XtVkzBeTx34w0eUmAVnrM6t+kSSGHaWlauT15sOty1jg0WSVEjcX8rm+eUk7eo6DFhR1Q
b5YBCSyrhrHyxv7Sk3eAtnpk+MKlhLJsHu6+/21lig6uuEQfWpqP4SFneU3ZyAZEzlvl71kTpwfr
KTsjOzyUsMSz2Df7n005PLXQ+pWtnhGDAtRcyR2GPlkJvvreux5ZVPqobgobReG3mSmNicfubO43
U5TTd2KMslJYyXNXk0Hk15kJbDVcVj0BjKaUlIBx+zXO6G05SO4KPfzddYf0myAPBBOwgLaJQ58h
1QoSEM1YUjeBDcGprKb4kgvpnP66/C2Ix5O4fTmqB1xVkjB2MKm6XwAcAqdSCW/fb/i3Pj5ifDGl
ylXNnhEe4dAjxPTkaD7qgP6D+zGN8ufFuyhtefnyQSrcIWOtkmeZx5Y65jHizM0h1bPmlnp/Yl8s
JZ15ddaa6gRnQxhNGKb5dhLYJO7kDv3Vpm5p1JEeDjdGRVt/nC0jHOPmRq6cn8tT13rCDqmd8jsz
0vkqwM30A9m8dKSlaXe1hEpGP4N2fIBPaoxk15eAq4PPnUC7XkqTgbTa+3EuTxpvMWV4YATVk0WP
QBhoCcLReA3SCRtENW5yvRHYCyi4vgs8IBX+/gEdpSfGHUHwdovSjg1YUYDcjcQ8q9+E74q0jC5R
jBd/OPqMmRVvKss/UUeJLmqm1jjZLKCc4kjOhuPavh6AIAwbJpKt5gYBl6MSHC8VeTG/BOGhfsGi
b6yu5mwU1Va76YlIhWYfAjchUOdCjnbueOD1Gun4pSK/6gbIozOwG1/4UxD/06i3RY5wCqLdujgV
pkpVVYMbSXT1WOY5g8St3PDhGaxuIWHHB6zTMSE5TbhMqHWqtwaD7VxtC3wYLb/Vln9GQyS4a0Ww
IhWACZ4Y03i7mnyekO80GCIzJepRwHCyhxDXWi1AUloOJntjqerH5sk40ePAGm8ZtT7ymY/jNdrS
OkSqUGRFQvpQtV9tOAy3tYrk9y8MPAhXgrZt9503ANXQF67MEUUYjqXPbi8RTlZgND5Fd5Dbg4Jn
3UKreM1tBFptXgNlPnYvlNbsDusYMFlJb389dnBq13t7F0QJD6roCpbQikWve7KYq6xLRYJDTz0N
h15qevouIRUmGgibC7Z8/eLKmcVzHB1wT3hF4ewflsudA0bXb5bdXhefSU/p8egELtgUETGwZqcH
cC1gCaw3ajCZPU5VXfEZcIWptXSXWClTklWOY6/ZncjLFODw/aZBTyDEbN0RYT7wHGetd3JbwN8+
pbk6nxv1rnSLWUtXQobNrYXuCO80beeXrE/oCs929t2Rhoca1y7WDGcSMnvSIRCuh+5WaaRoQgiB
yKFrdxsxJ3lj2c3iqN27/Cff4YS1kCABvDO9r0gtCsHcKeeqkFpBbTxKB9+aQlX38qY4efm99R5f
JjL7FngwpTJJvgYL+pVsTEVwiv86rVItqd1w6EgD5ovZNgiapDmfnQK+hsMhLmLCdXkWhcgwel4s
2w9QpohDiNHbD/+YXd+9Rsw4GkBS4NbS7Aq8qrj+DBYjMy3mi8vT2mQ0qYaqGwj665E2W9/Afq31
+UAVmtclNF1T3SyvRGyQxUxzgI+oQ1+b+MrQCkegYK1pOeYewi2bjSkMfdV8adh2x5cVYQkGRcED
7r1G0/dbG4Ck5HM/dfCMsAvPHmXLKcwkCaZumkCk0hZPwyWElea/KiQe8hbHqld/yxBf808VsxZy
j+jSZYwzCGq58SL0oIFXq0zYb8Zt2v/T/Xyv0m8fZs++xFbEnMoj0E2BNX/g79lwQePXP2DJqIo0
0ovzorRJAw8fWuWpEOBBerLnOEHRqBzPwk9ZVbSKnj1/m7kyvncYD8Sns1pcRtcoFWiz/ziwqYyt
XQoJkEnvfnqwy2dAC2OaXBcJZovA9u+7dMKc9+0fpWNPsUvkgtUWaSbiekLr8bgm3hmoaI+orSBh
8yRQj8/i0HCIj5psHPspaw0/PnHsY2LRO6bMbletV5aeSgo+4/+daCWqIZ4PLCJt34shmW8dOXPs
u6bYpZs5s3NR1g0rH1gZv1lw9ENztAjuY1oLrwUHPxcXxyVPrPE9+UbIksM3y4NxCovl4sc+u33y
lvTLREUWbLMAjfmGHGBCpmnYW0aNZSlNJcqc2QTiWsOjJhbv4BcuURT8EGIHcjmilAa+XsltHc9d
O8lmouKHxX0iB1z9NJUTLzgaaJS+h28nnbCBbfMzL7K3977qZBXyjfz5Cj2Shi1Ib4JRMwO0bnPN
Yj5mU4KmjmGwirUaR7YfJRzpw4GDaifeLvdbP5fvsco3KkQzjL1a7aVqaEY2g2XGZnhfx60ZuSHH
PDGycTj41PAOE6kxgXAo38Otw/o8nn9bfMscV+lmZXATPCvunIIvtcPoaoN86Ake25elGcIoeMix
nIEoQV+jYhkxWzaT
`protect end_protected




`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KMVw0FCOv34cWOupKA05LIFbQSQzhdC7cNx6tCC7Npkh6sezaILAhlbFmH18n8IdW398pPD6Glkh
nmMHOn6obA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
r2Vofo4ESYu6AQRP7OJMqj48QN1X+bTn4JEjmARwD+qhEKSRQmyGOUq1t8l0qg8qo/ZIs5VwKYwK
blMPD6vM/uEwnk5Wez0Hq/jPY0aEpB1pCERAX2X6smsXJzU2JpDb8Bv4jaiPQ9/mgDegydcxJcW4
WBwS5KXFO7Gsz3oKPK0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pAbtnX8wMTjyj7ktuU7kB3OsG4J3geGiLG/iiwFlNsW8S9qlZpamsi0d4sQtTqmPOjyAT23RYI03
3eJflbWyfGtfT0plGK6bngtMyTN/jf3W4syLadA6h7j9E8mOIobqiQmTamY9g0KJUU+ANrgjfOeN
szhoWM9qDRgcJaJU+Cx+nAY3VB4tTyv43oIrirLgR86OBanyXXakWvhEt54DbM0vCZ60t/V6QWMM
5AfcUu990jo+nQDtAof4C+iUq0lq5HXoPve30kHeLheDubNTRgn2Av6hPjPsQ5Qz0j2WAarM6KDn
7cHfTFTSgsr/E7X2uEKIN/4lJWHSxKUq7PDxUw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rPYRq8HUEihuLW+Cu/YM2rG8TnDS0/Gq3OuS7DyesuYUbl7NRmqXiLHKzc9+77PQjmWHaU9ZJY3w
N6YcIOiMSkWEQLpbLg/pbpfex+DdzHHsSFs08kLH0Aeoi6wEMuwmutXxMSWf8pv2siWUaPA+NGwt
ziAvFi/n69rNrniM8mNc01TDuU6TvFPBierNczf7TfHf/MJ0sVVYEoNF80pmcX5wvnwy8yXBKI0h
aARNqp8ky5v7QanJDB0j6CtBvpVG6YZ2Cm249wygZ8h9+3OgBMbaZZew8UY3M34veYOSjAxxnJQw
/3/KId/WU24TWBYnFoEwhShGNnpuhsluwktCvA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
H+vRkXrzIAXQKMevF01F0iWGRI6js2UlE0nDAE6dXjzlLvq3M3TgTAh1S5uwJFclzk5LaWErpkdd
bbGl6vqhScAbxp8N6yS+iKPZmIQgQybWc2aK6E5OT0qBcrXeLI9rd8c/FZH1E3d1/n4Ejgqjikka
Zri/Blr7vecUvt9ENOfmv8I2IwEibXrh+G+e6zXmAsiml/ciKeDtM4i+Ep7eUoVnlGB/uOC8buAq
eddIDAHqIu49VqNwin/vaacuHNEK0yjtupoIsxB8Fq4F8Wxk1tYNf80IQzD3C54Iz+D1ZmCe9IHQ
FU9XI2HrbdiAqeZMEgaa1bJs210sN9JTZGjtFw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
j2xQg2iDFbFFI7+dDRrAxN59y4jd3S1Zvtd25yqSjv9nr/Fw2RraTH8/F2fUIIHYeeg2Wby5LkJ2
CgWtYUuRfFFrqGhr7jf8OGrKjgf2FYM2Xn6Ltu9TuJNNkSLA2uR1ibWyQm3uIN98tYI9tyOskioh
MJOMCB7MiE3RwcNOta0=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XpqrVh5QI3WGWXCuXjnC9FYqu4ZL7+4Kk3kZlGgM/OdNMMdHTEE+gPHVGUx3Rt2e3mpY35HZ2V9r
iPS63FtPGbct+LA3iXsM8a26Sz1cR3DkQE/0Y7FY6mH9bqFXfJtntPHOz5eKls4LZH/lsg+59CjB
+WIVFVBGt455y8OplHxSSGYHCaWt0qT8zehnOZIx8jz3rxqduAMXu00jSfT3adACc+zTodb96KUD
xqOE3iNnyc0nU2JtLHvtKOuVLitKfLKEzKarbNEZ6kLp3bHG4da6dXCzxwe1GJ+OnfQYqkgJSU/b
hUOKvViAdP+Zre00Dm6xQdH/XIUwmpbDM9wlFw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 214080)
`protect data_block
kjWOEb06IAmTO195SUJaV7oq7SD/iUZvlFFDyvYX1X8Z24E9mxWj9/dOWA/GmBQD3YUNjWHzscXh
JlcVWSiYUd3XBgPmfu6PJXDBNaeHqfyhixiChosvthOpJBWkZuSeFCXwkiCC9XRsDsLK8sbNyF4O
fsKGEZACstnbeTOWMzgziWO7cUMKaNVWCAgZjaxaMjpm5LsyUBN/nym4VvvzNtAZ0rwEToByRKqa
Uvr7X/+3+S0id4pDtaNeTf9QzSduiE7ewX/om8JQhVlAigsqzPKiUDTpthHx9n1dqfyS+uYNEbJ9
pjUjluRCA+aHHc+FB0+xepRE5CPhoGTGO8wFsgHH+qWlwSUBhYBGb3t9hPzRaFwvJtrDGCRBp6/i
lTyWREea2PvBgn2tUtpZoMgo+ykVvd/mcBvh/2bG1WZXTd/FEhXtaCCjdZpso/Wm6o8wZHSf/8Gi
0Lpqxl1Gf9517mEeswvMVOyUbTg7Pq8WYIGcuRiylkBvZzM8U1GIk4FjjSEGHLN1ZF/0qJcvG2IZ
vJTHNgEE0qN5UgbSLe/IK+DdhtfVj/m/WNKEUyAAUXDkBffQaiT/OsHyOsRRlT6nRAxE2TC1SoY0
PIDqtVYp0p6WjLamS4BbWrmjqH7dqKZhAuM2kWbarhWJFUUjLAo4wnUwwHyuwCQgpkjuuWT4+oNm
1MbCpBSzXhX+ONPeJQ7sPY3wH42TzXF7GJhirFdnyMrg8X2nYeWZGWeYf5UDxG1WEzfP+mR4yhG/
/NNohR2dMS18Me0YVNKkQZ1L5yt9soO6nZN4tXyJRVTAwtMmbeg/P8YBXkwjps/h30u9pKJ1Frai
ezHQRRAI4Bq+rP4HgYBKhB4DXwiUD5GGtQU/CRYnVnOJCd0xFlheFxl4QEnBtb37yNWRrFADA6Cg
zFZ5P22+gGrEivChDK9jTUtdRtliMSzUeaGJL7b7m7RiMsOIBG2rzvpbbbi+A1/4EH7EqucEu0kU
8ucpfT5qEa6jKVM4JAaRfIbEAF1plloSqZyw9lR9iH94s4MFJ2ylFfbuupY8UgtSHtiauDuyRLkV
rwVfwPPUC9xdFcSfMPyuQO9WEuYoZHdCPSUQaR0HDdB3C2aiEXsm+kENZ6Q3UX+YzmMGtgQ97Wz1
ZFxilswjlALb5mXeoIdJ0axF0EINSUtBg8zxjIIyBQn45kkD7GWqe9tcueC8qExRCkqaQyTaZT0i
zTzNqMQdtCnaqY4a4Ze55RRikjMO1YpbM7osp+vx+aSclZGo9GvAFN45j7GUm9qvHE4pG86bqyWG
J6nbZ0ZPJMY0QsGnO3mv8ezRNEJUWJLYVBMXRhcD7XGFjV+BNyJBYM5BvtNZ27zrwwcX6K8bLWL6
+uS/fCUIyWYVFGB7Lf63m8HIa1/S2hmQT2I1ue0r5fVaV476XxS4bNr7ZGjQw/WPMQoKQ0DLaE6n
Hmrg4ujXk2ivzgZ6xaSRTZ2imK7re/yz3PF2WGH2lU5qU7aLtemm8ntzGcv/xzPhEJ8nK403wegQ
RY8HcEU1QlbeDN/tEbzDaIrLRzYuIkm0/JYz/6J6b+/zFWNYzZBjhtW9ZyKGbES+DovzCwZoXeQ4
sFMI4UOmWptQw043/uNuXAd/lwoQJTNhQY1c8UpImxH9uamq04JBDnHVVdV7OdMM3mIYbUmXI5Zb
wh25K+fEVeIhU/enXE3hE1awbz34fPSlp30glbUpCg1EEMt7iA2odpZdsnKLr3qiDCGY0ieo6MQH
dAn7ZqCPmzqj8SfQSvbBDPswvFUAPkkmNR/kHrCaIJCEr8vn8II2KejnoUHJwXTkARBGgupsNGiM
0CB8xYWSC4YJ4KIRA2rQW8T9v3LbxNqx9skYot5U5GdBJihnhj0qtUKFLCVykBGsZmVgV6y3LZiX
KDAurTur3She4DFrgnSZeMTTpHu/Z+xg5KNLDp0IX9MXmTvJjOGE0ivCSP1rb21+oJaa8PkL+DYm
H863cVqyy6YcKKSUEkgoCg60afZXUquzTc6BiPbIR9itdqIbxWkgxzkjx8W95/3URIODO8As0XHR
yiYwYK2YTA+zGUKJjce+41d7kMuJwoimJYZeMFUOClC8UzlIHC24X2CHOXKRpX79qLAGxLcZr2US
5gvwIyeAL0/dx8ngpzardqo8CDoo1zNECIe/BpZLglB+DkZRjZH5awmWJGXTvCyzCZcOed+DgStk
2D/RfK+BA0DrUB+JKoIuxD4JYtFbjJPA9DJuVVO2bw1HgCD3XnuT/L/eiwPH6mLVmxYWoi/AyL3p
dlmG+IdgRj8YpS4YPvAWWXNZfqWA2uOJsGUZF8d/+pnh3VcMKEX2cUjuIPcPmUUsPBWTneiuXSrJ
kWkOVaFLciSSs3VetQBwrjSGZO7EW50Q97y9rOK7a8C10ok6w8qVioZuKLhwDnv+O4lJFeDARLQ9
2RPkN9K9OrYtAXc3SWZXj9fgT5Hk/VbTG1jjGK5wPuBj/DthduSQ8eI2URX0/RrMbERGbmIwgtXF
UYF+OxZvo6Wp1zA95Czf5uvjh2AeMtcc+Xahbl8mbQTkdzdMgYKGvYWBDUICKUFVJG12U7I68BL1
CkBFnTIoYLyn4ONaXx+ZJXUqSuS340+uE8ccXfS81mtv7lvRiVPtUsCUkKE7/PBGa2r3wbqASEkO
K9z8s9Ud64rTXkITA2lGIuRLBaoghslZQ9A/9XDi7ftlDne4EZoYAbFcoueucnGJ+2JGyhHL+l2z
oHn+bQqsuZfOTrdmlgMJanUdUN3ITrcnedQtkgNrECpmxtBI0a+AxjlIGzNVpl2JpfSdoDxJ9r9T
dR7YoPxkj7L0LfIXfrAJwQ8F0m0Fh0fOmxnyVQJL9rijmTj2wgyrama8KYD/rsgxhgneF8B6STIA
ihGBZqxLGFOSXlrNv8Kv++JzqzqeaPqfCaxgPOwFt9brvfj7nsFIsNIVrbHRSirKtlHpjCLPx3mI
2i+IGuVrB7cWwHy4xroCMXnUTfj5moX8GLja4ZV/E1ZN4CbaTYw+9Den/9HSraY0ugn9TlS+uD0T
CoETyawUpbWEgdG4rygH4IH9MZ8TKI4l67Pn3isC2nlV+buABcaencP3jQfF+H67Jvga0zBMT8Xh
KevqAwnjK42yjSdVcaUHSEoAed3zit6bB0AFd+VAne9bBJaIynaNfRtB9H/y2nOP4uBy59QAErGY
P0SWpPUUBA+sGYCt3Y4PuVL15MTuwJTBaT7DixCQQ521om69OT71vQJP/mgWa87FBNTOHJLu5yhC
GYmjbJXTCSR0RjvwHgo7zTUFmfmPMYsqqQhEsRj3puvHsDuMWjcp4r57mGAYkMtpsFw5JT6+TcjI
Ws6A/9lpV+lH3PsXG3DnYcGh37rf27miOc9xjsPBawra7t0KvTyKpwFMUBHJheZeDCa32YbPxsov
MaozmGahZ80LVS7F7+7nEEUgzmTOW8er7+DwYS6EtUNqauAKiNFy/OP8j5wSiX7tKg4BjCZbl5N1
Ph26s3YiVuJP/rQp9qQMoj8FgxE+s+kTu2MBZ4JzVTbbAxGcwD9Qzt1gXrhwX+GusaBsK8FnQt+S
Qv67/ew4tCqbJgFZchLFWIqHeuyq1QwNUWme07dN5/6SRaOZR3PxgNp6ocPDru5GkrRp93KnovJd
QdxrPURIbl8xEDgfP68abiPnMvsQW3IvGw7zkBt57ZM1NuvsvWhEL/OHBGK9X22DdlaxbEz/YquA
FuH1A2dIlUcVdwB7SeetXbru9x9kwzXLZDdwIcW6HlAxl7M9wJk9dmL5ozMYuvdsDzTzWugVz5jD
lW7H9F9ouXMQtFm5XHuS+Au81Mflho0SLru0NV1Cmg8Z+bH0MHcN+c9iFG3Ey4RiSrr3OJTcSOgh
BW7bw+VpEQPpTLRqkHcag6z6O/QPlmDnY7v+DCVpa27M3Ic0ddJDU1tmBXH9mCujnPGpE4Nc1ua/
tWzQbEBagYg31wjoXYawbBjbvx3Ba16aMVRBPJ89gGP80gmhBy6yr3KiYPokwxmanYIBnfRnpxCc
77xWQkP3EKYN972X96wBhCA5Sdn0q0ZWJ2rOTkM+W/oFITxzyz0vQfD4cOwh6TVY/ufj6WcYeUTW
XIYwDG8FjSMk1hv9930iXjobkQgalK3Dz5axpRMI52udI6uJYWeaJK+enMniKx6mGbFcj9PIKE2I
X9szBJh/emo3jfCsDOsgtBuptn2v03UQDifnbDneKri2HX7x72d/SveQ6wJ3wLU+kt0zYjvAHAu2
0S7zjnSJKuQZ/wgQ+3mojHTczjGO2j4SiveVO5cwjHISrcoezDq3Y5MqaaUBqvbVWsdD7tiDvG13
MGJs4cmgLl0ZZPdCWinWekWw/oyuiGmTuto84Nc8ryXxDMduS8onFBPT/+t6fT7ismC++MiXQ+BJ
g7XiPGnDj78K7m4ct52RgSQ3Cbjx1L4jffT0h012NBLPJpsDMK4vCUkYlVgRglDwNRr4VBzuQ5hA
xhhhYupvPt7VBWptqHSRc5JbRgFseoILmxgOMekPO4WHCKo2mIZVM/OXGf9bDUcWWLrY6BrKNgdR
t3MuHyov5y1PXbYYHVamaIkJodWlLh0byFcZYPTk3ODiYzYW0Jeo4cIE6LgZQn8NhjIvzTgdrf4N
b8M9LDDP8V5vGpl+C1415x/jUhIvfBAMfPVAj9tMxYOMBw1YkmxeJkHuNtcuA2Kv4XWRCu5hT9tr
30MtfHkEARNldlfuVPTDaHLX2icb+bqLlG5J6bVcfvm1qnW14R/lze+Irtqhoc9rrTbEbEk1zrd5
/P84RP/hEk8YYBzTdcnlB429NJPlFlwNC9TPwmf2t31YVgQyFcGE0PjABQ2S5/Rb0y1kRZJ3nnmi
Pg1yz9hKi3uzwZE1IU9wMxIYJP3+P+kQGOtTRI5vhrYcX8UbsbGd3Ut7vuIEJxbcp3/r/T+CeEcQ
5KG3LVQfMysQFA4/IdHB/U/sJgyIGN0gjQfcnctxBjcBiZlPR17Qb7ouq7xvi3fI4KxktXY7WbDr
RNly6XybNab+FLPwThhfL4zikXPnuP6Ojf0KYlCLM5ebNVEQy0ixOPyQW96LiRO76MdtVw24nVJN
mffmCTnmb9K/WLl4iHrOP3VdmXiP1WiqNfIJv6dkPVClCNVDP9bDauIsA/NI4iHdMCWBq6f5CAdL
s+T24jh0/vp30ObJ0Zkewl2fJVi8y4bI6waYaBRX1+VfqQrEZYg/GknDqjeof43kD5mdkWITugmd
rHgtzewo3VpF+77+2IZnKonqP0i60z/GVqkBRfdeq3GD7hxCdf5FMYB3FS1rKi/1tDQq+cJMm6Ty
rffwhZOAZMDMYn7sWCLHrMGF8FDWZkU/isMVDPdyY972548t6iSsS5OKYc/Lqvr/jpBsuXCwC5Xg
zQ2YK95xnTfaFXgjQ241gnubmOebEh+vTY5wnqDyWpM7+t0oSGwHOLYsun4AYH+jc1uZMI1qHR+U
sLJ8UcuvAVP4fPypa+kAb5mHqSAbxTjQ8euO9uR4hBriWdPzcy7KKb3AaK+QQeZQFnfyhiIdd+FJ
uoSZLbdNoa9EF2E/ZXAS2hvGF+f+gsmXxN83xDqe77MixHVhv87til074dhtFRzf16nml6NVNw+/
i3oEDL+Fqf3IVn2Y2WDqcYSFaGix/ba/MaoylheXYF1ATo5SYUTktzarXG+ZfU1aIgVPPsMKwcaa
pyS++QT32W6ui2HokxYFbwVWZ1joWGGkzf7HwgP0EbyMoi6Vmm6dYO/kDixSn1diTuX2oryjwYs6
hYtcnGuPanrHlVkAgB2J1dSr+FeGaQ8Eq9gGHTiennq+oRNySHeX1GNOG+ej19je6paEyL/LfBib
/JDFrg2RlerQZHs1/1kqmUcaTboAIGhmvo+6hehjbnnmTy4H0XyPeBNtTZyg4FMBfR20bf/Rmn3W
ebesdukJ8wuEufvOzIRC+tq9bSIy1pBipeynASGN0DJIdT3nHenm6ViGKRMCur+xn/gv2PoeGn4W
x3GQKStMi4jc+TuNd45EJ9JchpRnEbgN33E9eMNyRPzf6TGJDlWOLL+9AaEdUzveeK0ErDuAsy5v
3zLC9CVWZLUqfRntZKXl5xw1FH1wOTSrXo5hV5mQrMPpbfISeP276noHbd+yrWJ6THPrHhugX9Uf
Yzf6Z1FQSOiQ713oVNdNw3S9k737ELialCiQQvbIhudmt10BUAwVLMcfIgtS76pJilJ6e21j+SjF
8dnO+tlbpmI4NJTdXqg0TLVEMuQe7AKnCceXyE8+NiAnGFMxGcG/6dWBVfnx2W7DjMnt3ige3Z/K
nPKfTy1L90ZLspztRLCvjxaH/4tuvM33WDmIsbjVce2G7p35737+UL+iV79cEI0/Ofp8DTHakZMZ
h32wpPsdOofr1sCtd8hT7jhJdTMuER48I1axW2B8PdNFXVLuMGjRNcNllmlDX6MLAeoiSeV0zdpi
9Tgn0tY2mB1ogFgkSX1+GKVz3tFUeBGaxxk5BkzhEnz8GlhpvAjK7jG667MXhislLLi0jRAAG5C0
uSvRuaYgrGyDt6QtVCu4VkUbFBae+W8D3keG6VazWiKi0WMai0z98RqHEU74cSOvMGCh4AoRo620
NQdwSn9+qGeGuYshhCDwonf8UxL0WknjsybY7gl8O8XD+42wAs5aeXOQEaxpm02KDKa+ibiyPEVl
DIzqpaQ66SKTRga557ptNphcBlCWBNJ9gM38RE1tq0bb8IYwpyjlqXmK12U0C+tG7se3gVsENPmy
h324XqJ3ysvlGKouwOQZaArR/eoUcrzy1dO0iekKjax54Rv5nAyeQ6pPz0dIDL6rdHOQbdkpmJ7g
h9fZ8/FlQlQSF37cUFffWjYITOFHu8FF2M0DZmF2wDTploBcyEPCB6/N1PwgStOaXlJ8aK2j2Iec
RJPYyTUh9JLMfOxrsMHWf7yPM9dL/CNDf1MgsOciSV9KRyDBjAH1H0fl7XHb26kCNSeyJLFS+Pqt
KDWhjM7ItERA7jabzj7EqdW9AYCpP902DA0d2Jv4hRiWpLrlfdoqPJPtydHBhoAv90WYH9db8s/F
6T2HqSYiHqA8za9u1dFE4wIdLjPEaLnG9Gcp9Tn2JqzJ+yQHpj4hTHcCIiM6oeT/7HR3JPTOJUiM
Mf/K4z6g9khdWlnvVDe4VaOspCxxLcWEoTk6xLblAXhtLYd6OzFdJLT7KJDKAU5N5eedWgN8DA24
8C0WVJB+Jh5zMzxcVsDW9TRkJ4u2M2FwtsRnMCaWFcm4CbFostc72FpxuZQVRUyIMTcdb6dZxTmm
ZCztrEEexidtfffjGDbpB9AhxD+DMsMJxy5lef02WapGDlVhRVwa1O4xkJkQgGeV6TGkl9/NMKo+
F/gk45zBSv1Hv7/Xr5y1rH2j9a3fExzIsMe8B5M8Wzb8CYs++bvTH14h4QNiLr4HksHCjYPXsUY1
LQ/BytdlU0twnBNMwbQRLzZzcdaAXShHcCATN6NfQJS+cuO2Pznf7V3rArRlQEhC0PmdP2GBOXN3
03GJL7W6A//5qU6kNfpttIwV05Y0HyN/6P73GwrjfESXR9pMJ5RZP30Rr+LLGYp3zJM16wVzs6UT
HdT1q+E0cPMA8yiI8uhEXNngq1BPzI49wY7aNrJ94N9pKEUbOhwNhJhcNI6GzprbzH9XWPYJqaSh
K+xSK/niJYP/kVxuaV95zA0FyGok2F1hMi4ypVTEkhpdMWcTltI4r5GdRslteq+cNHZEpJZIKZ3h
7Dejqju38VGE5C+ocaFcT00L5a2jANztIxhXYCdWdg4KIVGcZX+vYmY7qpToJ+OX9QMO2bmf4Uwl
EPji1iZb4LGNCur/SLpixHa0nNWQCqDE6ryEfvvtJ/07J261KMY1RIBiToLGfzWI5pJEgPNPnFDu
VelJk53phHB6WV834q0dqGyTfh2/dYCIuZPuoV6O+ygQmfQE0b4xkTrshb0DSGuvT7r3uShjsaNc
cTNzba8QCULRhpfyPy2gF8J3ZcMz0+VuOhLEYuhXot3SUj5grqqKh6cHBDALq3TpN3ff64xsAvbR
ESzaI+t60srq/GfeHWdepr9/vsZ6tyc1DfKmUOXZ1eAy2YJ5TqGu55OzF3uHAVyR++iTS2IteKoL
xOrMONUht8RrBkcdkRUh5kChA1gca5hnsM3BGIWnEKA9cjy9RT/BE7eiB0/TuRKVwaqdJuQSMPU+
QXHIp35Dohhzc9N5StWtbK0LmJ5x2xQSgTX586Xs5TBsB7jlJnYYAEY1yusaMrz1JlhgNnJ7NtpP
6bQjKCItxC8wFRihKr9ECWePSFefEtT+yn4yknkaqfEObhMK+HPXWNcQxXV3jWO5D9ySVzkVSV6N
6Sp8VfVmmdFuegt3iGz470SjjDJcCmB3PlM+b1MtRmf/OoOsYy6YquwoA0FObxWDcY6alY9s/buF
zoKEddywrMw1Yu5VQK/ODnb6LHRfCe6RjnKYEJ7xMmd41nZteJOlxpMkpD9t3l9877FvjMqfn0ph
guj3JP5d86KK6EHcSTna4ZlqgPtZzx2S160YSYRmQr8CzxCKP6fqdqyrve6VdqQFziD6/dH7dxo5
IyvIHGhf6RJYbZMJXE3jaWx+EKmjMP1P6Q4pa7LcUIn7Ao1G3KZITXWIrB96fv62NgfAqTBIXHbd
QWjdKa1lReS6KePk48gUotZ1BHyNVcKsuH4I7xSTazTqfhuNo4Zq8rAC6u97M/vstLlo/MMsT+79
6sXrxOK4aogfWA8Mv/qlEgaGrDBF2uI9DAZydbG670prJGThjkY+jnY6k55ipQ76/NDQANCECK+f
ZEaYfuvlomFTH1pQ1hbF2Ol/rj27g4V+CKR40isxQTNJKkspZ0hB3Kvo1W/VbdzjBFVzNk2Kgkqp
I3B86ZSDtowabF0w9NVt8097d4a7APQdhmmnUVuEaUD7b5pYU1JFLiapNIaTkhCY8tp4RNfy48Zp
l46PwYj0ACLszZYOVrS+fR768K+7URT9Gjg7dasAvPTWEiVLAPpim1dMCKDmonrfqRbb3glEV4n0
7JU/MOlL0y78qG2USv23KjIo+Nk8esWAL3/rDGr7gYpgxmKwsTimy1o3o/IHlHYZIazhc4D91rW3
pkIj6gr2YVmEK7Leo/uCnNSn09tDEydasX5lalj6TN4B/pgmO9JPCu0QRakWKEO6aWDQuarf2H8h
Y2EqTu0kxCMQBUv3FfYJ6FobVa6V5c3YUBLQgVdFWNGNq438iFQfESbDGnehkGjGENaA/nNFjcL0
13PbcNsVZ+7AlSVtannstwJfI4y8yvYhJuXWkADisdVGA58inWC7cq28Az6ucXR7bt2aR1kUxduA
+SnBGuQDNE67YyBrebN6VqQKuRaykK557Nr7gQ4ujC89ig7z+v+jZ1S0jGa5apRbaF4X2heXY6oB
vsHoFGknsyBdwY2TL7+/FZ/ueh2ebYt3vIPpMpMfJIEHoMVTc6gUbK8xAhP9dMcLIzgBpV5xKxGG
vJW/r1OfWZOCfakwi8NRfaWrER1yIB3IO1r1e+5h3GxxL4hlKkivthxDQaglcZ6lsYgvSZnGZgL7
x4vRGG4KCLLEcLdZTSURn+GrwKDtF2gMwbZ1EeUjLofKiEcSpHM/tH9MlB8SXAdH3+b0i2w7TlKm
KbANgns1Po4GUEOwBs7uWHP/uzgkGOoyVyWv2PCvfMJ/VNhXU7r+9tkxiYCsdXKIBbZqZ5LRSTU9
aK78g4KUWOHDnI+u58MPj/OxDz3mcDAybJXZMrQWPIRhNec/EfjggnPETGh9wDZNJUKswrji4ZSx
hahkSyj4dajHC8pADmsa99UoSVVvKqVsa5ShGg2QNxtkJfHelOdnl8Rj3S+CeshtwPW7bN1T+6j8
CEINH3WenPgU3HyAJWW9ZT6CFi3Pj5Fla0p3U9Fp1+HQhpLCCdAIIkV4fRRdc8bUSDbOwZhi5xEF
B05bMw1QBb2f509SBNkwPrDBn3sxjLlccLRN6tQBPjMigxCjiOEqdvgxyH4lj0diTDZlvF52lO35
z4eN7oWti2lgosRxY1zA42fSEkN+tPHME0Tcd2xu52Sz1lDArqYu8DsuAtoIQxjdHvHrMW98NO8s
D5e5Ot3y6CqDyLbko+cGHXKCzYJHiQYgdjE8tE5jmKBBtAG4ldj/0pHSc0V7bp8xtalXuEDc641h
/cTbESD0CfQKWF1BHzEwHbvz5rVPErpklgsr3yru46QM6mVEvquw8QgETmnJJo0m1ep+7OEx2Ugs
TTFvC0XqNr7n41wnce4IuH+PcX1wuRfS4TEsMrbpScidsyfPZYfOmmZxLsO87vLXxkHnZYkr1YEU
S6BOauBDGXXa5623h1Cshp57t4s8DC0QbBOM2M+b2EYbYAnw8InOfz/UQa699ZB+JeladAQpf4Pq
eKHP/nmFPbMOfXYXS1NVkOVJVtWDU71UZarmrKGE8w7du0/tg0hieawMt+/0JZajMe/r5o9BqDbK
XCrieIk1kfP57wkl8qGgapyJQzkqD20+lzg75yUZWcc7g1uKXiH6yLKmisR0Q4YGnzNo8KsJ+h20
Nez93w09GgMuTZE2DdDjFv19aLyK7QgCOLAJjahCP1SJguPOAWFKgEY04dUjZyFSsH1WkxZwwBF3
PXDIWFXlto1SdrFjfN0m7KLBqgqGC6uCLtbmgf+S8c6qrujA3kcrm2aDMYS8WJSUvXNCAdfj3r8B
0Jng49VyqeAQc5RZsT97RE2VMSDjFphh6yegeXLWDIPmpAWLhbbzlHVHlM6VCW0tcq2WQ5qVq26F
M6TX1/+4DWkstEf+LvU44wwEtEOWVNwxSmrsH1puZimP33U3/nCJ/GcK4Hkhx5c5088oCak7Gq9w
Nzy/4YWn/Ajer9ciXAYhLunoGvYIor/+poXy2+BqFdyCkEaJdo9bEKJ7jeGdNp8ipR/be0vIQ6ew
1iscc0r8z5pvlCeFeeZje+auyWhnM7pwwoc3qEYcaONyZ8mhjd0gw6FF0UC4hL8pmlG9s5OyorTO
cGVczyA378aIHfV32vDGpLGDo2/hK/VJyB/xBpDKlW5IlwxUQJNCGdkBHxeXn2AGiqaiCq18WZvi
MFuXzwY/ICbWz4++mu2HebqnvjTMtfxAEzdFeVKOb7YR9TyFHoO36aaVP2wkXfYqLEWMJ5gkLzmx
bM3Fv0VyIqmQwnzrRmfAIoJOT+nm8HiPFr2+/OqOZwCt9XK7pLuVCS/Rs4McBMZNQOiOi/4k1MH0
UFuQonIXMsX660aIeg2XFobYUQvakCXE6eyf+EMTgYOiyj5kEl6k8z14p7aLmMTkT4+p64FQOKkl
Ql4o6DdGIW0IfVtzwo32vrdadLVMjnTN4NnE6rD4oBgczRBP6n92NyvWhHex8fIv/tEj+xjZlfXl
7bS0TftOiqH9kd0nngr+/ZVd2B5rMqc5KCluL5r1qUteFCa68sVfRmn9+V1jVhtAJ/qigmiIX2N5
tev0t5emdXKHI/IIU1RcErVA+kjCw8zqhfxLyjvYQc20zMaDQLK66+BU/urLsPrSeAVzCzc47m91
pYnBGJQI9me/6hcYZ+/v9UjWhM5wcLVj1VqtYJdgzXc0g2Vz6A1c9Bv8Yjf758hSf/lIlTYiBmB1
mGaAPPYyx1w/nOwvxqSYa2JPAJ2q6xFelDyD6XQKD4xW9toPZkTbU8km/EP24UeDx14+28Vl8vXP
Dr6UNQagbQDteo4znuFEOcJZWVmuLgz76yOXuHtOgUpPQLw03YrYTSs50DhDb3zQV0VNN8rNhBuO
lCo3ahuXNiD0i0l6JogVAjUj/RiljJXIPR9rPlxW264qte3qbkbFtpdMzi3HoEQtVuHfMwTsSBIX
hGdCQ3TMfMUrNilWIo+DuxtNRKvEN1FpDgVUaiM6PKzqAxA6XI1ih63m9SqDZy+xGsM9s5GG9Peu
7hHgygx0c3SGCKNVPeLTwkXTieFFKETDMejIJqwJH5xzNEli8FQoPr0IdibcffyLw8REO+BdWDbE
FQeEkjG5QPoQ9cOxTzPugttJBx843NCzs17wsEAx0PDR0x6B6o7SUHoe0PJoLBY7YJD9XDolp8v/
yTs+ZZUHwVg71j4nTPbk06V1toJY5d/izDwrNYwnBpRJshYCIf7fvDl5VML4vpC3hiRLF7VmlPro
eJRHexI0BKQlEsMDCqrZ3Rrz3ZAWodIAjqrUm6CgifTB3tGbyR4gDgoU3M/J5cf4qUg/D23mCIO9
qBk+csjEExEMKWmUyw4/FGzQdtJKu1HWwt0BjSfPoj2c14kKHUaoKxV9fAuqEzIAjgyliP1dzvwL
4y/YUhO/EGFZsDrqUd8to74DRuHF7FU0TgejmMAyhUpGYNvTv/9UOi/Mjy2aFRqqeArIBrghQGtu
kjIMHyaRqhKlg5LAE7cOtwMKRcfLmTAuBpIfxLoOVccprnNfd4K4/MGSdWfBSsNbgCeYpofwBOxH
64ejtPX8zTzAaqA0rlOXqSjWayBNvyiBen9wr0S/Roj/i/6PpiZoZW4a87bK9jOqZbiwKulxOXvb
E0oDT5whpeWl0haCimUbdkj20Fm/CFi5gVxFFZzC03jz4HO/9i5nbm3P/Wwak6KONkRRXCnOqb7y
h0UKrChtBOG5CGLY4Ttn4elin51tuXmcDLnAOEI+TFDHZIkl1vuXG1tr2X9W/CWyf8tD0TLA5/hW
JREK0IxGuh9Qem2t+wV9/ExS58yYfqrSAc7PdtX1hO1igjSWXNYl2ObJGSbyLZXwF9q8LAPF5XL8
LEeCuOsaTNMURb4EdoU/PNSWNgFMiIUMZ53YwG2deQU+ZyJkldx6jHp1QOIRKPUIHsAP5YEH4sPs
lIxyKE9JkWv6x4R4EYRr2OsMmy1bQ5vUW78VUwNSStzsO8YK7MODt/mzZUwy9z9Mzfze3CPnbpdv
cuXsbeDW/K3OSRLGdXplEaozZPcY/tumtIoFV6FjNYt00pmG9LCfP249H7k2XfwlO+jrJLLuIAfu
RWd33Mph/GhWxnRzHS8eoIy7B/63m8POwdqXkthrjkDa9ChM8kpSHRRZ+N7HQq/A+m5AB/5nHE4h
UyQ0Tsyitc5sb02zhIyF6Sfvqv64vhMI5Ugkc3i8ak+Ix6rUIdZELvUHUzBxAlePCgv9c0Xiv8FW
l3pjLx6sOoXp1l/bTEhlbf5wZA4Wdx59k7XibEQXV4++wRig92L8/I7HhqGvQpOCGm3addud6Hsl
FLkrVeemDUAzIJtbj98P4C3gbY70skB/d1FQ5fUTDLiyglW+NtWAuRoIkaVuk56KJydZFhPLjq4o
5+K6ag8+sZSt0MJ3LlX7p6tTUEoNq+JCbwLM5CtGjfZWmPWco8FmyyjnAYL6NGnff8YQzhF+KvZ7
qJcfAcpeS2UppTD7vQvo85dgp8FtfAsw8gXAp73niaweJrKuQNtIQyFhFazgfCpI2f7L7lHF+jxy
RoAq8rdREA8yZ7Kf+CyCIkvuwaCnWHobieufVaQhSNbXQl86KZ8Relonu4ke+dSszYH46IGEgfu1
WRSxjZPJa24e1c1IshfQEhtjwSTeqFf1xXArrJjUctpgRvKa9BH3ueJZFMh+f8CLgrJyLH2MBMei
LIArPN9ZO8SFkHk/5q4yzR2ohGqqWgxT86JZ1ba3iBP/FNkHrdbYNRib0j+3Z2dGFy26E8DT44Qo
oZxZhIxaNqY1KtzoPa1/3Tg8/DByFb715lIZ3d/rWyyGld54oWGmmkHAbzWa3wgXuRIzpXoIzNPk
k+L3Vk65ovZkLWXE2UkDZ6BtZnwBQVnvtWLBaq/kmyIdViXXt8nmJe0K7Z18jttGeqanpMSRlOL+
CQqent79UgXnICpb4aHdDAwlss1xCtPDu34gWWMKoh3eXuazoDOeB/3tBahhwz8pqmgKHOym1/H9
mIOKSl4YmbucXBiAR/qy/GLL4fQxx6fVVTR0kVbNA8ROtoXI1z9T+ENRYp7N+lQEHJ1jLFt8teoY
uJVdzdO2vKgkCTJSxh+d6AAiu82Q0pv3tPOZ685EPd7Mli1LugOuCh9l0MzIULMryeyrpePx3AVV
+mADl/dHOjDpDpHBcCvQHBtCvONVjdUREAefoRUOTP1mjB94ZAkVVfQXoO608FXOO3wnkYU+1w2U
7Zt8e74kXiPsqDGVAv55dHXkiYhDHkJ+uSVvkSVkxJf3GnYRwJ9TbI/UfJJdGqeIJt2crdT9Q8N0
YeLU/12/JH9IKjmHvPiwrrla2R2WkHK9qdO7GFpqPXGba7pptI2dOeda2dkuKXZx1VIS/xdCxrcA
KRdXi0smmz0/CMT513vN0UngX4lyvtRLBHkU+e9onlX8/3QUDc4hsoeJp6RKOohU2L5Cp6IXPOa5
udCOhr6KnV3LJHLrQLVfxmkoG1idYeeBrvA7sv5YJYqviS/vSWFYRiBJCR2af/zyrh02M/iRir/c
i688M0U7XDZ8zKKanWXerIip9HfnDLy4NQuWtwRjA9xj7+CKbMTJ75+nXXl/5fXM52k6ynstOyW/
NpkHni/WjEzQctefnjwLuw1Tg855IZs9SpTWwtR0HWbbiTNZPIiykvl8NuSco33l6by3eGQlK6cX
43/4v9Ll+8NSM7wxF58xXxlxOFAC/WydyJXSAVzenGe+GGpvluqgpJ8Iu2ac6so22oCfNMCcza1Y
W0WSQ1tgUOPrNXStnREMMdCcBARJ37/bPTZkr2LzTQiNpjCjEQqi0pWlx+ThADOVoXMftx93m2P4
AW1s6/uVhqwfXjrEAGoyuP5O0gJg3/KiJDq1KLt8q0yhgaVF4yBSuak4fnMpoWhTcQqNdXjNy9Ty
KzRggw9n5u9yjRmqGGLTijpgvrTpTeocSlr8PZjfPtqxZh3kpC7V7wS96AHK4k2WkktnIp0d8U5N
nJmJiM54dkLbqXCHtyK1cbOH0JgRblOhGmlu24sqpFaIMCyuu7AVJfvZv0iWRjZE4a6eAvwAHpU8
WdjzNZbb4cK2SzIACXdZqBs3LKOhQ8O02O5jSB3JqFNdLRPPhXXq7S1XdKL1AxzTiLYyHJ15ALy8
HpQvC+UFERbXgejBXrV2AMxbezEnbox4gHwhhYTLHagJMnIO6qWDj56hNIGuvrorv/IFjmTZp62D
Oot7aPUAXjqTtR8dDOGGigsCQjVY+S7eaGgSeCUkPLWHeXNuG+NJKtH98Zdiy4/PvFTzRorXmeX5
CxeF9ahUnCfLERJuAECB3a4Bzte06qOdNVXJeAXzngF0RV9hirXVH6KuJRHH54Nn6l24yE6nETWf
Cd08IYHSTXa4GIx9tjbGrWsMQ/XflASw4PiiImXVLJGnIker15e12nzl3fCpBs7yz2zGI66WlW2t
Ye4XqShQIfwp5NFDU2z9wcEIpEyUDCW8geKd2zeoTBLgNe8K3P+aZJyhsVIBhCDVNyOx8chHHP+V
PIRHpETzRnK7pkYKFhRZzUEUeYFvhRTjXseA7bQMbB6mnJ6noMPRyBYYZWp+5LArsreLXqSeNvxv
Xdf/s+Dfklxfbt0BSdI8hjZfNzjAJ47VFXvss5nig96kQLBbCC8ZNQgUA98IskZsgbhlGtnyd115
1rubr7bElLgwVQppMdXNrjb877sW9D4wNIima2a7YE0clqT8cKHK3DCb6BAfNRjmIV0HgNAOoOiQ
4JE/+8+4oCPy42T7GgCC5VhyrVPU/0iXVPdHjA9H8IUmOxb1L1PUcZgQ89A6V2wD+45so4RiS+Qx
nqKXOXVMtDUIrXQQGjkcv2nuSDAi0MDy6a4czs4Vab3uGnS0pEsbLiLcV+1RuUCJcPar8SKUlVbp
1GyBPF+pfYHk5JjpRvvyVpnzqYtrRbRRpTxfaoOi6JddFh7cKNYgHItAZ6qagL4u6WREDjkN8l9l
jOwwamxDFp5PXJHLUcTzgLrpqdukzpfKcnNRdTLbqT5VQrCWWr0a0R2Nemu5Hi3Dgaw/vnsNhElR
Hf+AaM0HoT0TlJ5CRFtAnHngLcvLnUu1yupR3RyW2bRiK/uc9SdByvERtdJG+MTW96XlVWaCHEWB
0aEQB4TTJoB8lS0NPL46EkpYYTribWzycwRIg4HtCCZ5qUGhFcBS8fYZDKpU0eKoEUR2gzwW7tJn
qeFT7fMn5wHYcrpgVcPJ7m+0MpHFU4OtiGwduM85eAX2Ky+xirY73l6Uad6Rp9H+MkmaMI0bg8D8
/gjacv+YzuuRhOVPiX5pcb8ET3XrqGfgAW0lzzXWkr+RVwA0CCcErHrtdoaImIy6wtxpM1ht2LSa
RxkmEqSFgTfPLVI0K2bMUSEXyvuP9FfqLdjqqSVN+DojozfHu2tvJhJ8idE7wARMJpdU53IPhviH
20TiWjxp59ObcgC1WNxSyZS34/QxYVU2qUX7CH+CzHwUCV5PhZLlL9xz4viFo+HpjXP/L6JBqBSB
tzTa+YXC6PgV+Kwke7nVrJ4dErsYV/gJGI54qo53StxFPHU0KL+yieyU4mkBK7aSKNO6KiCHwezP
zA3PEToUTQUOqQ25pNiZs8b+y4nfFhOdsP+iGmLo4P+F7MqNUifFM+60TnFenrjHYKFnnot5jUR0
sHrCnqwVVfoceolKPwL55NkQVST9okT0wOO/rJgDk8c6E9ku+smkdjBUuNfLDPPshjmuGKOWHeYi
393JUUO2kYwyDfc0aAgbxrJzUo915OJ9pIucnKZifQhUrLt5gDUavMC5U1FJ+mVO+yiQEhptwElQ
3uGE/lcMcS0mQhfdoouu9CdkmDxLIX/gA9MwgzjRIkLEXwY25YCl4LWfKLsgZfjClkaw9V8ncWVY
LKxLUJC7k1l4vNV2As7BqQDAI6I0Zj81PmONAta/zEWH+bl3EAQtM+0IUYCd5X6pWzjqWoN/7UN7
5d/SuQ2C/vSG+By+LhmX8KsowdCPq8Hy8U2ihWtgD9zrtue/DG08RIELxVOBLcStC94K1fWC9IM/
6zcru/sNEnFQF2dE4NJKxJwJKbNTCJpzDi31V225CE56ype1m3PcLKQymW2uketPaQm3VKOwR1Ce
zqC9hyqO975s3rl6grDV4U1PJHLBAtRVwRk+ylLIks7TiiyrNSjw++bfKnPgsRXGOvSgKQ+XiVs9
LErbm6Bu2IZh51YZAw0A5Y0Auvzoa0N1fu3Waq5s7nCcGO9TQMnGuJGc8f7qaCVtiAA/rHLBw46h
vlMNQ/yLANDc8SCu/SEyq9flShZMgeeIsM3dW4k9h6pTqHbZ1pbMb/CDr7K75jzO+3GWFnEmMeJw
Z2fyhNw2nxxxBBxE4hbsPQLAAcl5n+v19G0zQ2m6Ekr+wIKTGpI4XxAbooVmZmuLRD5BXVMB2aRC
Hukd9EkY1ysc4f0cqTJmOO9dqimH6FQ7bHKPefQbHVzKmi9MWaX13KFOZffX6Bk0/g3Q+QONLoij
bJuY3KE4zeF0B5TvAoPZwtkCYrU8k3FKdCvFbmNsEV8Ce1WLgrXbFhFesiU8+nHVrDIaow6Ri+p1
AymaDra0hSPP4Qk1veC4v6rskr2riJ5PcWH1uBium0zk2/j4HNjlHEZwPyC7O6RKQs69hySV7BOv
gELyRbErPO1bQF+Gp2lFCVmD6Fl7Y/wI6tMQimlM3figiY7PHN/NJbrfqENStqAGDPHC8276G3IF
baFQOnKFTiocwoAYHS61G+LTcV8w09RZxtk/rUnyYDKxPZUrpEH5gxbgvCX7ZC/JIQIWYxTpP15+
yfPZdFiESfzztxeri3fzIxcMp3AJgd37W2zSeppdOOrRiVhNyGJNFAx2/GANCIPl7/74mn3k5qpg
i4mUFmc8fBylmQCgP+a3iz8k58RNPg7QGCsgRMGzq+wo2uRjtJLaWqEDWQbC2DNUGTQPZ16tURru
RKKgNvHkuE8nOawYKaWJH7ZsMdLpqZSbZ9EhRUjdjeuEcb09pTF7+mPwU1h5Pu0/iIz1IwiyexH6
X1eadNdOFxxXKvB8ITja+X50HlBVRl8c4y93W9+wgQWnP+9raT4HU2aZhYu/coXyMtMoFAiZ2EMf
Yw2IZAbiqo8FBGmScTmG/Nt7W/2vT6jfi/Fq/T8+NQ4r8gaX6WAub2s1Zz0V6XImOvPJLCJ7HrhN
gfZmH/xDTPtSrQMjhTWg4vl68cX6wS1JrD50jNEtwcmMTH60n2IeK1zT7WNPRm5o0MvVYR5YVSRF
m0bltdU74ds5tORmPTIkcH/y+5BlOjOhOjqiog14M7wKzvg57bIeJAlLIPSoPCH5uDO9xKbu+tn6
TTlzvN67IXlNCEptz2qUUCiW5rFdv6eDibBqCb+CP5yq5YkA//8Is655e9cXBxgS9zDi4OPM2nvc
CEQUJ2n3eQlt82s1MEsvM1mIVb0zanGDCSH5ojR4K9GgFhPzRWKNiUtCyeNK5+5IBuwrJA5K5ZHB
T8XX8JB8N4q9OZ8t2LzaHUOHJrRO1RCIHYlbAQpoZUZzzYKsjDfuTWyLuYcFUH9ZqKYtD5PSyVU4
lPlASe8tBMyrlA4FHxBzFLMB3UulDsfyVeYTCB4syfD7tH/DPA9h4I7TANl1M17oYKLwuTKfADo8
XWl2NItbD8252u3pHCUBIhl9Bnj+fWDm5vVFaRFFLlFaB2iUBZU7CFVe5wy/squDS/YPTcKWmFlW
tJajKP8b0jCvtI2S/dIqM4NQmLzjemDkPAYuH4ePz+hLlq2yWN7ce3Dc1WGcDPB7DPec3f2Bn3xL
aqOMIC6HiRdl80TF8+gvu47pTt0KN/3zMASSUg6LfgRsgtnHnLj+2EpxCGZNh7NirHb+D8Y+IBnY
wNi+QZV/MTtPKkkbSHk5Sx0xQYAbXfqYe/tQSdtZHP+MOyZ1/kwjp3dQrkQzL0YZiZ9UIi1JEG+2
0vcSKv608VETAP2WAZD/A8hKKjV+hSg6POY5hBVf/khTiqB7yXeZnCThseJqD/nHmlcCvz59NU0B
M26VbF672tn3zSmNmdcRCGbtFzDWXutCJpqjt3GuuH3WL8dDwHP4PMrPGCpQYD8i8nNyXRU5G/c/
xOYTYrQdc5Z8AxSc6EywzcEGyBSJGfJwbBa6P7thfZUAKAlE5+BXlv9joMcBcN7kt2Nuo1hKqx9S
xEd9nUzmo/PkAtoEpRKhLBD3sIP7WQibnjm0fbarZNcQB2xP95iL+3LGifLagXdW835NSZgKRcyu
ALm5JmHnlAtt93YFguWveTKToGDpga7P3DOopKv+oB714tK97pAEXTwjRV07p89j9nTwipNknPJd
/CZ8qx+CyyWT/efzlCIx5lflaTyvstmSHc70bdICNUVK9paMaP4osnPvd59zDAj+kcqjssSkR6o9
2IMOUMMGrQ7s0UZART3QZ5dagym4XBHmRe6o3SafDud5vCQy5uoqssM0oVkbMjHnhgnN/N4IY4Ri
pGRqiB+QX9FHD5EdsVu9n5q0mRdmWv0aIkInCDD9eo5mFl/yKim6jwCiFAUu6AFOY4kMRKuBBKTT
YbzGnDD7jH+IKzOHTTF/nZ+WhX9DbdXbl4j8WGv8Ak4VVcZ+9caV3uX+saM9Rsy7+JypJZV/tHkz
MKqEGThaWySsrDNLqd7DYVeyuufmbmMOoCPkUZQ2wibcNzwKVPCkzD6FaK5HowM6C3F7ETtTpUKN
XHDH9Wx570sD0ZYtjXDyCyQcG4EG/okTPVii/89kaZvoW+KNyb7xiXOPKEqe5SjIQO5MIrRAD7fw
K2kCJ61bmnhIP/MX3o6/SmdgFtx3EBDOsJDVfoduaILTZqUZgm/WukhYw5mr2Gq5/nUrw+P2hbjJ
eZ9W7n3aBbP57Tao1COoFBL0XE4zscI5nYd7q4inWMXC7t7KwMDz+bofD+Eh/22Gp8/0N1f+dU7T
8//fkcplwqfLLlVTS429B8bOsMWYukHePxEkIbxByIMxFtKfnM8cIpDjf8x7vCdousvi0nn3sxNc
315erYCtPM11BHoWUuLaoSw/NOEtKO8t8FiFUpJm/DICcKihijUQenE2ioCaZK/9Epje/HojKxTj
ypS8Sd5Bza6eMiunEKyFkcujTFxyqoFuT4I+ZgGoJwYETUvuSv6B2D74hpiG5BbsZiUB3uti3sJb
bm0HhacFPA64ShylXCRH7L+CcOqkpTGPHhMxoUjkDWEdTqRkBXbpm/jsrvINwz3qayxvsEpcnn4Z
UzrDXbFmdvjBsLGSe98ONgikQxelaBHmsbDGsG8aER3KbZbzuUhiNcfUMHd7XLIJJh0D0O85MuCT
HKUCGm5DTBou5VhRUM6GE/DAewXmyTA41nUdIBvD4IRE8+Fp/l4exYshxa4V+X2lSoijdxxBGiBy
1WtjuaPi8QBNG+Bo7DiXksEB6BHERmTXMjMfqsewqZ56sApkH7hmYKnyStFJu2enldDG9EP1pP6P
kEHhSbyMbUD9ufOdtC5T4Gza1vgpZ918G2Hr5lC9cC5MhHDvPzuuy2sI0AQN57kG3KzmTl1d3FKA
vJVORAX+IZmou4n6XpcrtELlJHZFFFM5gYNxx7067/l8fpPcgxoQVZGZo6mtmdzsOdh0XEOi1c4h
Ot/MJytIfGsEkUVwDqksBCTQxyTAoR1FjwkhnhrkyOz1FS8lDefUOFKMDijWKyWf5R7XurZrRAbV
DEkS/zxaSbHUZ2D3Fu5GryrZ2/2whnI2rJht8U6LcfCghCvKLvudckUZvGg4ya32998JZdCfzIyO
BvXaN1c6bRIjr2Thbc5XfQkQgPRX3fws94WSiG9mISqnsK74iQwKSNZXz9dxlKLEw2+wEMIapS7V
Sqt2Sn61Tst8MW3xibM6ixiXEdKx2dh1RBFhDkt6RkUVheY7HAb9Z+ZGEV8sNc45kgxBq1ghWIoP
HxuVfuLokARRoYeJfHABF2t4+z0e0AjAS3xtD+H2xd2zZ7gdQ+LHNkjAHd5E4claxYZ8uXOU65Ml
QBjOQBNdcSKgG9PZL0OxiaxbeEZr1s47fm2X/VvrMne90L2VJ3GOHijkSu1BVCRNlnzzFCVZkDRx
ROVKboc1VXgCSiWGNrKH/QDM5grFXMq39/AlUoA7jWzvBikIwBzKb5GHp1XlxjCM2ZSTzbaN5tL5
vXTNohk8qUNPqwQ6fhvrc6QYEpmQiQm6DzuzCEHb9BDsvHhn2g/szMWPkVmsf+oxxpVPoUx4KnsR
bkp+/2c4qJS4B3sVdgZi0UjIe7hpiC0zogF2giDQlQIBN8xITHTk0oimULKhicshr5iOr3nOZcsf
h+T92/imG3FEtecuJXFHnwQocrbVaQUXiQu3aECHMjBt0E8fgpy40TffnKKtOV8pQr89iPT+XNtc
zv2pZkfAQCqivgVvidcpGETyBmt4Yhtju6J72Yry7B1yatNnIrzOH9ZZseAOAwehJdDGLY0RBuwB
1E7ulz9dTj9FymsVuNwxxADFpsae6Rauket/BmJSwjWGspAKeobiiiKDEkbxmAaA8ErJgLSPLm6Z
amEI2sxAF0JZpQgFdHLDR0ZQh6hlGEhfXP8DL6rT3UG06EMoluXPXawOd88LJwDWxwwy301gksVR
B3/7vmEnLfXAXW5wxgwPgAulhOo3pHKj5aLCfA1G6TPjQB1fIMdLCFD0oZyunPjy32qfIHrTC1mw
766U4bp8C4f2Si3NmfKGu0clfYEyPKVaCS960sB3Z/mcPQWZXbGUhArMT2gVq9iRTxJcmmay4o0X
rT03xYOpuKPhmt8VAn7QcbeGQcewR/fy/btyY6ntqP9sf1yxpNkFjiU7NSgJgYJp/1vRTxGswmv8
vluhV9ohUaLKyirHbakQSHkfRMK2C/WDM7Vof+FZ3fUHOzDS5g0o3bOGlHbCW61KkegSoKtOWKTB
ywtuTrvKsw9zBbBi5TszjPGC96Es1bdvR8OHZOcnxZpAPuWqe7DCC8KI+9ke5lyj6wm5ZUDVZpVq
2X/bA2nKaGXoXkIUl/RplW/Xv62HD4VBI2F/pnISPYiuICKPPTKcaG1nDvT0IJFJHvOAL80aCuqM
4+QB2RV71e6x2kqIXmPtCz6+S5+fdB1/1VEtV/+vgowNoO7Xi+tYdz55kDVKQ6qodCzFqX30mfdO
gZfo04ZtQ4biVCnzPPGcfkcSsWrYLexjTmJ6SHRO8XBV30vUbjelbN+gYIfr2yjV977t3diamQ0V
sxrGlchi6Dw9RcS+fyNKA5o8lreJeNqPolZIyHNR/hihcr2Uue6d7ZqWX/RZvdKMLBNVZwvSfQS+
km1J+m+jmZFYL5+eTDbRLYw8uJ4drT8v2XeCo5pttOddMWPMTiCdnbbkhaQahg1yRAgqdgge+ybL
iiED0SvCOk2Efr4T7yOdty8fJoqsNrzrrlNZYwoMksQA8S23IhBB2Hsj8qEcTxBS6dD7RYsaVo2T
oY2WN0Nik43nTA0oBLStTv4JzxRcFVpuB5WblvdoabYE2zsJbJozmy1TguXkV6hwoen5r44batBL
EmqxWiDw9joTHplV8u3dBCpwDGoM52t35BNnuom5oXQ9sTiT9C/EmPzXYY5D2Nsot3Jf7aBM4Unm
fFrZBiwZ5KL0pSNtjSpyvKl18ZS8hgFiIFD9aZ+gNcXxsCx9EVCORqpIwBe6smQmtaF2ozSVELUV
/p+0BcE28jpSvu+3AXhv4PcRzvpf0CcEzzHVqECx5M//h4eHwOvto7HFMunCvlXKitqEGCqkMFkb
DN95ON+WAOW+Uiiops8MWVSufajdxOVmXwh0uIoZpAy7sniWZZehdN8MgOVCYQyg3nTZp0Yrs3cH
Pe/koqK7BuV3NreYzWbrq4zhXIAKFwsJzRlduAhRuPNVdStxmjsZq7u370s7JneHc7ZVf/TPF4aJ
choQ2HrIvhLOIdJ5Z0mcutR94ri/RcGttorytQ6IjHGPOjX0fYmnlubxKfCoSH/o8dHwjEf5Xkjr
t1pPQpqDyBWkJ7jN27U1vD5T9bRoI21oRo/G5J2ckPDG9O5ptwJrZ1vfhy2C6rDkIW3CEPN1CvNv
ifH2eew1qYuTnmOl+Z2DoZTeXP32wFu3enY9C2W4/+jg9rXvuIKzlX7/TH1JW8MgQ/opV7siTZdM
jvP0r6dEw1oVDmup5hh4peB3km92Tj8pXYkuorJLqLkcYO/VkquSpdDsp9aANqxil1jFSReu4yX+
n+DgPy/ChHgH+mKU2SohnTNiqcaWp7R8BD6P+Bx9LU7Sm6vjdejiWRcNFMiFqEicaGpZoXlLD6hy
LMnWhvDYk0Q3TxQi66oAG3Py9NePjP4fxEapMASFMqN/fOJv/1kAyfFtWNHRtX7YZVqLwq06nf7o
J/vU19ReC2obqB2a907AEbDfga9Elft+W7Yh+d8yGTdtfOgGVqzSBS3Ia4NHxkfDtS6svXEgtZS5
lbxfzdUF4RvwY1iAqhYmAgfzpY2hV/AEIyA8LwI2mos+c3xz9qhVv6X9lCoOHi1npvZY1IF440et
vwz7f8L3Aek5EDO5DMcYBYFUVLj9vwUvIACKUAcLnLsp8wWNuEElrETXEF9hRiKSKRecqXIGHASY
cBtt80PA3HDFdC95SDpjxt0cbS0UizCnFLsPwmLGWTKIzRudLRo8LXPkDRla72YKH3rKjI1BQass
cGxmEaa6SsFd4vQkK4F4Q5UOey8eYZI+KSVAMLh/CAcq6Y+cDRY1WAiqwgOilHhBevuVkxc0o/14
sb6N4WV/SMMp1O94akU0PCDiMbjsv/afBjmaw4UOKY5PQfKII+imP27K99OjYG+5t6BmmCloIruh
O4JDRNnu5X6FsMBHGfqykgDeG6cs7TzrMBTRH3gbQjV1AGRxPUZSOg4sRyKC+HKw0FJNifsMJuBH
uYmvjj+K0hJK5rkACva5kWpdIeizRgoDpCyPsVit5OmosptrpUmzd4xH+Sm9AmK9/ZLzCZgNw1JO
tMRur4Hsx6RoXPtcxGbBwf1o82BbLWhGoJb+UfV1/4nHpKqr9kQTeqQ9tAEW2QlFzC2T0WWp7vw+
wGXj/yHyJ9FCKmSZ7k7E1QrT5WEVtUbw1AFPvDt95RU0FEi+KQOv1cVGsx60kbYVXtNUxv6NToHG
0gc20BPTrNoxtphKmLla8PHfsuIUiKMayd3Zp1/ZhiDFMhQFVqEE/WJ42K2lZRVQVf+R8TD5yRLb
5m6fJL+PPpwGMTxO1jFI8jPuvyIp0N8sbmTBCjK/oKrieHg424r3OF7uSMYcLOLa+tz7h9p+jAYc
jeT5/klFz8lXEwBNuRRSmIjQLyxmjsndblcobFKOaJ2u+WOSqnLbh8rpaR63X1iL3za8L5oT9hit
Bkwvnhzzx0UFr/Y7+4EFZ3aErwXTyv1J09flmI/FC7spu7oYC2yYqqJXtwJHwVDJK+n2/GpkMj1F
1CpHHv48E+Xp+XeIvXjDdolX1fBxXlY1MC3/Z9jVDWVzr6LzoC8mqZpJ25G2CV7bOT8k6gFcFuCS
KIzmrC3YTl3IbIYZjopakZ0O4mJHSQcUx7yp9kCU4iF98JlgYS1AQQIBLVrhIbRGbGBUfrBWFlGI
l06p53tsOCBv+dfVvU0wos83e9T2MtiEsUl0XQLe0D6A8VEA6QLy3gEboy39WfIzIahuh6fMQwWt
UFcZQ92XraSXjlQVVeL09zM/pQXDfKLQeXMrn0wDMvmhYbwDm7tsWZLRtA3sv9Kk/WOCkqWg6YA/
XBHERiV/rBxJnHwCR1lJtRfCIrBQGBEqnNwjcfyJOsRLfLH5WX25u+kv/LYNOavBodynL32pKzKl
dayeBq0/+R3CFh0mzYA01ttX5/qinUjZxP/oXqVjNVkA1h33Btni57XFsmRNukCeO7tO9Y8AfRT/
xET8Lyzj7ni11adiWrP5DQViNSJ8Bocb+eSZyWgEjMs68HhfZyRjvITuNYkx+IPe48Gjn4aECR72
eyJqx4wzQJo1on2Yv1ZXkgPHkNjNXRN+dMd8+gm9uitMBmD83+SEqM7PjS6hJZ5rBAA5diG6U4fZ
d/ixRx7LNrYIjQxo9aBlA3KhV46Z9GonSJgfckQLOQkpmffUfOrqcVXXxg8p+RkzP3Agp+kQf5Gs
XuZYTLH6JXqZaxyYmBc3dHQiQ0+Dzns0CdMfGfIMeKmNWrQ2hsVOmA9rRjbyhho6naBG+D3fncIF
+GJ1RKK3R7qSi+ZLOTMgGXsunvwWsuBVoxx6jrS/XLbjzZwE7GHAgI0I6P1DykUS4I5iwlTatQa1
VSVD5opfgwfJTFLfMcwU7+bqgStntyi91XfQ5gy0fSaBJcRXAoPhHqBgMmMy7xOOcoAguyfA8nLd
OsXWx2mEMJM2kiyB2Y8rR+8/RVN2C77OooHXcnDRykuqv5CM+PPoYqJoAHH8YZzT6MixROSaVuVG
J0StAxWHckt0JVRPVu0b/drDyMHqtp/eEnw6ZJ4AZgIrsD2dG49pBrEQAvXER1f5X/XtuoQFwlpt
nBEbQTyyh5dEc9yuqLODrJn3YJ7MdYioWsr1/DSbcuk1uoRw1SNzf3YvS9Pc83XIeU0W5qtvnsBk
sclhqZHx2b0MGb+MfxrvNOr0l1oSTaf4Ahcshwbm+1jro4kYmKMHdCLJWPWxdZNYPqlREQ//EPGm
A9ygI3fyPGAMfY04NOIpWcO35gOyYT6Gjo5QC6iO1hjraUarUt43trr22NF5dk3rBDRvGnddPqHl
w2+i5S/KC8RE2WkrJzPnEvhOROYZdUa8CVNBhaDP2UCCOMwV8LpzJpwmA2BsUI62pntvG3R1nsTC
gbvP64MrMGhta2f4kFmWlABHPjUEHH7aY8WUJPXeF9rXM/ywnAAfgvRW1+g1MxyULH+nawyyQZtt
spx/Sy4ejwXckCakQZK0woXg7rvvplWhG9f5pHKz388CUVNa+OI0eRCjhzyAnhyDPkSYJHyQlm6/
Z4xiTEFh+ohqVrrc+3QQMJHLwNQHLRHT+x//k84PKzYPTzKlqmyyxTKSJmSVTq9K4H8v2aHo8R7c
D9U3WfXILRaDH1aYGB7UDflQJQyBwWCYTOGN5nlrV82dv12P6jU58MYdDHQuJl8epMiu5psm6Y0+
sGf3H2LOOpG2leJV3kXFp7xyc8LEF/zWXvBdNxX2z8mmYDJVZl+B5FcKWRk1v4LOSFJJIOZce51T
GzzOyyoYpwogJeHzQXwFAWWPAO9f8yHWPfCzSIRw5NdB2qcJ5cp4bFVPBuPE9VwMYoJ6mZBYZZvE
qQBS4rOVaUA43GWmUVQp4wjSCpIR0NwNc5HN+k0+eqhORsvu4j830GMZP6ltFtgUV+TqmM+iChB9
wSEJ0aiHxGq8Z5/ff5pOMQpgo0+4fSq9k0v43WgElMw2MQyrMVLAFIwfdWesrJVPOYvKMQCKk6Yz
lsb3vKaN4TjvkcxutQXfS6vwyJjlQQf7ccV/pCrNZAYEFPgVkDoQbQ9Qm0WCvfxncFQ/7aXxXYg0
hphnzo+Tl6Wr5D+UuT7dx+VTazofxOVY+HVlqDYcV5J7uowDS+sweZpwmr66M2m8D3nrZYxkL3aa
QvV6UtFYqy97H22nIhuwx7rYVZ41uTeDtfeyCQLooffR61+HiZ9F9GD0EyiTQqUYFIemlfx2r8ju
ej+bhtQ7NMhzJ1x2b2b/9oczuZLEw+UJMWoTiC1gS/LUZCo69pL30SyPiET9o5bCQFrhwODi8TG9
z2djh6jWuy78YxfTXhPBaD3NmGxBf+QOaPojOReyaXWgKT/FnfvhpzVnbwDNiO7c/ug9R1ZlcK0Q
wg4VoOGUoTqMicKEWaoaWZxKjeuekF5qMdEmBIBAH2AfJueqJgtKEjDxxSgGFJJh2VhPqK/y1JwN
Goz7ev78djGvLir0v9UNmeax1RqoWElVwd1T4V+Peq1YkG+HokYtWXUv8SFobKG87tj5YTLXsZkq
D2ia7E37+bU2a9norEkVpXHwcoJL1xRhTzmzdeyxO+Q6VKQu7dNgmnKbc1MGCHqHwfLqkR0Vg+w9
HCKBjG7w7r4wsSYnn7ktY0gIneNDn18YtdVVhmwrStK1P0LDqdYsIklbkKpvtORlp49uCPlp6zOM
dD/Qzf5uJeqQmggG++Mt0oWJ7yMlDSmzWIjbv2ODco1MlFRRuhZDj843ekq0NTHTORJ9NTIkmgph
GBP4Bd10ggFgmIMgIMyB0SUUQ33kxyEhtZ/23knqJlz+mp+7UVrEZclfRkRt9uf1KOQiVl2QUemF
3fFGVCGoRvuurrWMc/JHuDMSk/M34uecfnMx9EzEnOIONKbMQqhbotZ+hqht/eEIUfZlHjpyFsRS
TI2HG+zyNh/vBaKng6QkKOUbKF9ANVZGxoEab1ZhOJV8lXm7WDdIN0tRs3vmMJQSX3hqXGl6Vh2M
BJKr9Wi9lrtphuJ0X3RW6UwTEbLQ/5MkF7BnD5D31S6zgoyKMCtmIaGDdM9tzwLBmEBXA/qLX0AH
1Z7ddOBsQxwbf6/gQzSI7LjHXJHM7EyICstwaZEPyhDYpD03UxShvbXGei/35xs2ZA4iILcp8vGM
6y5AlZVff5+k+UNgp++ik9Zqu5mirhdfYcBKYqx6DAMIvJvuf+JwmDPLcRabRiyogVw2SweOU+QA
nHvu2HpR/5k9GBcjv2htS3lYtd746/3cCQaNxXOxSCy77CwCGCULnXX6ZxDJZYUgcvcnQLTv+sJM
ashzJeYAgJE0WuMvR8Y7VKXGsLbh1bDpuMrazcx8FqRhSU6Oa51jjVPwMl8gE9MZWHQNrp8pTLjQ
qJihEQpFgjSFuGxhATuG4TuujH5BbtigzpeZ+PSO/mGgOMB/ZtKAwmVQOElMaJSGic0VB0zXN3KZ
bfh39xPt8yiyMDl+LmtQQmCI+Vh7IZ9kcn7oRmyyoRxj/Oh2s+j2YtRugOH5KYyyRPi0q89PZXEd
QL2QW07hp2eAkMDvmazT20n/GxKLj+H+/psm96xwWbDS9AhWhSzXQW9tI/9YTR1iXTKf/T2UjME2
WnqMSPu+SRON6+uIdM9yqaK+4JyJOBvEDMHqoZZOy+bfSmgaJawBBnw+BUu2yuHiZlfn42D4TE5v
RJQmG13wWDyxzYF5Pe8G9fC6VRIm5XPaahVhzbeg3yTpWF0CUZLZbSeg+ZV6yiT6eMzo0jGl10V3
GlNGxHP7KA4Mie/jaaWFFI/rC1id9wG3Vr7qRL26DomFXvhThkdiPFZtrnG11C/5E7rEL4nGwIa7
88FJdj8GV+plvFF2OYJEDxPA4RJHlP2gWlHeUKQQjD7/6Ow9jp8XNhVKFU7AG+SlQjeGJMpUpjQ+
INLzwfzHZyoyka31JpPj/iygHyj5soOr3kb+av/s5INF8cvZTnorG0HEuMMS3BZ7I54/fGFLHOsz
5L8yUKM4WpwjfJNDZWZk2I1x2oOMs7xDp17cy2Ecb4BkWvriqgBNWYioTvoHeRWL9JAxb9kS2Cwx
3eLJUa4vlU9fnV6xGwRBnAgWFBuWCiux9+yz2oD6Meh4gH5I/B8QyA41OMnE8+0RHaQl2v54l45o
/ZFMF7WD+oONE/whKWS111foLdwYhDRLkcndEc99I1XcEXC+sHpvoPcHSKknC3g/LiTU6Nwb2Dcd
4zA5ttkHjWYmC/v/lZsscjv1g3DXR+IMlDmb3Gx1lElSLmY1bbQQg6NdrWBTQIkyC45Bd0ASA5Jt
TpqV4CZWOIYzZLpgD7Np3bv/Qg/LTFPWzivEEpMAZfzfFh15UblWDWLIHfaVp/In84rbMC1Ivt/I
HELT/LlMQ33vYRqKxbEv14W+IFrMECrZ1K5TwiZGkrBMELgS5luFVa7FHznT5PNQXy4ukcEtbHXY
Anufb9mxIrpIDKEhlmWUvb22gOPf7PDaSqVQk49BXygsK2s2LDQh+BBdbTY1sUL3NMw1A4nDYr+A
hRgaXQwMb4OoMYToNvpea1iLobqwGUdGhRsq13V3ebChGtG2JBqPLVE+6E8bvBTDqNfC3GWW7ieU
ZM3aiBMyaaCuN0liRpIKCGOBq2TETY91NxWN+WC7ENb6B4FVbDa/jPwI8e9Hyth4ZnYisKDvdtqX
AXPmXaNyszDsZSDUhOqBnM6IlKE2HUdgF/lQ4mTJlIDSnSxQbTn81adl/SpA1bfc5Jo1nflQ4s8H
mrCiPjNFkV0KAhDf2FXbxdyANzpuaU6jWgAGjSsEH81YXfCvwCH1q0TgFVVXZuFf+tkXM/1kXSS2
FBG058P6TcddW/NTucMr/1o9C3mdC8qBoyJMegSQPtOUnrN77JsSVIATtV16dbQOgFXy9TNPQZxT
v+1/t2Ws9w+oQUit5lW2BWgpFWUKMindxllGeAtAEOWQ+FHDHpjkZVwT0jEFQhxVCuK35ilDTi/+
/oVSMkB1p4/HronG7WgOB+17oWb1o9NDXe53QhAC4PUriSkfsjD7ri5TvGXrfPbCfImDL/6LRpyO
o2e8TS/+Vv6Z2IfZSisTEsBAllxlVidrAiptouMppoBIPssO5ihvh95v1i6Sb+nE/MhEwog9fANV
VHwp0UkyFIaSign4Cysbf4fYVtquj+lUZ96GUsGb6m4ZTYj2msF8TXEeCzjcBqtxvPPIqQ66pyLN
HIEs8TtnWHGIgtwmlWrsrDcZWDrCpK4dP73GMS5M8KdSYC/RCXHBTG7zMztoyg1gZSS3e5OGJg8Y
VV8yLYmOzg1Q/k1AOvf5nq0BYkJ9Fs54x8BONzbTFVK+xW5F2CH0hjNdBNnOAAuaGl4fehf87NPy
fUhkY9ClGbYhSoWnILO0aLL9QouthV1A03xaqvuL4BW/MCSnF7O0N0Nzwtfi/Z7hU183Rg+cmSAp
JTxijYasUKzVWiNOHN15OrwX/GnMJUAcEmG+ZTf03gOfVnDTQQjLWKLcVKNV5wkV99rxL9ll7t69
BZe7Ke5wGJFETxOI4Qk+873jjZnHVhQG/knppVC2YR4J9Cy4Zo1vGwHlAEkSkdlqmH+obz3C3N1F
BaMBcl07GSauwcVyVjdvHSs9qcd08LWWeysGdUHYPq7v7MHv0UUQSGPkgNKZxoRK8Amf6+WkRWCk
WrYKQIMZeQ86W0WslfdQP5FG1LkUuK45pO+BcUpV4MdTEcCK3Hd4n4bcXcEDubEu3m/I5abBeReg
msUHlnSqyAXu40nN4OmAhQwu/xPXaAZ+jtvxnmCkJQ5rX0lr963kLq/eBlt0kKc1kg1U6BBLKnrp
qbSYJpEjqZOyKmaYoJlcNDyg2r0BJf6xO3MHqhtx31PriFFZr7RHaNCmWABuCHmTBGEPALWDuyQO
G4+NySOdo8uWFMnBaFcuzPNDbyaOilfA7CQFWzaIP0w0YXZOWpsOu6cNiSM1q1/wxyYlqG5oWj3v
C541cFJBv0SCsN7vTi/DJv7UCxijjOXjxZu/SDqHSUOWqD610qLnl61Qvuo+WDij9YXY4/8muT+O
jXyzwNoOWNIafpO+dFD4ATaBkWIiy61nqfoskOt+PwR3Y+8kuN7xbUhG9+fI4lgXBXf5U3MM1C4p
+iZWymEn3aimAs5w5FGp8+lO19uEfyd1DmyCT7WjF2TTj0/zDt1usIUUOVBZmKd/hU9WDoHi7Q4d
3RAOZ4fifam/+Q2L2EBqLnntZYJuJP+pGIXDpjquJA6TZeRWnRcQ2+TRaOf+HrQ038/wQV/P3Gx/
9atIq0VDVWpuThHlq4SHxSAI8jR/oTvEX+HkAiT+3MEcZonxEQxgdlTyOplM8TS6BaNeHD7zLmVk
v9rQrRtY60c5uE2b6JnoG48uvxZRjZGwivFDjUTn2MTfQOeEJAq6rwoqHkpNJpEk0UgMXuPQTdgv
PX+QXAoL8soBhBtIYQ51Ialgd59denNb9OTafE5HPkPzJZualwJZtfXksCpWnvqPBxhVrHRfo8TU
p8cN1Q4x5ZV63ZnlrRYfgx5fYbtTmmhgfhuwGtm2ES5/SvxdMFcPIDgNikfFwYYOP3QAl9IIC9iL
2TMGM4BL6Pfssoq9lRYiZru4N2BSjjC6bGic6c7AbzNgqY+tABte3kCpVcCRdFOD4dZ/6s4dymvG
Kox5kGZGqWtSgGb4Qh+RGnWFF69iOZRIX2PJ1KvYBi3KL5GUTGSOxtr7PX7kfbtnMMCoXp8VqLY9
i5PtZwu4R0GtdKtwqaZ+M4v5LQV2i/7iHZh63dj91wJ9p2WoiXMqSEvTbwbDknspadtiulHLEBsI
i70Xa3f2RKmyAYFG8VSWi0EXrV5QCWShlrvUBtMYQIqApH0sFnDfyhyaUKFHhj1tehgx2THEqibb
9TW92ZBXueuMOOe3PHeCR27WpwmpxyqUi+4WKZaLysOyGa3N/UV/OpLRM3eAjQpDldpmY4NSdQSz
CluCHeOAh1w+ap3Jt+gRhTl77ixSu+t8R2Q6lCKRZvXHiTLDeBMLcJFT1ErH4loK8dwQbQ/xe1Es
3MX97d7nqeuic9js+wUp4TVP6/4TyWD8zDlOLwfDjML2eRgSjaB6DZz9y0dojLZyjWc1oGosRkwN
E66+Ekc2fUD9YKUGtUBvCHKwsqIkk7uq5Kbcz9wPgU7Dkzv5G+JWiNgJpWyp7vrCJgHHgggTbibg
/O9NToEqrcx1mbNTsptsgxemR8RxFtY7GKuHBCubL4YORr2f3MTsB7NGeGDL6N7qNYAdz36F8WC2
zFj+FthOKP+dj6ag1QxjNAA2m6YFfZBzi00R9ez2dJf5P7+6v2X3ytq99gOjCFK7rr/FL5BscDjD
udyEHP0tSO8Gi2atnbPkFR1HCs4WIUT2+CKCjFgaCT32UY5E9crN65Z/nq6MZLUDmNCLCTghVCWR
VUEYO3JkAhFyEmpseYtdPIfCjWFnHrlMLAIbicC73XUAHquVVqUtm4Cncr6dOpHA/ljWQjjeWmwC
WOzhAumC5CAMTwRbLR06StI+yP+go2Rk3kn76pQ78c1zU0/6hyLHcRM3SAdeg6dc4NwmfmRzEToR
bgh4DdNnAUjXipwMCsNRZgQr7ZwvFAPDG7Tev4h8RKPfytXLd7cXpXlV0kFZOC0TeTGZlTS3I6td
g3EbCISFGVvqp84yqByA9tXeqerw/PMd+6fGhUQ/8ewtbG0zgYcGT1NZwMKjDFLqjj0NLewjpmo0
17mPPXtWT+z6vaLgFEGEcd/CVnqE5tS1GBqVNqkfDAr5NaDZLO2MbjdGTkI/x3piVn3FqkgNzsJz
fFCrO1TpYiWs0SZYY289Ln9nqfOhXxKqLr9gjiIUqz005P8D99zo5b/9d4tnJnHp1Qjb4FU1Zhxm
/XnbjNAQ7LCWDhVB7YAFmAbAFmcDEWPz3gqTC8cvckN8EqB5MRXz6qjA9HzqQGzDt/hHu0Ykpvr1
nwkd8H6pRMan8RohfnbqqdeHjDcLBOH41SqbZaJA6gnoHtNtNoMnpEVjBRiIVEGwPQ1W0DXJGCZx
ECqngWc5ktYSl6kHGEuxiGqbaQumySlZL470WPc7rKJEk5oSpv3lqKfn25qxWJf4wGFf53bkWWpt
aorWqOJmJVQCndy+CfVeTZIz/IsSWsr/XrorfYBIzR3OCCM0qb5VZc9FTcWoWMTtlDGBxuLUQCuO
56MsLxYBCipqKfa1n8mOD+ZjNrA0ff911bVRkEVbWGOSPkMLoVFhvFPyEegHfQ+Q3SewzT5LlBOJ
PViGig5FeZBq3wwOnhKQ9rXw6npxifsfzAl3EtKWLn7zh7qvr5hDvRxvC2qi6AdfjBtsCqfgFkkf
CVShm4LevHHux8p93DRsNbtGeAxr+ktSdW1vdsMScJ5BQGO0C3W5kYbWVRDa09wRSU3G4klE9EFR
8jNvOxJP/VcrYsJq5aVW4Lrh72vvrZwjIrkrepSjNmcKRQA3tYytbxY7U6vZBIKBIz4tYPz+ncG8
40RJf0X4xiePdea+2PlItQvclPLYB52VnIRRBppNxgxrkgzo04nbhhYLDnCsPCRV2e3EeRqHB842
dXWYI9RBSuQRfqeF6zxpvE9z8UiRayOURdTx/iNgr49vE7dzsaOjGn5EijWbkGj4saU4n++7AgQT
sCKjH5br2rPMBPpTR3sqghhjpl92oInxAcpNfVZYrfBBzpqhmhg5VOP7rrfIZ1AhiiU3HaZvcfm9
OwctyrziX9qxLfLzi1tiBLrHXwk7AuutxWhPTsbSKPq6Iu8VEEsEBoqKhq9+s/veTwk+dPU1sePw
W9I59OHWX7U/Xg1RDsaGRWGnjB/zj//KmKsmmaCidvtpzLbUYRsPDaBlFpoR8W6B+Cby3o/9wJSB
XPtKAs6dOxEVTAn1KnR1ZD3GVckCvv7AG8ktr98peu0UhxjJSfE4rzsbN//eCKXhsPbKdWAqhLsL
0zO3Y2Qihutx5BtItv1O7usZU07LIsFzeoL87Sg76PtqirnB5f4QnDyLZiwdblf5g43Ogmcfc02+
kzSKY+62+u4A8KecRjv/aIw6WQK43u9Po3I9KEuVHx2TMRCSLcazdflAOPU6fZij4QoVoyppbetC
F/GCwk9sEp3qpTQwn047LYUZ+q3WLzhUxlPOn50YRXdCTSNublpNpky4mct/LabCzNmsDIXSSnmp
UvoIUrj89wpHYcuALNVL76o6L9lex//9vQeAWu9I3KV+X+YP+pwDMTW5eO7oenCp5AyYG3GZslkp
3NEZ7JdSLUhhJtWm+m/mGhS7f4TeJ1EwnANdRIsUt1XsofGi0HOGUOm1K5onY8AsolwMnqtkzGem
U/5PGsqbdCoLZ+Ks8UBIltAnoj3cWkFSTIY3fx3hg51tbukhwprRGjD04SxAXFdFp0fIz/Tcl21N
wB7xvGdN3eTZajWpiC9ppECOsk10Vhaxr3r+6k7IUbk9Thvlcwv+mRgUND2VYPCANhHZHooGgJs/
RGjBEDpAgQkJuTm/xbLHxeh07zVD4yN9lmxtytqupGz3bsU3s4Ti865e3mnlYxn9cGx/+6KKbkTA
vMYOO0WJ5HZyLdetjRvLEwyyCs4n/nCUp1XB5KVIaxAEwbcFtHiVr6TQ4EywOLBAIMiCCjl6/eKT
l/3mXbomnKamv/6f4vLGRkxfto/d3WGTYqMpjxV/4YUqj7lPpEyaVQBB8IawOLtptkWg/ksSe8og
d0FFwPb3wKcSR1foTxJE/obebPAskZ+lF30QVPUthf6qwCCygB2Z9Pi8IAe/eLeSMnyMOF3TTz9z
KyfumhB0FFF7sDU4L5hj/6aHlHA3+YM2LgwHLooASNCW91PV5gg5YWxkhxsVkDxJoz4DHv+js93X
pcSDaT3uYJM8FT667703VGc0rEazmt5cvB+vNYw1Gv5GSdz+RC8H/Ld1DsTL/bn0Yxe46lpdmIJs
8boozLULz6Mavi7L1+uF2e2pIkc0C95KwLltQ3eAnRsLx4WNQOTdwV7+00L9ezAaAWWXyngkiRjD
YPFb7Ih/cec+IaktzfcJyj7guigrN7gKq/SNPtjnu/uxMAVjIyq2To/0Sz7LFmlQgc+q10OIw9TV
6gQ991m9Fows0gMQvgK/9GDVq5+xy47ab0C4wNQDu/QvEfevK/iJR0Ng70Dbb6sGAU1KNR462Rt9
H0rW5IvzrAVFHd+CeG92vzuVPqinD2SjWlPJXbp4Uu6wu8h0O+0HeFpvtHEb+QE9TiwELsbSsqWi
BbcQluVhxbVtxG7KVBE5aKsWp9C7mwRk7AOhEnmshZ/3dpuYXNyqzcb2pXdQlTNPDtTpwBhFHeRL
vnoIfdXzZHh3K6ISW2wPKkjKBMF0UltS1a0PvtUO3YkIPMJgowdn2jOqURYgv1n8CSBBkK89Zb2T
/ydlKI8YF4wdiEu3OrPrJNWXd5zojoLni7mxjLk7EV3n6VjpgrfQ7daCUwhnDu9QUv3Ty3eCo09u
BJvrjgVmTlecOebwCFtq//kVLC9HhbWA4CqSv8xZz1lRQdSn9v0t4xPIriFMM+Hze4Rctb/gKAYV
WmHBvBCswl+tr2GmfIfnnKUQz1jnm94rlG1A/OxdTrIm8DHCitelqAoRcZkWVKMUb4fEROeOVZCC
wwMmU6rybCnr7e2Xrmjbi3Fkbm9IVy4RsOjmgB8fQ/xRUJzwRv/bhuC4wPRoOsAlSzcAaVcJTGOF
nmHR9kCyPFKMgn+rT4LAt/o2s4CuP8XcT5RMkt3kYT1cepjexZ02OXmqzFXVphwi7QRwjxNAZcRp
MIMqB4PE/MWgPrNnOwZXUJRFFXZiI+Y+iHrVeJT17QjgUnP5dOxwxqVSbDKIl9zwNOJJPPAaWyrc
+9wMteILnKXppQP/f7oyb9ctLlu0LiTZheO728T1VE+gN8cCd9kftZNJfZ4jug0VvhuEG3oN2D8/
MyRFTsDBQxNXQKBDrstpnlu7a2vXyj7+baELdRBCdQk8w2ZDXdHq4+XPnBj968YV0Idw9JXuMDBu
VMt9b9bH/+l3tia5uaEv8XiTLiBaKQQggaOV67EkL6qr58hfgCpNLGRNjBZuGWKQMqu4e3p40YE2
EqrwB6/kQCCebKNvTeDzCb/Yj7eZAzCth/nqBUeo0Ap4LKeHvqasxDZcaoUSQsPh0E+USEj7y0cC
XaHAdE62r3M8iion7rGDZbb896bDvizUrxVTLYg8nDJZxsImkB/t5Z+AGaHSI/qw7gWGWmfuLQT6
VNiOt3hLglapyYzuGiQKV107ckLs4IyWY9fCMIfixBptMF+FEm3P8vNQR2MuOb70HK5FhULUycwa
PWQv8RyT/p8xpa6/Ie71G6M08DbV8FxteKcUDQgx7jeFpBB9yZ0OOG+ZbRwCALqO0w2G+TebddVz
S3SwPIF7re/JMjIeuw0lWwlAxDhmbylYQnULWdVxYAiN+H/gXIe16VhVv0gn1FHS/UvzBmD8xNQG
yZwTS0KYtHsx796LlPQClizJr5k6JvvDm7EMqkWNi5ehOzZtd/mLIr4qbsChil9w93AtMjBVGbRe
gdgQMokDPxhEj73+IDVfHyx44I8H5mRgn1FLmzscKhh6BeamsEWk8fQv/gHPbCouyOKx5HwgBq3V
TS34AKxfl/d+fSdkJTHnJsIgl736OoComXpzVlCbVrM6s3fqvMt3wBm7eynPPnA5peaeFXX1lxbA
fdQO6pCLPMWweupaIkBVEzveCQwgJFkxbv92nOqJYyqAU3fmKt5CzO2XLzamn6dd5MdlIGc1R/dE
RY/5kLcuJX98y8LnB2yiZ+RT9MCEa1/937dRruFtQ5CE+INUMm4zXGpqLIpi4O8XQsF2MfdLK+6v
mI8oTnRKeaIG+34f1if86KSPG2Z8NAQ9gNELHg5MskjYIDPX+JOKw2VmDtTmdKarvCr7BXaKY1IK
6i3W4Y3+V0C3lGC6xUYT7kEHVoezoeAXpQCwTrx/qyWm50Y8lMZTHtBk7+tuGO/M4epH/XhcPBUv
uFkJdo87AuJVB5e/ZXO1/3w3+G6DXSyU6BxzlRYcMY1UjTSYvPYa9DcDCglCDPYxMe+MbMKX5MZA
TF5E4kHmuod3j6gzPvEn/PiTwok5BO72v35WoCbjE8fQLhep1M0Q/6/ZOsOKsAsQ01JZoDpZ9PEw
PeEFvjuUm7jHr3YV+BabgCjns+l2seDptYWl/qBVgpo8PGKDMyslKEjhqdrbadHTTub+fuPl6i2U
8UlWkUwZFXvwpCHuKU3RaeXl7yFhmesfI548liFDDDW7DQzLeWhSD3E5iFtF6dnG6nx7pV6jEY5M
42C1/9ngIT/1y/mOZaMCbKzGwvXFd33Y4eW+xZhHWbcIvvq94+IL1/WgVn4dd0G7w0bdXwQ3KGMX
/M3K8Zp4TMliZDYIdSOI8/BSQswZaVY4c4hGI+6hyPIaQS4aOhbBVi8knwey5KlKWiCNfYj2KQrP
N3SqJLBv++lZWaz5HeWtdLK/eTGtctrexWrwdt4UpM1/DRRBkI938CKCHF5itBqxAzY1HZkxkaaa
7Kq6ssbeQ5efzRPiBSVtyJADPhxOY5D6Qqv/hMf9BWoHHPZd25e7CMDcUsvO9yJVt/EofWP89jTA
7gudNJbF/52PPk51ylyUHZY6SDIxSBEf8S79CkwGMJD8MNBKRGbuB74Id5HrHN908xy3YcWtfZix
RGNOr2JnghkuXKBtOqRYCZnMeolM7zjaA4D2PSAw/C/bEKkBa0o9rhHZDAQYYl3kKk1LwpzEAx98
pgjl+eIrz0ji7JrcSPsQ2goAfQw/ILkkRnwpKFo/+q5Hx3sSTHbDXfbMp7xtRyKVXh5+drDvA2mb
egntoPWW5xyffsG0IVP6ibqg22IRw7CZ97MT8GfSByGiFjJUddD4QpS78n/iAQPhJGIPoYuEZyBA
ur7Dj44Ju2K0fMf446EH/Vcuu94WJuDG2KsxRdjtulwoCMC9Ms+I4XaerrKSgYxcWwFv41+PNxU+
83DjryHxRpHsZibX5giL1RPw4BFEFnNLg0F8Sp6fFuzhJVY7MgrugjS38hatVkUl5I/YlbWvGkVQ
FMLtA6VCoC4U0nB8VEWSOs2YcIpmikkd7d00LpU4qunwpTh35vWse72Ucb9o86y2EPd0inU7sdQX
9ZWCBARDQ2dEKLOZ0tzjh54JR+WUv3WIGIp8lFMQDzXX3SdzN30fyucxYEZNxiUulRNI++zoK/8F
CI/weHFEV+Y4WgPakeXNfS0TBdxKi1vwYfulBKwCS72If/MI82MeRxp9C9S0DYhPsz1CcDgVAxJJ
/IW5RjFwimdCVOcPq/BrFOVPOUgUN6o8YKdtCBU9HY2/3AmFswFRyU9I5OB0RFDzpcITiGCTYwz4
BplmaPM+X/83NpEUAT3yYKxhktLN1GzkM3zBLLf4fODJ0M30lBGuR565kZwNAZqT9kT58c3F9v/y
gu94Q2cKavdXEzcv24fx8w1IHgsSChFRlneC9qE4yErE48/M0Jy8At2o5RVkc07d18Re+AVJB8Aq
QS5pPQVKlhMJgOLep/LYDh8LLnV3djIQ3T1/1IrnpWifFD9Lr8wZ8H6qkRGANTS1hWfawLrN1vV9
3aMGghkEi51qQKE7VSjRq5DaHff2taOBkZtD/GRbA+DlNwz/wUUc4xKeBUo9Rx+oSO3+20wKF1Ll
W0Ocu+qhtKabKXD4haW/MkvThjG7w9XPpvmAUTSmFAKL4/H9z2pTigp4Yjw1pcyaG1BuiDzc2+Z7
rvUa7HSZjQwR448Woy4BNIB7sLKKc4eXQgpXy6uUOLze2dOwOfQIFg8DMlrtTK7qTEWr9r8k5UtR
YfYbhGlSZ61xUmcz4+7KXBnKRMdtHuxuW/pZAfkjMq6ULAFxHiZQwdNh3yUV8MhwMDgiXQ6IrY4m
hKjUJU6luJguyFnrrucW3tdbK268cn618AJC+YmBfSwfOsP5+Lf8El/f7oPwLlpvIkORN52NWhIv
qzIxFYgIbPn1NIaFfYlVBq+rilHr5GBZYo3peJUTg61QE+P7jDnudA+5UxZcJRxHmGaCmkgsk3I8
TXh971VOV7T/7WIvRBnxIzcn1S55ydatvnBsrK0oGIUxlOON3wIFRIepb2k6f5FiAoXHditVkNR7
oc8DG/aRWX09OfZbvwVv18cIsxaDRqaS/0W3sAs5LhrYe9ZOw3d4lLnLrTQ6dHJzB4KbpC7rK/Lz
LKfQzXzUNwync9OJy4dMnb02aEXqpc8u95LB8XzSnuZB7lSzzq8j1AOMh6AAgxV1hsYTXbFmWasB
EsfP90iRJEbbgzSHomJlmhDdz8AREWZAAzZvgz56w66RBe6vJPhvb6wBbhelezzloBwUvFbGkFNn
yIYcEPApgCVYIdUjGnpU9NAm1QM0pwaZREpTic5LQjBV8g7M1UA+CMmR84482ligBrqCw195uaUp
WJhXmzUmcmGHlfGenc7haiej5wV3N6u3IDePH8k8U56yoQtxB8QkrcV1s1842VY8nKCEFexVoTMw
0Uy/8PSX/VQERq6n1kCHx/4k5iVFpMOwoO6BpcsqN/5PwUpgRiIPE+BYRKV1P3jmRz65H+RFJqEc
ahrDrNuVVjc8W4Ls6tgZrh8VMBfJqsOo6DYnmPuwRLW053wf3Ic0hpB5+B5QXa51lTdSHb6HGgNH
eV1h19KTmsyNJvdT0n0pHP/DnfJSriTmueW4pE6GxZX1PTOiAb8cNvt3wn0l6IUzgYnmaGv/Mxl/
DpVHk3zffO02AplnsUi401GMHvWnG1YakBG1xHUw3nPlplXZDyPyJNjBHN/CRQ3Bvf2FRUwoJ28H
83MYLPhyRSe2Z/YL2sHD/qLqUorvvkfaMZnBfxwj/qyjJoyKxbamkg5oQnwU7HhYOHIzNc/B7BVd
SOHULbhTuhQ0F2WZfe/QHGOr+He2Uv7KPR9T8oGKpxGJEtleAcfhuvaIaDuAJg/iJcXr1adhLEhg
I5OLiigUgUzVzG5pScH/AQ+IEV57M5kEBSpkwcY83nhtRjSbAGi+AlEWsPW1Vea12uVHh4rc5PMb
Rb2Y2T80czHz1mwoXXeomyag6NYU9sBCtP2bir53LyPNOz+5FK73HTfr5J6cPZdCTJ191p/xbxvq
ejDPsDBEb+5ApYy+H0c0qvM4WNEjxGrfeec9DoXV8l2BuPk6or28bcB6/NmtAIn5TQVg0cAeOXb0
X+o0hgmHbG4RvG/HqqdUzJTSM0vyNBgWh7MHiFqTvvL3RQz9GPP7lISe8Btnh/1BePJ/4cYcxmOF
qqC1VVhE9io6bwQyQNIXDZco8ayP0EjwNf/JnqumyJS0MNIl8lJ8HaUB8soBikrTRpOw4cGcQvTa
2ju1WWc/uhec8z+QNKlnkU2UdBYymO02HJ9/FFbEUgy0hQlBX4yjFVFdS2Sy8E0mbbw9UDdJIGux
TBDxiJ7HGVyJDzFYShsk4J/Y3gDkOekv3oLX9isKeRSpX7z7IV1u2+ocoMFnpVGPNB1FfPbWxelx
tRSGhYOMStOu4OI8XRSbB8OMEHtiwQtWrP0MdofbUdbzeAvhRrrhRjQ8h6M+GmX5Lr9a4+B7Ry3N
mbiG32+v8kKDN1MdPmW9dreyzV6u6X+4cFqQJ0r022GX2vHyFanAOIICiRmrbz7ikq7G5MvSKuMv
k5//whWyzTL2fD6wXsM+zB2lJD6gz4T6edkGbbofVDKIddYeiq3WXEHC4DtuzEKfLuOzzpREyihX
aTiUm4hTFcSc4JNXAZ/AyKzOq6w39H9ri46s+/o2B9Rp0+9d7CWXettK1OM44HNrUAU1sJTp6Klb
0yfsJMt0uGSSw0YHnh7uKbuRassN1g7ctSaBsupz67A85YZBwpjULxGmFcbtvQf9SrDvq1kr/1t9
AcEZbDdPDV+fwzGb5l+eS/9YOvqB5gBqR47kPMeHLXGOUQcFQfI4sBAQlh5yV4ZG7+6RFB2S9XkS
btYQNs/YhbaSLaxn7hmjMezA/r7igZJrPrH/X9fVWnUZ0B6BE2pDgiGPXaAHbzRLZy2T0olbCen0
vEFWt5/TFwZkSgUs/x0Cog/qEz/GXpbhG6hlYvQgmpfvaSdIFUxCCZrfb2jGe7GXqrkIK9OLmME+
Bcl4wHpfOapY29MdGXrHETu37SfsPqDCiyXjHTu5jaff7G/AhoGwpZBpyhUO27OkbX+z1a7QLVVQ
jhf4rPqWoTgDcIbMpKLPKueJiCvAGTpH8hvPwvQDOwnhK4rxjHpbdCgSuzS/5+e28zTCc6esr/CH
xKgNGoCY4POK061JAjVkWrbGqK8gkXKLPnCpjw1FKh50creJEbOBNpbYkkrkTCuM0C4CItVvTbcD
Hpx6aGcB3vmx3V19SET1Jz3xS8wHTuUx56CCeiZP9Nz9ETZcfKN/aP/UYG7UXr8qrGqReuwqk9r1
w2dSS1U5M/xb0ci3SjR1qXdfs/KF5PbMkCX4Gqqg/u33kk+XIGzJ7XADy/z1o7zhtY31PoSGY84E
vmREb4r94WKxXA4oJvewe5X1SA1ubvbJcZA1T3S8N/u9unsBGN579fN+dtlr5M+CgWajGjyUVK4E
lvcGtEOFG4SfiRXxe0Z996gFblR+45Y6l8Mz0kt3DfZXtpwMqN8MaLG8+Z/HNl5uSDiLyrTI3Xqv
ETVqJjWlNBpTOI1+tAgsa4C/3v2FZZ032ElHtm6OQq77r8IJMo3Tm9YdaRBHueO6/XuCK6uVCgnI
U2d7Ipi66V8KJZZKAUpX/LqODqa5bhLJIlSNjY0K1rBy50riPPTCngPEkapGCvqVQjqr3LKKdVvm
FT2qZaCZqvA9yTYmoDVKtL89Yw+U+kn6kTC6AZi2UjdcdmfBtBSfvtZQCaiio/MaWvalVCU/N1Mt
PTabB8WBZnYQnDG+u+bVcyrI7g86C4NGEsf81bXsfVfgn4yO0qzenKRPOrJg12IV3TYgcndXW8XS
X4kSrft+OXBOWNmLBgIp4EfBzQP29GpihMBqYcXhNKhkm66rda9vsT79zDH4BfgmFUks64DYqekq
y+fD5wGi1ntnVNKCKgqo3hWl2vo+ge4WaG5s8+WqNa0UNKSbzcRd2v95kQ481I1DBLdhSn6Krinj
4Up0hJqfUEuQWzSeenwkMPGYsBRksP8pTF64n41pmF0sf0O46bJJFLd6D2ccDzs4iSo8YCax/O5o
ET0y2ksWnxkYmYlf9mLyaDMeRYia83J0LWnl0xnbvG7OoAh2hXg43PsE+6lwwGVfB0F4QYqXSVob
F9u2Cc1yeWAOSEfN5HQGgYUTNJeW6yTWw8+u/oRvjoo3l7UoPnNy3YFxRVfrYw74N6ugeJU2I/vH
azIG7QfnKM+OnF80U91vEZRrqZZTWN+InquSiS9Y8migtCaALRMEspSelg3b0AkE5ZundS7u57wG
Wx9gWMNYKgU0U+3xmh7rHFuLTg22LqU5WWCNhS3miCQSpACCZ1r/1Gm7O9YIENEmnrhw0qcMEu5Y
dQcVCyuuIr7XQtvAZi0Y+BqMcSAVdQBHFfIvDlBaUjnTuSZ8agwP/rGOwrDVpvONist6CKEP4cF/
8RTt7A9HxXw61mgKm0YubXzwKYUk1HI53tfwdnCR9tPK8AYMNKa4zgPStxv0xWaObTMVUW1y6bEF
pGoyA+Iy+qRq5HMfpUKR1tMf8ZbdmVYrHgvEXB9/dL4WPBsBoAQNKxfWplQXwf2PYD0GearDl4GC
SEZI1FSry/nYpv2ZBHQokdLovsWjZICD0PlJg7OUQMAlfBU0p9SikIZSQzxJNhRjRL2fUxdU5ADm
f5fay2RTWgJgX38mYvWeqh0AxV0KR0icgMKGqE9VYlRySv7vOqHKU0xnKtdoJRmfTVbkwnpLc6NF
/3bHBuIdlexETcIo8BgNGyKE88oktoHNs3AoCSNFqCQdIABNUs9pIPnt4aNuI2rJ9qj+xRxir1gp
cLtX0HUZ2xeyfpybGl7c+X2e9wTPFFe6MPX5gqG0pkZUVToolEXashvEUGGv+KZ5cpaZBB8eKZiW
QoNZEQrXlVkEyxoso/ZnwMwG2C5whQGfpeonbD6eMJtuYrguaase/crKapd9CMvnbzuUMSxurkSV
Qttv12g/v7IGs7nmKWh4JhjEwoKKUWlliPrSjUoZI+Qcn1Qmy6SJIT5rGDjNUlw8GBaZTYKw76NL
O4aabQLBMz9zbODFyiendUs8u+Z26bKkqkFRi57O18PFiiOdSIKcsH5vu+7qBYxSl6DJl5OLqNtd
0+0s658VyhEdI3Ad+U7i/4uhS7lwMxfUuhDzQUrsHVXzqy5tdf8Jv7UXKZ6UhpMGzrL+U983r5CZ
niohtNtQu/3/wwYjMJ6jd2ojMBUiS6uC/u/TWN6Ro6lb5crC2EJy0XZbnDF5nFV3DLgMfzYR06JJ
89qx3VL9yFmT3D7yAreLDEhrJThAHhG2nQF3Agbz/FLCGHj0AI9TzoPaZanlHVg7ewpZBZfO8SQh
HQZ6fbMDtPVTpLF+KBKsv5QxpkV2XMpsZSuThRLUUDnsKUCDigCdR+jS1QKQMZxfZdG4Q6jTpTey
3b1XbQQCPic4B0Ttf9pt8MLdp1EP/eXr51rWELY8RHoa3DFevG8/SFaciBhNiyYI+7GzOdkRWdsR
zEiOF7Nf+ckU6tS8FGvDx3KYd9hnfQo89eF/JXYeyytjcJ+8JqP5naNS/avnkbNK5ADCTifkJerM
Rp46Ydcd6V++IKWYG2Atd8aBRwj2oFybnKU9B5+wp5WpvOjSAatDp64RoVrTVX5w33LaGAAMzAMP
6lFy3P2rHPACfiI2BjJX007WkiXns8g0WX1ymjsrWoz6Whsr7i5Fb7I68kpFaWhkUeP9gKWePmxb
cK3EJGtZhzPb2YPsr9Yf3BSNkgay7JZN0McQQ6MjL1Quvcx3YgZkGC6uj/oCxMRDxa/kBE75BD72
/pgCBdM1iszozKC6kfBlVQpolrukPzqnw9tMpsXSIpSyXBZlGLVyMiErbjLK3NFAo91i+81MyNBY
5jczw8fsus0ni9JMWqLjoAbfd+do5lRthJ1ogS0J3DAr+qfv5kUVoQe131O5gMNl8meWj1qP6owN
TrKYmBwGuOzInPdhH3jzv3TckrmSVRD100nv6HkGI5WDHIB1LJAupbhsr68N9Lhhg/R/ow1uSENR
DZwOUHD6GW8HUnrpaWiHL2A7A7+toHRkrHQNIWJeKPLWZMWrWTlHHKkkBA7Oky9v5JCo4qJZiOkT
7g+nu/LQM8zyS31iW8zKBl4j+tG1TLVkwU0yF+sagCFMzsgncnxW4CkAhJO9LD4CIko9KjN+NbKX
xiPkFiQsbgaCkGRAjL6UvZtWmuSCDrpPUpXwzJ1RgQKsOWJSxdcbP22qaekbgruWWN4jKUv9LhsC
01jqWigfbAn3x4Hn/ucAcx/InfCyf24s2poafC3bpzpkuqZJSV9EfczdKIMEHoF3ER1OqACHr8v0
1N7OIytfuMH+jbgHUw/XOCRuofldf5Aa/b5hZ3BPLHn1RwD0ts49vC27dejyK70ofiLJZXLozs9y
G+/2L9TR2CbepHEQE3iwWDipzL3ht5P9qQcBDS3CHxYwKeo1euEwup68eCKd5/5AOxMcCHV3WqzI
f5IT860PeDQFWL2qOt7IC1akaPQ34naXwJP09KydoJ/KIXsMmJDbeqiYZaqIU06WwTbS0y/Ioes3
5ZXpLPRTS5JqDayfkZST9CjL0/QJHRdKXPnleeSW8Bb5MTVebz/G+9XpxI0LRYC8DCsiqfwwvnpX
Oeg46KTeBmvyOMB3lK+K11ycKbLtAHdZ88iuVN3WL3RRcThljylu5i/cvl2bpAfsGcvuNlegfd/B
2YThPsv1X6POoFXPIVIvI6ZW8qCcqhpHg/aSTnkZTlSKLbRUZzzq7axXY+Qks16DR2aXOTlTvznQ
OcVqCfc4+9hPUAi1MIMilyx6RpFnOzGORDH1Hxk3Nbyu0F0hdSx+KNEwAAEKdYzgo+8jFHnovpdR
BDvh2pipYB6xeqdBDtvbbMXjhlEYOzNWWGarZ0XrYyHKxxbBhBg9VbyhfvwKcaV5/PsybG9Iu66E
jwh3UDP5xOgKbTKrH4KJWKnrpxbdASt4cWtMr/SYg6omfbVrMdpY9ThRDkrGuCNgHCQ3hU69gDum
U7S/dTVWhWhvm0Xsv3828iUZv45uIc7kyt5ahcnetMgOcsYMQYCgYA053wDcTPHkiCYQXNRSkS1N
92G9K8YPqlVcJwNyCIyzHunIHYM1bPN32OCd1ZvL19a8dKOX5L+4Pl08h/k9IVxMXN7Q3hrBYDh5
WgyH7WFZZGLHTXX6Hmccp7fHuSdb8EjdpgQBhUafnvFHsJPfSxhDfuI5aaYRiqvqEKYsiyBGk+ei
+wiVfE01KiHO+uXmbcCQCqiC1e+t9RbcZcODmqfTPlku340rCR8PDgUfBaEKf7d1ckhYGF4ajpGU
yCoXnYM27g3Y85rd24SfyKP98V/03OQrQ8oHXvT9jE++x7dLqIbPh84BvFUNkwhynBqTfFR+TVBb
T96W3irnE9XXmVTmL4LxqTQLO/lAm34gouo6Xqj34HAZRPisLseWlCQG4+u1yT0tYbeDQ7O/1xAY
c9vHT0a3dkzplBuJ1cWB0lVSk9aUYEC4K2oz2VdDxYFqBZXsXluaRRmyV/ErgPj1t3ZnddlSkyqV
natR95gUujF3/V6OuKBkNnGdQ558mIlc/aD67wLeyc+KGuI5xPLg5KHeDNtPSZAt1P0Pr7iwxJvm
xaCFXFU6ybWlfdhVIeaY2YY3cW7DcCeohuOmuDmL0bYJNNG/6aYV4iyrJyf1XCZ0oPb99QwKxpm4
5Meorzldcg072fHdt4HxNqxkSgCt0L63K375zEj0HNPtH8b7fXnYNh7VSMpinS6zPXDkErbrTxDy
YXs3omieaIoLlKzPJLohHAff7wcrLSb6QZFlt2D1smJusePiFlczoTAEglKCn0w0xg1Tt7Ga/908
fVy8JYTqXYJav3QRxwJ8hLiR5yKtxymKc/3GTAY3bsUp4wBS4Jk550yqbTact2MWGfOL1eUJmfTW
9kaFabUF1iYETepNeowkNagzWrk/Wj/wGjx6QR+CQ3uVt9ATlUT25Eb8DM1Oq39HV/4DTlqfLsK7
mFdhICr1oFcT8otjMQT3EVHh03V210oJX8HbHS5G4CFaLkUPI3hft/gV4WhGRuAX13s2PvONaLGe
cPiXwkguHDLLkqw5vIiLD7hp1XuPQoYZTD8cj4EBig7+72wOa2VpPpN5B7I7tP9esgJHSLcQGXaT
5Tgl3xiRnPN3x68Ue+YY/l79us6U/3Xv4zg78gNEaR1UbycW1jdfAB9ic2EY2+e15T46XHNuyTXj
lUf3y2K1K/Bwdcp5i28X2HT/5FhOPykQIf8hSLCgt9GF5l2setgjvqu7qS/HQZtaTNHXGERu97aq
cMZ0a4VqtTpMm/Me2v7nzA0ZX+fm4WiKgAXdq0f0i+J0b9YoU/+amZc1oVyNBFJYwYo6t0/RBqyx
VCZCc3VUaUK0gwk2sSDr4XDw4GM3EvvzACy6EXpLQvIeF3jf5J517PhphrTYMg0Ob93x8QMnMk9n
wFlsHnTd9F0TJ8DDAbqsBGOydEG1sl1qib9XeQcJwzUzB3SI0VTRJmglYg04Sq0/cqNCfLhEWkQu
E+LNAc3tiOMDKoJACc09mdXqifwSEF0qYWf7+/mWf2SabmNodLQXlX0N/orZsJ8GOQrSsDJYjUMX
DUfjbpvLR06Dc2gf48PrpibG9z4BstJoaNAkgjXn9zvxbrJhz0nUG9eysmUy3KJ8r0rMRjUEELVQ
S1R/uk0/BG4NxSpRjc+hvVUihGTCBVGts4QdjN2FzLpK+lGPHF6i6BGvCzrjZO5+Gl1RIipeUQoF
YxOAddKcoTRSjNDRhayjC4p0kZswQv0PksqzbQforruRn5RcKBx2HTKuRy6qw/WwGddJpRix/M80
PmFkepplkcviY2Tw04FRzuXvqISpsCF8PgtE7sbSm1hK7Vi1/zxQEwiHACtlFvqz2QrsGOl88M2S
QLf2rtWfpaZUFkprDJGGF9dz5I56lcVdT7dQiGd7xJVWxVW+BTCPkfyzD2ZKxzlSkkluLFMQVLVZ
z6QiKVrTbVUFsFfuiyJek+w47Vap5ijqRRijuO8PyqyuWckXTwFdiiEa/5zw64yoiiXhOUXP6JQw
IoHHoYXHtnwUVJGUfIIu2BrwD7TSca/rM0VyhDAD5AsHqQgmFuSX6pEWSS38vcKe1d3tsOu6Utkx
NEXurgHKLTFbmMLiRX1U0QkxeX0TE5IzS2mv9gsezIRPt4u8AZXKbZbrtPmbCQF//gVsfC7q0/h/
rUqFIS1hIyrCg6mmiX7naYxG3rOntQc8EPsy342f8QjGdngtMCjnUDv41968zYNaA6H9g1/7zovG
+LSwGL7KB0xL+mtSzMZ0hl4uZ3/6xYKTibOMn8eDyl9i9v2Cimo0z5Oke8T74Q/SK4Fu0dTfIMZ8
xxfj3J7ZUQSZmdXfqEc1XXkcFZFG1NPQHfGPtpNyBPspWe8mM6sgL5sG6i28wC9AV2vbhFG3lJ3q
T6nVHHX57CrCWUXpjkvmgqM+mdHo8H3krNihR2NFt9aw8C6XDIkyda4aaTGgYlq00RJvcSS42mVK
XS/FCMVMKpv1uyLfn14w32shfUoykDNPTTonVMSq/7jWcAd0MubArL5YEnvyaOhaLNSQZ7enaqta
OuhYZ+8rEILPwACU/Em4m5X21G2On8APNW06FMqC6a3KxJDyndXmFgdW9DREzQDCdaFa1myBtAzR
olhX70uOgH7e0MHN70a/H4fBdWyJDRqkG3+Nf+BtkIkL9HwV+GgmbCeXwUoE0wWWOteHylZX4cgE
LSoZ3wqjLZTK9oK/ilfBU9x3jD+smk/VfhG4ZSvZ2MONbx2fJf4aYP1NdfBz2W3ulZI2JbN3C15X
YuMEL9AZAk2BBHF8wOb++3wioW3aODYcykT1MILV2Xwfr0z1fVEHd9g5fk+WpGZD/dA4P7fSuPKg
iid70/yAr/3HJcRHcvzqOaSw5bY5JNGzG50o7gdhabCKNv4DmYY/RHQTljFaeez2EEQXYUmMY1r1
o3TLEvw13CJAl4zU9RbPr+mSPc9PkZAYuXD4WFY9+ICA4E7iL0rFvfYCF6HkM9uv+f4Dh37Azu5r
ijl9biKiYFOFgyRJEeVpFfx23TqVhRpP0k1W320l7KSvKR5H80WH37V8SsO+CJh5CSJqTe6iHlkn
l1gSOHsJ5fulF5qSOhEFoaZihbVBP/9ARmSSGP02DSf3jbTmMSX+D666CpxHER6F/y+so2y7aQ55
IOkCcvHmPfaZ0ooE57ezkCCAz0bUnFHbLYTibtlqzgkkl+ZsRrGbB2idA/J/CDZRiLyrvKfa6SmO
2baHjKAE5YSAkKWKp/zPxWgB5rDQtzuIo7/hciqvAHedzYO0vnSaY7gf1Kcy4cygwOYHz9Va48Cy
AJrhhDLJl3OI8jZSUn6lu7osIOst6ABd7nVbMCZtutqxs43rQrSYoKA5tWMyMEV3sAEuB8aKaT9W
cG1T20wnSyyo3QHzhj0bmsrFHHaIR1sV9bXsPBLCg5KCR3c35pLbKbeKlLYAfcz+1SDHR48gs0wN
1KlFrlFfkDqK/2FAt/VxLKPQzGrxTUukuKm/E/ugtfvgBkd4xpWPv+0MvwU4oXYoZ9xFrXktqmUO
R30jCR/EWuyXFK4KOxBd00JFnt58QS0whMo8ld8UU5Tx7JW23uCLxEtReR/3qRjImUzX9yl1oi0q
hyEfknAfshQIORMZhqUdZRexQjOZyw3flBiuAWziP6OOiuuUBLbH9MfCWnxgF1Gd42FTwEnLmOyH
xJzhrcOSNDhSvgneVsfX0VNh+5/VBIiMt/uYf++MFOeWlWwzRsYaT/VqrG+kNjTPJnLYXyfr5Atp
bR24Y4kivI88Xu4Cds5Rtimqwg18AanJ62OcWxS7is11CzmS1pifj+b9SzHO2fQ6+wL60wGN4xFk
0MsdvBRDRPvKT9mWA5WKXHrGImZEPWIsrP+HxA6kyjOO4IuKWVD6yB2Taz8Er+vrJsRedb/OoY9S
kzLQ/uuEyOKYG8uRLtVaKAvWwrGng6ZFyC8/o2/U7a6kZzevf2PYm089fhW1+5n4mqaiv++MzbdC
J02W0dcT8Bw+h1FMnAomA614Z8kyh5JhPvojFyAsUyjjEwKsVHzRVBIgy6f+S9myfwrDc2apMoVr
DxVYkymhKHFE28JRbHpmyMw+n1KoyTgddtxledFIKQ/FNDmdxf+4aG/4bj58gMkRVJdFBg/taDdx
8c1BSNKNbXhlbZCmxjdP7+X2sLy9vx3PY4FplSBs+pdFG5WMS4lIlNf+sNPVswRCIGw1M9jG0arY
r9U/lA/1dJPhVxS+swgbMG6+vj/rq9RfuLpFzs8BGDLDqeNi8rk+RPz6SkYCtl2kWTM/fjHtu/Fx
B5TJLXHeCZxAIWjWdEeUGyQG1SLCDIkQ60XCWoEM1oaSvX4tRjZxLVU6zENKr4t0D4mKpE8rut/P
JQHA5KhdEI+nJUkAN5o0tqjLfpllil34h0Pyc2zYjD5r8i+xe5lVwHI+z4zfAWkYt1n7PLWQrdO2
XeGtKCa3YfEkdNNqhLuKn/R64EEZyZ1IR4m3xeuI3bpcweoxJdGEk6PodhDz4SRugn5wuoSCFGrr
aQin42pHMNAYr/noqM4zivccF7OAwpAmXxtzGHFwq5GGNUmtxqV6PqZHPHUStK4nDVbv6l8lLrY4
vx+rSAtFBvdG0M2xE4hbPSwyRdCGiwrHr7IaOdeuZ5fhxSL18URaYVMfd+8SSBWOCvl68fktRNHf
RmKeCHFrXJuQSe+muex0V43/O8RVaEy6ayXch1RbwjxqTzjPshZ68Um7LnKmOL0Dy3jNpZlGzicc
FoPpy97Kev3GDHi70wStK+RDGvJGHlguD4Vir8aJQVjUhQgplZ16nS4aYCVMWPYFSbSMpjAjSh9v
JKsD2uREWFUB7Bo2MJ9uFjswBnKyamCXW2Eh/a1DhuRL9DEeMmZz/Zqg9tl/gf3pD6EPe6jKgmyp
Bpv08WTTOQlc4dhnLiyymSffiJ3gh3AV2lt26tSwDDWbnxJVGlXO/6ssvqsobwhXKBLAbO8RYDcP
tXWCXj/tnWmQBaNEIBGNJ0HThaElJNoFOls/BPVFMcQPIPtVZm5Ef4IFZq9TJucOaEGdsN867TSF
Un5e3mZr76kLL/scUOyiedV04rgZzvoQBEOtkMN6u/cy0dYdHrKsdINsAU6LuKd45xTFBGnohA/I
riQP/CnylS1XyWx+YgMXWzvG8dFrpOwFEpH73iK6igocnSUyFfev/NuwAdeK/pJm4XmQl2YVcnYK
uUDzzlpS3tBFPFE9mboA1UApTNYeXGXRACi/0L3qWEQfR64suXq1V70fqomhJX/0fyjuQVXyyYr3
Kmee55JTFJ0siW+RM2w5CrqzHvxZddfOJRRxG9ExHV+Yjiv18f6MqTIf1M5dUow1M7dA4ABrpSt5
Qbu448XiJQanM3jPsAiy4EX5SE6oMWMtlKqs9ZIoB7WiVnNN7zeYaf2diy0B6auzVGiq8P2ajUkU
AmGVwZlrSdZS100mAh21DmWBgc8Eux6nCC7cFqwLSnY2IX33eRvjQDhbvtKAZFVF3DwB4O+smCQ+
GNWVfwK5esSn0yeE/HhZntneyjjr9Tw1dj0MsHiqB1z5n9bomA0RWuMDfBeVQ/dTbimCgud3NqJ+
hf6K+oNoi0DNr0Q5qTdoisKx30mbmr23FKu5fPUqPhngpXSNDZDjtPORaDx90AMjnk7d0s8hzpyr
OzT7259HkQDVzH8AKIw/S1oVe6h971EEGUMkLUfimpSMyXm1K9ZRiwtMinOzG2G1BL4fHch7iwrF
E1MTSCYQHnt2O1+m/7l7IKXM7hVx8nV4ok64gycayqTZTy7I+pHwCK4jbkhpTlEaPp2Y0gHhlaio
YGDfgvpVEZIE/h1qd/y1lgSbQIkOhXrUMB53/fxL7uZxfkqcANOjCeYF7Bhs8gupqPYT9x0Y6KuD
d4vnfXYQe5P1Jx1g9k7Wgv0g3HqL9wzEl22uj6gd0JFVppuoCsXBZCpYFPK94xOZVqYEBNtTDxID
PyZk2v8qg/8qDAfcSeZq1v2fTaBETloH87pE0Rz1/ortTx7zcmjgy/ZaYHOinjn8OIKy4H50wH6Q
8XfRHAEsTxBidAGLf78Qi7kzz4a2J+bOwtS4+HGr+XwJqJdsll646luq44mZ6tD05upj9i5WH5A3
1G3F7Kn0fWs21JWf8UP65mGVf4OF+zijEUeRYQcramK5azKb2KSxysCBqMC4BxsxcGqjMZ30jzvN
wbwb6C7INJOQ3h3k3MAXalCi6SxfuvNUQEjz1D5IBY3yT7PH0YmuZBt5+1QXBmdtfVErWwlSn/RP
T8McDxSVCtV3m8N2K8HGb49B4Vcgdk2ebfk127dde9Jk4CVliAIkLFliLKRmxPGFtQdsLfd+OuTh
qWtkGK4chWgaRKETCBUTiD0qLaL8xSpBM0TVn5A+hqqJeBgEH4R8Y0ssu56/TIi8FDCIo93prPBu
ixJruh96Z6DSgw5oe3bTxXBTDEaa2c4IjOY0BIlbjwiyELX5G/4HioTY3b/QJnPXIy2wOB63MT1i
QCFHkLGF0jLZbbgQS6Xlb65uBGItMBZ42DaIoi99CiGptQi0FEUMftPz+etGyV4tWKj6Xs8g6Oqw
u4GZ1gtDZpK9dpahBjOXexTNm0w9zI79NnepfHuy+pAlxipS8AO86d3WK2FB64pmYW7wZaomDIvT
CpFSIwMsLhAa+dEd1vrkoF1iXM7hDLu33LHUSINgHKkLnF97UCCBghxPEf7eRHxag6oGwdhjPAN2
btTGwFd1TB4+z+CGTFM2Spq1YKanyjlaixEW+axLfryYXestvDMuuXhsKxZQ+ng60O98xq9Vn3pl
CRT9QzPfjNuLzvdwVP/h9lQzlWTJZi6CNu+cOvGF+TRG2eoERxLIVvD24XTdWPFuJIxUncHs7Zjk
VHMDrP4hJBiY0WNtLDi/oak6fxPAru5i5U2C5biYpE5hhwJojYZnvlY3FDfkhXS+fwUB9g66u4vh
C4DWAyArqzzlt2Z3s5/FAEilqileJbFF8Z5OdNAzIwr7cb5FgA+LxhYQbb9MSuSnCW0N1VIFrJlW
DK1YM8Sb5nkQ9hgfYNeUbiFgxglcRZuVw6d42H+B+5iulx9HxhP2peC7bk6cDK5PQnAfZo3XS/ix
1WDA9bENBEKa1mSliE0dIsMfUfIRxqh+tEVBk64eXefZZy7olnKfUXTtGM5Y9uAIgkY0515zUSEI
gzFYLcvuCpAuDKLiIq0q1COpBkqQI1yhPxSRf54mYaqc1qB8nJza2IZbYlSGWh9gQcCsSp+mPlJh
0zKFhyG5fLNWSIAFCsDPtt5CT5Veqaqw+VzdwBmEJNyPucmkJSgfUI+QPHcZCrRR16l50vozQN4y
FWx6eHSeT96svzGKUOzI0jdEnKPPQPfJxxzJLjAXp5qxN3RGeDpN2JwEA+YxBTZxlXmYVhaHmI02
9lFNKK5lXzT58xgJg2JTmR95KQpy9EPHNyiKTDmfDVwVSiGPUAtbtxJvHYilbllmYXUuYeRvoqvS
q+p8HrMOEzptknM551S0hjXGrUvCM6gy9OIaUStoEDaabmBSu2Sbjfij4VCTzRtAK9nEvuhuXysR
eq3z+OAF+om6IeMiysbPZ/vM7yq9cyqEyfGezTSWU6a7jImXRvU7gZnY/VueVinZq+yBIssWNNe1
9AEXyOFwK103bQf/J7UJFKlKl4wzQ7eScEEeAtrFRwhC8oeB/3VFBaKKKEKh451rLQtISgLQZlfR
r9h+13J+pGK6OjBMWc9DIYGcPjcOzZLpw91CRXzSrkJJCiH/X/1NcEVlY0w6VZM1nvp6jZTYoDnQ
CZI8ZZ55eHdIfm6iWvr1zb50eZo95WVxvnmz0E03LIrHCidSpoUt7aFLFb+VXPgqARF59orP998q
bmbJrZDX5neN0vBi2XalHW9/4iEbd0pWosQXP1WFywAFHq/l79E/CHNgMyhVI91rEOtnKaM/h9Al
+HE/IuIUZt97jUYhKpSLmLXqOuMOygF21moq+6ioO7+RKcMWOa9JUTcLoXtYxWqyF5FURy32eZGN
DFMQm106Uk7dwtyvz+XRuidNTP1wyU69x3ZlwdUyqh1+XbH8H73PlilGp6/VhRCYv296f0LsQNcT
xY/GeiZfTChUBjYSg/36hUqftpRV8DKgySojsbPl5X8LAcp9/aDTW9t2H6bAc2kV2AK+TsJAxwVl
TFfXtYiOBFmNgjHVSjRYUCyzcqaUHKBxCXHgGypIYWczaJsi3HeT/myaH5JqkoLnLFYYeJ0qwjD4
/QZXx1ofVDbAzvcN1JBaem5+li9K88fnz70QSd4Rczu5ZiwKWl3Ev0VFmf2l5YB/uat0MRGQtYhn
edgRU+BESjFiJKbAAskaafIY0r4SwSkMvRHquW/q8c/t9oFdjaHDUZTdmcyeY88wDRx+Mqjk4o7x
bRVkHnwMZwtb+7m62NWZTbPMNGD+wUVLGq5zyUFYMb123UtKl5K1+3nJ8krmbQHb1K1hZRQAApRL
SsSOo7DTzNaAobbbnIcNK8nmoNQ/4T45KqARLHYDTMxJWkS/ZQB3wJaWRyKdL81BXwVYiPVMNxoo
VW2O19ekpx6sVTMrS96SwFWTPaXu6lP0N/JO1aeMsG8J+ykX3BQTrPzSwW83JE5BoML8OkhP2VG5
4m8YTohU2EABcD5ZcvRezJjwspgau6UyUs6JXlHmSPTs1Xpi+2sEP2AwkETQHQTh1Zi9iW2p0sbW
dD+4lp9M0FJnd9TasBAplxn6az5/2ZdZk0nnzMSAUi0voSA06kbOE9mNLQ0uSu5N7y5ro4y4zPuj
nc73z7Q3uUw4Copp337zDNhQDfG2u1KlA5psfBozQawLi43AvIvFPr12f4ihTvyx9/7i3wkfCS7R
wJgFYf8wRrujRG9zRika3xtCRnCREdHvvYoljSFGINzl1vUHqu1sIQNstRfWMuNCv2JJj6dtrfQ1
AzT1iPfjhlE3j21Igm/wq8yam+WoA09hV/7am3GiDDj6YrVzteN9X/UluX4WMlyM5awi69KIPucn
Cmj1LTGfPKsvVL1Aymfh1k4BbwSrrCBEbjanHmYWfMs+Kgryh2n4GuFnmsjO5FErrstQPx38v1Xr
r1UjBTUr88eAqOoJab3Yjh+Ns4fCMBkPD9DVyd8HsVjwpRSla9ZQJpBKnseBgJ1kZuy843CHUF+w
aln4gm9TO7jDLVH/4wTTNp18Er+7xxnYp2RtJrHlgAalILBZSYbb9TpjOuBgjXsszpD7F8pSz7Vq
Lkcc6ZHYjxIMGxozzHED9bgsuIYPq2qyUGPbaRAvMfsDWzHQCARIpNyGdjZmY2hIQrFEWYn+HwBs
wukSXj3JVQcD7d2K/t9HSH0bXDhsPpg0eQ6bi84sPUgatKZEAfM658O+oxtijyGNdoZmnp0Nl4RF
6qbMx2Qb/5etzr3gdZxaEudDlWT7khJVFwarUvmRy//ul5zk52vm8RHMS9ZDhui+lzqhPGiXu0hB
n9c1rv4q5uJxLwQTGaDflUJ0PB1QEbNIpb/V6JHnJ9tXoQRTRv6EFJZ5fu7MQH+hfRwfMqht8yYs
oJ2uw3XgBFDNppAXGLUmsi1t6BjJAD6BV2WCDIWiAxhNWLsPNDk6WOj6Qg6M5WCzvJkW3Q16hyvj
dm69EdkR33GoRHawuvCAsNSb36yimQOVdQ3a8Bk2ZJXlYKRpqid/0FqwTpbex7KBdqggMSs5GfS4
+IhRyE8ka+k4IBiZWEjkYP/EAoqFC9i+LQ7fG690hBHyDjPa3H5eb+fKAo/AjhPii563BofAlX1f
S5k3efUROYp5gaSecNT/gSK05yA4TGAcDFTBeoYNUNpFwjQF03C2NqmcyrnHUz78zpgapD6EuyA6
NJ4ujzEmTxvlo9R0BSxf33x7OOwLlgN1vnGG2omiEOT+DWRsMKwPUlaF/ptWnBbg+owrV/r6setz
fcbN2TiXxGjIl9axaatMMiRt2OgZK0NaA8fBRfTTFd6Y/cJ0a6d7q2AYQvLlSS388g4QJf4kK7WP
jz9Xc1irt8OiRTsyT2GzOTn/8xh4kygmrdiMlksL9+Hx5PhBdbX4j91xZbxWKycMljhdlK1XD+mH
1WiLkmOp07rclZvBjzGxwS4/aIV4QYEcl/ocHMTP2mVPZj0r977o3AqxSdHA5ECLpA4tPk9/gWtw
LI9za8MEqxFY0/rgsScH5rZQ+KFlmzwVwTAPDOfijnyFw2sgb481Kb8FITzDZ3SNyX2oRwjnAeAw
7UuUWkTHcMPuF6rseMWMTBlDSrrNOxn0rm9WKFwb6mIvhx6itVMsJz+HYZ9V6FxCkffhpQ0IBvmo
nJaqZLim9kFqyM1G9D5Lv1N1vdzPa7IQP3RkBjMhdjzs6b026d3IyL0nsE1BJBQfYvILPqmzpIxQ
fZ6vt4sWiQkAcc8qnvmlCYX/tj9PaBjlhTe8RtDRBY5ntSYp8zRQSzNw6xSrjxRNESDkUkMxjV1F
dKhXjVnr9vE6P2AUPoiOLiAcAfOo+7YKisXxRmjE4juGOlxTPlkkIM0PLQPvT8pZGuc8bzZXHFQv
u9ke15O7Ri8E2vTCJVIVeQWb+PlshHjerM5ToGMcBr086WU8dvMgV+cBEoQgcQb9Z7R1Rl335mHm
8kzSE1d9DBOoMCya0kZdwwSceUrj6joGJ/s3qOl2oYtFNs+8bCNYFl4WBTCd3LuurPvhW+SE0nOE
eDJXpxq3HVSoERZOvBqEUKtFcpC/5XR3KhQatjB7CbB5Asah/igfK5ox+//NqY3cbpDufPqdrEyn
eQ6182oXDoKugZsA5NfZRZzqL7hT4M3Ue+mSY+Fy3vcVVjWVdwhFjRFyy+SR5DUcohr92wRsn+P0
prUldvWR1GNHKWGgFC7FtlI0hUdtul/sNbRR22Gxr05EC2/GypmnsmhHj7G8sptymKYY2/lVE3Sj
tEunERtL717+sBiNzVe6/MRGpfbfQO+mzzb8Hs0tCvY71KhhG43q9ns/j79XYhjePxZtjNrpPAG4
rgqP+vzsPI6S437E/6PIhRXCriwXZ8vwSznp+MqtHhEiA4kzrLuRJ5xgzAJsEAbkXs6f0kE4Wh2n
nshnlIjaw2p4hLPt5g+deDOX9V6slP8oyaGuetYZ6641ZPam9d7RAAvGOZHHIrbqUbGwtucoImJ1
Jt4jiGiZhBoMgBIKNxLqq7IZTriMdLokNHxkBeyXkwgTas25rbxqXDrXnpYfpimQNjDESsk3HtC/
qzA1EM+jASQbS+qodN/V/aG1D0q/79CTybjqu5DVb6zgEyPzdos8PJuKJySYmVEh0IGE7fCUc4ll
JAZMD656wMNKnpdY9zfxsZ8eFo4N9pQ5IFVRDqHCcKnFy0qg/hlLq2xN+zABC1VVS4DTx1LhFoem
h0fisMp9gc16PyhuqG6n6w8WsQzbQQg3ZgRDy77f9U/43mGZgm4coj4rSf9OA6OiNKXBngZjLbav
CwoDKek72QAdzLUSwYHL6hhDRJRvmXLR65+wGVE1+JU0FvkLt5w+Qympmc2nunA0RihuDunmAe/O
zJZDhVWSfEi6TFxKOuPyXGR8+NARR8xVG/iyinKN5zhk1p4q9gNxhcFQle0VPHVtL3whx6HdboLY
iM8DyajUyA7zkVlmAeEA5QrrVK1132Mb3OnvP/owx3naTLOBDhgxAwusRZlwXEcfYLcwlYk2O896
UywT5gSOB7tfM/v+HAR3AOWnsv7Z5MRBIFb32MjPuSIdxAsgcwei+KPhx69HrTpgcSQ+O2Ha8uI+
6CTLE6+GJT+qZ0Nz6z/gYK/a5umhQ3CgME0arHPkwvscyhRdKMFoh1r4Xzc5z+Qx2gQiKLCnAtyP
RDxnX+hw1ShPySUy+WbYDrPDOYYAzodtzYP3HJl3hJGwWLy574FlFyO7BbAFRk1rnZkn4ze5PFR5
Grx0QeZhb0u8jQpWNX35OSSbCdQtVgUrseh0hs64oajDh/5EFjhf6C0+OyS14rDhQqhjfqkhu0Pc
qT8sMaAYWqlx5VKnVBporEyFtEW2bisVkzApzW4iRBifkKNgN/O8lDN0fTXXA67y+pL72lpN0z5a
CajZ0qOWwi9qwNLe4H5X6AeDsMYxXmdV11QChHl+VVMFRLgPJ1c6PknMHtju2QiPnJHpwWudvimE
1lUFlcjSDwpVUXyL7zHQCInhNtXm5QM+7WNi892bprwPySjnBchOyyJoyhy2lI6RwMgxRgy8ln2A
6rP25IhkFfEQEkWMx8FAAoP4wpPE9csCiDlqgRTnOGGYAH07WSMURGEcM0NB7+ID0z26QbsjsKfN
EpiE3QcXzsd/0exbtjaK/akQtDMwi6dgMhB/IuiaT+Pkh8hZCBPnAZRjlzNeFJCQShQ4IgxVCggR
GeFfY6OVdxHW4O/K+Swqj3hIJJs8PgrAKfRY6Lw+UpWj/Gkg6pXjqUtc5DLsx8kQwtDjDDiu1vzq
97ObaHAiTxZk90NzXVEChXOPK2k370EV1RO5no67jHcowbRGW1IwnWEPfXWKaJTDj9W/Wl2NEAC9
tZWfgvQ2gtZCggX3MJaN/HhHHWtVjdbbCTt4Nh9lloAdwAW1+26PgbrkhQ9L05fYAgZ0g5oE3Sru
xUF177zx7SFvmLwfo1uf/tYG5aeHHw3Kh8C9iIqrmTktKdwfRzQOv1efacvGpWRA0AO0xrRlmA90
Az9O6B59DgHe4iqGzdIjNBe+bcVrkPKgO2z+JWROqd5IstKkwDZPSw/NCY8KOTI92qzwJOoOjilj
f2gnv4a88zz6MYjniFt6l7lO/yWTqjGVGP4QseIcV097H0HYonts3eq2jjixNEqidyYRPVccjt9e
uTB7JQdHKFwlMv26/j0mpIzTBj2gl2iy2vvyJSyMUieKRTXbOZkyFWXWAEK7TsvSIiuQIOSt4aWS
yqOQKGc1TP91AXOMfkEXoCDHlLuJlSMb0SYG7ymFqupWBWtP11gcm+gXvQLh/xM7lPFmn0Rofrt5
iI56vk8DLum8YsmhYN0jAMUMXJuEvkW1g2FMCZ8QXdfOM+Ozaj40JyG8R4tRzsE1+wmt2lCBKFi1
5EBTEGJ1zUlTV7MwvjSrGCDnEWC/BMxwdd9Q6eDoS64OjvtcTbGb4iFx9e556A9+tDT1O2ibCRow
20GtF/9SW2AFUhdkqcic1xXIOgyVaES+PXhJUvEHr7/HhOr2zh7UVGl2kZ2Z6uNjt5pxtQhsAzT+
OKBeZ8iLZHicNlBVMKKFJOGsJOd0iBn/XlM9+E08rw9shxjv8p3iRiQTr6qO5NRej51ite5mSuld
OKle3U8PJkrl65Di0Csz9trkp7bG4YqYd9Gcgi7H/Q+BkPIk++TpNTiA+O8VDWFZhQEWMtgurSzh
j1cIxmegzom0zPHqjPFj4VJotelNf0MMgdWDdOsJFvC2V1/h2JEDC7dMlguqaDwGugEEfOz7g30k
QYS2vJPjoWR3jvyOlfBCMCxR/pdcp7qgeQfdS3TBAlBf52OJMO5DLKzOAyel72qCIq5DwtzHtvNY
fVXr6qFZKmlAq/GZ6QZU05if1EOC1AhDfzmioQ6d0x9fD0m1hufYRYxG/Gc7Us/FuteN9p+7x6K0
0O77hTYFDoCU6Izs9Il01wBE3FJnmWrOMX0kBCxNTRaDHEVFinvMqfEQJ1qDzdwL1GXrtGOXL95t
VR3nX+O+bimq0P3wKtuYT5ZEBNCc9qUBfiGQR72aoVX6oYMHe9o4J32GYYb9/sJtDGDLRBPpCBMk
ZV6Q2Rt4OH1QWBzVOnBUHvGdOtsPr0NcxNVaL+Wof/DpozD3QtvgCFCM0hnbkVPuLmmrZPOFIWHe
jccQrnG3baX9NoBhbCvKEvli2+DEqStxJSxWY7i14g8SlfWfAImcHbIUo5U09wdLdTfbfz6O7vJN
zBEvF09W6RN3KPoJ7XA5PlDknhwSpA1dZfdmJ8QBu/XumH8YzfHJTEf8RqpdpLKkuRrIIM9bGI0I
3HVGocOJzPPtc+zNn8BaIv//elAIsbn/FDhlfJeUSySjwf7EKxs4blNXiD4kyuhXH22JhJfcbsDU
Q8XyxWotPGurDGKoKNaQg2ED+MVbAwfbp4fb+yjWNLOy09nR8vV4toyW+cUgkI8Mj027DvU9Q2GC
OzDtQIgFsFC62tf1Af4oC8i8vYd2ZFI2x5Sf21rduFF1DPQ3XjWfax+UQgiuuyaAEqoS+DF/zvx/
3erxHPRtUlTYWty4BzEEE9IfP2yUnAyeQuFimXzzfHYyl86wvbuDk4hgly6x560Hk6XgWyfmDV/U
LKoxAVKfR2f7BuHBgzSOgLM3MUqBMbSqHaHY077TygXt0CENdjn3t1etiVJMRGYFMCRPDhd94G6C
/RNwZ9XGHrliry9oZf94c4axN1oHLr1uCsHPqdCnIc0C6EagR8gKg8ywM9iu/84Ai3eNvQTqcW1e
uZJJ8O8z5G+JOhEV0oBrhrLFyp2TrdywgKm+YhxlrcQT7TUlNE+SMwzCv1YkrVWWii8cDhq8jQSS
34br5X6hzYwm1UXXxJbFZD0X5+r3CBVzE1trscZ8sbsFD+qPw73GbRL/0Y+rMl9ceXoCqK/mNs3F
qw2hakXU/zuPg19Rda1d2QaX0lLhOOv9g+T2hRr/TzesJuaAJzpo+Q7Pcy18GsOKpnnFLQsPAhQP
dhg8zPnTCYik2txL4j67gZOTlkryHrMnoQZx30ojWeHcXFv4q1MIrsrCeerq4+Bh96lrIsBAKlsC
dH3TwXNMzWqjiJKJ9pXcXwavkSZEWNma0jZeLKgebfZ72O0h/F8VpxxtrSKLJE6s2Ub26VWsQfWU
/UV3dE98lgCPr3EZwESiOkzhZomHM2S3dsAVBoX24zuaqBx87PfxmmQ+TJlPNNB/p8p2DjcnT18Q
Drgv6GXx4rFrbEoDR3/izNybgZPkfxpKUJnN1BEJqaMDzTiPIA/yaPDrRpE9cURsQOvNdsroBRch
uRq+Fb6ViA/atmX7u/ps0qPMIROb55taUvu206QtpSQ7rD2/WtbaRyT96bmCc3Htoe1CEM6rkFRP
G/xNLqRvX+2WQYBSEaxaep/pS2a24k42kmT2GTcQtoDDxSnmBjabK8UQqQl2ngve921HPnQ0JifK
J8aDY+pQttk3CGeUi6+p1Nteesnunu6k5UA65V0rKKXB20CEtDv1mWzB3Sz/DSQUbrwVSXMs7YSJ
QJQARXmcTS4YeHdD+weGUz0meEnbVPbW0pKb0dp5KgsIXtudOTnKNNuInoxhWxqJqbNljvuV/rUG
zdso/9cr0zFIEfm96k1GSjuqxeJTAbIt4Nw/oeudyxbiK1i0tFWlKrxVffPStclIGdmLE3wIzjdR
PI3EpXLzpF5YJUr0+LbFk84zndPdcOJWminE/M1lsG8sgoosjZBmMQw5faBZscqHwvppNmy6Wqlx
JBM+7Ve/bdnkOwid7K0ZH17guZKoe9pwSawuM3FzkrtyqJqVIO6rDJyqx1UW5Pyq3Jwhz/O7E801
tZnAklzVTgr1o7b6VOSuJFWTTKO6S9x8OWzh6X7VGw5DF+HcVr78mvTE1KF/o+S1+rsVlxwYZc+4
XwhCgUrjKAa7mxlVccheKpdl02eqhcJ+OjkKKnADkfbFN+CTn3v+e0JiTB0/YKAqHYKbK42/VOm2
BWqow4ogyqBsQdHUHC58hBU3Wht2zTCbg6XiEaj6PKF16Bgqn6dCd15xz1rHtXduht+TuVX/Qj08
WZwzwReYyNoAH1qKbLIsJgP94TmMaNt8poyTUBA/wL+sM96vNXtC2nWZd0g7XYl3FF75niOrEfH/
kC6q7Z3LfRPAAs2fRIaCMlP91wLXU6O0rxKhGvnSmzTsFSMRMukY9xASbsGp7AUSIjJ/TuFPq7yP
9uBeWS5zzTxhGyDsotGO3VUO3gkssbgYqlRT8IBLYpcJOoww0u/qCyA6K25hojInTwxAcD0OyI98
QqQFbSBiQ13H+iq1yeM7yuSZKQNCSew3cdObqn/n2kCTMVdXT2tCJdl7CqYG3Jcc+yIUVY/I1CWR
lnqcHQCDmY+ShL0+sfAtF3w5XN1QOZ3K4ki9RmgbGiBijbTtracgikf23a3KA6lFvNX0w2FM2Z5x
Y5eWZxyw0yOhGHYt+YXEu41Csa7tVO+9H/AQVVN0HPuKMgrItGBmYXQKv/rP9C5s+5D2fyhfr4lg
4xFfY+p7o5ne/u4+dMkEECN7LamH/p9ZhFkXpq2oHpGUV39CMiOK1oNvj1Lo97G9Ks1itYowWFkz
lA6XKOnToqkudX+5ecayF6VcZRODLDWAxhPKxrhPgK/mGUnCYsUgfYZa3rT14CrVCAkykk1t6GXY
dmvj5e87TYrgG8ck/j4RCxpaNgXPUyZzbb8YBkXlUKEQ1KmHF18i9W9AnKDZnNwOG8/Z5XI+3KJ4
JoO+IUMbhoK7nG13Q3lyIHUVC1RgNGcyPWf0ztcJwnrAkuiKFSoJ3luaGqkd4Q66tExBj6t2masn
NSJtOIvcEs307HYsERcNTCLcgI2LskCV/yrYhLfOX736fGA2FgesEbADeDY0MygfW2OM7elIyUUh
w2Nu0NNfTW2nm+cRdU8NqFW9jbaXJo4YODyYa+GtW0aL/73KANZmXo3kRLvel18BCj81BE7joNqu
InQ5Y67XfDORpoh1A23JWiaPipvGydlqY6t20k0AbFTyA5mGSS5V6kmr5cYfOCq6P0z2QZqAhszA
ijBe2I/asGVLzHu8n8EiaZs7zfQ2Hn/bsOZLfCdqepNCunD+MQPOLdPVRIAVQsGR5DeeIkBrGmkW
L5KLtIZa/Yj6zHFV4Hluv1fsCNV8ainxRd78CW6qk55QeIvnlZNU014rorUSTgX1eve+hdFZ9Iol
WPVlH4JcZSWbdhuYmwU0t44RSzuwlL0yhU/wpNkyzCP8964ZflDliGI8kNcbHbkXvs0b+d1CI3JJ
6HDc2+9EIgHVL6nDMn/T8HkQSSkL+rhdnCoLfog0i9IEnon55KhZFZ/Rsa6G4MI/qQWImjwQ3rhm
RXbfffjTFa/vFg+qBNaid82NGAf9v/UGQf3B0i3HTOHkdLkKSRNCMkKwV0IT9QG8WLJV68lQ7N/p
3an0ThdPEf/Gi9hCis+PsCw//LhxSWpCV607+kmaO0yPvRdRgFjY8GCRmaMnHogEpMvoqABHW8n7
GM2Aq2Ad9n0/FN4pSKVEt+EOuGeMeoHl+GssInziyiNwuVpJi0EFQq490YAeJMqJCNLXNRA1Dybw
13S1u/qzr6tn1gPyAKP5z/ppMYfWs4t+K9wiZk5oIHsbU+fB1iurVdfHt/xPzLXiNXB7nUj+jz42
sAPS5vhkWXKet8HKp2Wc8LG6JLV2VEH7T67YvAQX8MKWMOJVXUjTU1TXssTH3iFWx3YrAzP17tbf
ZoZqozLCQiRRicxWtGypVc9MJMtiPqepbNqKsMk8V3l2E228Kgj8cauMOAkikR6qm5hZYoo+flgu
nn1ckpzqLmrg5nFGUKQU4cbEy5xqZXf63JvP8fSDYNSHJ9XmE9xpYxrRJTQC/drv6ZmGyaOFJ7Dt
/Dq8yTm7eInhlT4j1AAuv030oMq+td1gHte5oZP6gYzqR2J86pZuMA2jdi7z7jRAS0lWzoXKGY2O
X5U3JEVAT2roW3Aeu3symi6R4hNcWNM5hnafp5vgsm/sw0a04oUcjKOyyRbk5UXDlZRlqKBfiuU/
BzSS73jflazcZNQy1MBCNLP7+9b/ZprZlbN/fq8M6/4NRTsFg5GSPMMBfAZ2dn83lSRxnuWVpimq
E+u3Q9sqcYQZM5Ax62suR+md90aO+t9TAgpCGcCXVszWwLauZASLeaPL4LICJgzyG7RId1HR0mjK
//BQaiJvCOvZPmN5rEXsQ8PcUE1dl/OTPxr9FgNp5H9veM8MOPKnPILJrD7VZRV7VxR4Ei0ro3X0
YctGzY0sdlWhcD3tRnCNRHCyGYJm2c0HCD0UVgDBnc9SXKOEIpOQ8UMGHvMCyTyZj4hCf51VaFsP
JIBZMFj5REJntzYQzLC0MuYinatBAAxCixg1h7jYs5ad81NdTIFXq/+KQ2Gn4/gEoQO6hwwKtwKZ
x8mubkUOli39KOkzayhyDUGc/m67pN5CVg5jhcTqWPZLsCGwpub1OF7la55R/fTaINHI9lVtdRTZ
Aa/v0kpm5ADDodPxwFqKwBLiI2piMQMmIKkrtAfLmp65Il4IW8YHHc2mvu31fYh0UNkC5hQewuXu
o/CuSvClhguPegwBQXeEe0SnjAj8rL1xVZOpycVMnJrt46XD99TZGhsNPYIhWR3JOS5s85Xyzp2i
gfT21YB124biyFJYX5MzGEHancRN0+WsWOvstXUw3IZiNkGnBg0yWXIgABLrrTF3lyyj1eK4nDSL
OlmL6PUWfNSJufkBL2a6AB8T1Yhh5O5FgxT9y+wvVqN7UimrDAj/a97KKxfg31lEKBDgTavgLtVS
+CC6xveehdu0T/5bQLUpOGZlxhWTY7Gszu4oZM+3Ll1KSl7Nyl17XIjvJQuYxK9AIWYOB8yYkTsD
3BW5IO4dVLaWyLHrqGY4W+kxL60y/g83kIx5No0qMZeP2CfOtAZgDLK7dYyUrA7j9hB3hBNL9nog
MDHM2xAFzVgfUbtrnhzASsua0LBDoLkcjfj2Z6VF686uAnC4RlKuAgqTP7XDZ6aTVksaONWRR9qm
WRizu3LlSl5B3vEo+QZxBCIOtdq3cU9nwNhzO7Jifo53HpFwlCVInzcHzfvPA6/Lv8DWDuQ3lzmG
gENh2XKONnUOfgHBQZ4fROPn9RjS2C5vSi2c8ddee5j71i/Oz6eMpmQJYxEaG5RmmE75ZZuu2zzc
7anx+/k1bM/6xmDVZq5NJilLfbHmPHq+GbaT9RrateBMXv5T47aAVgbZ3wrgLYsCVRYCjKR3W6Ax
0mSCvc47zjO23LyI25m5fEAdSueN7FhIcVK0bcRf4pkHpdDC9iGKz54ithFAhiNQv2sE/g66BZ4F
9Mpf6H48v0n1sDvzUEdeCS0uTHjcrpplCD3CgFjWZ+EF6DC8aqumqoXBEGZzadKLaKAOzboI3tRj
h2U0GRRmMeaDPBvMOuMPwNqjRGULyXrm4xnYGmY6VKA9dUw+naOYxNO572f3aqD9t4GoHTJfDeuw
cEp3iWFeKTMsILjXDDNAOhaPORQL1i8b24xnbr1B7m9+8wi4JI8Jj0RDde5oWEhl5MBYakvHRRfx
bHjUEFYUKjJAEviIT+3EbVdVsvtve32SPWuHUxyWYDIecFAgsgIBDqbfOgSBPKWulyWwv792srMb
2utGR5jc/PlpluDNhQQnRUc9BVrzTPqTW57mMlZWTqYmNy1uZl3Bvv4H7QsdE+jaPoBE+dxk8FWa
tkGtXmh1BZG1sf5j0pPnUx3cJnD9WpnUdIrNpydYIPNtygBCmDNrFgY6m/XHmOLxdKXsD2QhzFop
s7h9xzfbh6ccG3VyaAPxcmWaIYqw78hGV9y/Wigm3n/06Em+HWw1teyVjvUzt367eTJtgoPWqsmA
sjWo/m1pKClkODMgnhYFSsibq+4LqZasWqBIY6ChVY8ZdYUpkcI1+AFGDeO8kXTDaSP3fL5HQdLK
aURq7X7Rt4GtQ2ZxPyb+CKKkmxUi5UB821Iw5pPB+3SsyPzM1BUXvI9zwsdnc206jHx6+412fEft
N3xF3D2ORBv6yb+XJdyxzUoK4kMDUaadaDowFypB4BhuEHIt/L1R/cj+LDwNXz6QLe25DsNIsU2j
vs0Qk3CLwbtNAR6gDfWnyxjCSy8bhCm5vOczU3thzzbtHaWqi406KnU2giF4+WF6qHaLNwfprEB0
Rb/NneFcJUml03bykdoiDQnyj2Rcj5hxAlfOkbZKvKPNhQUui8j56WABJ7FXrru2GNsZVS4a5zm1
aqLWOBb17jIremEHZTAefkIAoNVfOH+UF3aWpKjXTXBDYsxHVVjed+nFMoIVlze665mRhWuvqB5V
2+MkaKPMmJnNnres4xjpwxQf6MNDlWsuVcvuZiqyOYg1eEV2fV98fmj534aLPFnV6ztJ55xSvAJ2
VW4/y9/UV1z100SSHXmX6T/HrxqHrc+nxWJuJrYqPdAisfFqpr53IUYtqLa8SKKSlksBDIJmTCGm
M2J5idLoXFxwkdfz6wvKJh4mCAm7mrk/ixyuutgLxA9QbUY/8MbmuJym2dsnb/rFIx57y3B6PSOS
LEXXwavqbDgG1E3q5IARREhibHvHsNb9rkU9zpojDYclOSo+N8fTv2puxHeUcokY33nMRIWaI+zF
Gd3aZW4O1l5pfvLCwbzTZGKHxlac7ghLQkDkY0uk8BJ++8nV3jaUqN67uNj74AjEZk/bapUOsFiL
dd8W6vFHl4Af8JBcZGKOBPtU4KRNLyxdBFSMDwfc71NVTbOxTbZ67xXOgbcJru8G55tc4/h+7jyg
zEvglfdCpQvvuuyYMxdrVsfygfcZ4t1E1KEGDar2D0xRAcmrFYWB3kXyUZg0CW7UhEBtaOxZ79xs
szCHyYt/nZ3X5VkCeRNpjtIHiC+G6M786mfwVTj9gc/5UvfUySZymrH30zBzsGNfiTd4BV1/yVY0
nPRN76ILvenIFITHiWMwweiyPKcjwXzsHrJ2nW3CDY9MOYBvmHWtgfHE6i/VJKNGzvV+Ib7J5/zb
7lPxu3biC8Jgepdxyg02bOBq0ZWBGTJN3dODGRsCoA2hdbokEXqJzMviDx6gme8Ey8tXvjX7bOWx
O0YZvA72f2x+TwHcjdfIdwaaOGROfK7UakNwFgfFTqDUU4WAFSXvQmUq0lZ3CDntn4YwWxjTIIJe
a1IMoPI8lpLWC8EjsxkvUh5/GqdJJc9TRpGDkELSdrVjZeaxGAJt4j5lh8O9USedL4T1FGU1H6Ky
45RkVckLB4R+frWpDnqA7jJkqJOU6o2w/fTJfdtw7O8m3c0cJY8ejQPX2yaJxgYP/Xrl8yqbkp/j
/y4cAWfmKH5UOw7NgHNvJY7lurEIIHSkHOoV0/8dj8UCcHpglWeRbM/qlE1va+idlX6M1gac0Fbn
TV76COS5REG3vevWJVA0lrN6iOpNXdZYjA6H6LddgkvVeHGCixodyKyTqC2x+WLY+I71+1MgSjXV
wz0oiiPGhP7YZmvYZQ6/X3WFKYhgb9psCFuSnNRLCI+SADwnhl9CKV8Kl6UiKr6U3eGuOSXNtllr
sgJx1JSGY4wuLexySJnajeiKdO+NJZn8iWB0NiJ9YZtztX4EfJuPGwOnGi/SW3M2ZV+sah37ThCo
TLWTaeL2shNOJ7Q29QZQ8RbQotw9zVk51suRx3rbzvArSUOel5do87jswS0Pusd95WDhbG2RHQZ/
mAyF7QiZNWLkkzGCHYjizrUpu0erKFqmBVP05DL6KEdw2GRWhLBfr1uZbbTevwg2pV4NCKFpDha8
ShWuiUIrXhDHbaU7Sf9T6q85zPuAMpBWA4VFxj1b71NeZsS71HICBih3S8nPJtGfk4IrZTK7a+Ri
UsKvrk2TiUO/gLdczkXaQ2vbQQewSydpeVmkTPQA+KtvMe3GC13ZvI9gAWEU9cMDWkBceYqW1izC
Q5LDh4FOWPj1TG9iv+R9cLVCboYtrarGTvAbU1GH1hCzIHo9ohnJO1ZkJUM9aEG5Ys75qVaM0arU
G3b2G/1HE6KjNU7tnvzU8/iwzdgXIpz4eUNf3BWfqLG3auEjEVnWM4bCmr7kw1JKp98MGrDNl4G0
p54Epr4+EUNUcvVLWfEOAWyuMoROrJbOQunZjRglabCJwxh7U5xHTyLlg/wrDAhtnSzmVtyjUzwz
29d6X0f1yizJ/3Gz7K2ZPmr2qqHee3ZDEyjK9hn58ddSRvuYAUI0GTUlRe/WH9lmWR8RyotWop6u
afGhoia3mXqoB0jY19CYmet3qHc+mCfh+CsbdJk6jeOtlGJI7CqtH+YE7+eHyysZPG5tFEtgpqP0
Gefse1q0IL+TQlYMsTJaXpRsiLZ6CAbPj0YmaoLdmS0/ifddlWwAnKCol3ZDV+ItVtvaJ8OJHCuS
CAp1/YCJ00DXZqzC4bCJZVGoO5NF7ef8ucSQGsqxC9dmQJKqn5bwVx3aqHPefDriuLereWn8+nBJ
QaF4B6BfqiF6VDCqLp3m16E3ySvVMDp2NRX5OkR7sPiwAk6VlWdgkfhJ9YpmszxA16bbePSd/vNe
4IeFkqSCz3Oe/tX78FlFGkJYTt1HRfYmrhhPT2QgyBobs7+APi1b64hyVmOji7bwRD7brIjl8LPX
qfNwiGnKxOgmrKwAzH20v0xLw0ROiKNBuI1AuP5wkMS8B5dmaE37DxktcXoIbzaYSrEub1oBCQuT
5hr3PvykYA7CRAzY368TueOZDqkxPjJfJa9I6nQSEHTEhNd231CKTk+8gp7NJP7AxlrfAvQY0RWE
hQu+baqug2Iaq7lrn57yeL/9aXqZ6IUP8OkUDP20nchh3KQUqGBlk6YBH0VRLU3uSrEEglDyqUB4
sleTIOBJHbQC42aBJQkx4oM5esKDV1VFWXZOHkPsR4xu7kmB0NbUWjHo+CHRz45+AUu+UMhfo2JD
Df1FiV6AeI3LypBjYgQX+f27E1RBB40E1BNVqZpLdqu+N5fOHPFKSpBS3ORQTI6fCqmoQ2Ln/V+U
jnxO1p7wMo3XdKM21HyYVeQpvew73wuGSmtSp17kLVocf+Y1tJilqq5nLnTY8tlC3614XH7sLNFC
9HeELENcUUfawTzhKLX9e7jQIZ4G+7bwXkF5pdO1Y9IKN6SZYGJcJ+XFGHncZ40PhZLMn0oXYec5
yGIcjs420tv4EYAyxt0XEjUs2pOcWEuxWEozPRACod7Ct1LCR2/FydFb67ddp04hKTfqCKRD70La
Qiq0Jw6r83FdDTQOB42F8la/wQJ7Dd2VZiJgtaSG8xSE6FGVXVCOtX9e0unkqyVArxVMoSwwFSCh
YbBRkkCzQ/080RJ/cI59n59iz32kgu8nyKGS0m4u+whK3TFD5Pw9EsNtMYr6BRkG5dd2HotSqulu
YMmcaIasnj3cArzU6/ZCpmdVvOn4T+GOVKoesmPYK95kALtrvElBLCATDSXmdUveEL3NxnNMLXUg
HUlrlarjPvxDAjR9OVbkrnOj65JN9sc0tTAQECuoo3EvNlUtUXpu1CpYHjuJ1YJUmmjOxs558jdm
WsyZ/tTK054JJnDQA42bNBWYU+GYQfx+q+/z9uRQ3VSwmqtMP77qPUt3I0A+CeJ+GShc6YVY/Crv
BEUSzVCxwgkI7FFDu0PbRxPHIweZm9lQlYIfP+kaSjfOj/DclKelxecr0P8CSpUqqQ+UyO+wquo/
p8hO+4xf6plQUu+idKJ4x9Ne8/acnrmh9QqtCqp4EVVYdzju1kP5R0ieUGwN+pfnm/d6rP6s/nIm
Blkm4VeHZHwypyvyAnP/+BOQaGlVHVuq0fqKa8v3qUFyhrevpHo097fKxV8vSH7GZM4YwV2kJVe5
gneFQJ38C6i/KO81wQAquZ6jtHZjB2h0ua9Hy5vON2uRBI0Dq71eX+zJxMUKUniE0Eru3XDqETEc
HAqjU6HhBzqtEs9SG1GKE4Sp1a9C/3BRX7BJi/5AKkLbDNusrNtorA2Xf8Yo8QmrW4jSqBitZz9I
OsfUa6rytsS0leDKt4aVih0T7+wqbUFT+cYN+UHAxCIfM3m0m7mYSB46yLok4KCFjIqYcir9rFLd
9YpdnQvPgp4bvssv4g9HBuHZSrc/6d3O/7ptrOevtAiEr27R7r6chcYc1o4VVPYVU9RkbEeMhpmZ
7VBkrNIOegOPIq7mQd5Uwqc7fJQgZ898yNfE1tJMnaUV8m+9C8hZfe5NjeP13fXt6PeRZPSolfkI
2fwc9SPHmoZrqA0eggzou7y3YFXCsZKEhL+PabtAqEGudfsAzF8U1IzUnlMMPILPFn5i38V/2+Xc
OITGvW3KXPl0LxJsPvekvdQI/lFzyrh7yceUmbGhirPBokOMlQoVjY0+BLG80bTo/laDlWpdMtbi
zW7ZszLb5kWpHC1ELcJg/bpNu6qI3EMBNCSAk+a5aWAc3XDpTNZBZ4lrACmnRQOuXSgDE/rKhc4e
TtlErhe3mwNMTKwb+fk6ag/dznaH/kJX1MiiiDjznqoc1g4+//sWZVZpzERnI9jfDGacoDsZFI0Z
/KkaF1PPpzUzfP6aiKOlIM9UG5D+GpJ4bMfMtPQkfx8K7hG4PC86fNwO6vvEa2js+IAshoNJhuE6
ULSSMt4fWnmXDOMW9Enw+P5bibu2rAe1oTxX69kA6esRKp4MrMMC5EtEKZFGi/pUaG2wLf8sYAX+
sR2kFgtnijZXCZ8vRLARs8LHfvmtlMXPFI9LuimfKjdRebrAUr8Ft4dzvlUdL8S1EaRLkWdQoDem
EuonwWzM8mAWsyyqWWqgGU5RdSmQ+CiUmvxh65NgXA/J4W4QfXXWpb3eMYAZcNd/Pxla+RgU3uMZ
8BhCngR3FPG9HpVlZYlPqYGly0PKitR4niwFnWXzHXQ9KbKs4fFEQVk2DuStqNXnPsNlH9vPlnhG
3zFBXvDuUQHJ2TK70W5wkY8LoR7Tu0LvaPSBcY+eANIDUOSvd67FNDsJeZMI7agHoRduqRba8JI9
Usc4PLe014rsQ55wOutzwyVARlfBpxH6vysKMN9yprW0ouu3x3UgLaKcWpDDo1PokcpWCHEiXU+T
h9yRSqV2qn09UWv4NWR8GcCih+s2cWOLEpkBQ0Lk7DCPWvFYFoaqWuFlPZkOcQoAZ9I7QqWqcZQK
M9x1jUVqTWFfJBc8Cim1gWa713MtTXfK/lE+ZC/+QqypbMCJeaHhECvazHGov7WYLQixL56/SMhz
jdtLZ1yGKGAVcD40aQ+qAS7fWpywynADp2APK43404hvjDq1dWVswdZHTkI/uQn9ZPx1wc01tZZ7
Ml0J5rubP3oK0jbp+Ezv8I9FbWihz+W8WH6WsNHeHAFpodfhw0w6f1WZyMwK3ZJqZiNlKcB1EBzq
iR44OuIrsMaRmOARlkdDGRfOo1aZK57M8+SIP1lJcxlQlQ8GlV6zPMCwWbHQJi6JieTkBqn+J/NJ
ORyN/GiOs3BYA6uScV3f/JEj3+mdqfqeHccxn33ta1mjtN1tfCBBGjZwnka0XoxHVz7rXXYYcKxS
bD7EwQjobW0SqNQA6ZOB49Me8XUAm91MiTHtE1v94oXjVEflRTTlFBNaEPaxq3XJLtClYXGuKbXN
aHOWEhH7yZthtOnrVnBUXmx+72+i+xH0CIFde00PXVBeNy2fwSRo905Od4vl6KArEHG6irhQ49l+
rBF3RX5EPNRXuJLGI3rwQhwb2DsMs1DN68ABsRJXbolsDMFi2ThqQLy385Io50/XtMS5hzyQAqhZ
CvKULtEwc0ZEJ9JeiIKtZk927I3S8ptZR/a9asbF24rvWW5yhQaNsr9Dyqlvb9Iw0GtsVf/YOttl
CaqL3e3gJ0uErSD7bXiRSFZOvNhk3AdbybzkAptNdneBLqQAzBi76XKXAjf1U4+5Mo1I/14z5iHM
EWbHn8FmG1LUX6ZVRXhng4mlsG2naqaG9CvIlL5cLE+rWlcKoODd9fyVNPTMtLUdcwjdbm4B+g7v
vsIFkr8kAQtlmIQcbk4Yj0YULT1VfarZKGlF+RJ3Ya2X0a+0/VsWURjVsf8llH+uZMsSrlZQTiQH
BvFyrMfwFrYQHFgaKE3Y8BbyvV2SK8g7tKcYVHuzEsokuXwwiVR9OTBwxJnntzg4OtQNATTlTdXS
12XwV1l6cCY2+va/aYerWnw6uHCEDLxg89dOJzX1NHsm4IKd6dSOdnZi8Ja4YsGwsI0gIYD5+HtY
T4SOEgu3UsuAQZasmNSkZqwaYwAk4sV494zl4C/yZPOd1apUaySQq03tb/6bFuE0jACQPm+PqTGS
nLiGtDnbZiXbg6AnqNNNCxvFT4NdrbpbGOMWaIMBhOPCIVLJZbJU++FwmH/2HkB5E4YHuQokRS5Y
NGHduxoLjdyeOyyZLECYgEbCz53L6lQNkfAwtbA8o6VRH2ugAjXEgguH+G78e7vBzAfxp5/8CLKU
oUjaLaj1xV7DVc7+7neWUAnm+FklrLjvZ4QP1VJl5Yem9IGSmwVNzk1lCRDx2q22w1ebPzjLIu06
gAZQsFQiEf89Gz4yw1fCZGLWBu8qrsvaorIKP2sIk/kJz6BY9nYF5Ys1Qm04ls1uLC5CSLhOL6cR
TTo29NdWxCz96A6ljtJBguQSQOyu+h6S+rYlIRdTFT27VVsHOWo2v3aEEfSzMz3YXDOVeEYyzYbq
Jb0N88LkwjE6RhigJ8O18zExguG/ObBNcjybqgB+gs7e+DPyQmNAubHxgQqaV464f+jmYIdjyg0Z
LaUxeMNH6kbNwr4XDFVucRvf+zfPwsWqO81HTU2U9llxCc/7thNtGuIqQc6P0G58mfYzV1k+7efb
z5rWDEZCjECftcRL+M+XBoDoIyagSJ9xFVPaGS+hREpYdjIBwNRyU4TPg95ADIBAKvPcoAWWTTpl
236LosUDhdKxlOGz5TSEdSRUI8rpwQ1Z+Lnx2Xa/jvoHA3vFmCnc005IfFK4PjZgcEOw8I5U+bBp
5iQGkRAycfjX0r5ga1dYXB6cAUPPypyGtukoq5AnDhtyS4dJbNFLXqn/m2bzPLnMR4OIE5UUrPwR
dMbUnKtGNJRTwQoDRC/dnoI2oFMmC6Omr98bHOvGt4OgmSdsagEul7MoKt0vYiK9m8VQKbKOF7md
rP7+JHgJKAPeN8EY4Bhh/4r187FciewbLyUEtSm5DMhmv3kg2Yv4A6YF+ZZqENL/isnaV/Tn4mm0
pL6L8uZcn6/FMLQs4fLWw+VHF7a02w3k4J9LHUGSyALRGZ09JnNw8II56yCTM180vBwUTOKTojV8
sWul/TOkT/x67VEc+AuahFcwpNx0XmTFiW/g36+pDfmosB0E82qug/RpwMK3rimBwjwTpnWl5sUo
BbYjG8BQHVemGVXd8IKZRa/1gWmFVCBGgDcHR1bYbl8zhfpWUyhzirVvkiye7wIGCv9rzw2N5VRl
VBycaOwrK+ABdFZZDvLVYB9cy8/V/ZgX/ywcQWlI+Ffl96G8hiw1ilba7jEgkRmxRSQjnL/8yYKF
jU2D/ZhoNF1ve1GOEqZxBTVTS3gBkruTlpMNm2D7IMNZ8CXvUPJHmSbckrxSWtB8eqkK08SDWjEE
gMvJO8gMSdC95lWETsnl9wqoiRLT5cT90gIQ0K2GBmQpoLF1SaR25MGXhvNrgO+xEY5f5VNqp7zZ
deg4vpRiEO24CTRRtpM21RoAW2+DX0V+yWw/dLIzGLJl86NjuxhD5Zf7R2n/v4kj/IEFmlupCmGK
BQ5ny1ykyxww8y7CTH4IoItsGVPTNUO+NTytcaj3kePkHVCyuxRqo2DxsMG3KjglXclGp+tkDVfH
j3g0HAr+r3pIRHQcN9MHrL2Kc3eqqCKrajSbZsFY0nzBG7MLourfzGRtkfClBLjatcAISpGDfLPa
GTzUSE6HcSZnZKWVfFYFcIz8dyz2BnICIcLtM8o06ywngWJUd0uJ1v6B3RAzmTs34N3LXEpSdngi
fC1aOdbOvQJFx4d3Vjcdw1sjD8oIpKKG0FtAw61yNJ4DWIKf4X7qJnrqcEpkmVomyFPFWy4QTiuZ
ryLWO2AtAYUmbRktTeoixzqz8FW4D/ne0gh/VVnfbS7ZqznLWJL37AFB/fLLD5cEan3emWITyA4j
FuNlBM8SwX04Y9GhdNP7+hWpJgQdAIKisB//awc8uqp1dh/UPeqt1IhxJuqyCd0hrH6wpMrtMBsg
Wp5dS2H5GjeArVaD7NBS72/9AliwXnF9YWzi8/8UHZVbDUcNsXnAcBuRtxhaFOr8aEI80LnRXWuY
FmrxlZ5UMBGr+q0F7s4PfYC1Z+QCoqSEaJOfQzGad4PXyYN4DXA60uI1qEqZiPQAcob0X/e04L6E
oy6osRa6nDbdZHwboXSTg71pD+TuyYczLp0wgnPU0Hc3jcj8FY+sNjfxSlyzSj+jPZJaG0jmI5KS
kj0N1mND176SPXoTOd98hGOnO6OEaoMjrCAi1DRd3vz0y1mz6ICRmskjG3CXlyoWjgUjFryiKu9N
WWbU5B0G9hB50xDv/DpRSMIS4Ab7Daf1fV+TQwsBnEO3049V/nSaIBiUPxJVM8AFp0e2LqeM6Vjn
/hvV+ev5RkfpvWLpX7YuGKEBjMMqxfx7pnQLgkV85Vx6iPTpHmlBrhlenMUCH1aopITnd17901iI
ANx8THCNn1NPPScyc6XzztaTDu3OasK9zGD3A+jWdzV/cRqvw2plQ5OGwSuq4IMEoNR0f5yqDAZR
MQqysTcvsQ0r7Bqsy4k838kPB+HJ7RVF2yGdOiLJ7cFX1f4hgDsq2etQdZbX7Yvdnc12mdxRsmI1
LiAZRLaYvXkFLr4s/VCKnrqZfAlSrUi6oK5PSa9CGP9vwnOI0PMTeDrT1poJZFgqKAxoFzsx4OZF
DRp9BKonkHbyf8kuQXSQNyECrpJuYmLVaww4e/ezqAl6Z1tufhcSXekhrd65sok7UhM+xfu0fMqO
hrGEnmS99+b/cS+l2flCqUERYKtpxmw6aSO3/2cjieQXAfIlIrGluzocRVc8blQO0FEfJY8NSx+A
o6j2ALQYgtxqAQ6xKbxWxXVWJ0DnjAUDCX+3+RuEQRm/YdGfYhFx2aBt4pQsvAtxsPO8Dw5Nf/HU
K+E2Uqgt+d5PFPfiS+afOi+kF7t6/rVXodCKsqWmkBoS9pbLcnukf/HQ58uzGUw73c85Ta89H1zX
NwjN1xa84uRVteMErixUVPSqWXHTHBtD4jeV+gts/VYOG/B0dEOW1DE97GbwqFGlZjXY1S/Zfj8o
ZraeV/K5F8BeLbAlWnd6w0z4NxkGD8id5SokTervTzvxOJL8FLALUks54alyqz0jEdsIKFndJc5V
2mNUSpHlMGJXN76PqLQbv/h9l8BbxB4J4UbRvdS6t893W2ovywKDH2yRxgUn1zY2m24+nQGD371V
HWQn62QzMFZUpZ8CePJyxayWWgX8fAk7bVK3QmsobwVZx9eR8RK64p7Ko2caYYHcddZfDC/OOTKG
HqXs/U2ZM/MsGBFOLcIsVMDRJviU/d/oEWeKdbNzTFfrLIlG2Nnq7u7fdH/qZx9o6y4EyO5vULiO
jw3accVUNt3L0m8L/r55aE7Q8VaKbxPBi5oIgOPb/Iz7mqX/W0Hx3yzTbImDulYZJVDa4kRsDe7f
/9AU5Wl68cLPVnXNV01clmShls6l73jVWDC1DHQkVOqAwUedgggbNxWL3axIZ3WMkZd7EvuspzRj
2LJHgnCMhH4vm/xB7AjnCZw1rDfulkN6JrSjwyEGBiUi40wh6ofHIJr8iOaa9rfzVhzCVDm0Hy3f
CbuomLPv3g4vwc1Dd9Bz6dT7YRhiuE/1l6GtVQRqLVah4mvBC1L9N8NTY0bYsZatSzQDLShICD7o
C/qTTD9lxykwM8Z/Mv8ALaVPW6C4aBQQy5uurzAzBl9j5gPOXLYTsss7XsStfqlbVWJBMG+Q6oNc
RKUTJ7V9WfzeelLRcPXJVW3nqiQjg82TYvYr5r3roJgxsNxtRMLm6SPlNXylR/Lio/V6Fhfov4Vx
hi7JjAY+M9GSaVeUs3PliioQKxZPrsHUZ9rIx2w12B9/oU/5amz/Jb1REaSqwMZykRw63LRnKlgT
UQFte19iHNzjlzlVKOuIdrpcDzTqCdhzxG/dJ2vfqhSvfT7VKU58bF/AYKGCLpcy6cuNuI2EEPuf
nSYe25o6RL9GTKdZPYtGySTOoMfbKL8xE/BcxgeblY4htKQIaz7pGe0zEd6TW9dLIumFcpqcpr/f
6z+QhNXNnC8tcExdYI9rCiBKpwpZNOym7B6GWI/4Lb1SM88NbLF7RiV9mifMze6vX1/367s5nb6E
UlS4sr6oY/3p18bWGEl5UUoj08BDaw1JRl1/+vPMRDFh1fBuVGLiEABptHhcqzIZWp/dDjiP0XiH
/TY04tgbCYckY09qac6QhW1hDQXM1fs8Oyl0qAO10giwy/Lbr4nHShu/0afkLMZ2E4RnFLr9zxV+
or+GHVvFj9BckzgQInXDfn/qbVHv+aD+mFuqpHZuNkNThW2qh5zVEkRG4/FIGq4hXbncHGCBo/Av
uJvxOeHc/w29Pc3nuDU17BBefL9hz4ukVS+dcLBaT3lDK4eZhDKYZ189hJgiuI0GaOVUoP3yRcxh
M0vMjamBMYKyvofdX6Dg+6etX29y/gQ64DBrPVoED+lHxBEKQe7j2MwpeiIfdiWYjsuAMyeXYcAc
GJlCWtg+lsYhvWub4Hu4GTE/VG2fxL7WQxIKwXK5C1V62r9sy8CMqYaGwTxWNef6PG5mabwBs6eV
oqml3kLr4t55WJP8p6d8VFO6+yyVTtin1CcKooGpOWXP7weZY7/BZIz0T820ObQoJpPC5hevfYtP
9Gj9/scPCUhS0jyP8jvNDtjop6fsf5QqyUcKizAhsZqdRLLByIMoxI1vjQkw7Hyvly4/RgSlrhHy
TnModxX2wve8rNzzSIbqJv4DDOmnM+qZSXBr+UqZBvHQ3W3d5VvxRqSWC84P7vU9gy8UTlgMYFkY
8cyVNedMRJJLTWZJ0n3zZUzVIp75dMCgJ5MmFlcnnhpUzVprCScueWVkdSyDiP+YmMTWhm3mXRSX
w1SFCb6256g0I4vHakmeokaq/HOaFY6HNeWi9T0FBTtRcShqMETK1Emu2+/Y7Wi3OV+j5W7qJ95D
GlbrSO/cBb3u92RLG5IyIkC2FoX1avKrR3KmbMnxm4gwvrMz9JbR2xPnoqrdaDuKdIzznKei4j8T
P1A/qrD3HYYKo15hwlqvu3hrVRiTnv3hwPHlaWyLmIkbfqpsWe7eVSVQtBkvLFrYDX9wiH/DBHhb
NPz2pHBrZolsq6y2zEr3utK5QLtsApjjI3HeN9JXQ4w2l8KzfZOF77T3kT6COd5nYZaRgMauND+5
N0dW/4w6vVgvEXgmHctZiWohnd52jRkMTVZTSsRSHCV9Cin0q3fnmBmQxq571FkQ+mWU8ENTEeF5
dlnnlp7w9aSIEXzXyYKllHsJkX59zcDxE4jnyu+82aUWGAqZskj5r/9/ZEVD+kmeBrYleSHcnKFA
9nBTOHLJ79MHXkyHlntNWMKue0nVynbIj/Fh5fCeUKkpU32ZvpCnPS6zEb4gTabKgvjinkLjawCs
Tw0FSGLA6YounKuqt1/I0okG1Jjuz+WJkYgjq5R7bENx8EL8CIC0n5NWmphQitn7UJuRHIdwX/M+
quN3UW7ELxqQ18dveL6J7sw2Z+kQdB4ed+5uCMn0KQMwf0hpp5+zOIIlmzK2xTD1aj/OjtNuNkiw
KxMCg+SiI1C8B6k90l8Jq8y3Vfs2Yw8WSNbqqErGRQjYxZq2vuHrnvU/qh4rnnWvNHcMLTT5S7YQ
Wx0BG+ctcURh72te5CbbJAboTbL/az0c9c0OLrqZj01XAvob3iMRQBLfIGAVoHs24yacvSxfP61V
0I6uIfWgpruu9OHripc7zB0+60Ff5rG+LysKDMkYPMYYGr6QUAH8ia9+JVWF+QczkuN/oOFUwk8t
5SvGBA89UqXnr6zEgs/KUbuq3bmxvXFjGu0bq62fWpdyWxXjACRcpAS9WU4WBzwW4ob9hX0Zo99l
spd5TDLNWADn2+VjVKtgYQAvFcP2PBv9izZAld/hkSlSeXAB03cuyehcZJeGZ0ZQVAks5J1sy3Wv
c9UJDXTwsak69YylMSuE099TSPmOAnlqpSzbYNyTWINkx4+YRw0lJc6+L4OexVLFo2UBSEiKkrXI
MF13DLmJQriYFaOp/Tw1nNaUQSphiCmQYF1ZKBaqcAAY6Xa0FSyOdFsQHdlEUhqv8WAuiPg7lhZX
IR6hV9tX2d2yFHKB6bAG+6mhzpEJ5Jj3W/07hX80d1oQ2yPI8+5Vy0YkQvIXkTRBjOeQycEygzVK
N9kAwUVEUcewIbFUTwtIS8M4M++lCaJodZiHVUIZKh+1rfcsS8z9LUiDamrOdRKx4nwTGhOv8gKc
FwllFeNxs15ZHiV9zBJd6lvzEWnoZQixchv1GPUCwerTSaolqrvMPsFmMXrRHpa/RCaO/4uOTPVj
YXqGwD24f4GgSFv2hjz3etY9Grvd0LoI1Kp06ObN4ffuKcjHNZDmJWrshmcEE29KN7g1hELcOA47
hDQC4J7XMj7vusfpDYZ84mqLZrB9R7cke+VMKlolDvipsCIo8Z2p8n10kD9znr9yBmeuCMidRQ5J
4YTyybvIIt627Mg6IEYFsukICsstp4hnJKcqnga6477dTdXAkqAlucw1fZHbbhOCCrCyFKsevl2r
IDTbnXcMHrUxFF4URHTNhsA+X5z4SjPSHd+qTshko+kat22rAGPb1au3WvyAJQQw6kAXxpLIghdP
f5pZU4dZNducu3Udyes2lQbfMN7kWstTaossxoBOcyVB3g4brIA+/UMnJcbQEdu91Hj/u4ShJBXk
akOVmfi4yYpxDioM/8j++cpOAPpFXUc4SgZr4uvYNe5NCQ0zZeqF2Wy1sN3L/WUJEuMQxtcSMAfw
qA3CA+KsfgIHipXUPlHmtwKpAquwp9wKbD99bUdAG49bh1XvyVxvrlu0ns4SezLvlzPv5KGo3A8Z
FLlWmtkNqMTjeo4Mcxjo6xeqjdDQLA0Sz/oAMdqQjFX2kDBkxreSdZiTbvQXHLZ6e8nT79DRx47i
LpXWh0X4nGafNMDZa7EGFPerO+ouyT7FgI8L6VTOw02+PpGMH1fDImXjbTq2D5dWyc7n/uTA7V9Y
JqBGZ5nUo6JoRMhLf3q2yOz58sdX+4xDSrnaWgvzQ99Ukg7S7zGW4UsGdL6Q2l2tuz6u79cU1Gn0
TFGudf6k7B+ZT5H8eBDwqAgAsael1pn2u+bcEPOmGGEqSiFeWgbjbpzx67Dpa7LrzzK+WIVsgTx8
BRyG9TxpbB3AcQ9e7/MhB6W8vbvvPC3UAeJv5rspuVtL1xr+7wfz+RZ8N+hBlY2hItq1uWSSRp3p
s5DDszNL5Fb8vP6jH1lYowGyTlCfjXU0uwxw9RdYk4z3SHUDdKmAFCAgs3e/zRmv+FHp6l/1Kt7j
wE1HkHPYGcj63gdPEjI2VoFqisdGP+QWgA82Dy6eG2RaW43SgLiKIuSuYL/BURCBbnozfi8MRdZB
pngJL8Gsd8g/zl+QBYqJ6GujoqLZikhv9m3sL8btZrpEy+3aWAyRgEOD4lXBwlE/U0rFZGJnfRKu
GAD/Vn3cX1A/bESU9WLcrVfHFSSBddudSQovZz//2A39Bfn6RDjCf6gVPOGws+wlHCtF685ABJ8M
e87x0wn9NkUJfsTJC/7IVkKKa3q1FwhJS67tcKc+Fd5ySn3KGLBaA+QEc/5pQOQjV1NxVTLdVcdZ
DIpKnM+a9oUIlA8EhpQ2IMBDQXu39x0p1PoQM199GtVFNKl7sVxJojpQybheC2JNTv81mRA3NsIw
DyQSVZp675hmnZYxgZVXNrkq3FRIUehWaJUFeJZ6OpG3OuMe23lkYwVhNpZbiXPP5gJtc5Dk68Bx
GlBWpuRNEjNS2/XUGabmEq6i88kyUy+2xZ9dE3SBMp6twGgkhVqi3jRXjeX+30U2ZvIHIFJ4A2D2
WNexJ+Xb5kyoTALo47TmtsBlz0FeNUOACK+RR1/v8U2qempIejy9vR+aMMkLKfZgbBCAFVxM5qjt
qtKG673tutywiVPr9c7rZMbtAvHxIQYLpQTmLSR6r+rQcwi6JDG55eIV+yZGwUkaGVrm7eKFcTJc
TnoEHbxT7KvPTTzVZ4tmz+Y2XTy0ZceNYlSrpiZHGU3tZzVXPEVDoemQPsBqvwMIqn4lme7ez9da
O2t34dfgnOfiLuecrxkssNAPkdVyWawr08l9O98kL745ih46cnEMnYu+ev30iFnbV3JgzH3gDFGd
xJadTYQ0O+ra1qAs19VkTIlYCHW72Pv4gpKzsNE7acBFhyFt3i+Td4d3q/N8ssYC+ptXlg3PREE5
4Y1VETilY3I1Be2iHfKOISu/cYM8GPfCPBfq3veH72mPY0s7NGaf+Igd/3xD2OD5oSzyA1XRs03q
zqKBMXaAv0NGlT6/sw7NvbUChkNj7ygBbnGGX9lXklzLn8SuxnUUFPrHfcnpVU3p6NES3Fu+JcBW
P2q3HI1qvw5KVCzO9AFGeEzi2l1vUVXoHDZaxiSJb+AbMjMh4lms+2PvoA7aqJBC+0yOkC2y+ZC5
IccIKKlI16U89cWSn2m9JiKPYsBqy1g1M3pbT1OYbmT10dmMop+Qof0neeo3lBMH8Iv3aNIeL5U8
SAUmC8AtHz/hFbUs3EnLRmW8DjCqLZTw1ZaQUsDTAfivGVLhIsf1etBtMFsWtnWnSA92yhNcMe94
BAJqz7exdov6WY51rfKdxdaVK9OyYil7rbQL6FL0bJvtn1uYN5WEoMK/+IYnlrHZKvKmKWHPxu8H
ZrhTR5kCtW+ar/MmBXK8g4uMEJi4MO0sFmxkT+R1J0X/5h6L7U5gQH0xmUQcZy+g38RQwhxd0Ocr
Np0EkbPgNoZ+qQPTs19kzHyS6p35xaP6BkdUSzAqxs4voyn3b1BrGJ/mDnwwAlRsaX9nX76WI1yA
Vt78hUC11WY8O8dDviW6TtCpM1kbFXCDU+VAZHS0xp/nPfn9O5q/BLKrTPfiPT6lBU4GQkJqaghx
NPELQw11lyOIIOn5k4Y885rTprfFCbKQXirtbmd85kWFfhRjtCNV900bNHJ8vQ8ef6JBlweQ1B+M
vg5pwqQTEewmrp+LZ4sHEqfkHT2Ce1JsEsIz9Ilhy6BlZGEFM4/vwgHxheqrbup9BEfs4p1mvCGA
AVS272E9YxU4Df1tXaoDmzsUM/3pWlDENVGwPug3UlEcG/uaRrTNiKv0C80RccYZMwApVj79M+Qo
VPNcOZVkwyUOQrFe/v0TnGDfvPOmDyKY6vd5EeGEkpvnJIDw+raK3EaaaYXJg3wAYMHk+4JzX60r
hLnXB2I9NU61ktikQg3GqHQ+V8N6OptHAQtDjE77GKxx/iXDxn+INYDYKpldH/BNobpQm6Zx28E7
phD3Ee1zJVt+JjigaI+sTyIpURRPv48NzIqGCTRfdlgPGqTQGDX5jOYEZh8U3h17c1aw+NNi+i23
YO4VvFrs7pWRsRiUoRXP7aaR/+oyBvSytR1TK0LOR1S983ACYf3Gm5Ig4Up+D6SqTfzM8mX9f2JW
fSwhCYtJCefDXHusfMEraKcnn3OSxvHn3ivsoNfQDWBGPwzyR1PZKYl0o+eqLiaXsRn1ZJ+ysZFB
CXiVBm0d9dSVJ8t94UPnsEIcX47HkoWC/+16sbRLV9SCJKH3OpoFesMo3i5yH8J2pymJwNw8bHOM
BCPob+op7gJW7aLzMyKizVDd6ZXz7MyP1Uxh3NIwAKnDGMSadYYmjDpJ8TXYtdiGs1aitOtXeWsl
+lo1NcCeJYk0wH0YSaY0Y68NSbOJHlfr+lHtFJUxA/Bk2JQ/PxMqBxqsnhyV3QxIiy/irGT6xAMX
RBEim+PXHCBvTCHMTJm0JM5k5b7vSzyVY6LqVuQgScu/+HoXVBL5xdqCeFDFS1nl8iGE3avv4Zhz
iqh4kfW6nBEnEAVVYwASUbaLqGPMfFafyrDuKvPwWDJENLQYbkMalaHYqFj4njUYB149TGBEdQ7s
KJ5gQEpPdgldoSxM8tQZY1UwlRGPsoqh6S/ky7zhCWY3NrmfukJxs44LyU1eN1M6Eabz80o8Djs4
fU8dscgZ2jcN2NpngFOyS5vDzK3Mn1tlFRZVpf9VGDHEPaI3QEzdO5blQdWCTS/NVN8EDZ84xvjQ
AfJDpUjOpBQB0hMj7QrTSUSwpkFZ9wvUjNUmxhGyGwvCb/ZD9JwI96UEwhptfDIKBQMSXrc0fpWN
jAU7asTVcuYcW8kqY43aM6g+ALMDPG25maK2uS0h+LQh5X+3aI+PhePP9edYD5OmoUdHhBDNwtae
HTq2VY5dgccOnFeDkMOP5kd/vhYiDQiacxPjqW3qnsuh0gNk1oW8G1WqA0Vn+gDDGIgUE2gg1zat
w/GKJubsl64Oynx/pWgDp1mfq5LcDSwSyWw9F9y+kmeQ6BY2eYNY+BqSF36jf9shHHffeobC7NEN
GBKTecyrb0A+nwdqqA87L+2n3rXKcl7sjd7jtNZN7xmtUTJQKxhvHDDH3NsWyt1hYMeNBkBd6slC
x78IKhtUfhCH1KJevEFjR8/gS1wNLbuJHDoGAqv3RDapDy/RGbkkFawoIYfiwR654wIy66vNNic7
ASyFjNOyNQv8bLp5The9caRJdKDYpOzrS+UWeNf7TQjxXEYgV4zXro/rQ9R/o0ThMydiYr2wncgM
p3DvRtXY0TRE5zhjc07Lc49xrT0JsKG2f6qp3HyA+wCG/O6OlriGZhqSSQXVpxwFvWlitzxSq4CX
lOprcuI4xLH5Cqd/qcw8ysiRqOwWgaWvNOqr9VHItAYJeiuR1Z1xL907if6vc5PVC33JZGrRduQ8
ZEdk9wu8wh0rVxcG62SFZQqzsqyB/zNPugSmRsJrVuwkt180n8bSGTFd9uizREPwpR4qZZYKxJnp
e9CRSePbt7UBSHioXKNtez5YL4nnbySsb9vB26WwxYfAGqha/WEH5Un/LBlEQuBeMhb+pip5sP6n
TMwKZiKZ5ATZic5zvwnlgJqOo4aqr1Wnk73NubwcFrZiaZ48V8vbQM1/qCAXKuN/EnC30ceoE8J2
Cn0Wlygz++NDjOU4pBFz+5oZw+sJ4tBp93nmHFoKDD+tidQYxSklJtBDcpvUtn2H/5qSy2F3RB2A
NPsy8adE1lmkw4zWlSd4C1ZwcsRUFR6d2H6QR4jEGNtOS3xZTCPZnqPO7aRwUJA3DycSvfq9WMMx
wz73bMHzRqOWynYcIcwvE5l364xqwkusScS7uOZuoQZaH2ajRA5M6lX1Zk46MyzmBCqTI/2uxVq3
gs2Zf/zWTCYINefiodZBAzmtkdpn6wat/SA1w2d9g4msDV8obxJc/YUdeR0Vx0ZznW0VJxxVtbVm
9EruoMq3J6KPmJggIBKCQruohbOjmVT5AONnaojRfYZS45kwfuPSa9BnQ8irOfEsOMraF98jAdFS
ZHqMdrH8cJ699iZEb25eVjDfBRuoyDF7VFw7bpABAPthEA+Ws69tuKUWbr82hVKCmiptr5K0mWgS
XlgJMCWGFN9339AxIQGmc9szAYUCeQc4ra/7o/Mbc6qFpB74LLsSKmnQtFcMFM71CVmsEVJuxC0M
/vvJ7SrJZrsxGJxixy7ToqAajTPd1UCS9Lh8oIUS6Qmj4QWukL1HrB42tsaRI1faxNa9RrNaO6fQ
ZNzoFkPyaUh9XLOCW8joqv8S5yqm7uDNF2M0wZkBZZ/FYbwKQR6eUsLk8MyP+bWqWbyfTe4sKKiN
uC2TySIYaK1vTVWxS/oFjvZ9KLsXqbVS5ToofCVfNrD0LLlZ06YgvIFs341stqN5zkDR9ewKVdms
EG2gYK3VfIuY8bIJkRlE2qddnDBUz4HeF4yMg2Achfp1erPv4sxd3R6Bn10ASFnG4C7+LTB5VJWi
GC57IbhPu0hTTCPZrdhOExKuRtmnhSYerVJOUSvP7qviZ04w91cG+XHDhWM214KJbRR2VnTpCr18
AT0VPJmuoX7aNct4Q5LacrLA1rScMdK7xkvr2UjFojoFo4ZcAr4bIU15bCKoLGvh267H1m5rwEc1
aAwqZHVWoCdg0B+oCxgH1+z8MBtVCiLPvv2c11J1nFmwVD85LfSlzMqGnbwdK470yLnwquJXnQl8
v/4yAPoVc0VUHgINt8wxEl1G12kkI3zKRWAWyyHyVRfEPeGJC2QmPbLFwPrFK9hkvLTCPLhYeZl1
OcgV2gZZL9jEeM5wQXPCb3FTfJmjjP3K4KsEJTXX7WgKYSisDTJfyKdeMT+QtLvaG52XZsm6PjtE
Wtud/gb+ykeIOkDm+0XtGKujj2SUWB2Qaho8tGOO1McbaKC4wYmDEu7tZVl3zkxXFsRM/LajQcdJ
+KGZ4O2ZHyDL7QXz3ufbgEH1uprJo4iIWUPnEdJ0K6IHBmZpXXT7FDAFKHGQZQ6nlB716tU/i7y9
+ABbt25hDZStRZJiT9i5ABmZIW9RVCKCrIYJP8TtJkbwN/NND+eHMXgTn0gA1b2sWQJbYM7/Bb6Q
uhdd+X1rG1jdHCO1ftYPvG9VUd16XZt0t1Syli5Iud7eO9RQZI/Z3GH8whJj6juKDyz74D0gPdjt
OGMdYgfXjSrzlxge/NdgH7soUaWm4CC3zSqbDUdhAZjThiiQfR7gACsFR3ubt6sjlLYKo4R2jRYB
xwOTRjWH6CwUNtkwJgXduDChtn3H4/KPNvJe1h7uwTUP1PhT3FpSYkE4vQgppLD1j01ME2S3ijv0
fHCom4DAzCRRJXsrLqMysX+/LQiZx6q6aJrb6LU9Q+0QEhR56ukVAB6H/DeEE1JmvSB5brLDdB8r
E6ZtF34LSsN3b6FljjINIk+geVZgxkYcagRM/w/Ogoi4byMzJo2NuOsOsRp402+qwRHKSO6XZhHU
4Klvq66oxFLW9dCRoCptOwce4htWrzxmZCCF3sWAtxw9SloQX/h9C5qZjxqv6jNlFVGa7x/DvzeQ
Zs+V2smbBQg/OB138teFT3iwV/SSFGLrEjX9DuXe+XMZ7DBf8A4cPKFhYa5A2bwx88+tQlE85Cut
W+Ivsi17Qq2G9HX3lJp1EjS82Pr8V4GmGBP8Jne2QNZs7n0mIw8gXRkJgP6KE3R22BIZylrMag7y
4dI52Bmh8PzVWLYdPxZY4JhhWsjIkDMC9qoYOGtBCYsjzXOoOuDBGkX33TwSgBOzZmbj1gQLSA/b
JssYM9tpaWDUvU92JRe3Stw37CBTCFdgq97wqz3pcuUGRTO9kIlsQ/DdGdoNsCphD+RYHtPGPPcW
jh5QHUIUQq/YDiKO+moNLxs2Wu6jsN8XF3MrohPJg4tXPRS+Y9stJRic6k2nnivy3R3ipwnrglS0
26QDUR0B2+Ly4OwjRn9q1FIng5cH7dDWdMpcVzibRaXA0MX1NEAH3XIdby9/Rxx37OsVKs160hVJ
Usia29OQ7p5DunmXDA/L7f6fliqly8ihaG/0mkbTbEhNG+WgbbvL2Rx2nWiqf64+QRNRTskZJ8IY
ZAlNIkokX5+esn/9320KFAMSjpsPYWRhkbdpSJ8RSeZ33ZbJ1x/f8lXkFiLJu8Cf4JwaJLQWjy5h
wwo2muESqQ1Aig4brlEsW8ErwozAyJ4Xp8HxaT7CjPUeOnJNGJ+KPL1+vHi1Q5YoCQv5rj1pZ5SD
H6TSByATmhJovmwCrWl09LS78CydTNbZW4K+es0apKjcqyW8HZDQH1GVzkWnFP5jlbIXxVKa5Y2g
w2fA3aIM08VCNI9NRtqO6E37a0M8cBw9PfiFOk+QAhxlVdN178QhGyUX/c1+H03S5mlY00vKtBd6
DjIoPrMBmiv0g+3MH8iwdKP2saLXxiRfRutHf81qkYGzkERjIdl0mc2gy8GlRuwE0WNhsANFiRE4
+xTNdfIa4uhnc2GV3zH0P5VTUeZ+90TRKFuhsm34FmCu++ru7sFLoKbsG23GH7UJMZssSrJBm9vj
yAVt66OMdqTxwkNT+/3qbuxFVT5M049sR81WctP9/fUZbpWrrNTsUBZZSiCxjlqtqP05z136fM1O
8n8OiKv4xa0kdNQjWjIqSQWcZ5zmyN07vmREVEeUevOyBqvglY9avesMc1ztGgCQmexiftLckhKY
+ex/nAlWLRVjjub6Z0N09VKsy7wTC/h2hjKghS55qR6+E2YAbyggWZdZCzJU6szExaKRU1Bo9YBi
6PthzOeoJ8TfbCxtZY1VIWppKSa08HQX6i82nXMSgm+9CP2rM79SpYOHpUL83HjG6MGrvuDLj5sU
aVmwJlkqdAmBzjRShufvuEY03ppIGkrBLs254B6ktIJkoKM70uESK0AFiyvfOWctOuX6qg4NXeng
Z+u0nJs6b0rPmrVOjkEVeoAQz6dnHBpaaJzhTD6Eecc7u1/Pxgzw12zRGjfEinZ61nXl/wySgBbQ
5hnjq9nBLpnWpVmCy5ogzTKFJqqGCi9XUoGoDS1yX+yYkq64FoorheFYi0zH/sRH8o7uJRMSWHCm
pH5Gl7aOo1YY4nRqwhIMhZ9bSSD6bQCV0mVrGumsc18qXSjzaDBEuwMFuGVRiLAms/BlMVt9kWm5
rhhF+wzMjlrpXdDfHWbp/nehfEaFxp1Z4entyCwORc84c2oGHZ42RffW4QN9iZ5B1jEZRfOtqGpU
NPt4AMYysk4M7W9dZGFjNPuon9OO8RDS5ZRc38/C/rfHun2ddVBaWZ5rme7RalTS2MF9vUYS+wFv
j8in9KjrNS+oSinKMK8MpcohOumdTFi2YLVvnXMKHw+t4ldFMwFOZg4cWQ/egSEpZo3SagrD2orV
QhLsKqM8tHNge1Nv3Fg1HktM0FGB2pSIbmMru804bKnnGY2mrS+etTSha4Z/70PkOrrG0WT61GOx
XejeVVraSyVbVmjxVLSmYqaVFA+5JoQbkCordhqidThyN4E165uZEqdKN2e1Bj19GMDX5Y9opOkb
syb4zV8HKsomM+p4wiPm8NB3GXVqTqg6rMRTl8p/Er5eylnPwR5KR8QtwZ1uNDtTGwk+Y/JhsI0b
VT0+IC8LeRj7KLmLa3LLMIgxM+cmF4/tztWohzULT55hODZV6Nja7/vOnPF0t2Z0wvm5F6S/990k
6Bm0FC4x3v6XgTXPqwuSYV8Kdhb+1CgVgNlNKpt/4X8NjwIXNzINrCrwPqN6+SVduqCaYSK9OiKn
m8v7zcXh5bb1B/o74EvPD/1wfESuFmOfqy4IetfClm+/VcQLKQVUTwd3HdRvoCBR92t24q+VbJQF
A8gOm9oSqEWgYTtqXSnamkNqrBlxEJdH4r4Y77zANdLLRKeRvjK+B+8zf0tRAO3rNp5s0CzdkYMS
OAeCQqAH+5y7Gie28gme924REhxqlRanGoOAb4xf4aPkFI+hHODs5BwwI1HQfzrhonELrsZBz+e6
f+B1wTplQqB+NkrwZiNmd+L7jGoTHewplSTTW4hI9BKNoWuQ5dd1whIoJQ5MG+veEckTs8n30M91
hohQwyNjC1UFe0ec4hCbbGSD6HkwwiodrRJ1tYr0DKdhBetJa7zB10uOFjEdAqu2DfVlQRAHNrOd
UtWbXeMxnWVx3SFQpvsHqn6+LNwzt9GBUnUk8YZ82Q8NwFE+UQ2rjI4noNpje8Zukd3JPpjWnmAv
mw4sBO/AAd5VMlaZ823WVmjg1gxwtI8aOa7ZuHiXsMHRGj9IwIFZ63eBQxgxaMJzj+k9aFA6WA/s
X1U6fuRK6kTt+Dd7UF7jTZcZoUgKM1t9XHrx+Lp10Vp/rwdLIx5t3w5fY33vH4gtys9nNOA9SqD5
wQimRGi9Mzev1tm/VpW9SzAoqpYmxc5KDrY9wqPFVt1osfyITbKZzQxCDNPMIx+gnilRJYyeHYx0
rNq1xcQHd3pbCflP6v/Vetkvs/gCucMP4tXjiyylnmfOvJmMrcmDhF3OFkGGWZ7qYl3f8SeakrU4
NsJ6fAcitc8Y1jI+fhSyfl+AKq5yYOGZSGEW4DL1pBgyL7RxLiySCZkiTSILk778wrQfWSpb41vV
WY6bv12FNibyJiG31ftDP5noaKfeeiTxQolgIstWH1XD3Zaxau3YJ3lRM1cwEeXyowR8wp/Fm+Iw
oNS1Tk2ZUzNfJdNtePOK8YLKrJNqUum9MhWbZIlnctw1D1C+dNGwIyGunbBngQ3B6dKddO3Jh5A4
aGkpwghNGHMGETj9I+ZIviZ1JSYBmU/P7pA79cW3BethNtXOORldt+s+p1x+qrT3SxoA3OkpbKW/
c/FR6joH9tPLcNPPbUizrWS+lMyhxXTwk/3+u/HMW/2oIDf52y+6/M6ksvI9lmS4hp3246E001Vf
zmxX0Lx0tTe2LJXZ4+RbGjQJwKfdXHa+wLCq64H9g+yVHb7ZZ3FVdxt7wjeAeSmLCb4tNj0JgMlt
Hd08yED1x1FCLq97guC7os04IBzgR9yWeQjT70hKTUjdhBhfWlKXA3o/OoqNfiq1JWlf2xImhYhc
CbKgi4odulhHM5OWeGRZz/mDSYGgL5wncUoJuP+u3Cc18MMAIgLbeBUu3/aKg1O6vpTVmj0RHOhm
dtAotLOeJZTEVkCOXjhmLiEnhZJ46Atwz3Qk95vul8DjfWB1RNygxKzASXtt99tOGVkecmqLWQS8
HDyFW2F+MsC6IwoqLQghFfYeTo4PyG7guzqdJYgIvEr6xBLS72tVSDHQL7IG2KNOSdjtBnpSAIry
8V5sOoSpbwwI7sHdiS5K98vGfgwAmK0V+56iZoxhOuOMz3YbHCFm0qOwfCCFsB/spCNO2O0LAAEX
/QzB4AmsvT28jTGCUKoCX6ZsPESraAEFuZWF3rDTbDqkRDkKV5EldF/VVTTeAHSzFnyDjMoop9df
rBuPLz53UmZeuoSNcDwCrfTCDQxxl4ckV2jFGdU4GI4+esm1abtkFrIU5A7rjKfEbDOHMEvBb5pm
pfvm2SFJ3q/BUM7G7+ZQVp51w0nKU5xxwJN2MLcgZljqxaR4YH7YiNpVcct1eXZcfAyiZbTbrvzx
LHcQC038+T4wTMsTHSgkdFuWWP373HB80S0/bFK/NTPPmbYo6/LaymSc91rkQup5+njZihX63VgN
rlav+tyeRCvwXYSiNoiUVgPqZ8uw05z0M3GznMcmrQ4+RKDXA5tYPIaHRmfZzIBqKYng4Cnp3zHL
hfL1gl4eDF8hZ+cmjhCSCrHjOd6MCEprUa/4BSrYfsl0Blj8MKiiPzzIUXPVsitikbuPS/NBQRWA
va64oYRedabQqe/U1+3hst3UEw/cX7WFqpcCMJQ0xPq8c3JT8dtzsa/fLR2daQs1LIVGPh3RX8oZ
VRQ9OqFobTbSMMbrDkWopgz0p9vIYfxN+zjjHBDL3rQCHyRTXGb2nblwZAHdCCQVd5/2DOPN8WcF
go+S/8/+PLPt9VI0Nl6ncHH8iaNAfUXUZ/w1xpoAXkKwAL0AHDhUHw33hFpciKdQoz7nuffZtmqn
qMrpKpbz5zc4TyJAdwfwmolIKtqqsgy1oonUkHH8/mPvuL+ADtZRtycE13BMqSRiT1BjjzviOPo3
I0iIpkjuY0OaJXwO0BOcuLBN6pBj/utX07kJCwoDViDPtyD29qUXfyh2QSKZqHKL+V8y0a2Q8Yc5
spNjN9ct0mBj/vaUuHO34mvQ293scaz0IcbwcTntgE27RQH68OfzizO2JBCC9l2eDSV+wHtmegKA
fzZJZXgmwzDmfQ23iU/3vKedblbHj+3Y+nq1Aff140Cxp+PQC6g5ekeMG5KZFtZeae1ctSlx/Elw
/5dEAb+Wtbc3Ds6M8D6HumFCnbeOpQMZlidbvVmqx/3NgIEkt79Izo1x5fSiJReLmmpQ3T02ZoOy
C0mSEkkzVZPqLJpKclXGG3szagXMZWlsTNx2t9iSK+35aD2QHZJtSKJzjvS66DHm1L/XqnZEBZNz
4n+gBiVXxF8ZzcIz8suiZ4FYiABQxw6BAI7Xz2DnE6tfTWNcSYj2UlqFD2ZuFNpQSfNYflBQDIQr
tuvAwXCwJwgZ4UJjI8IvS4Usci7FuBgN/iNvOw9idanNZUWw7BNTtASEygMB7sHwZ9NksPB5EbAu
zMOKfWVwz/vyhWoYHxaIqXeV6GNKLPNlI0Ae8ktL+y1uhob7r4+5lH+f/fNWA3fKUvQbPcynA7E0
CIWZjVBJaggKiRAWemKI6XNbMhrxbXoLdN3tvjCsgyrdlpmBGNyu8uUP7svn/Ahq8MS5G9wcrXFD
Bk39iuSQma1qFyh8TrA5J6Jy5yD80eA/1p6l2nuQ4NhxJfog/NMuQVKn959jpJHIZIEC5fzxjcfn
aomFzWtCKTiDrOzg7+FKAQi+VYwStExUK4ld0TZA3gs4+K3VIL9rHJQeUN4pl3u0773YAMMDSCk8
y9iHFdZQj4MBLhQSPgKRMMAcyVUweN9ElI8dT5f6qEvuTF+eNvJk5I+rk9rL7a81Z8AqKVrv+f9L
pfdi66ujQ5Zl8f4gDzeZ3HnHG+Bc0k1ba72S0zk2nLQy/DAlAkjdoOJfwbcV5KJAC5zwxWuJZfmj
52GHKjRtKbZl6Rvj388AM8QCMgUNusn+TX9kIQixlmTobIcJ02IRz53UWU2vT4AnkYVq+9/cTZLi
EaVjvk/j1QocC2qYnoHMELmlzsr93pRbazX2qoeTDM6kUn8mdM/3nrMrNePp/yNAUQtTxCXgir4h
H6zTknt3oyrm1DSUj1iguSL86mEMOdsY1NUSMMNtEeX90qr/6nbpZSMEdPGvH4p016mlju/IMfP9
KUtGddxyV24eovj+MSLJTv/m0cGpmJQTgUJtXk1wASFUVLKmz6R0h3y2P9XSYNn21sGdbcgjHTto
4ef5vMgbzn65A0zg8J/hwnroj6rJIjithlnOOvW111abffut6A7YKCMPjHkH9vTrAb+uV7Juecii
bM5ic5mpCYltp62tRt+2C2p7fXf0fvp/fND4EDYUjMUlDRtQOfotC90Ma2Dgxokm9JlRvdGH6saw
Uu7wXbUnbZLspIlM9t8Xb7r+cuPIrvAskjwcSY3qGa68LTgxIhriD6adnF5S0pM9rab9FRnp6cxd
ooxFIDnOJd5Ex3rOGf9gCCqR9wME3xQ7xZb4pbga+pQBWBLXL1Z+5JTmaA6/UZIdzfk2n+skffty
C3KOAaM9GO4WR9lDya4Bx5zsQ9CCK26xWkAQw2sL1t+KP61323lWQ/C6VQQ1OCNS3fhuq224Cs4T
DLe7cqX7B7h85aJe1AhiBFdJ05Ri10Zpn10YS3Xf/2BU6a9iaN5GO9zcLIfiRnxg0c6HevFpFUxf
rCtXvb07nf6dAxEtlZXevI0TaBYAOjqIxwdhn73OQXzucjMxzF/VTOljFw6CfvnCPtez/eMIxiMh
p+IA6HF9dZQfBlNVBwfYL3XqCgFCKT+K6PpRHRafIzSPokPx1L4b0lhTA+t3QYZRGFu/Ql4Q88Fl
iVVpWGkcMhvVEXtVHMYHL8RK7b6vodGj2DYqWIdquf6KPEMedSeMCaB6lswnQMzhxuyp0y0CkFLY
/NHrzNSutWPO8cME55PlPpSUfbE3L4ZlhrbP+rA15vXTri1ZA0jIerOwKxuFt96bMyExurZLiamR
mUj4vHMyozfdHV/Xk0cMtH6fDhMos+ZT3G5g1OQp+hkBb1yKAbF7hgdpYDRoebOxptWbVq+L8Jw5
tWAHK3mrrvi6Yl91pXqOFpNSW3xwYmx7yTJGMoM1CSggQq504mgu+WoLe9ypvucu/rrO1jjTn9/i
9JYqxN4F3EUPVoEVtJFXfUV3grWKFwQu6WMhYOMYHbnHB3J1UEFkLiwq7746SxA3tBV2owGLxva+
dScLYeY+O674RFoSmzDCToVQBwyyJAbCYJj516K9nPrUVfyPZq1fPALd8K8+rg+z7LAzxLieUsx0
zyPCBUDLggCqb/nxk69ShzkA4qiBmAe9urgTqFNWka6rDqcQAw3oEl4YmTsfZ/EUT3BGdwDnCmbk
DHvdi1uGAgdgPFQ5kFWN1oxH8rOF5NQAAxLQHxJkR7Lo6fmGRZrPUOUaCCOzFEG6EPrZBCU+CgkN
K1rsFSZ52C+aW0z4H0SStu1ROVTLqZraD5L3SEZ7/4U2Mec1UqK0/DKrQAmCP/KpGYNNKnUQkeJi
yxmnR3QmuqmypEGMrLH9UqtfmJ9tB8deausXVeB7jAqkcMBcSUqxEmKHKt/KA/hRwIVlATZ4pbcV
8E/a7xPqsaoRcm1/HLTG+ZSpEG4I24tkvGtRFVhArdckCx2rwZubEHVOR/pIU0qbo9+NDLgxum2h
49eIfllnVKAwjOJuM1Ef1U/AOPSc3YU86lcpTyf0tDNAt/Gwbo0KN4OT8T/2GurFic/MydLSkeWj
9rAkCipRZ3eUT3pSrO/fSX94TyncSR9JlYBsGE6dQPYYvWsiENbaSUQN+t5yDVXe/A6ZEdf4Y+j2
VWlEsDtR8qwVb6CSiGo4Jc0BWVrC7I7xT7TBrtw/20M+6w1W5LECGZ8+2Jck01+0ODiGgotiOhAW
/3yepmgAl9dFiRofTB4zIbvstLxdyXxbIDxSWkBU+/jYbtcEJGU1dbbyEAc9+KnPZBDD39bbPZlR
QpwQQSoLI4jtC/Humk0dCv1rSHmYWlU8bn34mwTZ/TBbooJj2s0JU1Liqol2BQ1k+6NeE71xtW7w
nEoodrU5YSj03Ifyzgn2ucXG2/JSvYDWF0n6IhXdYn5QLbqmuW/SMXL2400KRC+HEeFnShAGWK0r
MCpW0PRBUxZpsNdDLl/iUZ7Ne0oD6wZX5G4+bkW/QyIlhzUwbqtWrzVpep4b5whQfcZZVED1Mfp0
JucY4uH6GcYr+4vkh22qhpwuTinUo+Y35qJEYckw7AL5qnt8RXj1Aiq0UDKLPc64PXG7qtzJo+ih
+2qKPfJ5ZaOKYSkC89d7YdBFWh5ZyBqUeh0Q+qTPHxKTGTuLf0Rs4JG60NQwEOFL7PQwSL5pUs/3
rx9+CVVSkSa4yvwZWb6kCMiblKo7gVyL4HprUNbRWxJ2OL6CXK8MTg6QKmnYhaJr2j/AH3ScIjLh
nx0BLw+2/yfVM29nU/fUYj5d9ESsoKl7Vy5SsyzCZhvgxpnXeeQS4di3tCk+QlX9kKVq0lhcLKg0
PuK6YZYhMbtJbwn9emDUXWjU3CoVbbVYenJ15lN14JbDSoZe64jIG6QRv/yHw+enb+XTQFM+RlTu
SSsOc909ukJhL9JUWOdKB6zBXnrUm+kVPr8vZdka52cHsluj7BQsF0SL1byjYbs09d8qu7yhproI
G6QysemX/U0NbSgEoCpZp9TQG7hRmMg+JoHzEIR/dftfmvBQGRWqvNX/TrcPneXPOO0P99v2SWei
0nDaXV2AtU+wrqleWKW+i0g8FjLfxOnU0IdBTGhFk1XKr1XQnfbxMFz/NcJhVMZY4EKq3zI43pzy
tnZm+wlgo8FIuF131MKoXLkZ0C8I5rwEOYoGgqE0IIxFjRaF29IgMn6iCQAUt3allieLuk4eGyh4
Q44NhVXP7ySkF7na3ypTnv2rfNOgjaqAAJIB/0vcVnfKGLUjbm49emGSOeWxh83oCpvzrUuu7Puj
TaRMqhRCFilXoRXvTDGXST0UG/KBUxHSyU0KqXPfSZOVNQpO0spDvmxmHo/z3esFhxHuFQ3+necQ
IxhVcVvnjkpk2vyHwtv1cihp7l1qTbwLIboZe7bhwD4Qv7K4YhzbqfhLKLXwz4vwOEcZPufptTq8
CkW9O1Cf+cGnSuW0AqatJVGfuHxFLH2RwjsNtz2aLl/H865XfOJBwVY4Wg+l11zVTNmPg3DISm5O
5u9mEh721uCCLz2TJ6sb3Eyab3OL51eMkuEYl15czWolq9KrAUbj+3GdR4vY27l5JhQ3kvZJkM8g
51fliJ57twwCuxUfdjvqJj0oXFcbkMKalw00Y0BJ38yvTiWUwk9Wr+olOGXdN6/v0ExwgHKgQF3z
xM3kq72UIKMWkjYE2DzCoOGqWCyGZrNji5vz25o+NOhGdViH21xzI/EMHo/8cY2y+4n+LY3NQ+EP
t5PAYmbmM4AIhHAAIo2M+XxMhmaYIhdnokb6+nXrhVH/kA9g543OgFOjPBOYlhbXM+pmMeGJQh4v
PSWSZ8HFPUgDebQfhWm1R88pJCoxXapjACLNomby2v4qRyql6BkcetIGbTNQdArlmr9wMScAYd3B
Xo5fmTLWJ1V9RWqmsPWlivw4p5pdR9QsDJ9AyVJH//iqKqH8472rPNm9Hr+Ts2I9Fb7/8Bg63dBg
gZS/N2RtSIVhez7W18ftkedCNDbHhr0A0S+U+85fpfK+b+wW4uj1PK84y8HQsdPBD1sRp4H29/e5
tocSBOKsQdvNMu+NeVftw5MKBx9/ZnO+x/Tz9xogZfhx7s+1NGlZu4aWwPLGGzNv19kPGx3JL/69
4jpMKFVY/BJpxBwXmkRkk/Y9OfsWSgNQGAFzmsixlE7eQNATJmwJGUnGSPAoNRcaFlTlEelrjk5f
zG1bQri9kExXmwKGBMqOj61dDFbsdOtgXb7ZdsHE9e5uSuct94WQz4I908LEs24ON6F3DW7f1k1i
KYQCLBp4WXMsmRBpohYf/EVY6BpbvJ8vcU6ZM/TN7vrnOg2xN1+nPShZ6DkvQ57mfGadRTh8pdr3
XInYi40TY4w9kB82J4VAv5p29hPrwzbmvMfaZCZ1JtpBzuwM+5h9yDdg4/eO8HarhILLI4qyBdGy
iwMFM2MuL3pmK7JwLfGRHfXd49I0TSnMaAA3Qzsr94g5U2f6Up8ZcmTGPvzPdWqyAet62UVSfbWm
g5lQfzwCXFUWXGn8ZiP+uBfI6SWdwK+ENhDEs/4W8YG+2dgUfpNAdSsRUtVQrKYM8QiS82LZW8tn
8sm3l5tKZ2/xrJNicy5C5JCykG6glY3oYgdSDgwCrsbPjlqyAnyf+ew26kthk54NqER1PJ/eQjG3
1/H0UOjvmrT6HNbfI7tXHClYPIdjNSKm17S7jdGc+rkx3uZz2fq4bGofMSS6cltrk0bVO3VrdAMe
tb5lC1/mgit0CSLWiDQnJjMDckSNQrNr/Cu7h4mnV1SMY5g8P3SghjF/Hg6fNT0YmxhXiRHF2GqH
zmEBB9HOkhdBGmQihxJXLVNFYNelIRzuOkt5kmg7LHkfdk+sI6+lxUYOHcD4VjWJylbx+HRvglzi
M1Npg0WldJmFE6ijuXv9n4PSQOpD34yukLli7bOVf0MHzxavvnvRpD/Mr9yts8RXglu+wW9ljRDQ
euttMBubrP/LMSKmlN/inrpgqaLlLISd/DhW05WgQow5WgJ8vSOG1DxJX+xgYZaZIrth6RX+HVQz
LUSSIfrhhNjltXV2iqZKcxTeRz8j45MYv9YKrMoAUzmL5jpbEleelMMC2qYkP5x3f+XuT0o3n2nI
vpSYlH2owh8sapE5SGa7OfWg+j+mTUhFu4TCGgi27eaHVwpX7x9GO9JF+YYgV9/UwQxwr89Ru9EN
ncXkH4k7/xUQ6UVikcBxowiVUMgNbhOw68CVt6HGwUc6N75hP9jICGstkA/SMe0wjqGaS34Jjbdx
uo95iLuRGkcaPedTzxiJZdseQkUbX2RJminHjLiaMcKa9meCT2p3rDDs8tyGr0MZmVTYwsHr2hwx
DktSPjVy4J9Z0zYHHmBDX7fXhJ5otX6CIREDQJu92CM4s39tQrndTt5LPFuchUkD82JoQl92gt8t
LkdnAh2cJt1SpOeKLUNC+MPMddsEtgQdHLOE7vASDtG0s255qu5TsgaViEFYX/lZWCJ0WOkyvDc/
4aFWjaB6+vZi9Myygav7bXaf3GgjIyac2Rk191owjPmCyY5upfInf8ePCwxeNvHtJYpjQEQA86pP
J1B4SL9xh6bVwq0g6wE80/VFkPPmXD13Ecan9y3VhYZg1v0l7DikEFY9FXdM8KCPXg1o+tjJy51O
qQl5RpimTsigBGzc4m9F6QGr+6GDrpWCX//Gre9bBTzQmGTZqOgquR/71Jiuv4eg+W0vFxZivQ2+
Ou8FY3O5We7AK7SY7lLC25aJdSlBtJLBAnbJgxhVQ4Ux1pGAHj+FMP1OXFollxHrxzfwua7ZhUBJ
hM1H7OGI/oiE0QuHGUqpNpC53+oM9c7N5oelzwfbqdOzNXXa7J+mcQ3X9ZN8QHychlVdnVfmO0O8
MbMd0ofc3AFbl6wqcREJhopzg/nsRQEXFN3ggJnJC8wanhMSqVGz5Lqyrc+ybO7X6jorW29aWHOQ
a+lPk0T0ChOvXBsUQzDNu+V+3tFBk5ZaGC4WF3YNRdHQXkUozzMJyo4diS4vmeBajzuEWfw1tB3q
kLBAssR0VP/RakL57aiB5IsvDvZO1no18+IizUXqHhsOpscqGxt0z8VUajf6LgWYfk4usiZ8foIK
eyAO+0/XCZ3zKof20zwzhRtNLIuOfvSdtGKt20heWSGuaOo3TNKVALCUMvUYl/NIaxx0zm4tp8Ok
GnLdDJaxix89Q4cGPqXxifrKRPxZQp7ih+X5zVUA46TeiuStAlix8r7K4D39F7TWUVZHSMlg2td+
G+E/H2ecGmjB95AK0G4gi9f4ArBnwNVGBiLurvy6tTUePYed9SbBxtutf9w3ULsYrlq6aK3cNYKF
7Hb9HvJO6LldyhM8dVh1KcczEF/5h65QdLz6K1WXGQpV0bIqMPnXz7/X1/E70jprfPLMOGoxmrVg
FdBwlCztU0r0YSY04zDkPcdLa0AOR6zQBDy5RbE5WFPGRuRe+7QDtzOiBsLOkLA26uTmNZcXCHzb
5wNgHcYcpCjrZTztsY6Q7TzuzfoFQtk+nwjWnNF2q8orjmUTvfFgQwjyjKpa0y0Q7kj6Y8wADeIz
wPCW5ca5o0QcyaVGBFUYVvu1XdB2/3hCoTHqP/r8TWrqKSoyUi5OrhmxcBrPYWNgPLgPPDf9kg/b
+CTwuqYlIcBJsYiwJyzGzVSfrtzb7YM5dBYfL60suZhRhXJsluXvwDzb2tLWZKlWJoRgltEJxbn0
zxp/WepNKyqKjd1NFa/ZeFDJCV7QAVCOHqAGPAukeUUjkm742JkslAKMNITDyZ0FRd7/O8RsC37Q
Cm9KRgWkKIMIPJEXdwpblSDHDubMFfZEk6q/UbOi06usauduDEPKSBeWrYqDo6HQuOApHIdwyGd/
pzwcZOg6ncxmhSfmfvwflK5GFpFkOg9obbRZZ27w8FJC9ItSNgzSSjPKfShJEqRZp7dN2A94borP
gmTrlmIjdvBLf4aQ5FGJxjPMofc4UVA48InKEMUlZi7KWuvCFpnRdfZ1VoPslDLPPBvUlD/UitmG
NK99YDk/o2hYBT6PlMju+VVdpZqM4ZE+3CXxcgo0q7PrFYVNmPu0zqbasY1uT0ynHJCsbm55WaA0
/AMyVFF+sghzkJ6WKPyPfQx0xSLu8vJRJD3U4lvYPin+uLzD1xohssxjWp42K1VN61ZUGoZ80XUw
ofkKr/f41KjvKVkeYan7qfcEWUjd/qJMvil1Lyqx5VzAGl4Sw6h+MFQNaj2FtYlaurHt5TX8Oi2q
jZdV5mUNt8CuDSYkoXkt/zVtyE6bfascVoRVMCzCiNW9Z/c3Ymxph6zmH1+0uuCcnpTtqhB0NSXC
GlKtMn+wiICJOttEVd5dbJpFn2toQp6yW+Yd8y3jJRP8cV7k2LfBjnVvJyLfMHIwO68+BUEgPTMp
YptgDBj/+Xrd5djPnjkLfWSI6HG85ERQdcxFTPYTPSfOmxvQoF9NBN457bvU+N4BfLgXKH7l47Hu
+rOHrzBS4FA6SYTmKV7TBOFaTLNYBS/OGngFnLwt2ZpsHj2o/ZjpL0Ya4+r+yNKeO8re0ZKG/Rk+
4iLsxvvj0yv5iH2kOMf0RPrDfy6wEIUppplAbuoSZhGTYjrDg808pWmTF+AdK8WRX3zMmRyixGgD
yFbiLNrMonf1oOMvREzrzedIMYkaDViU8S9WAzRO2hppzoCBncEcum4WH3rtbWHGqPSfghcPdzLA
KeKaejnK6dbFXIf3HTfKBlYfNte8iwC4PyL4xNmoqzU0rMxUXqXYXyTwzRV5ghAoU86ifqOL+EI3
DH8JEVKEf3OsO28hSaN8ELldLJIVqajCHYRunz5ab92046y27G6a74qnKPqZeqTAx0FAeoKXzunx
uGZfEg+jNAuUy8B3poEQOcCVZyPl4lJ/gZa6v89zAQSRawCFd5kdWPChJvEO7QCjo+DNPH3QXr8i
/w5ultJgJp8FAANJlcG26gYukxXmgw1x40/4L3eXAXyjLenIxR4dyC6kcXacTpeOTMdwotqTF+bQ
dqWcdY+x5DPr4nhDgFfe+XS1acQ7DTnOZGzbGkCr3BkGt7IeTgNYDxXNQcSMWCts+b83UWgUJBC4
GduZzO27FXGTy2CnSFnO30t19h6lgQOm6J8sY7hMq2hD1R2Loz5v0ROMFK49d0z8UsrcnzbPJ3W3
kJY3iOFS592e5Tp6ZBieH7dv34OQED71YBT2sDd6XaU1nyKwb/ZbObxpt6rO5lMPzxMDqFfMDKaR
dDj7pxRjhJC5nAn9JLgvQSALUTGRSAHjPspbRMuoyM+wQdEzGlfYu2/438gtvicT2+ZRdMZX9v38
ndrL74wfiBafRHRj4w0mOdU/DiWvCkyZpzXdfs15M5kDikBJ9ClMinToPGuAREJlcZM9nzSyznRU
ObjY795Ond3nnFIepWqNtuHgwgJiinGaoxWUdI7VVmPQ4VS6BixoiBYV8FCGzut79yp7m82m7a40
m7CUnw2/SUX3bggqKSOf1olHOLIiSdOQf/8HAgZRGVn21094p44VroQf9vjIgfiIli9MojbgwUMk
ihlePXKkLt5kWgGixqNzrDpxSTIa6BaXN7tCVhp3jF4kZMQpWWYJrpcOyU82B4vXh4qCLrS2Hrje
ta6nHlcz6+wnTMnnzp2+0D69x5AwF/a8S1B24o6ZkbHFzjVon77qNXv6Ju7tR9Wb25m308OEAoi8
S+EIrmTk2/zCZyM8OjlaatNWn/CesOyjE8cCac1LVZrtpsAB40YcCTeFn2K1NvBETEOoVffyUHT9
YjJW+Tb068qiWwZeyFJ6+97imBuqrqiYr3WL4lcxZO6mZV8LXYKFLRlD4N+6BPVaKCpVkVzc7g32
ZIHzgkufWrpjeakuZKkbGrmx4rm+yhuwkfjb8dtrJN0wHhXNew0+Giaxys8MzgnDQ5rn4s0WpKP8
xHWYje3ScVf+4XxZOYiTcnyEX8dOKVBTpnyu3liILmksZHwiG5vjqU5t8YKfDQuFYnTLlA1WSuY3
27WvBVIdNuJW6nGeD8D2EzPgKl4Ri8Ruiz3y6eiDKn0k2XfGJaoozjfeOAxw5JJllJa91/xqdVPu
ZaIRlsXS9E2bPQM2Mi+EBPjGge81CDDNaKnTtE8WwzWBa62xBRXSvPOWmH96geeIsy2KtCVfB7gY
vH1w58QYYfJsp2qY1PV8GWjdmsle3TowA1KdJzdA8+w8o8kBB19gWmXtVgEYTAOnayrf+OqzfLty
9EJyw+xF3dS2Pv0t663KP8RUGZSx1VlZP4WzU9G+VQxI8lQDrqR1s5hVyjbKHz+oU3nqNEMrAsdb
4uWf0pucybNb8s4ZcBIR7YhCC12u0l0fFPxvBSdsl3tNnXd6NP64DbDo3M5oZQNOENerwBMDQoUG
ftR0fyqMSeEnWJUBP6OKTkrXC2Qp1ohHJd9lYU3RSXorHZRqt/LexXx9BWZJl2TdOUCxgtwt3zk4
wDus6OVpjrAHWR1nI4r0aLtffThz5HJXTu6zjGHD0DsSC3TU4b8uXD4ky/Zl4izAmwUQPxMvqf9J
ngyycJ7nRPTyjOS0c5iYZyID9Ec2Wcl4mqI/g3/QjtTVK3Db8fgGU6dvNITBMFxoEMlhCU4EX/Mp
qD7e4YaE2E40/A8eJlwmsZP5H1cR4Bs0mYGwB31t76qAQ+o/TQejhe6bQ6+vTIh+OElvqPiIF9GO
lc4qKN4tKn/Z2VGGXiDq08+OjvjVbH9q1HWBpoXGnguFOMBa52nDIHFYomgJI7kvKolND9ONqk9K
tCWB0f107+cxt2dzKihMo4nNurauJyO88BQdq7Gpd2oFSHAkFJbU4+EK0z4fv/0xQgXxj657lohr
bxnHlD6eR5bj3Osou6I7WRNJ5cdfRsJ9mK1zZEkI/Dq71SYEPJ8NNNvqW9kmODaTZbqe0tplWOjK
aQ1g2Fdt/LjJBXT1ZqP50Piy3HfJPD/Cj55Ad3K2YL5M5wd7tbNomswZ3/jI208i/pES8QE1Sdu9
wd5koFu43nIOeJ2k48vWRDdtxq30XUv+QCHnCAttyJOBq3yr4dlXQm9N3zUENQ3wsanLtqswh331
HJM37h1ewiXSTlFwTJrB1QTNOpEJMMRcLBzq9DGPCylaqGX7JJrKVt4/ryYotrdxNR0VPRhsl9vf
dtMTq1xTDlCN8GeTMLv22Ld+dadYwcqcrB0XAOzUIAwbFPOpM7hh4bdO28gFnGkc0NBHcGJ2BNgH
whU3OfzwhE3ztuxNtobI8aAcxBsQ3vpzshnuex39QeZbnUWgosm39XEKIw0kmlknC5EoPVYUa3Sp
0b5d7fBFBNq9QG3stsKvhrgaTUu8mhLPxLemQ6o80xBGVGyQNLhjtHpSGgq/9ZAdMWfeskWRIqbT
F9R3Ohgmy+Mk0CipAaYL/6yXCYq8vFOiXq1HWAlxV3R7ofmTWjagYYCPVUbCwSk/7UoTUS4RD1ab
eyaKaO4RwRm73dR6YMtOpmrO4ZyUc85BKs6pl4z8H6uEuwtSbMfp+li6D1tk3AKTO7MUYPB8eRAH
Su9jXOC6zLqY2KB4DbhmrcIubtAQ/POj9XEzj2hzvbuZ1lDjX82FXgp/gHKspEctIF9n0SQhYIyU
+PNY+c2nVa9W9WcjKEuNlbH1g1akxV3stAM0ihwLuhys/WN085GewJoTGnXJhjdJAw9EaI7F6Sj5
zfE3ukDlNmeptsdITKmlCO5s21wlxxtkdyYjFu/yNADgjMONOb4s3c9pntQOhVyvXzA3/t3vbrO/
UTITHuzK5VhdLm2TN/qA380jKiv3sC4KgAo60tiGuHyd9gspzyvTgvS4UYxAN/+NfQ1uG310h9ET
K4ERgIa61BXCkAKgm9VHkbmVHaVQ+pUd2QYUOFAkdrAKDFBwqDjULcsdFlSBkGt10ETI9Q8ZUNAl
pZ4QHdBB1MYS+jOmuTAuYybytYJcOhahDuCMsHytYEaaxAmpGZQdq58SaLhhIAVTLVdkOnmHs1aO
cBSNTSKbz5/pDZpTahgcct3SVzv01BQMroG/phNzVR9IwDNfpLFAJUPEOCAC/VuLmGbmV8VzkY7m
1E+HBzc+xqOzQvmTmub03GuSm1pGMyyF/Z8n3LB4Rx0PzukuPmaH0VArrSgv+O/c1SeyxMr2Lla6
Rp2JNP/raCyg01zUbImLYB8fNMofvE90pfBymErhjwjkXJKP0uBDPsa3FNQeZiPEGAs+IABqURYf
FSUnJij8riJ19wKbYBm3/yZC5/ba4tG1KmT/jRAbAkNrCZM9AbcybYbbHJMEUEykbAEjxOI43C5t
7erVIsoTYP3iircN2fQbpBn+3m+KVb3LCaHS1LF93hJHqJ3/Uo2Ix9vt4rquuPgaumd6F0IC6BW7
KyZD8ez32GozsU0/ONRoL67XX+i5P7kVQXG3pLbK1jHZx8bdp52/YtW+2cPXBIlzohezEOnkdvxt
lofR97RGsZWvFlXOVGg4Cwhpu0PX/on/KXyUo6TcF/P8BTMGLB7a3D0jI22NmOifOvQslFsWvlWl
PADBh09Vwjy74229dgM8XHjEEZczeDEeMXG+e/8ftwISnIyBMxgigujxCZTIIhTAYOOPbtpL6Rri
we6F28R6Fs3n9tLwktrTZML/LOaXKFkUT7PD4/HNh3Z9MT+Wc3l2HpBYcn0GGsKQiKM43Qjo7ETT
0MSYX5t0YuwJNqXoQ97gfuFTdY+KN2r2ahNqst5bUxflatkQ/ElJoyhw9OkpOGURq8D8jAxo1lWZ
oinA6fbL1NrIV3G23sIeOJBNDTAPXGVCXho1i5A5VymQUPJLapJKkQF1Z6H9P88ECtXmeolRlnZt
RKNRdr6HRfjlO+vSbjHMv52yRi1pNoAmN6gXkzmyj7Oug/0Ak4DUAKvGASq6p18pHcoOiNIcapa/
xrxKbtgGtOlFJXmdkMNtoqwfzS7EglO2yKcCDY1XBaGVfYNZ7wpB20YyXnATbR6HBBh3qixbrTmh
lp+nysEI4ErFtvPleDRa9cRuzzEidPsmvHWPCE2i/FI1ikBguwvdhrAxukygTeJvO8908aYRX46z
D8859DKoycnWXAXNYcc0GxI9CCyAPqiXo5/MTmc81FX61RBGXqJ+SJk7nfol/wML3XudKfRuAeWu
pxRQi/P4Sw/+/caMoDcOjPqlFsXB/Q0t9YtcYVNraGozOlpQkzZ49WcWxVH3I2NGUadyi8PDMJJi
6ra764OTUnj7CR43V4up5wtQ4vToi8WzMgdN8TLnnsOYiqVq99Q0QC1dXjxCDHHMjsAN1f3PfHj7
dv2/XYfLVSDbYz2yeUYGdt6EsBD6cwoEgLLlgA7yJbsClHrMyNvdXgMQ/oiQHu7sRDW+eIcsvZhx
Oh8X1PVU97Iq/Pw10R0Kk774LvtRN4q/s8bts04udep/Wq/9suz3UWh+IIicxQijyepivUtB651A
7DMYLfxh5WNyj/0SA36jcEzUH/c+uswk8O9P3r8UI54Ocui845CKO4/97YSWQE5bFRo9k+PQ5jX8
7wb8pT+8OKsjCDW65AcQnrQCcQ/Qr/XNqHd1fmBNc0VKAcgXFloxXPnf8jTR9RpvlW+okezWsAHH
AI5+WwVBvIp43+j220GkzpY4ikzpec20MDoTkgdK3xAbqwXZ6j40eO7yN0Z0wP6ImtBk2OgERyGo
RS/lfFBK8UTuuZNgiHAZAAilIGHqsTD4UBhKJ1b5rvWDN3z5MvYo8zC49D5sujnKQzX+DKr7szEL
e1nphxztzs/Il79wS97xvNZ5JpJ7V61nbAdrplZrQFz7pPAlW+UiqOk4WeFDsLTU9ZNZqYY03gGh
qKLhQ0sPuKahXaRS1Q7TjtjlUH++08e7pIRd67ZtbesrRAFV9ybvEWFEePXnusPJVOAqUlQfHvlF
MBahmWnx13KPTi4fHn3Y/++CXOZnI7Nk7djRsdrL/WjnMs8irETU+GODP5JVljuuWsnMFC4CdMZf
kuAEf05yYB3EGSsq+WgswPBhjb2xih6mnfe68teiKkt2+jQdJGSQoAqA2II3h2r29A5WQUM+RsDB
l38e6PGi0FG20y+QNcFyOE2SFxekx7NOdcEfu4j/kLNV4qygoWbLDSTi9WgJGFHcKatx7ouc8o2k
EvCrckD6GLHe29O9tqy4TomkBr9R4Ko2DwAHeYckzOBYHslXaMpiu4sI0Rr9sWnbD3u30hk6EkXy
RsL/Ii91TMJbVP7Fg6/+Cw7/KkjL49xzwZpZZuX+7h2Wu4kZc0FkidVL97Qm+35WDykVAOn6cIVd
J6w24Rb6ONAuYCgpQaeEIwm+ROr9IiuvQaO44+4rhzA7QD4rFn0YvYWu2u/ahqFrAwk7/Bamvfy3
OUJ+msmWas7WKLVi42QMCnx57SzNAMW5Ln+9Jl97yciMvR2eAY27/CZnVMcD60mHz7gUkpmj3Ko9
m8JVtKB4JCUNclASYiCUIsXr7IJEWkE4mdU5W/miQAbrqGdI3ok+CyTnEN0zT2qnA+1WOSGvTfG1
aNwGJt1mM40CLCgRtv56LdOc7I2twXGWTdL9R1JGYi2Zs3V08FfZk7H0jL/1HRYEFGF+MgDd0vaA
WSNi69IWtIouJdtrFXlE+l055faTvpmWocljQCdM6OFOVCPqzROiHqU33acP4vp4OWOYBxnPDI2e
HrM00YeUC4lc/iBNEBEy6E6iy8aeIH+JxCM6Qf0D+6nmL8SrGwUk8KxiodXzrmRy4wLurXYYS6Ii
MAX7/Ge1Uo/5a1B0X3DLz58oyTOSf5qJ520jEts1OegfeWaJ3nah5J9AYghZ+zLN3TBGfE1e8NLc
/Fr079HxQY1nia/e8fn5r6V6CWbzV/P2c3csSJcipy9NHRlXGVVUmZq8MZfrJfjCbxGcQ6Z0cwyx
s8D/2JWDa+IVhCXjl3zcq8EOutg7Nzg6a3jZV6zv/emRO0OdvYr80MVRCgs+PiokFFqQH40rJSOY
0tBba11EZp5YRqp+i1yl10X/0u7x32WGpzcOPnlS3pk2+lEKJ3D2IfsePomgammoTJj8feltdOax
QY7FCmHybvQsosaVqg0HTyhlSljZ4rXCYpJrrXcM5+UXQHfu168Q+CseATdpIHeoZD1fVspPDjTF
HWpDJ8W9niummyYyJvpCDgfM2q0OQje2yw6RwgF/q/jnY3ZU2iVQbphQK0uVEaDwVaC/LcROX6Cw
9fOrechBkI0MNpd+KaUVUnpok73dA7MPJefB4wEBEqnCPxUG6y6ohsF6Mtsq/toC1Hhm5K1Hw9Km
WgX+YJdgOXWC7eorc7sjHERj+fNHPw3/CUdadfJ4GxeRDerbQDkpShep90GmX8rZ2a559kqq48tR
sW/XEhUcxe4ycD13eVYvFC1opXiLLtFkBNTPhiCz4VwYKx8gw3LzKL6N3Lsy+uZshdTOeRqSf4Sv
JVytOX4ONt41LVAoO1hZBlxeE/FPI5hPIzcXe/cbc7TkrDET+0/oMQ4JOTrOvX0UpXTZEwkJxLf0
u8Sa32yb7XS7qfVvvkyOtFpoG2iru/u9AOjA/lsOTyec4Zrd1dX41gI+7uyCJIMsrhXYssVWRKXS
SDe0+yD90rdbPrIuVVwTHEunpncNs5Ctp2E1cEQHseS1xh98hAxBPLu/CMgzFp7+LgxrNM45vtG8
jTbHOpBkSJ57TFq8cesFTkYYIqD1/WsiLlOAgYipNSKJgil0Nl5vVJncSwSDncDf8ButOsJkFsp/
HHxnDh7hc0pXLdEGCAYpJ4+0hxIj5q7e7G2j41iRKwHZHK7ougbr9UK5U6uWbbDGcAYu7hsNB4AT
W8ezAzaklySaQTD1m2Y6fLsvISoAkgPI9esxmkW/Re8xGQH0TLR2bmn1abh2B0ZFuN9wwJsoK4G7
J7AUhU68T7s60REkmhOxxyshwEGcG6V1SmUFHa6CORItfGXKH7Xw/UUx7qetDOky/SCLUnX0hI54
DLMQKzrxeh/29hOBBlshzFEkarAV2t4siu/wZN1BEdjwZFJVUcrdzX+9h+je7byymJQysImBMBG3
7aKHC4h0VWAbpN1WhenNUH904RrIUN4wLMDIg+9jg++mkIlhwa6Zq5tUPpbzAq2C0YAaCXr1s6Kt
9D97y9L6JyKCtMYbI/3k0l0gRDa/6xfWQaYLEsdc4w6tVSA+6dNyA4/cwHzrhdOVkh/ZI0oKWgog
etSuG6N7kq+ZAKJZ/VwCMxrqBD9KkZSm/edqSB6hzXKPmxXtWycM0xoZveyq6m9Vs2dxRcQfHmoP
1RFLmGOo2pKg9wexzsiJIgWWfoh2xPo9364Gk6d2IHdSgPEdovsGAovMtdgJzKbPZ0U+Ew3DEzak
zij4mr+euaZcqnxPPFt3u1Jo9MLDg4J8qv0gYAvxNKiRXAiqHWOU5B9YVZNjFSN3pgvYuMjNK0SF
A/phynaJZkhHErDflFqzMkSb6saWjhwh52RL293Svu9zjNXqfJ/OMKl0a18smmnceaLCTFsuJNal
GlWVLOCoTU/q2k2zE9Yq48KeD5QYD3TOzOR3PvCUR1QF5pQ+HquuccEsYRDtm0aMc1ibd32PnW2H
96iAzVD2+D/eDSDH88gck/ck3K7mgWhteBil6ilb7zZ4T2WVKdtqCtWhMjYXBxB/u6IX8tR4Tp7M
I1URu6ekHMRlb8N4vtW4LjZrcylraFTFFBdeNz5UGUl3JlwPHIlfQNOh4mWweLptoouhGqWKXnOB
zy6NaRPKXb5poCA1AjyI39tKdn1m+1H6YdgdZVNKDeje123X/tajrcQzMc27YVs4SelaCwcjlfC/
h+ikPmqBzaeDHwYcbRlwjpPbCCDufWocrI9ZBNQioK9DwigGI27a95WUmRg/rMJbEOVZSA8MmT/z
He6g7AZ9uReSLYOb3RjBacdQla1pazIaNLxEqicXKZiRhMdH6x+xV6Iedwq6l9QcogLaAHnwKqTy
whQ+cfqqJ2zPCGP10f3TicK7jH0a64+nqMVjFq9z/MwwaivBZ0qhk7alMeaiHjJncBTVr2Yq9Wdp
lEi9QCeFD3euBfhg1DsqQZwft5RSr7dg7bIba7/zBfh9nd+PJdSmKmtcyvqltFUCuO9AY2CFcWCT
nGVaG16s8Gd19EtFExLfr4i/LDN7Sigk8St2tiS0Ru7uvOExBfIK1Xb4r+Cu2qBG4NvQVSwX4ZGQ
/mHCDQC/Z9j0qhSzHqVNPF7p/3OVf8eylP0lbb6yrC/mvsuEQa+rin0tVuatGczyRfwF8TXddW31
MnT4Oj1YhSkpPLShE8KPvs/hTlijd7KZ1gBpYfnRn3LY+QWLIkQNzrpmW65E/BXY89WGWuW25qWH
apGrRxNeMuK16sxVqicD6s83O4vkJdGNvki5QNCWX1LOu/7BfY1iytJpREWHpO3IUuoVpDris9je
8fDoavu4rl6wM45h5ma+9EfYlGY7jO+xJgLEk8W2coVYXKDYoi5FErNuZcNwaVjgAG3UsPbSnjIS
NhzbpNhGdMTBjPOthkZoQFMjFlxTDL9amYiSbIDxvKlW+a+XzwJK7bMQgTIH9bpewJg2pb6S8PUG
lW16u03A7G+llOKhSrvchEoqyxHRBrY8/xhllfyXWNjb/z8EdOKVV+eSGoW5q+Sc5aDnv2t17mld
bTRSmL1CrbLMLExVAB7rgi3aw/dt339q2KvYfqP2DfIMPMbP8t+sd8SUEOsj7hzxSU6qFaN5xqTh
Py9mnovy1yyR9Lxd7VQq3kzVOmxPU4QYO0lnWk/WBEIGPYWrYuA46He7hbSbNg/qV7W5cYS89746
EryWk+a+QDfVFMLvgc3i5pkra7YvPQZOTOpVWLL1sS70yf0oeZANCSgY7uz0qH7YQKDcdO4aHTB1
VLH/i2oO7sbhn18QMb9od9ab5+M4DsSa8JP5S8xnweyX9Afc952mMXckLCURkCpTWwW6jHbplnuC
n5BQgdC4zCOTGs75A4E17TSMZ5SiNSPRK4f3D7OHt5xIvf0mLFWzPMP2DUt7kFar+mvkCiL2chTE
6fXhtSH+4FqDxQrvNpuz8upQrmJbbQApgmm0tKLVPgG1XWDoN23RHH2sI/Lpp6tbFrIbsyWg/d3T
AtzN8ZgZnNszA8czejxMcNQr7gB2FnvofDAzTjC3vdFQTufV01GjrFkv3zItBFgV8O2bUUn7U9YO
yfnaXTYZ0y4WGFDSDcbcBvdrCLGdsH/gphW5TYn8WeBPA6S2yummipPD9RYwuyjkxKYGCp70Whfl
abLkuYi0odrhrKsqOBqJqEJ9LD8F8NuFeDC/ZVdslre/hYbz7EpEwjELkvKkInphT/ErP9jMd1yO
OYtTnVcYKK5ZAfgqGiJwVg4frVAqAi94teOvbu4KpwLTEnMQ+r3ECrgG55iTHDslx1/ZEB0NAZiP
nX87d+7INgIbDX/CNhGzC3+axsCTRnf8DLbt2E1+OAziTzsMYN8ko0UXW+qQLBDMynRkKkPO78pl
9C4DA/7iUat7iQda1nTPMZTpUO4X0q838XBOYnuekAgVQ7VRRLdewrtfjfMWhj42eFZDpRcWSEm/
9MNt1DgfqYcLTaYnnMRzW8QLGDZ/j77GL7hDfRr2SU18M3Xvec9I/ImRvt9HTK78+zqEtq4eMBzM
QrYqeSzVp+b0L2dZkW496Z8htzS2gP1GlI7O6q4iAyGe6sGFlpP0u1Z1NbVsPi6/c3DiP2R9P2u+
f26T2cOWn0yEYm94A1Wsp9bXa5yPZg1GsSnavjh9wGew/yQzQhRcuQcctqIPS0UjshOA0RV/O59m
/qSW13zacwBYIACyf3VVzpDz6jcHD/K4IWeY/U7OKnZqEKG55IKLoRq4E+Fhb3ZB+LXxjV0hOQ/+
h96P02/6AsLBVHbkkAYR+CINWSaXdjXDcpimDobrLRxMqsrZxAoRE1nqyzbJMUAPuDlrTP/Mo+jr
+64G6i15N7cMjT5SA6w7krfu7jh+HsR8RtpXJ05k6oC3aP/SdGx3i4zoViXA/QInmi8ZJGCIITWB
9h/qmscm7xR9hOx0tmDUTTjeIoqYGbe8cXu8xKQyWRelGBsQIOeo/zxVgTpA+kxjLCN9QcNpLbCT
gqAY+1QOntiJ1lgyRLfTStq6zYUpYRwVNkn6k0jMWHF0lXjrY4ofR4puGMj6iM3hKuVyOZHkeAqC
YRaJPMaFzQsaVWmOZ5gEjje4L1zyBWo8LNhTNPA/FnOqflVXrEVuEcRwyPni62F9o4aTxR9go2Bh
7h+CIbCSYdHNwTNph2o36wMy7S0/Cs4BXegyzbhdghGmhEhoQxgCfij4Sh2n36m4Z3XGo8XNr7nA
CuFlhOQqjJ56qJqfBkPDMhdhl5Fx5NLWgfO2E1dHkSS2P8lPZrZktdu+Tl6n58da0/83aKGHOWa3
LijtLHaNCx9AJU1nC55gEXT1wM+Kg9NeWhmta+mXQU31m3RSzbIAbJMHQ0Um3ZBtUJuz7vuLDQQc
aiShtuWhayGwQUmFr5ZIKRo6dFRS8ikqfZVJPCkvoDE4eBGCtlWvtIHMbYXh8QWX4fRxzAmGPPNQ
AxVLao2ECLBxIYlZfL3NWgbEM49lPsACZF9pyUTgztWxXIoTNYmj3kU51lyv7ViB0VdwQGPQURq2
wbpCj3LC7MuEEZ6ZFtgXlZRRBshgEwvIjo+gU8nZuJA5FnJaHHQtRxOW7OP3/lAPgDFwYOfvhN4l
M8XKgWZV8z0eXbI0Fps3sWuxWltHzusJUUvX9Ywl6gR13b3cAr4FZsX7gVAKUi7UGqfy4cI4M+VI
bEsXtKbENGBTRxEctseNLgIeWIoCsIzUA3qrat0on4hx1Iv0GVMkMbK+cGgBWjaNlwxiXMNlK8rt
/jCh1AA6QkKEtvgaJx+WCLAd6V3Z2SC2suRk5u2oyEn5o4MWHqWN8l2Cf7lIZQaXKOBpGTyJ/3vt
lUtZaUUBVNbRrhmCivN2ZtXBposL2SMYOPR6QKYhfPYPNc25aX7OW0GLWDwrO6T2gxNkUY7zNAUO
qwf8zAz4fX8bPpnIarDOIdy2pb1+N0WijG9lIHcMy8Lrr5oXSxWp1+Iu6XzWnOnedP5EcvYKxLk3
Ny2w7zdmayYwTG/Wb2ZgNEn8hlkWDc1UTZ4CJ5cRXT6Zh4HUd7dNH4OdNlDTOHpQV+KD5K3hFbjV
YbwQY1CCMxBxaqN7IDPjXLmlLYO3L83yEYstSPuHtkG9zMB2hUHZj+NTAXGT4bnOFFrNJxB4yYAA
gBGOC5XweFrUM7dpusVnJvxcAgbHdPF8nvCCVdF/4PUfX0IRt7BdBDRaz9JXbY0dz52aWrAhjHKr
aQOJu+Vu5ylf8Sx3L3x1PtwO61sC1PETCSgqw01mGHIXsHE79k3iZOO3qODBGbAzKWg2/Q2UxEAH
r12QcXUss4F3y1bPI3tjkRU21Cxyz9lBwq9S3F2ZH/frBMpRq5ednRfooe6+0wvUen07jmEsCMww
y//9mCtnGl0e/xh5WCi1e613wXP+DJfR6XW802t4b9x/Pr73LPaVEnMKeAcujXRMrkCYegAF+O/c
IajrhZX8H+cb1kWaLR9lbW0sHqmzCphVQ/xIimT3JQeyExd3kokh4kdNbSLTnW8WLhs2MyG9NgmZ
FLlDv7+MOxQsVtB/OB0k3aXda2ISOkrwXXQkeZTqcpTAQo4hs07DpM680ue2poeQGNp8SW9013Hh
LpXWtbbmhhquwFnN9gHkJILOdqojHNfxM3I6jydLun+zMDg+8kjNhXEwdv/3Ms3v34sIcZKTw4uv
XoGgNt5JcHyFfLI00FNZUrETZcoJPwQQA2H2CgZpeVyqznYgEso32sNWtDyWTgIwDYdhAq5L3mjg
W2P3wd03Rdr0gfp7cW78zwplm6ntdegUMJ7zpVG/ghb0tgkGD2TZQmto+CnpArr3W26tHr+T48gS
HT79tLFritk52qvcalLd2VBIfob1uVgFrpFblIFj4nFBbS1v0pU9CZTXRrPXkWnwjmPKl+eS8Ffc
iJgjAsIa1Spa9WbBUwyUIu0IiwGoCps19Kp0EbYiaF50lH5htxfqd5A96OvLpDkhDVtQbFhy/bV5
iwHuJ79EjYIeYR84cB5qKNJ4Cr+yiBVzOqvQwGF9zwZemP9Wjvx8TfAnIYvwdCbioTgKWQ37Nhu0
zCa8k/LHO69sEC7aI2EVclPoheUTJFdph8yU6n22IIvz9xTlXC3QPt8ODNgGXGOAMqYsrtFGjap6
xcgfXHIk+539o6quLHOmlmgL9vc+xZ/Ylqjbz4Ako/RdtcaKF2YZuju8Af20mwhRNpx+N9ZpQv9s
Alh9qPNercH8IF6/gl/eHlN9reF/n+AQWqjBGQL+jSNoggbCinkloGfzCYAuGRf3pW5D3f9BsZrr
ncHE+3k3KhyDaUrZOeJzyCFUGe5LdGBfrexw4eLCGwdB0gM5V/SsfojcHhG0qhNcJLr4z7gyeEiE
n/MntTV5F6Ns4kK9T5+lnY+VwNaE+QdIl1iN/voTDR/7zaUFA2dPz0iLOlcyz1rwTyQKYkG23l9S
Yhy9rTDpKJ2QUUCbK42hmE0vEoWBVt24GaYDgHtTYFxBq7lfaUiZ3wPQKTWynSYCxL0ax8pNtK7B
mtlKBi+L4rpNnorNlqEP3UDfa6Or586vQVMMIrJeJuObUipBq5Dcan3jwTfSYaiaC2N6k4XDVSSq
W5Cvv3fFf+09QM4z8+CIzB2mxxZD8dBQJoZFvZ4gLMfOvbU/UJ0hO2R1OD9AuFxZCNZC4xRlb5Rg
P+68BSi+4yz9x649uWM27uSC5P20Op7AhQsmCYuEK5XwnjfMUR/YsTCa5rxWhtn2H+yyv5tyft1p
Z0jiQTOezcLeVyvpKvQgsGGGurTe9YG+qW63SPRqR35IcJ/KbSyzfr6BG2EZwG0ep3+WC+DqH6Ym
kcTy8+NaBScsSXDFEKw5zColP9W2BCNF9BHuzgV5xE6tVXM5MO62EbiIn5IOKiithg/A5boM7THN
jQWK/ehekI02sCDsW+kjDJaDrG9SLbUYTFJMcKHjkzPcwhEZG49lXnDx5dgEneA3t+Hoj2vHPbe2
69Xyq5sJPO76xO80dhtpusprBGfg1UZ4fhJViZ/vvxccFIusZtekKkHNZu4+Ld11yGht2+JRtB+B
SKv8wRWFuf5a5reORsaqIRlwpYRGE2tyj515CvkqFaB/9St5CO1CNXA2qLmMM8gmHD27+3rn7qIa
YKXzZu6oCPzcDqFmA2xELsUil5r2xC5HTYXh3AO9lfNkHkYQiy92+1WSadB43nq4cSSCuAnkb1AY
9JTfMG2Q6rVgtI/W8aN4LF9mGMihdOONu25AK0IDN+t+ouWGpKgBU7EhfZIZar7JGm59gDZyD9nL
akDI7AVXhgV5YsFA5qazIz57+8eqNhCYT4p5+xwAbwreLkIYMlelv0j1F1Nf5V19qomlzUXTwar+
hIW4QiESGpIi+vI4vhivj+Qq6jSI+sMO6R7DvC5ZbMrMs5XkrTOXaWc4xTnqTnW+7Hz4I+SosgqP
QicbbOY0qEEnc0VYpC7809TPxd4RIKXj8xkCJDEpa2IvvgwzbTRMLkUkAvvMat1n+RNliSojo/i9
pBLOh7XeKA7GE4PRw4b29u8oBibPNYq+E7O8KrkoGDC8wh4FhL7VOcoJtrfp4Mbb61r0XGUP0cvn
6VlMvDLKWuxq1n7G5FT8EM9huX6JSsEn3IzHU+TT6O96If2sgnbQfTo2PeC1lZpAAb3bGgS2gQMK
zUSK+AvczhdG9iN/fHhBtEfnTOCjUOB1Lip2xVvq084iNaY2gv5Vb/0v86eDotH5cMyEKYOfU4qt
daEmwuWRNVG1pad/cFgdyZuDTY6/sgx531gbBX2kxF2KyPklomcuiHTOZ5ayfUMVWzcq8xlESt5/
z+tB/pMP+fmZESeASYh3FqKN17IFMFa8Mb7WjZEJa3qjr+nAcGPGEIyYz7hlgDcKS2CoROMtxzvk
N7PUZ4opYKobJuJ3yqyIFDY7QbzmptGZDZJ8uc2EiRE9b2futCXlWsPM1pVyXVSNuGs9WhRfVZNY
IvJmS0h+gud+OIeQOldr2HkeLLUi9lzocDnOlyFIOXyCXciN4HA3d86PfgL/HjYDmsknfeH2QvXN
IgG56EaAwSxOS1QbLcUpYl/1Fam5NkQjcRwHcz+MuLGFfKxjHnms4UWGYjJ3rwmjfZy9/jzTy/qG
DYWr/85v/Nbug8clq44t4iYrq0kb+FWKgZffROu0alIjREpPhJkIepZ/XV3o7Vaq0CRP/qlDxx+g
lqL1u4VJqRhRTKonunqt1dGxtebYPnheHARP86qT6jr9lsqyVaopVmxK2Hcqr3kTreSNpGptQDX4
gBB9Yfs9eWYPJJc9pII7FPACOkTbCHP0Xu+MjbbieVPa84XaTiRlSWt8EuWkD0wy/0UkzDfH6AIM
3yYa6RpRjWGJ9EaMGeIakLOxgbwTFioiOnmacPfYDXmUfSxU23By6v7daUBINpgJTsmTz7NignUf
wbjRvtBGkLNlqzJ75bZP0dXE9GcWZ96XvLF+2OTkdv9uuIX8PKm2WDKBWp4BZYHWDsZ5g4EwgyJi
F7aVtXPVxhTWn3up8koZFhezARSHR+9+UKJ8iThvYt6rLYI4VLxwEC6akSVldXlRtSZRim4RYBjs
JHL8cq81cbDtIQkDl7ja/H/h19HBqC4e+UH9gVoK0ovF6pYIdNMt7f2Wn7yFiiQxOaDCLb+EpfWd
/3F5MK3uuqu+eL6KouW+XMEJ+wwgLKjEjFKnMP4qIykdkgsGtO/a5eNgOQlV2Xmv0vyIDjVXmXKn
mPkRHIyoOL+VCZDqwFK2MbJGbOXAONZsYSoVAA8YzFrT/XfEIk/VxYAUBdHlYOvk1L8fOFNJ4uTA
cI/VViq04U7rtyoDRgfiIOVeVX6WH11rch9l9aQgWcgXrSlz0HbFRK6UvDwHsgeAgDG5x9VucoYB
60Ad4+Exe/4fK0UJCrkE/C5XeJOvdRQA5gtbsRKT5wlso1MhEzUawJP0DDJ0cbrHNeNAnm2cNspg
whmO4pEIUMogx/kt5t5cTkEM52v8dIMlEvCAbe79I6DMM/Uv00r0jVVtl4ZB/A2tlD31F/ToPJWf
sqgHh6AEF+8ZSFtckFcFL+qJ7vG2qgJV46f9B5bSYerjIBh/w7Wx9xfbSw4DIbWwOZJCIjYTVOKG
ORxW/3OZrmx2pP6j/2N9hg/BVifVzQHzbN8hAIUQbR4HhWS3aOpdK00Bm/xKexetpAQSitRhLWoC
1odhI8l1ceNoN+MzhqB3/sn9nYpaU9rU5arOv3JqodX87i+7lSpNlRBKBatGwgT2b5XuNRsULizV
InrT+WJ8HO3M1ifRMp2CLwAbZA5vtmW2i85qwB7odvWwa255EBrfgbYMEnFJmsmQ9akMmo00Wsed
tWE9iyGgO7h+qtOFV/AqUmYsYWmmywx+Y0dgZwe4G7YH1Lt2C++7SctvJuj3mDRDpaxabUx/OaHT
T0j7ua+wTMVCyGdkwEPrXPVf/KtvvJgbbLHMShV1T/DywgCRD84lW9BFfE7zLQwiYEpec2T24wd8
oV6ZvuLqp0DB4d41ZyEcoZ9iMGGHU2aXw0NoWWzhOTvwwKNUx2UVvNl/2l5/dci+xbdWxRK4hU/Q
oY4Ro9xCLhrL9Jca+Rg6xIgMJrpRa9iR3nQ+LOinEObKTcwkZijqnrvZAItckqP8NnOo+hTeXcYX
qgTA3ydOg7y651Qmbbr4hMNlyLUYICJAQePG6EhSsVSy/dlyiJiqfBwjCBhD1EDF8vTFTCjkjO90
IBmbXVxYAPCaqhX3/gsHLkSzV2HjNjuz2RnG2iuCMGRPQNiC5F/oBPggZoUHkEnxxDZbEejow9PT
MSkQ/UUyh4A4XkED8e8as0P3rUapIKX/9WNx6aZIAX1tF8662r4uGfkyStxwZQ/XQ83tQGqvNiWx
Ha5R03YvQAPfbrZ3ClVuoB4eIGTBIBVR0BVVECA3BUV7donh7BK1FT1bhajVGTfImzlmo8xH0aJn
n4B++Aty9Evovw0v3X0tLe3cANWCEg0840HPU0tj/oARddxpV6RRMAipWF6fJ7nYIzNGSNi98UsZ
O2J0ON6HaaOYrzMMGCMN3RPpwacdsYWwDJwtHSWUMXbURJIKC+cxWjUJINyrEYBeztvPqduE6ZZG
nbC7CSPZ6zVZEe6ra78EBp31ww/fPq16j3m7F79MQFKF+C0GJdVH8d+/gKSY2lampuFPjmtxblDY
d/xQoqVOR/3IqWJ3dbx/Aq63XVxhv+Vp8QSAKQwG9pmts5juZ/1iEBtnQL196pftofScvNmJesS+
A+RQ/3WRZyZG3Q8qW7yYSZrHM4/8v/HplW3ELz8VFTiajRL+4CoSvSm+6fZ4iMb3FqTW5DUg/jjW
BPZOz+Yrs1a01f5eKpEySWzHYDDhBWVfjQPTCUd1oPj3NHKiPycDl4v0Xq357gGQ55/GFynLgbRm
enwELi21v7PybBdasuNUVyhrbyyyyQTE0JLDwRa0iuy47fpPFg4ZxSjFilpzRPr+2tJlNxgQo8Kz
8f19VmYxRZBezBsiAFn9iAI/B/cCb0hKMDX1JduQ/jVbMATd0gbkLK6iK+1dOn+BbVFOx0ktMqSJ
X4VUOHgYaT4t+LXu+hwfqnW7xPPnHqefJWoXg9J0WYBt8c1rBaHleEZEhAH+MSUyKA165r05PfjC
L6IQRX4+g6K/8Mz6jnT9fPSnSgB7L9MPhYSvWySYmco3RszNxgQ/TGYbv9wV7yhmg+mAt0AgvOQw
vOw5aGu5PkXTdYPDJcsVeUYTz48OAWp50QWPDO/SHDGZME7w10KRwgWW/g4fIIfEr4nq82Q0gWK2
f6w3WtX3MLMvX7mWJTUc7Uw6PamOyD4NKeOIF3S3HyzLPejImRZHBZx4izoXx5GIWFOR1yMtI3iB
FmF6XN7v7tO704TUimyRBAFulQHBZOHdJQTYFDN98SQ/DyblgRA32AxoqzG9/IoductciRMrauU6
KnT77mBW3vkIKyElI0QE5KpXWDCmS6RkadUeDLqryH/ZGjC/vty9elZPYv9co+drsc0MHv8atWM6
PyWIUhcffigGydXBlBiDmf+JR0yYxYfQE2NI28j4NVMof27S1WyFkfVfb5HXg5NwwIOxt6Xfgiw4
5EA1Rk4wRN4k/ayBYFp7t0uSlbABJdWK+U68NUvW8na8tkc54cZ0a4KS3dgzoaODt/SGE6nqlARQ
+G1Sb4n3x5ltEH76YiMcUVmeelOavCvHXRAkYlMhLaVQ4dwEwWDoN4lLZvL8hh0uSzGEZgvMts0A
dOHXg3HkCNA2s5KpO7/aq215Snmq5ps7w8N5t5BMfvmkfaURKww6ZwzIutsnWVZJYpviZCei+3YO
pUDOAjAU6Lz1+rsu6FA6YYlqQM5dJBvtuFA2qxFTwu7GFhuCVuNfF9HgqmAgEUkyzf8ckaLy7QkJ
rB/tl4gOfUVc5bjaFJWR6VwnvAvXL5hzNsEYlGCB6G+Q9VrcUN4ThBeaMnkETPUSoZ91DIpWQr1m
uSqmtGzl644VjBA4YIaTcvhJnnTq8B9S10cveVVDHiPe1xdXi2wOop/Uz4DYYgw0D2+n6VCLRE6z
9ra6e1HAtYmkeXE4T8bBEq28zn849Lyoz+280kpTCU+QwvWqT23xA0/NgEnfbn3x0jP+SqckuqgF
LsGITP+H97Ouk87xaU74XR8s8hVzov9XeE1KR177nHyXtOE5A+aMBGPKnE9BFLlQPGUEAFQbNKDC
sPYeXvTmjcG/bt9Xl8u3L3N2cHgdZD9Hz+WRjozxpEL0k3MSKxcleZzvfU8+8KP3n+DBEKQF8UsX
F2VTBELltKxBdrOsatX93OVBVlNH8s3yGaC+XmYdNRbHZIgB3w0F7rPZnRyqRpdOkjlTaVDAuvlh
+QfGxUcbTkZB7W5njee/wPTYAMT0oeKwQIIrICQE5I8bkJbvyXFaJlgGISRWBFmZq8x73PMMPYQ8
LY7XvOdCtkIJV0vw0qSdkD8kmGGceV4N7Fb+P8pOpPc073J2rsAaWQCR0ai5j4dRiM8UD1xsQ3f6
6NcCmiATdQEY0TRCJHYkM25jRrePt8jGLSxiKwq31Uzbdfv4uz1I5EwBeMDR5RYVvL1JLTFfB+8V
YMu615RICDGgTK26ahLfa5Z6sNtAC+ZoA43JcFzSxYDmPh00abLXKPi0KZz5CRh4iBKlQx9u125a
d+ENqUaiO0kxN609r2tAMUJU5L2Y0K3yjFU6nGHDQaG7MpqcMQCAp5hE9a8DMwk/pd6afvN+BHmr
rOPkJg6Yi6n/DWm8/Qi1jTiLBeCvZyy1Xh5FgS7I9VxCbXettixN/fqSAPFGjiDGrq8qizt4jB5i
gNncQ/A5NoACrGlJq/Kc9sy8LSyj1VV0bJAh2/QvtUa1A4rJjZ5qk0NAPv9oaQpl9HWcs6ws7TBZ
mdbEREWILmz4LybDfBg8u2it+KMhlNjrL2z+ICIuTkrlOwIrsAb23lwCX1LWclPUV9Qx9wGPW9BT
cLf7ddqRBwwQzVbngYEehSEwbYG2owWOA/ogeLwWhP+ijthIlmG1vCrGrFN4LxewrkNURHEpF4b6
L+ggccvDoz+vyLC1ZlO/+R3vhYq3176jgRO/iaED73Dc65RXSYWVCP2KLM2FTKgxNT4lhKtzX4ap
umrQeAavNyLFz3745AktBKzd+37GPUa8NLMdnrXz88B3BkGaumHm9OPNmAZbxSDTTaTlkgprZMCV
tn76PnpdJ5RLoaLbIwASKTIvl/g9tGVaNq4FVirIl4cz321YI1COtzM/sgAPbmP36YZiWIpJJOfE
AzKNFmxGMPF/5f1iSOs4J1/tGhRO6aTI/N78a2q1djf1CC1Y3iNvENLuuAY0HN2t5w2/VL4AG6jQ
BsgEOddR/vDVUyEO54nDqk7GwtgxL6b51VkqztQBq7OJxK6YqWj7SzY6D1GTkpHqxx4wmJFhAvTb
3NPXiCS/kTsb9N3xVdybFA4xIaPbfet7f2LZt8DwDfo/z7qPUtPmOrZsk3w51sBb7kT7OE5f5R9A
hKMk45Qv0Z3mS6KADBzk/1zEwn/NekEEtABNbm9DGzo1tWD6UmT0Et5fdTpWmc2yfz1XJ/9OEXuv
12JyCXj2Ylq66giHAI1NEfv6fkioS9XlUeBy1pY+Dey4gOBNpd7tu44hMBcA29pK6iTy68OAu1Cm
APuoGzJot/gg8sJAyQv8weDCiL6rBw2EAds2GZvubVe2eC1qv8eHx/vkBB10w5Dlt7MnLQ3LYfvI
pJUkJ+2dVyOhnliHnnLl2M9VgpZPNQ7eD5QizADyutw2sCVZPJuL9BGrViZ5ERX7U9Kqp1GkxF+l
s6U8kTRwgzDhCheoymUJ5B1F+S5IRQ516CtWKyteg2Flor3AsgL/Pgaj/0bJNkPag3muYGWKCefM
hsBO/cDGmmu4J6LuOtZJ0aa7rOMKq2Nb/a5jN0hzezF1clIBViasmyMtW6S6WK1QDJ3ydrZbyMZw
lE+FjXqfo1BDR/LoV/dIRyn5lrM9xeG2NjZv8dQHByAc3ghMK0/GcEDTDTa8wzYCmxTepnZ4u55r
nbUqx0eZChtk7m931TePm99bgwadXN6Ws+RJX82cDrb1FOdkpD7XDB58H/2PdYmWheBG6sATXYNH
ghIpIbXpy+i3ja1ZmyqpswyOB8jwX9nCPq6CK0W82+rXnEXj11hyxW4h9rlxa+2vj3YC6cOw9M2u
ArkR1HCiMJBHlHRfTfX+J801XLxk98m5BMHA4u/S+AmilFTePDiWrTUoWWBL9MIG5E0r5smKla8W
XOE0fssb5J+jNLtH3yhXLhGypiWSjUf9/3ynVF7jXm6ZA0gpK3LlNPnLipRrRBNtDdRkKIv98Zdo
g07sS++JS5mzB1zfhR1NGPatwsLkS+oLtRdJ9vnxUVldzszn31+oVsB/jLF/llu4LwLiOkrMJ1Er
4KNb1iN3xa39YS5ny8XNA/680jS5a788LthnRTh+3oYY5RmaV0uH5jukmhq5lAx1D3FO2l2UIJth
tv8/183C0hV9l4vTfJfFoto7QykqkZes0kUl7cj0L+yPWZTvuNftOf1DVuSJp3heqjzpG49mfxid
t/fDJJvcwiUi/CT1n2u33MSvtVMiVBn82YSLrcTd/dycYVLFA0b2M02/py361vprl6onSWph2Z9f
KahDkth4J9LoUgHwLw+/NcQDwYS7Y2T6ev0zZKi1SRHm/EVjbVChf6qfh1isNdJgstZSRue+0h0t
o6uSA4ZZ5Dcgf02DIoHkIOdo26CIj7Y73pjYVJYUQ5BcrrNfWuuxaBd+SRvIUZmsKNrVhAe8yZM8
gXSnPWA7RPwmgww44m3MEhxxDrpqXwssqtKebG60p8TvhcS4rtFA0+NW4RGh0nCo93VbTDHzm8mu
2upda7DlWaEcwFK6XYFMRh5lKYNGL04o4RiqWfjFSx+m8dgxcOp7kSnLR3h8sGDLzq4Q+/HHN+31
gz9EjTGgCAufVltuX/nH/vA8DOMsD3OFx9AmoxbhHKndWw35DC6Dv123sa7I+qmk2lg9SYm+s+JA
jRQt0sWh+1WHroqssWlUhSBNtepDhWNera+WzvUOw9eofNEULNd2beEtQ3rd1/x4htoWAGYT45AR
+QEnNE02kXvZ6vZEVnTRkAjdqIaFvBHr9lXlpXZJmgaS3H81oxkgMwjifPylqEWB24/NSFmkniAF
7yWhUJUzql1IoOEuqm7MtWP0ACfNx7SIiuru7M6VMbfLCsFM99JbVmeir0wzTq1eVfkdi9E07gIL
uVlEJcJtT5ussueMhxgmragtdja1929i6CauGe/oAOIphXaGyWpiw1hCkDKw0DF6faBLwpp28ZkF
Gvq1ZoaopxE4MS3wRpucHWauosG3nSRVPIFSiatqmdpllUcXjvy5Q5DnUerA3ORiAygdYstPbnK6
GTTkc8YS6lW7vIXi1sl8EFuVjqnVeeKDoGeiBxY730ZcS1BkUFz5qeG7H5/ywcRbnbxHrg4cEef5
sD0Q4ZgJ4L/UhZbU1xDRgTIOiTa7w08HuHJlQMhSu8cw8pgat9aCr+fGP+yStgay6lF0hhfYH5I9
v1bKQxY5yYGiqudgIbri5tsGdSn9OHzbkmP/NoFcI3ZUCEr1OvKjS1gr2qFfBcfOI/cnIzE9zXyF
VpkY7k9MDltn4ia08cgAERMqZ+hZWSi8odv3dZHa8LjC+Zu5JUz50pkgD+mVIfRhLlNJSuONZqQQ
qH0B3XZ8oWfVjDDaQ7RQnMivos3gUYY0sQIBVrl5MsGAG0/pb8M77fr8O7JbxK7w7J+61G5s1tlz
kdXvd/S6gcDy7E5gAnEyrCw8n4DdtWmrtZhjLYGEiUNQBx49+Rh9vjIUwV8wkHtzMiCh5wB5l3wQ
VvsXGLwIeSNukVF0JPYsPXOG06gLNZ0Fw60TdVTgfBfTE5NUR/Ab3bd7ZBd0V+ahZ+ICYqa09hWm
Q6FeAYlpWJDF4+Algeo/HdbSfXASs+PuPLZsd6VFK61UheevyZAmhj0MblrefIo0nznE7LAzLSJd
WQrZnT9dczNkO/rXEthv7sbu93JTDS9fvVm1QlVeMf5ZjPPGK4X/sH5KSmysAZyM5TRCHS8XTGHC
AvTpjpOapxNZUq/ER7bFMMHHO/uJEyvr2EESzlq1lX1qtzF1wxxOBkOeKCjIUUOgmCsqFJChK4ry
AIbjLz8+ASbiEdlBR3wu1pKYOwTGr6RDyis6dx2v+ZSRgU1nFBj5+D7vHVNSAfOwCJVYDbS9JnPG
smzPyVCmLoTq3JLJiIevhmezyikGaSOEVUhAw/VTCTjjQKN1iOZx9EQ0luvKLSoVmMmPohVsAhKn
Bbp9m+zMEaB7vG21azdlC78Fe9ZhblVSV9o422KGN3WJyvIatrlmFvCuHA/XrJXjpCLZna+S2vqF
TRUfSfsftdsLrhT5HRMBvMaS8QNY7R+gaIJBiKAV+HZrZy3FirQeSoHG9LycdC3IS1igUOApdOa+
IBhegwPA6ItMiDqpS7kc8fMYGOuETxW9zgc1Ivt8AVnUHdZxNR/xhcG7euO7zj6WPOzlg60jqVVQ
jOWAoH2i2VkBJocS3mAVu3ErbOfDk/7g6av6iftRE5WF5oO4sEbZ8Y+xed2RYgUJe1UVsCM+m4Wd
mEPwOrv5pxXJ/UshuwYvDmKV+trouTbPrYO4Q2vikEcsBcfQBqjFts/QzuKUxgUGIQnKxjdDiHFq
/oqoPObgEPmUTgoP4JLGA+/mKHN6/LaIJ45Feg+Ch/MA2IkeTwz5eYP40w67TEpNXaRfGavWNEdQ
/8gOApf1EzdkuBGMbquXNptIF2anK+3jWdHCEK9cOJORmWZfM12paEFFqkU5zQc5mTLrtuD211Zy
Px7RY/suBsp+voLRxcc9iqH/HtvcRIYEKjcqt3nSoVwayd+G86mT8R6yiEBD6rG8f16wiG6yMghi
mlAeeYFvCJZsUkgf1kPYy0R8AEdM6FdUiAPvSBXCjkAw2CTx3ucorgOG2BBSOSriqCTIR6cTfDOA
JUfaPi1LkP8BJ1LMjYnpipUoyw5eWc+oselMuoLuaOL53N8V9zVehmVynA7xDf4NBjc1iKoKcRUu
vo+lMFiEsczwQHUssJ+VBrIj/dbngvfw0OYd7t3Gbw0sbwdxHgMHT+qFiqehAXJLD7FkoXMvY25F
gS5OQg2QRP/jObkfxZGyg/5ARgXUq1VnBn77JmnBsgouc2mFZRXXSdGgnNQbr9Ge7m0ErNKmWbtE
jZao6k0id90s/3jSomWMGBD2C7DM9bZiDjvdYVRouwXlxo/v3Z6pZ6bvjo0xuVLQFCn6y8onkpaA
hw3UGKpaBislclSTeygBBEWQGmRieIHcrbgnMIgxqzr3REqBUg/1E9hK6KN77V5QyeAAT8r1CxTT
UvD3RzxNk4sjJ0Va3r6ua2MxZCiTp7/2eVPKBfKXORgh3Ifj6T50YCxBgZdTxH9HLVpxvOhnNFhv
D5ts8S9TKm+L+TGiMpce/Fp+MYRTlN0CKDUaWO+VuUnJ9exbmbwwpvqE/3vhPCE8V4SGe3hdC6Kb
ifSC7L62ME4onUvIj+yP2uTb4sIROSgkdh0VkYv1w3lENfRHUWQgLP7JiodoLQGhcZTX/jDJeipj
rVvrCwpSCJvm1lYWwdyajNLnS/mSNWw4i3vPrHf449VbfdrizNS3Q3w+K5Ua/xFoCT9X6bLUWnD7
6rUpGJnLHfwXHJqzRoptIBtWxShWqYE2coV3SAOfoOZtUO9cVKoB1DVqtD+qgsmfYjz4WTRn5uWB
min0wCZEudJkRE9nCm4erG6qHUi5WhrHnMqzNIKUEudIiY9DXmYvj1q3rpl1/MR8k+/30N5W0RyR
7eD//1NuB3VroA8YpGhO95h+Un8tfQi/eeEVkQKiV6Zx1s9/B+OzBwKqk3hKDAFOO/PydnL2T78p
QHswjPQXeFXIZMt70+As0VzDhROdER3G0X9fx7h5fmn1YLNaMpqpH0PmXAn7jIVVE99E+wVNGq0I
0QWDf1x5ObolJLB+dizjSLNeNjhLBPDoVWRQJgDtBQxYhSjdouSMMF4qyfjheyPiWH5FR1TiNMgs
4IxwCrulVx0dwYTKnxccsgypyulP0TCtU7q4E9MtK9C8arG/h2g9ttVgwjKjSYXTe7uOXl7ddL6b
/08sLg00HnfKbC11R9RRV6umS/sid/9T6FHPKtcylDI5MY777yKqbg5Yg5WzXy41Lx0gQZmj5+7j
NyCsAm+uAwY+cJBeiky/0IWz6/LjYIZeJ6QHtytfHKXaBGuV+euvmnI+nOysePE4EDneJdqTPA2U
Fi5iVZKxh8qAXUR5wVvFIFQ42xeUPIq41AJOlEM73CV4J0VgKS53FXAQ4GaNJKTDxNJhx3A113e7
htBJNG2TC1fgAAWOYAKcwf3I0wFI/gb0JMYvEQwiq8edfik4Hexo5hzPRSrGcvIbyGZOgIggdmim
5oEF8u/8W5zu9MoFWHHb+hzslapn91q/PxkYYLr2ZwNLtgdcaEOFQ5ch4iQR+uGcgEXIxcMn9qKk
KhbeKKJDKEn52Pm/pW/rMJMJ9AvCbSOD3qT9RoirNq9bZyqAJ220L7uueiZEubqPGnx+nDWzP6kN
J5XqSBUOAAFBl4ITIGd8KQWrASxAXVrtmWxfqeWqN9QBDL4loU2vCm0+yu3SRxd6j3HiOXqCyEkV
7RdKZoOnBJESH+E4cjEUKyGiNmkPhMIWaHiXZxKr5pzm71uYJsv4NpKNTpC4KUHeQSBG1lFu/Ol9
X8aZGUOs3GUGCxPU1IFTKhJueXJ771nOkleceKFof4Ox1b9tJOm3pOvHgMSQtGc9m7bLmDn/59hx
VFimE8C1UVKmZQqsMhLRSggmWrI/BboCKUkyIRRAjYdrcUWkBQvjLR8ntrAaVo9plF4iTtzNfdJX
jKz/uWHzZipdRWKYVIo2923eprJP/3n9h12+y/prdnyw9sG4x/StOtbFmdPPSX0bYtYQ9Hrj806C
2hs1u1TCui5YvM5sWDyvcG4vauTL0IJ4bNe1bKXcYbsJvGeQv+Zws5chRjxcb8jmJd6PYbcdNx+k
/vpPa3STEHKoWdKMkRd+MDmQO2WiELyV6xolAHC57MBkhxhiNZylIJe85cRaB9I5iImj1Xwa4Ibe
CLNUVYXEEyimt5nKppEO6sKQMxqse66IYQLK2ViuTMfBSFZo/Z5I1kASWm7yJZ1OodJxX+NXjv3H
zUFBQ8DtSDZZmdhYL4G2T7uZWm8V9fgflF2xw9LQf1XnQgaODFHvxUPuyMTurGKLFwBeU4gHNGRo
B6lPc4Wn/vFoonBM1woaxKCxeZXeKXDF2oxs7r0wSw0kQEaXYpZKwqkzSbUnAlATyYPEXQ2iIqoK
nAdOGhKNTY4RP1CjdQ8vm4Iz7+1CJYFaeOpPkJoHHjOaw1jiCQzkob4caoPeb83q/M3d7QtzYTxu
rG89Jd+oOxEDNe2zg6G6cVDVGRMAaec+2TE8nTHrlC54g6tqFFPIz9GUAa5uJvVs+tcGhrSMwYNX
yh1gjoQv6xMebx3tqy3CvwT1ZbFGNqwbuWKE8XlLJDG85MQy2zWkupSwAF6Ow/8csYakNQ2zuowW
e8Ky7/JOIsCIJJqQKnOVcLz/VY2IwQURHoLP2Myaj7jFgq2xeeKUa+gqmIEhNHkz8BtilSpGQZ5V
b63TqTNv00cym7DCdvh87jwb8QU9/JtymeURMq4zpN2henA6Fg1C8s8Ud+hr4sEdaTA19hRTk+Mn
5XTnCDdChIor/eCLhg1Vw6Vp9KwyCmifwe5/TXKUftcacg9RcEhcKB6gTGbGReKhPbU+L0b5GD5f
3ROBWKZGI/jpoTgCIq/o91XO1EOenMeJr9cOxApOzz7VFHnP11wqXSTf7OWHJps2IRsiQaptXovj
hqtQumV/vuiqD487KS1JYJeWDigFhCGVYzc+5OUBCeKobM8aGwjTfykxH5BGFFuIW3ShICamrcEM
tvjNTu48ufTa21MO1KOqg3EjfI1MtTgZiejNemyHSuSjQ8StCE8pO1yvOQza/RiuMCnA5AIVV4Yr
SIm6I7MQvh+RLgnXlGIoRXRpcjOAeZ3p4/4/MLfCNiTlz1e9fIyZVBOqGv22Z5MQJAWlUmfVqs21
iwlxJ3YLtaBeibUmW+D4tgDwuAUPp6PN34Jrch6rG2n/W580sPt8nSTxfV04SSkkHhMPJL5zN8Cw
KwwoHzb1oJXjTUjmseMianTUPM4e9v13Pk8GT70fX0HH7r1Hc0U+h1yEcr3wyKHmLCRNd/Ep1r+x
6ZDfbzTCIY9Mj42c+M9SMMYV8Ro6VEzLVNbHlJk8eCaZnxFXe6UF+A07mMCyRQtBylOznApr63UZ
TvU+Jj5PVef9UQRDbHKsCKP0niH4dOU3aA1HoGM0gMsr3zFHacaPfk5vV6/ZQKfoQFn2a/EZRLvh
MMP+iOx1HXMhRKjlxIIwCnqpm1LUSmk6ZMY4/4ShY21rmJqDk7pdEBESMhSBu5Lk+q9BeXJQJW8/
BhSwRwnWVs3FUIwyTqSUcmWkl/qsI9jmEA+2zjtg11ZesnXvFmn2cGVb0/NyUKHLr4rGcA2rxVKo
pTSxeCHRAjtHeV0ooaaaB9wOqwDGFO7SVIDSEDBudRuUgmWsL2uqhNejap6+gbgQlXzEfiIGpvjV
2C7CJr+0T5wELv4a0SCJJB9kIrxXpWcuFmPttzeU6a63tB0CAn3zuJkdiIXz/IB3tM/zkYe1jn6m
5pWp9zlvQwqRvYJRaLVtsS0MNl89YQ7J1qFj3dFU7iShbYJEsncMIOVxbvtj42Pazw036mJYgcCV
yDoqcVofONWWkQRQBmQR4XrKKFU8ZKJAkH5VgOCGhzm9uLJiA2+pSq7Qn6KJC1ijkDJrgaJGy6aF
ySAonnHODscs5Ar0mAF8bVDgAs62QgiCoWDyEDHNURRwgp5qiFCxXcXMYl2hCqIqmzTEINwAGrBU
vJkOfCdABrTA/0lZzhMO0tqRMGFMU8mN3XPW0jlxcUgHXN6DnavPSDZbPIBfim9+HQif6UxUXQ3M
Jl5+Uog+scrMs3ihkuzywSQ3owTzfmiiQ4uUELw0MjncUf3W0fVIZ6zklC8vM37GbfVvbN0njtZo
qAaIJUHfoulCp2BCoeFQbI4wOn821+lKY2BNThxH8STxMJCPt7tpwU+D/jXQ9KZ0R4JOMpnfMk3Y
RJSKfQJXJQ81DqWJ+mSHpF92P4LHT/EOJ4EIccxr6RQqmOovAfOVWaAk/Cn/BiINv/sKud+FsZCi
4mAAKS9Ou4jVnNjwhZLCKANz7BtxDu+iwH1F6AhqaexH0C76e/ZlJxO7VFkMht0eYMD799wevHRH
gEV4I/2JemQSqS4Nf2GpdbAsiJMd/VqZNiBechOauNd6C0qnO6qsk3la9v77qCWjyN/Gd5BMy8ip
wDBLlvFLI3brSnNs33hFSbtUND/iw/9fYDx8JXpRIhq2CuxICr5dWOi3mQvTPugT84gzvw3vY8ng
TQ2KkRXwybKU29QZqiFxaKC3MH18K2ros05vJHnpkmFh3UnurGwC4+7bcw0RC7G3oU5fxrRMRdvK
aaVnFNZCXwKw517Ue+dOJeqnm0iKbwmgW9AeHzDzsXQWgGKr0PNfiWYDv4ve4HS+rez0wZYZGAgh
1+Zy94yF7sBlU4byv5vM19sB8oZRrIPFEPTt+yRAk7vl8PwvYyZe6XHLiEfNHx38Wc9QKIzLTXpN
D91Q3gLKvVpEjgFZmuzhGc7GYlFMgsUappCnUJQpsr7kFGvA8Wyty64fa9b3y8na+wQsBjW7Y/9j
A5HN6eG0oxATeYlfXWxTDaxphMtQwiWThN1hhgZHy8PV0Z7gXAbo2I8aPvyWTHGxn94ia7q/cEPE
I5VI3qhnKsLSMntU6UHzs4MQXXVix1DTpoHJ86O5xbxSsoAHNYwhXAfOmzJpVcdz/YvDDFPRyNmd
EDDVimezkrst0QLCer7bkp6SmuI3hVu+oyvce93lwyNu/opruVVuVQu6ZsLoz3jS5hMkG4bbM0pk
C98C92CVXUgc9pBIEgviES4mKHuBu2HGAppeQVwb2q0x3EidSkUaXPVRCY50QD13VM4uzI8tKm4Z
9Ysw71u+fgMMfQ3iPPsrNzSvDMfw7DvjB1iG0pq9dybJuWj3hq4Vf4pTSeVjQvNB4Ze0jLOpW6DF
MH3kVQ5J1PRpvLRYaqoV9vRgFJnbFNyCyeDptFFRBxDz/efEG9gZ0IcBFW8OYeJzbuF/w+77rFtB
ECeTEeUMRm+YB3tTJsd7IAFz6tqcaLinMg4epUNOCBX8+sjbJzj3vp0ROnbefogTCQBCEVIoh0p0
U3bFiHYXpGGN2S9gih6DnnkEf5iKzbDdeUsqmPMh52aQtN7+v6RCUiUdZEBBfml+tvDA0y639TD6
NWFWE4vWThPTZcI8RCksxWD88KbmuRfKm9qKrtg0ZHbbbyzVseLCvkROBp9tkqkd9xVWOukWkgRz
0a5ww01BKgz8ocSExWwtadSBVRbR2axm7Y/TzGZY1kI9J0m32oKpSnh02GiOc4ALt1AwUmEamqOE
sD2XFb4ZgwTIqHpBf+eMLFef3mAur949qACn0sXMgCH50HAZp7G1QYZiHoisnuBXsJ0y5XUhrBCq
rIke+rbVLoqaZCkiKKoCCqljpgZvD4l6kJIMN1zquVibSdm6HklhJSPJ+oLBjR/v9FGsfh7SSi6U
0cJmvIrgikvlvBDzPvk0Z+Tiq/U/SaunOuNVZMpncyjzv5bdnCC+/IS0WwjQGPRQqPg8AGDTYxZi
Nk1yqO4IvzuBSa1NKC7XTW9aIdER7TAv3A9urZ6xWNRo5kO1s0/DzgO4eEORggqoeTVxeL5/eFb/
WpsOhLA+CcXKW8oc8fYIGkyrdDAnQnZwgBlZEwyWsp31b1UzcdlSZGH1PIkQV4e5QU9a/NhnpINL
H2+FOg1mRI5LqkYFJ+fNKv86I4yKuCUfmcwIG8Fzt/6LLQHG32HFUcR514nUXNqxncqVw1qhbUek
wkH0YdhANjs0057IKjgR701jws6vA9wJN11Uq3LnbhAn+hhn4fQCS2DejZ+QfXIXdjMPr+wTJUIA
B3CwD57EWw+Ey84hi5kjYN+FBY2ZKXnBcZgLTaehYkRWF8OR8WOr72clgU5yVvnVUEt3zh+ANyXt
hDdL0zSYaSzsdq0IYJGKEQ0bpYpNoNEsxisO+MERHS9XzsjeQucZbVOPJwSE/Mfv/E9iWvlMB6Y8
W6ubNFTYpQdFssQ5VPfOCTythqj5iH7udcdwdKrWEWDWmcslrL23dphvbfe8iKc6nbQUuXMjaYRz
toWslHwf4lOajgNQnr4zTuFNg+O2ifM0Yl5jsPhQsAJ1tXKNw3/cNX15mEi3RHOo0f7wTROXkrMl
QO8ATjvD4XB8zulHWjY5ZBEBl1JxIVEugGMeo5oFIaOGLwRQQAmggz40fPHh/Juzfptsp/y63y2U
Mb/tQ23YMuPBj8ATXG+EGpfiTuLhQHMd1IvcnbVy0X5j62fTCWWmPHIEUX3tKa8QTU0cA3931YrN
gefiXhWop98HXt8ih9jUTfYgAsUsdBDm0QOzYju8ynm1J5RLOFGfjA/B+s9wC2ecePceh94C1Lov
OGrlMN3QdsozRYxx1YkWUclkP9hlllpAmCdGZ23lfVotTDAIeCHhgrsh9bi0hx0CZw4d0+pWCCKQ
rjL3yi922CMSRkp/ZhU/JXmxwNkKbMx5Mvaf9LaLluNwO85FytWdx0th7TkYcUXPzOeBdx2rhiK1
Q+o9V0iVdgpQ05JJERCt81TYNn9v6gFL1aY/Peas5Fw4o34PwTwB6Qr0CzDpQ2X9HnwJepZC0Sd7
5c5CiSFDUyU17DVI7/3vR2BPP77Gd/J/kwHZ/l3ALHYm0a8xwnDxjYZIL9YywZz2sNVwyKq1TSyQ
wkiR1jXmvCYagiIXAJouEJi1RdF7AHvO5yIAvYsElEc7rReE7sS3WJWxZGiq5sRspSVz9FfCxVXP
qYA03VaIXPK4whfBTi4pQ8joXbDK5TNl6QdBjSTHwfqTn1leVo7nG1i/NYmkONeI1neE92SWGV4T
2/oTXB5hw0GfwCcrFR3Pe/V4SqJFAdnDGYbD0EWCTGQH+QfSymvdgR/dST3zZGWRkcmOZKP2URB4
D+txs7FQtJ/eR9TnJnfKkggw/Bg3wEH3g/hf2YPu5zZ/nIAZtBzsd5TJOX9vZNBFMI160ZqIZyCo
JCqbGLK5k4JZ65wsxz6Ghd4MvV8S2hWi4n/tiA+bk1xYaYq+pzdId4zZw4VKBvvTiw8l0iH4bB8+
XD43pZaVnkWzdx/NTPetGOq5c5El/4eeMFl83Lb9bKeqtMF7bfnoYPu7CQ2PwIZgvo2TVnoGqOAO
cfQbgoyWhAtKZwMkXJ5M+cOagr6GG1Ymk2YvyWLjf8N/QxSTwt8twbWgMBsqbSaQZUWIMsWjoSvw
Y3UQkYhySoy4RQxRtWH3qEDh2iTPsnlpLBSifCnb3itkjTSVaYYPTQcEdRTcgx7LoYuA+rRvxy0n
3cdM1vHyjmObfQ5Toximxm4QGc0kFWbRQjPMlnbY6BBOhqxz92GfS20ZLcUhqZEHKQx5XfrYcJFh
3ax26LAVw88BMgotuBKvZs1KtWLrTHf72LiIrIyTsm0sK6/sT0JM1eh3cWS/GNrBfFuznvCDFWNL
CeBtDs1XbkAPMMUU9i4RC4WLYb9JTnMe5WYZw2opu9C4qPPPgKUquB8mFGbMBrlN8X75oYMbRbW8
0JatbZAlKuwB7kokrTZhUKykEu0AqrzVUNSOlP7ia3p9CLKMN0NS0wTRBINND6/XqCg6TexzTUuf
F0Y0n8UzruOGSXYe+VBohycaUNCoFdDxeDSQX5H8ClJRw4Ud4BTXivAGfh9L8ovFsSmp4UWdO5u6
3XOi4xekQnlCsaTRKimXbkImq81tqFSd/TbbNbhkj0JZNqMRBEAJWDk4k3+j9rS1MP9t+DXepvMS
bwvS7KW9QBG20avOgPiXehYiauAXlDPsG9vaCK73VWaUplzj8clgSKi1yoV6z5fmvrXYEuihGg+9
njXIU7UINX25YkYbKEHq7kHsePOvVo3YoHSQdy3IDtrNLra0TOfMcrIjCIf9oPNnkJQt59JNdmPj
1QYDD0+jFxKk7pQ1bCaXXPgqLklybarIggPIfIMJPxmnvKVAYvNDGFgxwToH1wVqqFBDOL+xxRsU
6P7FQndzMsVrICV0G/wDFlMOsplN77eM92h96og6ASpO7k7UuVYHDG7lsrBvHal1dLlfTlqOZ9aw
jOBD2M5/j9WvzNQ912zxTd3lHmBEngxdSuYH4MfwvuJna4aCYmvrqXayTYAMRVh2Q5Lzg2hDWmwA
2a96sKddJycaXqpcwqi4FvlCwNAwNjLc3NtuM6+VPZ+5vmAZts5w4Dy86TlczZSVXL98CTSD/myu
IRVdGq/LxHRBJRZSqyEIeDve1UuBLXdEMqePIx45lM4tEnY5d1XNjN4lHqZk8U3Gd5e2fk0zkvbA
RMZ5c9QyelP3p4po4djWjlpuDOcOgC2y5A/5K+9eDzMwwitwnMmvJaEBS4+6IuPiUrI/GLxTjadH
mBFtEu2f11hFL8KmDXWUtk0IOxnWuy+yTSpb48HDy26FsMTdG3NWqPT+9zQeCbduxbeBn8cY8rmK
gvwIC8aoaJP2HL2Djpf+wDwOuIULSzLgT10TB7nsFUrTVstbhgzI46wko4E0liF1kWHpNJqswlx+
YfR4rZcYIPgRRYSG6ZXEiEVorACTbX+MO/CoBMw8JnAD2bnI9hg7oDMrRi4V2H1B0ZbmO0xRHbKB
JNjb+c4GtPnacLJRUQV4GHaEf3txlBKzuBTM0hK2RF/ElEGFipwKp7e4fDSmKOneEfZtQebpGW04
VSafex1tSJ7MRnGN74CoV6+QFo7w/7rBDz613JQI+ivInQdP9md/I6FL1d4n+QdP1ajM+Tvu8NRb
K1SRVIzDETKKLsKkTVK2KR7XmRbF89qtbHl3gOvLKgSHlUp5qcKknXTk2DpH4KOxYT/DQB0UENPe
ydral2zJOVInDaFEUxR6lf4TqdMFJLLStAQ5U8Bb1ExzB/wSK8MiBsGtx35I5OOqyeXLz98SvY+I
7GNQVeghFBDq5u06KW7nrV9UzWokslR6rre81vwZdAsUD9EKh4YH/X75IE5z7QxT/3fMDNEyibK1
aega4UrO2m5HBif0N/KbXS1/HgNIYd9eq6JdUi/nQHxKN84NtXZzJ1WYOP/bXqD+FGdWrsBVg122
YuDAwbono9PGwItBO0gflNSKfV0TlGVTob1Ik5eoTFPk0W7J1VifkeIxUNH3vLu9TvzHHZRzzcKk
rOvK6xiNLGPFBHJu62cGDrdhVto5lNKA6yjm+DYHo2JmdUygtuSUZZQafGwtjguSbc2RP9NbxKW6
Id8yYpJPhqRH72FAP5djEiC1HifoTxYUT6fHhUiAC7pkpG3V9ZBAehBkU4m9+V3m1rl03hZfp1gd
LZId4sBreDU2vUV8wVLQTT9kEBWlfAcEtuYaLxyQxtArGxyJ+HXWZwDh9FrfV3RUTjCnyaDQjy4F
D3xIyNj7NNx/Ra+hLl7W+AXyOsSf3CpqZjT6PqOrqv0+KlR+SpN2kg9/G8LrBjCJnS2qDenX4+N/
oMypQJdFhCxpUUndAVqfwiEawUqBdiGo/FAPEJKTObP1W8sqPZMehvefWPphy+xcmGXDkhbMnIqi
VAvLE0wjpHAnLt+Zd+eeE8SMGEQ7ZSViBDGON7psPnR8xqgg5SmyobAzCupiOdP8H3BhV7+v8BeD
R46aihHYSGiwm1/DnT7K0FdsaLBxa3XM8iFWkmaUlMOnW0NcBRy+wgqWVZQelSjmbWwh2WLL8MTW
6FV3muZ+wD/+qV7ZU12OojzrHK2EoALyqUN9NPvbPGKGnAg1r+UtX4rZR2KAUT6Vc4l7vzEOHLJP
n6PMnN3Z/5zCIId28KQXje363+MlJeQDO4k1aZEftI8dVYrv0fWlvtHZxJtAv38sjb/81+C6qdcH
TEOAi3jVMvKw/87+8VRu7I0OehEuKC+NJeRFbZCa2E5I6+Uz4xYk+J6pOzk+LhVVv841eYJfICFw
m3hxfOBNjqMp4JLbGSdcKR7URsJfN0o85tc2SP7H1Gab4q88HTMaotwL4oVm7b0HSI5N+s1/SvRO
fX9Uxx+Jgum2Zs43oIsWzbop8eYrf5ooOSplX6gaskQZTxVqBYGKUPL/j9pafI0UOfdBE1xOUi25
1cAMf0BgQ7R+8Hlm0o/IaHDA4u33IG6fjf1k+obyygMstsypiy908xm4kJFOwy4h/txBEc0EcOed
kuu9tkhRtBEtuuGXFa6vucfFz5GwwmkogbFJt7XwEt7/ji+kd2dERTV8MJFe4zFwroAeTrdD4+sr
gNRbbBkoc0ERDnRH3/bXFPjMlAEv6D9meqFSb8a2z7sy70cnVgMhKUThWv5T6iFBGvN4Swj8fHOE
O/J4TT0wejUZ9fyHiLbjo73etXUwZlADccVWmeM7SxQeVNu5bEDEw6wLUsX7AkTQqvRPeqXQGQ5T
VMR1CXMSG7RG6ndn+pAmHl9IfkEcpXJRAQ/tNasAH/gRrqj+EM6MZ0+Miq3c2qDGYOcaBFcrvSQo
4Fyv6wjy2m20z/GI9uUcqBPrAWtzvY9Z1q3E9NwkKWhLLbp1WSIP2MriijD6DDzsF2yqTWpDQR7i
yniEtGn/mROna75AZBtXvQ5QfvLNM945VjvcbtYdwePuPTVmmmDUgxvmXBJtMInkYv1baybas/0M
9lfInPS7Q68HJaNfJmRhGrEMkUoTOc3JvTjkRLS8/qPYjMd4RQ9yPEaKnoh21aLM5hIuPKTKS7eg
Vz/kK7kEiBNdB2htS1r4JZ/YqFl8qI8l5ADQxrXAvmUZTA+E1yBNu6b2JPGyesYVtN6v6fhbHQ31
iy0TPIZn1CBNQ/BaqcbAyxiEWBNXSyqJpgN9Pk/Ma5WQcwDhZ4zyJcEQmal11qOR9/DzXsJQXtQj
jBrFutObKIYvxZ+91HFYarhyQac8c/7PzI28WDyF+/WOkgUKjh3zYKtGK2+lMsiuIPcTrf8g7ukf
1xg/e3+zW+8w93xFBGghQ1oKxNao/enJ5OMSlW3sz6UeFjAVM5i0BPnamvU7GAzDy9SE9V8H67KY
SskQyheUuzMUs1hwuH4GN3bk6kHRYLEP2ZM1zLl46EqrJBsi/5vj3aGsv0vhQaN8y++WeKJRlo2A
EMaU52iX3bZU/OdWwjlUlan2X3ksofqUOfMkCIiCegPDGVEO+4QfXAc66Nhi02s044FhYv6P8vln
X9HQKhHqoDWkz6IZ3HisOnT8GvjXaR1g0euPvtaCAoFffFGfqj4rMg2QPQn/fwtW3YPEVxPjPLNi
K+R/E0MxRygtkOdvPwCo9oT9DZNOwG6wFKF3yui3Od5mlt+QeK/9OjiA7BIMgbJq79b0HM35Mwj0
MF8S8Nhfoa3V7Bbzwu9+dLSDmZtwAJSFQRJqjCP6Rbof+C7T4/kja987jB8LTcuF5p9CUwolZBm5
LfsfZbJbgimPpffnozixSpH/RB0kvnUAwPrEZVy2ILICbquXURGSHgdAuE4ttRUZcCIVZCwT95cd
8wT+rRLCwtjn2rRqBqDh5WdeEusaJVHeWz5lZVhx8CcjWVQmTp9WNN/NGtgF3ErgkFzjGriy9dTU
m4vgpraT/fwfnansbPQMs433+EXr6rtQW+uYwhSUdmou1s5x2nnEUDcpozbF6eueq3po18VAAiKp
qRPJDNZ8aF/vdkhtzF7AGE6YacdvvJ4a4C97u4w8uW0a/ByoK36R86gyA19zi5E579ZFZ7EYMkS/
/d0TxsEwK/vxpcKRyiBVr7873LSEn92m0z5HWnZIhlLLtB00nlv4ecYxMq7cSftkRMd74hPaW9YP
Ri3qQorOAP6SPskxE8oIK1+a8VEAxnU/1IoVseRf1z7XvUl4HqpiRUjcmL1hHoPJgdNIV1bAOrmm
fCPRE4byzK+pjyxYkJnDhUyNGT8g2YZqq0OBo40Xy9WLW20YfRoBYUVEUmckueWAjMUmlbgdrdIJ
6wNlKy48RWYbzYxErtq65xb+ZHjetEi2LMExraFxSg516OczCPzm0cu6gMMWYRWVTMwY47n8x1xB
Lg35jyRKegKfZNehjW8ngZ+kk5fNzozgb+GIfgHxJDI8pMm9CCQUEgYxbqMIefoW70da1oqBKIbW
9tXoKdzxHPJq9ATVANa+pzkajgg6lq1qlre9TtzCA1EbQp844YsTEX7dsJsEKhoJTo3r6pAxhIKV
ZYCPWxXm+41Erd8WqAgv/JDBznAvaHl72fqPZPd5HBs+AvIUoIevON7cqFkFi5XoUKBuq7hcdaiN
Z6TsuZZib/2vX7gqEcN8fFj5Pk3gv8Exe6PYB1iZMFeUpFVr7JHEfCLbx6P3fwM5d5TUAyryHztm
+OqaqFewGbeAkGaJHSNeSmqeSmnKNLmYu+sae0hMuOhoJ8SbCR9KUrdn/hp8IP1b2pXgW6cV62AE
SlBWrfS5J8mrdNnZs6NgZmTmJInoD8RN0dq5vuddbxHtWkMqYPBAZWoHyz+dC2XJB1X9kmyZrEgC
oxmZF+ZGOYDqJ0z+tiEPGxZkoA1LoeHamgbWFMd0kHctHv5QbD4Mxj+fxHhp0fhfx7kYh0lAnckS
clx3KOXtKZbtXXrnvMJjHM52FKfLoC1mTlxgPRv9EoOfsVM8UdMn4Cw3t+M1OW4Li9WKqusjr6+G
xUDscWlwH96/atCVf9mES1VgRwj6K3T1eUAutNekj29fDZTRnKf94QLG3AriiP2lh/2xDDC/dZ0n
pP53cgkJjnuZqghYvtEzy4bVZRn+Z3JhQB3KF8mqnlwN0WhxtAvHsdxJnSw3uSGfxXdomljLM00f
mBHMCPvgTC/M7baKkToThPzH66nERK7l/llprkWC5/279qdFBht/JAYfQXZDofG8oUjGLOY1jLVO
G01tfoY6PWbhUzTe20u7/xHgJoIuXx2stx+uGoCaQK+/Ha4iX8dwVhUfILlR2rlUE7sBOvNik/YB
q9iX9WuqOyW3XfkfyssrJmo085RJoLJWRwgoq1s31G0fSiPhpayIg8vkZSvs6Gjk0Cp9me5w+jeK
T1buSn9BT/3ktSLSttivaL/kkde6aRi+5gPY9pdRQEdwpN0hHlG4abf95wIuhSSmQnS8BbJxwA7y
A3uZnRMBsAnUENIffl982BdpFGlCAxGhjdQHnWKUP3TnDv5RqSMFk/xD3I3+ffNqeerLmNxeTZMR
MJMoMKHt1qAsd2j6e0Tn/iJQE7e/+8NYRfr0Rm8FX7giivmWGslyc0jJcYBPp07tgsAZtJw6yiYe
0j3AqfkD02zbKU0/fYqVkgfpsSoYTMVSO7WBTbHpAcrCRQTo7/ADqM44pm2SYv7hC5BIAV6XTPRn
ECd31GHhkRvTBJ0MfreuQOi7ApuJdZzntCPmuPtkfxZVQzOnZU6h1DIlwfJT4FpA7D+OaYehLtij
AKSponNIAOwnJsfnnE8a0h4S4x+0dLO4TG+Hw73cNswjSDmoz3aDXRqV6Rn/yL6k/Of5skSmUpRE
FdZ+YNBa4TfSr1ra0JCGhhMyo4Z0Oi7YN4U9mxVwxnsIaKqi6vur++gFr7cLa9YGk1I/1dG42+Bj
ALXL6X+vorAf8Uu2FtqoAuXKYzWSNdFfAHA6lRYYvOdwdAxKU2w0voN/dqivrbFpBRnhFT/Tl8MY
L0oOW3ItgnKvMBhaxeXAeBIJLNl+pzjs/u2LsJh5ueb7VmDVQk0XoP4QvyE2WIzr0kbidunc+zh7
xvSuamDD6k6PCdUTpp2sGqv8X3l87euuEOT7ESn5Se3tJlTAopbVXNkfOSRPu7PToUBODhM9kTtv
PS61dPVEq/InCwMxTTWu4W5udVBbMA2XvBJwZSBuoVK8KEXBgIcc0Wna8GOxzy6uDe5XTIo5BbS9
m+jQUSt9yFk4WtogmTlDN6yyWNhJSHnibjtlIKESTQLoyV6HHocluDGpFJFXECpxbimA58Wqkn3K
FslJWthvLxdAUUihfAH5tc9MhjIQ60eZI3ObQrdIL6VnoycN5dCB7/mAsits2S4uq5WFxEo7LG9N
fu9AuSUDwArHQa0oueAz+nDReIirjGEu+Lqix2l3A812PqS6y4DiehjcgQmfx1VzPIJRMfmDBMLS
8AHDBqvJSzuAmIVyqTZgMqzZxiYbAbMOvYTFT8Gawv9LTSvbrUGldeqvMeUB+cfTzR2zu4LYTBzI
XOl9oPs/Nl0v/M1Vug8IwhUVsQ7NMAE1fEQ2X5ATltKL0hBCneTIBT1EBg4939ANC01P5EAfsoo3
a3X9tHNGMEB+AVmgntTSB/yo0zLlYMkksL3oz0xU1bUKkPp9rfDjhoWa8JV8JreYsNnSeXsjb/kv
E3gyapfKJ37BdTOMukc7NmKDy/DJ8XZS4pb/kni4uX4w87fzadOhiyirw9oaLZ8dyMURafP+KBRB
X4sCnPfBmq2dZMY1NC9zYGYGFELxurle5fAJoOQjyg7h9rNtmw+GiZa9KExKNoYGRgE+ETj+GEDK
t7+q4E2eVJCy8Gn/6FjMfQaWiphwxikKsUuSBTobX2Q5OvmTemIv8t5WrfNMHk/rmZnjBL9kTVB7
FSvwOrYCBCBeDB0z+H/iDeY1jzPnI+3RO2xqy5DI/S8b3MtapVQQF30xN/Y/rfJ4YWpL+Z/+yELw
CF7VzASDsk+u9ZcOaE2LXKVJtwbn+eMgagPI4zcVDHU0NhhGyUTwg0uRrqEN/7jGHJ2GFeEuHRth
vc7oZau68ifcKY7HTdaHm2GW37ZddOtwxT8/uqHjj3ReNysveG9FKQOfN/5thUu9x3vSwlNd0hQY
GKoGl+0hIbhFuRWr9f6N+kcvKuUom7me1tTVIFcDrY7/bEEPwsfYaxyAp8AinIHr+sDQ0o9/8+cu
lM0EJTGboxe7tZ3s7PsWHj/SRSsEZJmNv1ooSnGGhpdXrALqWbW+BbpK/fyMCu9GqpS4y0J4l8YK
IiuLpbCvxqWsbNumYxiMhTYola3TFhpTC1w66u1FVyjztRruAFZtlCh4v9mgYLxOYCoJdcQbXJpK
Aazeg8xZrFW9QAKFcVleE53w7R/tsTCNa4G0A4x2Wq/wv9nMvSLLilxhJiRkVkb8oVtSXqZ9E6LV
hjfxk+XrSDpXAugKuoHIB79zPCCSevsbAvALJnqV7urUH+DD0JoPtG/aUWQgeq4GCJ28aejJdBlL
WijgtPfBwvnhUegr01LMX8MkDtNa3FmTXDXJJyzsXYQpdHCxcSgcor2inxdeAZXODwXFUi5XG0dl
3oSIl5LhGF96TMcv4hSDs4crIcTMRB0d3LvuVCM/Ekoh6eRhruvZ+F2EHpj59/CvmCnijMLNW/Xj
X/O0az42qhfg7WbzTjrn5c+dRIH8LJjU6l35qQz068UK9tmtpEuE3ycTfEneebfhnTNQ6IM0lvDL
VlcJX6+yGVdOalLvW9v1VkvXprpY55szT6TscvZLuuGMTINdvy2+v6UytWLLIF1BWitd70LkSqq+
JMeFV+85W0BLAGFiVib5KGpxn2h1LAliGu6H8G2/7Nopef9mRmtHc01DEME0MjhdMI6JNIwvLdbN
zAWKfkz/dgEaXAfnPckvD7UFlBUel9A4YNxZn9xCoWYizGS0s1CbCz9Ybr/pv/YrOxuSqlG1FuoX
behy5lAr3sBmN5nIivKA/zUPtATsZdFHpRWkvqMnv0II+wpOpkiC1sIANXc6IdsMlp3u7LOdbL0H
/wyKFI/W1ofWRDdtX0eHwta/LxlwaKKD9vLzVJeq3deI1Ip0GvXZv6R3uwTYZpHKIiu7CGyMTz5v
6Jt4OwUr2zxtXiBP7MnbrnrZZ5T83FLZzTHKtnzjX8eDV9iE0n65w7T2pV8qTLevv5SQYG3RCyAP
24Vbv2yrbwXYKyHBDffqdBIaTWK8BfB1tziwdnDPmwenJ5ngpZs1w8pMNgy/lSikt1V+K3gWTmFA
+tczSmxDeUq2vvSXShmTFIfCSenLbne04q0i4VudsH7w+dG1hU80T7ad4OVpx+koaWn8bvL90w3R
EysQrAlEdhz72hahUgCifyTyn0eJEmDilpWA0RNgTHRjTEH80doefd2vWCgE0mKavyEeu9xNoSnc
LjEFxr9X+qrC7NacrwwYHAugd6dO8IGi4rhlLxkOfu28Bib+K8o28NIj7wHGtu5Wtkabm+B0Imic
CMAbQEPOEErxF8x535F6QIjKDqZurGLsrtAXEBg/2yczNu2L4jEpwEgTGSY3J3X0Ncv64w8UlgU3
yzm+Ml4f7qBg/4wcqP65QzydfTN5jVnh6iyvFb4iyuny+rzCpbXMI4DMYdTk/n3YlS7Tx2NwsPIC
Sbt3rlOqqJS721q2WiEjvmh+vH+O6w5DKU1yfg3gXTCGb6JoZ3CvwY8Zws7y14fM+Gjv9w2/seLy
/Nawq7LLagfslxNa2MuCcy3mQVYuqEPcQ3WYpRYtZHpBvGpS8Rnl7cocbXRJvWQw4e5a3cnGDYEx
SSd8ZJok7fCh1vNQkLpRaBJCj+fU8vYaO1F+RRjisLXxXVIk7FELDItZugpHoVkEvSIGNQIiPhdL
2fWy0Fspat+FQirp7YLxPwzMl2U81DWJ/9eCbnIS+HsXduosmIFIEeVNYjeak1IzV3VVyN0fJZQe
JQi3QaO3reKTql+1qDjbAhVzUfUju1lpY+EK9rBTqd6wbFOnPL5szSKTgS9FBOhOFIeU2baenW89
uwkPS9SU91ctg8LGrKHkUvUkRIVhiFfeSrs/wAn5b4xQ1ALykQIGShYm0CBeczSTsziv+Xqw5sDl
8dDQcjxWlAwy0EOighvk+lDaPbV1fA9tPeYzQ+SSuwHG/a/5N669VpOB5liv4RriW0PgNiBRtXku
VYpTuatINDJbh3QkImyXVrFF/AsmCRxI9OBMg7f+dDoDi1vOUQ3XnpgebK2/513Kh3iOyFSjghRX
f+5p+YIIHR5kSagA2FZggd/XdZP+x8fLd23OSyohoAqGRqZAKsOAkZukofCkFSiaSZQfAvLWgp9Q
+elYUUFoSkCMi2Dv9mTU14nvuSxC2/xUTpQJ2q+fyR0STuBs9t0+tfahJF1akiRkCxpgPxeGiCTV
p3VQmPPI+BnJ4B6HQlP5OWslMKA1A7CDUVMzuhkNb+QEms8Cyg/WKq8NPcKyPoA3lG8cb+jVHml8
1hHcsm2WL6IMc4HPhkt7L9FRaSHnH65ytdIUEfGvQwYA4QVPKcZLLX9XcvhWWCGOAmDTW/LOizeW
J/jBcZyqnxZJxeGDk979C7jXCdP9+cYkI3PXt0ZeAigdKQ2WslGanuSY6eTvqVDPdynTi1W9UEel
MgUVaERdNbySe79usMHCUXiJ0N75JAaYoGqMoK0JYqD3W1WhbXU0ck7gatMXxSSCFXaMjNh5SqlR
wkic6XZX6Kwt5FVZZSkbjENy/0D8B3KH6trchexeffPf5F4nLJ/oUcaknJD9ha+6G1y6G/YOfqx7
pKlH6m6mGOCkyqFtgHRYcadmIEloer29rfHv4T9CyGrEhTLu9z8idtIawnYJrchbvWoqkwx06Msk
3cVNIZN5ZMd4na0iuPqux1w/yqGbir5x+NRI5jOyZ7RsLFyi0G4uyfg86CEklvJiMnpHxIXYFDU/
cPY+FQTo4B7+DiOyOAwEFJFQb/b5MTyb5coXO/u6+B15TTGcA/G0FLB0t/CAyBU8lwtTcXlRr+GZ
3+JGMR0oDlbXcjQ22FdtI3Q13ufgZ69M23TN8nbY8TOz1CmW0AwaHFqUS3QaqZrmKxcG82DffolR
MEe4latzWP/B+clJGkshbaUAOKiwGtbxouPMELRh8UM8Ur93WcL3pJh/kQF23+eOB5JAUxyYuBC9
R1HApx7yF5NQT9FqhmrMFL9x+XbOlw94+sHNB7nK1oqS2IJ/PASvRQAKIkYcCpI5pnVlPMjf4Z9Y
ccUYVhBL2Luz7K1OQd/ImVHHLN0wjm+L8FvcGOeOtdmhf4mOkzyvtgLZfVyw5Cmccj6HwQ+F5o+F
AOyQ3a1+Qc2ZYiGTRRyTONjrT+XWwsRFJRzV+0uH4o5wjIXvzaXsd5JV7o5PmQ6+ytAxDwJY0e8K
Om62AAXdXZ5CgEOY9VXpajnwANRwqlfn7ACc86Awpp6gWsPS4EvQoLSLwZq8/M1HPcnEnyVqq2Py
et9Ed4X7Vhbm+j215PaFGszJfSLrkm5KXhb5L5YOuDXp3mxQnH544VOeABwrEZufS0NCbkEUy7Eo
XocvqTIqpNaBqdnpo6MVz7teF3mmwGxHvUE9JrP422k1rgkil+f7YS2j88Soeo/yq4AmFvqcvh09
aGzcgSJbEDUmx+TqTFRkcHFxFCmIVC9eZw8qC+VPtjS7R3VkFisJsUPMHZ8G0jmHsrfXiKqIQXMM
BN1NuraKT7Glb+NVC6rSYIGjS9QBTUx3ZvL9NKcb+7iIDS4oAN5oPj7dh7KJqqkm7UWgcfyXlaFp
f7KLi/BYQI4kWC7AAJSt5sgypm96Yv//C9F76AiH9/vE2O5qHJ1H7l6hQUazusyH9DYKDPEpph/S
3UgKmu7oOuQWCyLj1UlljQCxfxNlB+VuHZsAj1Vzq5WBgWimGEY1eEZcDEqVwNN1DTOM1G/7alv1
qDicAK46kDPXHa812hgBjDX6T2qcBr5oMY/UE2v7QiaVLxOM72lrcfIEoXNmyibpm7NvqjCYrzCL
omKrzdPizmjRm9eHUfd1jSKGJz1M0kpK8I9N8Yib7kbBXXc67BdDCos1F7MDGOlhBDLxGuxJ2Sj1
+kt72jFjWM0g4jKoWOr48CALJXxy1UA3I1bKPCKz1tQJ2uih/BfdjF35yM/Ut6PfILj6bsO1il11
mL0SJ07pHQ/XrO1GGNNcX0+ckmLx4cwbIBPnLOKy+d3VW1tlxHMHWDfZlgjNp4XN/kQx2zcViAWn
ZcGo7xkleD36iQ7k3020mGGuP+Q+WhNPRGNbc/C3+XqSrR73jpPn3pDxnFfBR/pBwejn8YIOts8b
CV/aJg9Sa5W/+BAFvTtvVX3xdu3Kbo10I455L8xOkIkSrJLO4ieRpSDnv3ZGBxUfKePsspjBVgS9
NeQKwYf/TDMzpGvAMQ6Oq1eCFNQnnv/MKV7u4/IGx3vrG+nRCshRyD+/vSixizB2indmk2kXRwKM
RYWy2kWKV1b/4B005v3st0u8PysXEPODghgESSpBZIG77bTGqyJvrrnJJlRt4u34bFU5CLwlrzNf
6tTv6DC18myuu0LiK84ylovTRf61LAV0PMuDlHv271/0yplKuC1twvjPWq/9ufWoBRlzlTXuohxj
S+eL/vqe2UYww2jrW7gUQSo7VOXKjnylBdkrpXaie0EP9s0y5fDUW07IMbwxyu8gQAWD2Fy3/PM8
lfJydYLQkWZTogRogXzEUi+dFYqHauuT8lX/nfqny7o3O7zarHD88KXDpJAuY6rukzGKQ7YsF075
2KBMjQYuo2fAoVHY0fpznHvsyA3geCvV86wRWuiMY43GB9or5b8+mN30NfQ/u8hIHajNoolM4WSd
RZ5F55KQ5DseDY2UAp1dgICY9VQxyuNZoosdd8tbHuh002NIBMXcZIB5awcPUko32maH638lOEaj
owM+BICqY7x5wa3cmBa75SQCO4QpWkzT31nZnxyYItgXkUWFb7HE+Cc4vcSNwDxuCFlpd43pOIIE
WcFxB/FP4cJlYciO2GjQv8PryJiufQ1nwgT5h5wjIs1VuRx0DgqMQp1B5cCwIAiMyLEyDxerNqLc
RFU9HUxvXXemJcJzpAFF5JJCJUFO1kp7SqrFNhJ838BMw42Y1/3TAdzw6G9w80lEr2qu6hDQU2Hy
BTerV0B0RQdFdkc6QbGQZjpbL9sdHOdjimRnfT7tjab+m8P66IhZi32MORB6rqbjwlMnBhxfKY7K
FfWCusn53fDhMFbwZusZ3/A/6r6GBgJMhXMfRWAZXXGclNvEiWy/l9js6LJUypOfHRfeZlTvlQFW
4wnXI6ZPcYgjQeDWt/1bS8ejBNkwf1BdV/VH8/7B7+3ERQsm7jE9JbveHpOJhIHH2ub8PNJdMgXs
WMDvOrLe05eBtdof+VvvOiO/ZcFIdm+XddZfrLP+iEr2GAACF/MJxpesv1+GutCrT3ZFWhIVJGO+
Kqo9Si4y8MTCAhwgEnaHVM2WSRIhmUiwef2O2gPlSYEKBed5K9BKCVlSJ4/i1/zw72JoiRX8wN89
M6OfYU6JdPdidtqdg8uKL6/YD4gTcj+o6llRminb6W4vGyZgRyTqnmDkJExOwrDRryFSFr+fdoDB
qIftijT3JUPpFfvyUaWUrewc8bltXax30P1T69X07zD5BLdw8M4kO50JPi3QRSNA5/IQkEkH0rrj
zc3fVZkIJXltpm+eHxdo/GRlY904RiLEwTCFZqENQgwHORELpYlTX2qw9qNndFAUNiqSEs9k4sX9
i5uk0msXN66HJBeU0QcD05JJYLY4cqb4+cIYeSBVrymtqK1hpMdY+d7xTRvFnxQ8z/fSZcYhIPMb
rp4OoAZSttfKdqDcKMOyhdXa0E7E18dabVD///rmbVHd35ybas+3wv0fDV79LNf7DG0PKmONSXc2
R8ibRybIgbtJdUUy+siRBnQxMi82eLKggtvzsrPEmigFFmdAOKw5xgO1we8yd1rcqvVZ263VJM0A
AW5DIL4At/wYncF7N1k3mGj20Yiha43FbbU4K3K0SeMChvLqmTRjPnC59Q6urJqaUPe55KjyFfMn
v8T02w2KRu3Anne0mQxl62rPfLFp2NQR5tB94bGXFkknvp8YNiw2dYi7/X0wxpue2SbK/o2JRCCa
3oWe+ZS0wB/Gblc6h1pSqQkCTwPnCKmXpE1z9tDqdm9D9aDvKtWpi2OaKcRmLpaWtcUPK2FAgi//
MurN0YdLgwFL6AfL3HFsQGeYSvc39pBu8BmZqVT0TkyfVcQvO05VsSimx+bOUnUZH2JRNSh6HW6C
dR3UKR8tCpmJtFlYFCyhPQpPjmDXlpIZqw8PM90/xI/2hFWNIjgsBFCR1L4kKbs8jPfig944bJ/0
ck5iOC7bXfQMS6ucWCsZADxGtWEQlBLY8VTyO6kPmnpqwh58f2jRf4xqikW4UFRqzjDLtYkYztad
RXpwBEKkyuhbgeqk9GF5ag+YP75BsA4OlIz65YN14431lVHhhZA/UiMt6d7kNAcIHbNTKvx3fPDq
NGmjqQq39cgAGlouUpAca/rs9ZA7pl4Rpl1do138+Uiwacc5YISDHKJIzt2tIaJW6Gj61RlXyjzZ
20IAoym5wf/+jA7A05lM3ohh3cVVoafxsoaG/NT5SFgughHxqA2mknXOlvxPTV9NOeLCfqrU8MlA
TBiNYRkt23y/tXyZBo+F+ABuT3zQFXPNSFb5OLEfyaxfUar5AwwUmvMWK4nT4UO/858lnE+mAMD5
+F8JvCY6kpDKW0EaaryYupJOl2h7Lb+5OuWE2oOfHNh/CShKv1rU9KTp9g0vBGXFNyiUeoliGEoD
9v/yI1FcZ6tZg10Oaj63voefV0xT9T8e8fD/Ggwl0LH6jITHAETo+kMg9ycuIh+qHn31TbPdrc2D
wE89r5TbyGlDT1xhM0MCdQqIot3rkWb4o9ARCLI8mUSNe+2z7M88F4rbubu7vH31qdVrg2GOC5cM
cG/Bni7qhgXX3+8jTGzbHgA4bU0eLdcPuj9DbtHv1Sp5cccZX1d0D3dwRhUpP6PhyoO+I1cYu9jX
IIYsqBQ6r8VTaZ8yzi0VC18yt1W8UxwDhPunHyHMBPOfHKz9pV3oq1EYtgqBT2fazOSsnDVRI7rk
XilW9VSyJ9pxXiBdz/uQ3iZoXg4mxZXatolFhsXwDT944SloTOXc+ql+B4ZGy3ZYGQ+DiYSIgf6v
T0BBxc84s0asfR8TowDn/iU9tAuKcutW8fKoSfwtCtUVX5sPYF71K0d9CiM6VbnskXLwVPoYDG8M
ymrPZv8lNZ4aOLfguhO7HakeM2og/4J03Uhltwy3EqTYEUM0CP7FQT0wqGbxKgcsCiGiSs1Sc2Lw
4/mwuP3TOv8EKlEQBj09OAoQBmYEk18lJ9mEim3thoRG5Lu+WS7f7dIJ+jk4Z3cMDRomhXNZZcLG
s+58xo70xFqODt+uDWPIUYmj86sdtru2wyWwczjiDT51WebEzXywKSit5G/GfBeOYpCPPFSlMWLM
lBYfftpH+uYleJoTgp5SbmVyvetIfDxf/OryohaXhwnl/4wuxPK4Wk5bdbhN0t//rVDxIs7pT85Z
4goFT4d9m0ymTx8hMbm4e3rjxqG+keVYaqC08eOJo1P+dqOdF8VWZ1l/0PTB2taP96vp+lkySotH
1wpJWkXCNaeG/nJUBZ6+LpbAtrJRUZYz6AaZVdHtyzCTmbFUyyU9aoo+fkWabzRJtKUVopDPqtn0
SQy/hSIq+CM3RSmDu6/Z0wglQZEOevmucbGKT6phFn/xLe9DkUZ4zNo2UJGM01eKOINZyrmDY4hP
Oc2MHM4wOru/MWKIjYNWcU0QJ3R9k2qilWVpdXGh5q4anCUj4sW6IPkaODQAJTJ/RXWPKZNjFlpn
r2LGw8LZBs24HT043EhEmgxHP2pgsvqpVDtWl+m0a/Yz3zGl9CcfIQhFnI39G9JRnvd0A22boJ6y
Dz/+Q/Ek6gRZfrT7o4lRumiC/OS76LBiTLhQKeLFjr/wNrjsj9FlGzNj3wt7OBlVwdLQNLPlW50G
cr3JfjVESz0p5gZk8lFBNGV3bAfd1mtfuFX57cmJm5B55cEvAcuDKbuKfo5oMg+Fb0M+DdRXWV9h
9AGHub6gjhLa6+jwVsRAP5sj6TzIeNB3yIeNklOvVPqFccPoKneNcovjSOEWDoI8ChMiPzIYHFFf
4c4STm5bQPjAUEN0zve8ub8ToXf/+9+hVyUI2iPwBfe1sZXqWZLS1Zlru7jz4sXowVUTIUqIZJJY
vE376uNrHmbBOH+yQhGzeMOV+0ebgJcWr2+ZrkSCOCc2uEUPQXe+8HFw15uTlr96PajPXyahw2jG
JvRHKp2s2d+xU7iiqmru5DoVLALU0SNadiE2E7lCC66vfSDVb6H29HxImS6RdXGDKi2SfSs7goRd
cyl5MK/SrmT0Y+Cp8Je2oaHoyTbFNkKQQg9ff0kjIYGJosq0ngOcZ7KLQWXjELVT3AaG9sCQQb9E
TB1HeGNzNzg1Q2CDrZW7/osKKLeshdMl93Pbd0AgKwd4Cm+3llFBo2ZVd/pgHLSCzKPogC6LdWfh
LacZYmoZWYat+QOpRC2bK/cCSInfShavwMfjaFz18qe+/kTzhkzo2znnKt4BfWNfmNS5U+5f9s7c
TDTfNycU4SgToGUKRTs84UWKs9O0ZUC2u9yoQKKpg6I9jGY44eYstCpesAznya9Ixoemp2TkkTGD
h+S9Gv1CNPKGcnnAz559g+K9xpK3H0NY9Z3hU3FHvXr3+pOKV+PkN+52d/nu1OiF5+Zwv298pHhq
m7dxdKDZpfphliS9faGXVaHbA0gdNf+EHwU3Ey19zv2tsPszeVdVBWbb/oJM2lzmR8Uoh+2eeHlc
QK06PC+lxAxEYHI/RLe+2UZ+TG7eCkgWyM8sQ0oUO9/76ww7802axZ5egysEkPlbrpL5VmyzgWia
kcqNlx7NsoYjx+o7+2tMFmUJkPcFU0HnU5zj075NeXLClnC55D4djFR6Qa0C0mpzvbnQRsQ/WucG
lkv9sYvaK8yS85VU13lJgbddP7x1t9OsgQXTRca0S90hzdD+asnONtv0ai0TIHfRY+Nqrhul4bIA
1w0PIJuG7EW/EoxPMMWRuA3Zc28BEmyQprkt0NRkaE2+ztbHWVsETI/V1HBZecW44bHM8vM5/XYp
WkSmu+uvOlAf763D4hQlLVd2EjpyI1mt2QrxpkPdJ3cYKccTuYnLyMjKODKgo0KFEbivbs0DstIv
QYhZxfFtg71vhdqFA1Bs5VwDCJVQkfWpBgL9Ok4N8L78cFZmdxQAKo1zB2h5ux+WbUcgm6zjNGIs
hBapU58AHTn0IiU4zMVqXpzf5ePwm80f9lC7GqKUZK3upCuyOZ/IamBSFnmNqwC1mI9ajwKInVnY
c3Z7k+YggAGJB+P0o9XRvo1xBF3c56KpUg8w3uBkr1F4NTx9y0swtaPX0BiLlD0L0aH7/zj24Cz9
m/qRbmnakw3lvC9Yoq428CQFoJlP+crWf4R9jXHzubTodeqh7NmsbqVRoi2WAlng4zwtEJ6I6crB
ga7qj+y01SCMavUy62ofdZG+F8bWNbBZq433Dl9JPArLmaPOUfmOxuD69059GJhNh0/rUrtp/bFZ
vhfeA5aL2Efd1XbI3pchZ4cnSUPEpwSlfrjurx8BTapDmBU6BPQaloKmtoJskN7JB5jTkI/NQUsr
dqc/8JmgMRIFasw367Yhx7jIu4G4k+yAhI3UC2tRZ5dxHkp/HdTKotfP2pDngc2LN74jLa8Jz3+3
GpzCV7qbfT1jjjTg8IT99ng1KLJawIkwkDVKxKtjV66OPTOroQMbEcUuPJkAnuqkF42c6zQ2eRg2
o5LBM4wMZl114xcuJg4rPdqLIwgAmeyOeJsDDg5meC+vivewTDd1SVSip4/nilElsynjEITg7ifj
/8I1g3+eVOeXHYoah93uPu93prWfDJdm7Km0aiUUV0alwKY7Wi157VG4t6CS//FnDm6V27Az/3mE
bkeYK1liM21tMsUVTOnSSXglBtc0emEwTQ4COsSE4f+eZL7jixs+IfOT0/63GdQemghDnlLPBDY5
iRn6Cfyyhi7Sy+SChl4e6/EQ9HC4gCAVTINe1h/RuKG8gT3ifugm+/wtK8KpDI69ZWeeIOgq9VLj
qvNMecPiK5ViymM/YgKHpJJj0UcoCe/g6eYJOLUycxuUz57ocIh050KaIpfaJvpID5DgLoao+LZO
tbuM3evoju576R9zU9ok5gsFFKzSmGRSjXSRbCoLI8T2bPp0YD1lwSJHxRL30BgE6+0mIrcSt7Jv
DVwekmK5AJQsP2py1SkXTxsHu7M5ksrIcTin8k4znPoHcprTqJut9Jb4vsFSj1roIIGFBASWnoS2
rc8HK9B3efUqxvmxaHIh128TIaXB10QrOWWWXdmNutj3o7MnqIRCxTWx7D8v6lH0+hMWKm24pF4N
9DbGsgiA8m3VVA00EEPWtMkaNhBtRgzRw/DeZvimd5V32laP/IJdIZr1rBYSnE+Pup8tBLqOj9aE
XVuAMGzcSWgbPwGysld5pSfFJ/Kgx50NOjUFv9YQsSKgItsl57HBP257sMGIKiQZw7+ICS96slji
70pXqGNM9bFFEi7lYWwy3Hhd+4dS2nVj1HtgVFLajxsppylzeiIlrsOe1HmUGK0kGyF1hoi4BArt
53DCWg+xzHrW+K46ZI8/z08lr1RSltMmbopHedChdRKYtDUw50bLsKZkieCTrEnosoVYGdXd063X
G5qrh2N+oeUIVY64xVm9/DyBssMkO5iTxEmA8Fkzu5jHqhxEakwTUmDCQU52F0naniuF4lKqbc26
cifxDBTybHZwzozqX1epHYsLNPIpXBAivhUgIRblk0c5mwpGe7UeFOLZybGvdtKChuL4r9ZfTac2
GsR8swLw7vRZKbGl552BeqkoAi8EXbeiUKpnx7vGvYcSx/3YpHzX6iPvtsGNi9jqfVocTncIBpZP
lHIM2mbFNwgCWywdkUbVtaevkSeppRGh88Ok77wEp2USd8Xfk38TIfw8+vNZn7l/HwAPrShYzYrD
XcYQMo1MM/RslsRC/obvksij8SsntBGymEGUUOZhn4H2+W+oe98LZmGc1M8T0n0Tf8OotTeqI5Do
bR9/2pNDd2MH03Ch9OsN/hkqsD/LGXaYv6dDP9oz4xwpDd1mPvWE93SvV6+8d88O/FqbYU7vRVae
iJJgffs8L0qAppkDdwp4S0+tz9nNe+d2CBlwPQscNpRAJqKU2WpArufQEBdboJcRilrFoQVpN+cK
C95a6nayloSSzHTeRLuXhR9MrAtqR5W4gbcvqDBaw9rOFJgfg/Kjwe4e7L/v55KJ8ZtgEAuZiGQX
17gS4SPVaNoTm4W4YWyAba7IFZhtl+Tg/09Tl1BJXg84hED9TKLzvxJG9KYHvHE+H4IW2dGjXvVv
JKkX6CxOhLHfE95q2jynThkSlaF6L/ew5O3uC3WewGS6PWdN8Z32h93nE1V/s1yefXsqr5aRvCys
gggCxcGg/tETEQZ3eel+mba1ziegQjsUvOepHspWS2OzHbp7XFgporlcbq4VLkg7Q+M8LHqMmCYY
zHFZVLU5HzKNI/JJneGozQqIRNTkU/WEJnVsJ1Q7eZujLa7IDQkuOhIETF3QXp/P/mypviUGXsCW
u82o0LppnVA/lwU0/ygIW/nRobEMKYlIM0KaKp2RZwYFgdET2vVV/wcKUBYHxUulmjZPgzvxjnaP
ru2cpM5jc9U9sG7Xuyxop5DFpZ2B9lVUBkWTvHeya2+TESx85zU8EKKMT1iDKGQbl0MhFEYvT9J8
3RY/yoy4hcWGu6MW4dpJoAoOK4N3eMBVK0JAPpWJTu6auDzPBeQehUiNGCAv1P4N2W8y3sdKGgFK
WJG5/5m+xei6HzHMiIGkSi8Bj+vyqP6U9wL4J87956xLV/aJQXpWqp2WSe207nsdmOAdK1dOwEID
oXP7hywSgGYgVLlKCi91LBcavP3DCBgORp12/WaSFNQZNLKZEyHxzV4XOlqhh8ObhpPeD4zeCLkF
qzVRW3yt1oIf3DWc48zcm5D6KV4fzuaI/Gh/Fk3NHjk25vlG6gz9+sBAtwvga92GmSRV01dnhK9v
WmDZywfGj1atBpFWAZBWRQf+wkt6bbjiSZnfmlOIx7mXW4vHM41UGjlHeKCzdppg4xyeGsMRH1vs
DFQ1WYbMYWnS7R2XwzkY0Q0gyuCif622RFjrMFO9HNT1DBNM5qDLMs2VreRNproaywEUVMleEzBK
BRrrFri2xTGCmV7B1h/6Tl9i53DfZ0pEQjCKFzVWMWEowWTl+PDQ4S3k2t5VEFSyq5dLtwUJtKni
t1QLOlk2LaIeQ8uRODO1TbS9eSjmJmHmbOH9N+YDELmdxwpWfPGAo6aHlgW6pmSzjBYnWBzlgEzH
ROXRrGbQSyv7zUzBWIcTHgq9KUje88/dqnMB5p/DiwCdsLzUWWHD584sCMOfJtEwRnU9SO8LrEJf
LY4JutFtiF/V2WAXmKsRdjWzxHc5ZTEnNaZZsNnz2jBMWBHqp/5bHn5RNOQudhXRKV3sZW3qlupf
uBjZ6WzF8DIuMOw8InwPcYurhoJ+58aEBQPSEi/eNbRkrGGagSZVs0NdWlP++cer5uokhfqzwOMF
YkNm4sQo/kCMasnngjJ7c0L29AH4c+j7w+fXMDGnTRXyP4mY7hG1IiFHjJimb18uktyBU+DkYsvE
Ep9d2GRd/404XCuMyUzKB88JTPMkkeaBHCa7Uq1Hf7sK0ilTKRwiMBu9k4Xtn6azHwUtMgWgt1sB
/6iqXH5h7vDh9JmbxDGjV0wURSHZmkO6Cm3x1M6tVnVcGIKfe/tdGJBq2wvFuv3/HEVvWuArZo6b
fgCpUoEN5YGFzfYDgxxz43mj4oDOEXkxkPI/ycNNY95/HWunTqXk02snXRe4xJDW42DTssaBxY1m
Ds5b052SQKngIxbYUWga4mOz4BfrgPTdJaQYtJKAU/KUycxa+z8+0MCEjVZMNOAeMkqUG/w4yFWp
Exq9nxp6wAIe0noUw7rpflCTyu/G4GlbYrfJIoq+iQbs+f7M8fpaUnaXAszS8nYJoVbHFyx9vLHW
F+/+dG+yYuGostKjCD+QEZ5hi3JqiuYBiWQKKnjXNfNm2Ps0UIpJF/mkgHsjb3HEcbmENCzUw9pv
PL9nYjtmBqguBYymtZ9I910tumat+xbX3wp2DzCWrblh+7VAcGdVZN7kwllVti+v1bj9oIa6w3xP
zbhSmRYkxm9nTHPiHl4mVJS9itrNGTP759fp2eoPLiUFT948/OJV+6JgR8kjdotI0S6fUKyRY684
KqNvLv6zyyaNOaSh+mW6+ZQgAmxnaolY3Swjf2AC3XkvJw39fDNRk21MkWvaEIhelLs+IvX6DWJM
B3jPobw7e6IKEFJvBpUOZOLymbKGWMhnwT1WccSw0bx2fxtYeu+NcayYV15yY66m3YM7piYVpPzK
jk7Zz6dZckh+aRA+qXTYj0HYA/R6Hj5mgx1BT9mmKvcxGkVRVbL9+dXgmcTKrxzF+hrrNfLd8qYb
bZ+w5H69E4CfcKoaWAnvTDvVs5MMNKWKQClCXdeH+aSZ3ew1N9G3vF58gqGFG6seO1gtGLibZkCs
Yf8UP+5OnR+5ycsJRzZiNqoLqCIoJXfWKqVS/avIc3Rml84AQcCvYKwGRhNEnVNCg5ITcu93haOg
WTM8ViwcWWV2tkRIra6OIXP9k5kWeJA9IlfDMTYVgLjE5Yt0SCXO9Ys5mz66eA8K7m7aiDbg9vTD
Qm230juXJtjFvr6WVvPq7TwJXxUxSJ5hTdyX8suceQOPfD+VacJDRQNd3WvYRK66GYhXYRQSoJq/
aaeRRIHoV2lqEIo01R3kFpLaUR58Dt7W0R4nhSO2G+OCm5ovBg0TPMzx5vRaUCoiLTMV7rR5W//v
R9egA2LzrGxwSkkm23rSuiLY8cv8QPmkGeyKlGLfgAQBFu+zN/itIp2+uT9SfqAQdkEDYWMy6kBp
u7iYYgSzJJXXeQwNT4jDIMQXNgMX1ORSLucUpoH6j5d2jKAeKi1OvJ4Xs8hEdMz7x0Q6r7JNFNcU
Z0ctylE31SiBW3U6mkzAHuTMto5Di9xJ/oDGGetacJR5bG9Jlj694lU2pI19GSKuyXsBfFU2QVVF
VTjxzBYMJmZwY0mYr97505biwxYgE95gKix1sqRE1WpJ5n1yLrSPbLCmB52QacsBA7AcD4sD52px
DZPxLHKdNXzMLlTevW+1rBHk2XnykZ+DZ3iA6BeQz7C8/U6gmVBCThxvxHDx8YppfmBn53p3VLU9
QOJiNQsDyatCJDnkr4kCZZUVCKAzj7ZVwDFSn/931WaAcAUqhwqQm297msggtfAvwAkmZMt8wKnr
aEtXD+XhS8u8S6QwjpGzmb9OKsxHGQpAYyeUgVSHUSkZYcikvOw28tvg8hxaPJGyRE5VQPjT/zxz
fPbNnYFMoYXaULyh413uPOpzQ5U8Tf3zgK7rIs7b6affYVBQK63+Aaj9DZPIsXzSrCf1vUQe+/v9
o/zom9hIs+xesZk7f/hvFOQ02jxufAZyH6XbFVrt2p2Fka2Wg1UBw/oAOFNOJ5r91QVFM7H8eui3
lP6oGP0KwzbSBtROMHo0XIJK/8fgPXHqSbf+ui0ep1RCyzO7t7891j/X8tEB+CbaY9Yac8x57H/s
H9E0xG3JX3eRnLC2EDkrJ3npyJOvCr+t6TcGKGp6GAt7I5TFzKpBl0BH2nqPJ2DCuhdx4ml/iIB8
eHhXLoJFeWdA8TbvTEhv6snG13ycU8vDvJpsK61g/4fN4y+pXg2VMimfRi9ENTAICZ5aDx4vCo3y
UKNBNScHk6VDEFhJK+w34dnG7ctdPGoodfXAEftOZmbeXOhW/jOfDV7YBQdB5S92JCz6eBHOQ2Wv
nDNyYJp59BYiz+hB72G55daLQxttkieEdBRUQ11BIi1YPwrCYTrUyzxP4H+IZ/g04/5IgCDYAnBv
orB978olM/y/QVRhKYMW2sQ5Ri0YPF8TALLb1P8fPut94ZMQr39sMhd1+NASU/38edLnU2vEBzM9
7GT482yzCBBTeMxatlwFbTbe6dmbf7MfCk3zFflImjBcc3SXBW7GlyewZx2Y7fGjpP4AuGeWtWy4
gNRl8jtSW9TxwDt08/CcTluLsfi6dp5kWdm7w9zGQPqJxPXoB4AaJGtdFMQyzctQmCn1LWIRf7xZ
tyDylXvMcJDVif6NlXpFuzx4BIcEdQcZfc76+ZBobtM/N00z3xXnKPT1ApYTQbcQe2llWU/tAx5o
3l89UTbc/7mfiL67WMCVH0LUQ/OGUzOODBeJwu1BDIRrDwHdDW65qXGslbEhvkFtsNWA25kvXVWf
gQ2l+7vEsnonfTH6FN7ZDohWN2VenAqkbewZCIHaGJ1ppbnnEVWs7V95YbMXXqiw8/AdGu4M5I0D
fXnRsmwGCi2ItfrPTPZQacN1QHPqMAv0lsf2Mf6KLKx9DH8aw4Y7Yo5Q56P4NytkG1Ryjex83esp
m47hvxvjWCuRvUVaLhXYEbBXqQuw/9ukM9Yv54zU7hAYzN19rARK1+QllpUbyPPJA/k2HqnzbGsh
7eyvm6lP/p0rhPfJ1lbE/JTwVJA0A6OqcHGFi4fDouC1/F6IcibAPTtr7m+VTqhL84rzPWEb/ChQ
XV4dBcLOfUfx+ADMIeLYcWlssBX4PxHW7Gd359JHf3KjZnvrbycqafRXAwcGhHuTpSTRwbEzf8KY
7+fw3PZAVxCwqnXLsNIZ0y0HOExsoK2dzGYT4+T/ofnxv4NE/3nk5j4I8vFyenD9PYuIh+QyqqIZ
2ZkpNWFi422CXUNSYWMUZkgWKFHEaJ0zeGS05SZ5Scxo+KhfPkz7jvKt0tavdrqsg27zrvLnCCcb
52FjPPGT7k1ALT7s6nsDdiOCZ+X3WhY8673VhZGFNzZXPNhCVKpc1547gu6hEctpBchx5AKQaQNi
xHeeB0cz8F6D7GSO+0P+22ROWdiCKg8b841ln/LLd319ywUabfGJk48XrKMGgjvhWwbvFB+FP2Oc
wrCUwTRpypF0gRM5lwF0/vxr7JD58uEooZXwSVMGfge+ZqAD2vK2uMDFce/7Hy38eGBHolIugEho
zze5oot3uB10KBAAIO3rzfjQiHASLBnfVO/XbtTfLQi9ugBIv6Qc9hvODLmihzQ/bNfz/gjN13tN
kYzgkeysGVgG7VCMpv5LdIB8krbhTH88nK1cC3FaoxtZLPprnYxu1oFzvjhpgXoyG7X36/ME7t1z
71fkpVkuWpBQEGkPPojc4Oplhm62lfie4piagXKZoDsWqawTuhg9xCrVofPYWbWfIXpxQrSYob7G
bMT0jkeU56pgxbcONKaT/W1pIvk+p0aT7sLoD4IlCaK21vtEJqLPvShKNhvyDKdBEBXj3LZleHbD
60/yRpLMHdQ1CjbTirze/ouPlAUrIEu84F0Niy/Oem3WGooXhn/T0Oo7q4SVmXjWDafgpmpzkXbl
TmhFVcDvvCmEKwbQBnakAihDh/EB//SBoF6hbit+ULfY6+KbX5yMVbut/nwAnuKq0FEV+oO/QK2i
2CAn99FlfaMW0xhihzN6+gWU5hqDi9IBhcQAoSKA0rQ8O/H6CLk7AuqA/AYaOFsSd9fYJmYR82bU
10tZxvfOOb79BXDCVpFj0p+l5S6ic26u0pndGpD1vKf45hssg0nQPFHrD6vepDF/D2ciBaxEovnM
+D4BkTHL6iLe2R/J/BYAtxMkcDh36MbGsg89K9wcbDm0lTyVmt7XmRwbSLtYTMLtgl0FmZemEdIi
AOlh9zdWqAVqRNFstCwqinXaMoDIkzz/CuBSKwd8UE6TDOHGMBc1wXCZ8dpiwDiUcXVPr77Vze0A
ypkYiWEYzJP3XXJi7KgxympzRkQm77UUC8pRbSvWj0pey/l8CntWquSNH1qqUW/TwT8KVYb554hj
SmYkJEzop5k8OL1MKi5n/Mp7EULOSimCYpIxkrmyN5Jx3f+qYqYTq+/SeudnW9Zpbi8LSTrVZ2gj
p48qVzCGkHBZijhQwv8lVAqk3TQn4sfEw0oW2gF0Dy13tFqqULp//0eB83Ny2IK6On0J2UIBPiwU
X1hhrGUw88QBVo80Kim/HI36gVkeFHkUQBWp1Hmr79CchVWYbqgrgBg++1K00aTrjEWOgyC2AtFg
5Xj4pi1TgCYQmoP/kdZV2X8nL/v7h2yNsU5ENertbEyFRTN2sbV2CJ24pWf5MS3W2N7oUR1xcOeO
ti+AR1N4IiTVJEM2ppid42n3Jg/lkje3qA+hgKNw72rx7c1oExpjrsz+feZP81YWCYgSypq88Zbi
rEicZFpFbWbkzFmZ+Y8MQ5bk6IlNWng9qj1jiO+4liFj4DNqk7EmxI3sQvHInJ6aUU4DcAI7vITr
6vpb8tf/msTmDaU1jA1TrAXMLXk4f6FkZILH9XvXnKUahfbJguZomEb790acxaNNhLZsiKprfmbQ
xQctZOfI0zETxPctFzSHEHdkb0v1r7iMa+sNxzT5+32uc3kLFO/pSERNjvD7ho2T96MtVcz2NaAa
3HOkswhH0u8K1bEb6QGu0h4F0J2E93cBGmHSDVTo+N0jScjIiD/Q2S+xEuCdNaSr2SW3VrQxc+lt
nK04u+xNg0vfvnRQMvALwCD8x98jy59JzOR+Az2cMBy2XN6yEfeSUAJ4GNwwD2J/k+K6VHzXN1oW
MQkw4/DuKQoBO3f58Ev50vxTPeLDlQjncRnGXY6c+MpsNY/MvqsiUDXwRSts3ey2b1f0JA2Jn9h0
/F5pKx8+u/6U2W/EBGWIElG2b4T2ZUUqjHjv2LsNyIdvXOTQ6/+aevGikfNxXS0PfouZ8wSle07D
KGi9tO8E0WBJ7JTwoXwYTyVKLxJRy+A99iVWnR/AJCtO1auqVQbGk0KB8XZvDhlsZ3lQvODwwYvC
vPGkv8xZMSSGj2xuPGKPGIiaezIeugbm//CXI0P7Hc5Ct28aG2RN36osi+xTrnmpYg3cRH8u+nnz
Nm0QAt3enuD3rcBUJMlADM2kwwBQqVun1Vjw37GFiOcZgYnRpfEwzsnPRHlc/bAW3whhfdHnWNPT
EpJCZa+clHkgcxzWe0THfeGwDYutRyVqfP964ppjO2jnGipi1tMc0230FvZKpr56HiWE8fyBcQuO
qxCpKDAdbYl8LPYwjM56sXSedIUAu1z+UK/ezogBe+7yv8dQdj30o0kVNGqdT1Db1AILGUHhjEyA
BX2jCOmrs2l6BH+8+WCDjJ+8foxDWsRPkGUf2chQvL/luPB/9rfCXs6bMp+il5/CaeIqsp8zvgDB
Xfo8kn3Hhy/Qk8nFZuDoRQAfHOg9VMF8TiJna0Vy51PbRR8KIp0GWFoWY40CBxQXR9KPRcjw3mBK
icJ4OxX3sanuZ5cxEAk7uC47nhx/5d0gmWUlNLAxcyS2suCrM5ukpuF71EV+TkWZYY54laXrjMF3
aiTY5RVul7u+b87unN/uY2RVfSm6qQHh9HcTxA/tlkAdP5o3wNesi3Z6YOvQkg9WmRs4U5wd49cH
o/Vj1/gssKMeO7Lhxde4tZUD/58pBDbPPNG8w/K2A8mw0SVn3iyskwpLW3hqOnjsi0Z1PLJKE3u6
6GvCaFHNNByq6wmZ3Ye40Jyst8IZ+35y1+xfmCHSWQLcHbIOx+wpfIYXXRPyZoynht0g2SuZrW4n
h1jx01Hj4GYlTNEHB0uJwu9iq5obDd9H6I4/lWRmgKWPKKG87sXFWs2qXFRUkj+QONSRdKX2H0vV
WkSAI2sy/TagMUXvQfG732uHhPNtDQZ6t2ikkNMB0/L/tpvkMrRhm8k4DzvrNKRzFTN6kQmPEI92
6fSZ9C7WLJgcXMwj0QmaY0OEF3anqsj9OI4MXul7YXM+Gp+b8pyUgHQJNvDl8XVGFEPp/mz/tV7P
wPHYbe3LJjHpgKzQSPttbeqQr3LB0sh2TmMOMMM+AoGQ/qQjtyGYU9sgIegjs2ipR/oaUZmRpiDA
UEMH/onwFX5w0CJCIXKheyUWCgdZXfNHcu/hAmMZd+kO1Im84pB/XWCY6As/RtaZEpZErk/bU+fO
Rfo/hIRgTi0+pzIQxKjr1q6AUy7qD3/qZ09kZRDTSKGOKywYDqF/XT8tIH8Rnmu/2sG/xdig6WDe
TW6i0t0N2ivJO0Ncy98lWPPMAeaYg8vS1rFkEO8VdA6nvgyyamVFkwL2ppI5+DZAsh0bLXM6zmyZ
vIX1hHJXAhQSIFC0njtswe2Uqf4Y7HrNp6+SU5tejdrHIoDtPf/IObq0sTTcG69KBWZnFJsEZdjn
U9FrqEubhNqnwP40ItQXAKk6bvxRaRh5pHipuPJi+6mdQJrUWursdGRvjbDlSsIHbx7XqCrBX7vP
xw8mgfEMnYczD7QBX82Gb1UdUQZyEJycktC/Ul3R9PbeknHb+JmMXKTUAsG6Aj7UMIW5SeiPpT2O
loS7eOSlZ5LkhIjJoNEIQfeFnbz7xghyk8nKZZw4eBBpC/CCWY6c+PcL3VR+XXnYSODGHDQ2WG/o
G8lfAqc3VnbctaIWb+rqzFltrwP+pgWGTP8k7nVs+lyWOqJLNuGbEwvqzACxsPWZH6/RRxP3oRDd
S8nwIJIb9wRKpyRGq4OF3k08FbuwhDlkF3dMpgYEw+xjE1WTAQG9PqyxMzBM4rCdF3a3LvOVefOi
Y6rL3UAl6GaBqizl7NcI07IHnhFxuqoagp3m9PMFUJxZyXC0V/KSLL+idmDHj2Ktbl1UbnScH7OY
VQpPQY9zO5ogENZUPpd2Jp/ffdI/ND6wS5ZFTn9gVuuKnjRN22UN1hTTxQEn0KuBvUa3UyzSnVNF
mAbAkAb2gHst5sg0sJUnq1hVV1XXzIybwC/4xF0gFMMy4zxlklAQtx0QYinNfJcFsdnRLWkVQvG6
qVYqhfUPMMitIHgok64eJmVRZB7qetwK2Z+OxJyH+09mKH39Hotujq7IHtJ/ihvduieIo+HPheVz
cpo7K9gOvGjdFP92HafG2t8G9yGIgDif7rknJldYJn3f3bJCuR23APEpE4wK0O96c6fhEvP3ITOn
2mVrRcO42gZuoSDhcFKyq3v03HZu6UHwFQJYkWnjmM8lprTktrPohj9sPD8GWLFe0wfMHs5DYh3c
V7Fgxs0DDNQuUu01HXflxn06d/kiMGn5iiyRU1zFz7A9nuW81NAAIiKpyd28ZhAilkN7M8SrmOAh
45LoaoD5XsHpCjLIebzsPN9MBSytgnT7pdywZaVmbxXvZYJ1TI6FLFWCjqfcTH2YQS7tYxKu34OK
myRenLRaB2MYzAa23DBEA7BoX8M4v8bKy6h9z5ELP+LaAiDyRChXokLuqDja3tE3q3mrnGol+4sA
PqplHreExYpFI+PnLUoB9D8ec4GiVj5rzNn8oUS+Isg95WwCpdOP6IFJDKSz+px+q0GzW7qCtrk9
RRGdrDwnjlrBf1CxYEjDRIEYNh8FreUV9ow8VonION+zH7yohAnFbmOU6+ZuHxWWUhBevD9WCN/4
07avo+nwR65WIkEX97k5DP5ScJ+ZkZ0ThZPGFK5mt78hvy69DgjKfrMcERzZB9P8Niny38BEKq4x
oRttKROeNvYOPo6f/ikYFu76iWf+4Uvvj93jhXLsIPg55v9k19DolJpDmw5Y+JZhOhI5Hisi3CvW
mq8FAYwHn33RNGNpRAvJpVJDDY8bc3NuyjRw6uxlkABhcV+PRt8dIR7SZoSsubPDaNpRYkUP46Y2
8Me2ymWIjYHR/Lq2syzopunBM5ct7fQcws/3YM6tknGtFI29/blyJfA1aBSrbxbn5NzUMRmq1Kup
h+6m8UV4wHMZrUcAZ9tuChJ8WxofhYefn+zAKocUPIAY9S8GxFiHxPCkcOCyoyOusoKoA88HXLSy
nqvzTSmZ5gpGrwnpplYTp5U9IUordJB/msRTKu5CJyPXkS7ID0u0Oh2SbcJYhMqt07LSF55teoBh
n3a2krVKumYkt5tj8nexUhVbTrgCo9Lpx7EIsptj903iD6rIdH58ubJ1tDF+lMH/P34M1MgNOLfx
XWZE3XOyQrzEU/gcJJfhgPcEERXF0CAQyGLuVfOzxCybFsZCSNw0GeivLZ5GKWbwCMJnfOi39hzf
EIwFLzBdSF3WlJ66I5KLkAxYNxGBOjNAGjBhYuk6pMoJmvhXBD92uoppOqREgo1TBqkwiKo8UUK2
tDL/5MuEW+20nHRyyOmKKO/GQWgE/qgpAgTKSZV78o0jSLPt9ieWAABaQDThtjQLjuskMaSQB0qi
mx7VrDwsqzXJIBdAPmDmFfCrsg9tIGQoo7KgH+XApEV60C3XwrLTN3e1Qs39CheOTPEdY3O3M6aA
nUHoYA3DGHRhmltMq3T7t8OVW853SGnBgXSYi7QV3szp5b8z9uk+3yCC8KyBKPBVxKPHWSiKrIk3
ZTSJ9ryolHgfNM7bl+wIU2P7lonFciB7Y8Lw5SYnIZknW5NqvgRwaBssO14oQR7BtsaKjr+vjHec
pYnHo11gfWwExGmlZBS/1hQ5NNHB3ZDUk4M/da9xR9ubeH79R8ADtlHOa8oqjr3EXMTnx+6b2nUx
CEAJYaFCxru0mkWsigPYJabqROzsyTU2i9CW9I4foGhS4975/fO7G0GBAx3qpRLD0gNDCwsoaD+o
pMS5PZA6iis4Ke9Dyv5b2PuAvqzx31MapsX2dag88EnJ6QpfY387+vDXxosW3XKmgmBLd+0yj4hU
/kzd3B8qW7TlAdrK4moT98fUQ/Prz719hgDBMat7V6tHJImmkwBnyU+KrEN9whm8ZYEEnG9JJHBJ
sdurB6W0FeoTJCLhQq4mvp2ILYwB9mohGn5zK56k6qKv7TGzQVTjoVqdhB7zZSKEpXsXXNPvBfAb
I8tNC4UoMSmzYSIsGZKSvfhUJuHlZMcx2ENBR4PudA2BdHEOrh62lIw3uWQurG1WEKDYzxUx8BBf
d/7cIWR6bDnU/Rs4B0CggRpfK+6xwUdDZB41QUn8wDBWGyehwkxOjh0ObbF7OH2Vd0McgBQHMj0q
gt1MgaDRXmM+SDP3nXOo7V4yD/hWu7cH0GXkQrynl1Uv/MtEAAG+Qltj/SSUMDnqt3uUEsyeAV8w
iuOZ4faN/RPZl+dRWgl+kIObJ1kH3urEZPlUhN7oNwGilLafDf6HFqMumBoizTIQQ6CX3t5YxLOF
fD3jgNnLBUY4Y7d7VRtsmS0uPRRazHayb8eT32tQoFhUqvVf/DNyLsk1GyAWHHZIYAOKl8iLwb54
UvFuABR+zUSKPh35l0+P7kXHsN3oniYZzWnR6bV9/thdKbZJtrd6U67o06Z9qlQc/Ra86jJNIP7F
axEqpESw/e74NYMZIVhBeQk+v5lc2ItyDXBkzarXPBM6b+gdAdbOMg8BA3oXNojS+867OQzDnn9V
+c6O36bl4hWM4RQgxqGKu8mb1Ug25fFUXai2BoYcq2sUpmSYxMMGSjuMv8jOB8XfJ+LtbxNM0X+X
FetYjdWQ18NSL2wQZVFIAM0wShhFo3QSdqX1r4klZn9kaNmS/nvJElsNCiHswWep4+A8Zz2+R0Ah
p6ISln58gCmUeYPVnvuyiwD8wJzncmBH7AveWMzpHeHxuU9M8h9XJs2SL43cMgrKXMCLUG7/T7x+
kPvdYB3ps/7gOlMo19j8MmW4j3dBi5J1cRwT8C/zmps+DfqrHWoJi7wUUTYbLiK7dCQG6RAkNPUi
vOkQbVdpu0sjGaLAW7uExyLVsr+b/SDoyI3QLlD1jomA2WlTAc7IjsT0ts3MjofoRRd7bmISem3J
weX1IcRtXqNsQXnZSSIda0QV/S2WuIVKcoyDitliuaniaRl8tLtVghTqMnQuUZ3uksfHJMVdnwWk
oDikNsJkZwKoIJlTL75hIQzQC9x2yw8o+bTQL0GdsyiqKCF4r0/k3QElGURx6jCo7WXyWCdXQhdm
dJr/D4P/gt0uNsgtdXUdvBM9xsEkhT8vpsmMQ7Or/xrq0Us7drCOrzPaG7tfwP2rc2FMxPds2LBv
jaZ/ZNgsggvteuJASpN1z0UbmxOaUItqQbTbV/61sG2Fqn5xsSIsqdAxNgvVSMZ3jZJ3CJPycd9Q
8E4Sr7exeIShxOzrSJArBJ/KqT0ekUNa5TzA2RBIhAlygCSo3CPWJkqK8EK5xK+0Mm28557KhHmJ
q4st4kegnvGbqmHMa6k4CVIkfqrisukWsTvgF1UTVGoA0t5hp94wDO1xp2+UMOV7pv8kP1dXKmSr
digJN+iaIjmpIFWx101I8q6GdX9ezJbUErnwH7lXnk2UVzhK5G63xolAPGRDEpeJPz/YKeC09Dt2
b0YuWSrF2fi/MNRkqFqmtp47Dl14QPV7wHUMz+2C9EX7tWophDHl8Qn6gAAQ+BS0HrrzUPSy1NQP
7RKKkIolmFjCMVFUlGqXpjr3f/GtxiaI/EI9EPgoa7eSlK4RQJUImVcfSkpqGSSIN/p2bz724k2L
9aJr8OJ/PX3Ij0/2XhB04dwy4iAuhPe7zAjr9BanM5QD8oajYKHKBVVFvQKV94yKw8WYYElUV92P
G7DvlX75km3yWz8yJIguSVUdU5GTnntrAKMlbPTx08MoMwgKduHv9sGLAuxmJhkFSidBX5nq3FWr
4wYnexJT4V/liV7OaqnmGeowfN4k+f1QBTo0hLrJD/W81kEFDaZ5vo1F3BVgkfp00yLbqirTmLXH
KsAdHRC+m6+ugHjoR+Hk28MdBEQ/Bj6mNUwiXVJaAg6SqdVIFg86RPZ6eG1TPmnj/Qu5ocPmV4Aj
tVjSYFbgdiCy8NMBKpSADu5G3lV/AiXng+Atnxte9LPFYlTGt5/jjlNbmK+65Q8sQJfqlJLEkQr7
Wcv6T4aHdIZBnA7YyO5pShnvRkR/23p9g+9zBGXywN3qsbEYXAA//Kbj+Q9Ht1v7wXn7lWDx3dvX
TubACDnPQF+xUF0FcLOw1NPh344ymqWahQSb4JwLqHughffbVJ5olOu+OM/mvNqNhrDguMeWaCm+
CS2U6mD8Yv/EylgHfvKK+24vDN6X6jxmjh3vPsqyK0cPFLK/dpfDD75LANB27uy7mJoNo0W4qECT
MKt1I43mh8yvTzMjIfM8xF0lnRG7mTN0ntBSb15v9vOH8ptBZLdFqNbNiYydx9OrGw7a4/1W0zBi
XHTZI1i8z9YGkefgltONWd9DAkSYExXnh3Q6rAiaxG3RdL1JrqklzsqZ17XAKfBxIEJx81dr1NJE
4vj7ROtBzjyh3GKWIGkuatX2HXddH3SnPTjtALRygJkkozFB/m3QgCFe7D4zOSoHEIancQMleFje
G6j1/RYpbu+06RsMZ2qqMbhxQov815L/ryBbP8Q8pFFvvj2aRa/Cbtpr8RuHC1YFHT51qUY6og6C
lFs3K9gNTyLaWli4aTqNurhkoGnBO1qDYBuwlA2I/+/QoJgHDQyEjNps5ewsMsAabZyDpmQ0q44o
1YDdCtp4+r7tBEE4hbhsgdYHjhDjJU7IULklKXX+DIh8VQJT0nW6iB2yl6B8UmValLqjDoxzFxP7
RkqiTroOTOyDOP/e44gC6KrVCxue5HVi391birLMMt63eMtlsbduNtytZjLQf5jCAZvsy4X3Ydx5
U7Iga8PJUGmMA9cpkIdYS8ObyHM+vq5li9Qr0A4djhF+T3J/KGToyggY5jDUhqNPGdfeAoLbdmQi
I8sz/eTr7zpNKtCvX9ySgnYxVQTkeNTuF3lZTRxathRiuIqLMMS4YakR4vZLCyXO9Gapl5N8yOEw
XrxFqGodvzAQMnIbYJDEr+gA/YDLEPIG5zmS7L4arFiaigcP3HaIpbFxkNTwn3b5qpG/WKKAnRvG
4CUtJER6h3au0wJXEbqcWse/o5Fxktrnl2rKqL67TAN1ukJZN5gAwyE8e4DRVpJs0lz5uGO/yEZY
xDBRJP49SW5BEi9hOz64AuulPokwyYMTAiu5HwDyuUwOhO2Dtum7sLNnVeD6HVm+DED7doLVNf1K
zaH2B+16GUJmX4u63cfiW9i3U/yywwOjsr7veVusP0bbiGeZU/oJ6hIGifOdnK5Z8ZEbhMRaFn9s
fhUsiPk6gMOT8SYJ5hh8dQrQDAC4GpF1TR/Vi+jokGEiJZN4Zgf1TwnGKJu/xdJHcWuhW12nCQkM
Ro+QDDsXDbM1TWIuzhGao6gHjjBg9FtbaUIBjFjvhCni54pRUMcU2s7JxkrXesiqfG7q/WTST/fQ
Mx1Y+RWBEeqHcfdMuK13zECr+H1Jj5/3b7UoWoeMU5j65oPnbh7gyIkhV5hpP97cQnOltVsQj9t9
jmVrXyIUYrBiHqAPMooDRxS+IjcbdeCy4Q/9eRx/wZ72ooAR0/D8zCm3RQacVsDEtNIFZ7Sgj9sw
U88rz6fiwEEQ6QFvdIfvxbDFTxv9UH/n9BkVcbu88+TwufbmCfrwWKJ+P0hZK6A3yKcWMvlD9W80
+U2eyQ6U9Ab2wnztojY2+Xz5sNuX2Tge1tu+NCjueJfIeHkHQmvUh+kt3IM3E6PF+lV42GEBVCTH
GHunEsiL7jWR/gqotxcEPubcnFd19pXlgjrj9XtXeljeSDlTOtZF+msbIf5p7tWreZELWPDR2MyU
aAlwgcj9eUdWx6p2ON1ah0EZy6qkprC2eqbK27TCA3Hc/wEVXRmE7BPMeNdr9/dA68c+qlN5CL/C
8/z/G7h6QzBANsX7AQAgQICPEJ4oHtQf9DqoUgnPN6d7dR2XOxbGZqVBGbe+sKJrrLkzbCBFlEQm
hRUH4pknLnFArpJZb9qm98fZGCXizcpHcITD3rBOhkmf+DUMVGtA6kfaFRz8S4h53L4XlK3TvN9a
+NxKYjgsYjSFJs0rE6RuIzH7hgm3ktJuwicMZsb9H0BLBV65foQvd38iN/cbVtE+0uiU9MQA18H7
OAbNzTsMyJ95tctwccz5DkWtFHgiurvEn1vmKF/ucrsJtZ7uvvuODth1CGeU1VZIuqhKJ5IZCGtT
BgZYU7Etk4mlP9uqrD16CsoyNYZ9Ly0BSlXWSzr7evWO02f5AqZorFBq4dzOApDsUtCyY4X6kVM0
qG9GrU9dAwZWZvmeRabJq1J2wsvZkNWZmOxe+9eVnXIJbShwUapRuT041W5NCCP7G90HMJrpu4fc
5y58X3Mufcl1Pbi6qw1SWTEbRLn6URMJUAbSLfAIt2c9ukVDUuqw2E3Urrm8bunOKI66HdY5r2FQ
iA8CWBJF/U8A7aINDHOTqmHegEXHyzCdT7AxOZSCu3wpJ6iTClINVTsGGNzKX61NjLdo+OeWramg
XvFuSkMwvGyKeRMysf4PJqW5RiqumC5HLUJdvJKr+VLQja2MGB5tcpSCprp37g4Zxz14mRbhE1t7
TVL3YkOJbYoLH09whHMSvYIZ/wuNHNidyV7gHsSz0Eb8VQ+02M8C50c66r4ZlktrpxSevYxRz1+d
rWptzfArOPRKSVBiHQpt6nYiAZ1ayW2OAlhd81pJQL/6DqkPS0nghYvusxHBhEDd2qfjJsqrKu1N
FiAaTdAc4WXFQDjh8GmxV0SqcjG3YEgF8hMOiQCJMAibjJcPhUw/XzvMc5ZNi/Bg9lfuyRf6Uojo
f4fqQudG73nxNmsVEBJtbuZug0zpGC6BeIxI0ZtOerbYu2B9z+QdZMme//5jhF5jXQhgzkkBM137
5OCN/HRQNzY+RTRcy50KGcMhQJ3dPPPvQpVNeMEU01XTMmydMG5gPlnC5IkRyeChoJkNQTJygIgb
d26cZ7IYIhMB/1GrkwyIdbrDHzGVwwGpdO1Un0zwJg+SHcZgSryjOhkQDqJfx/gKYTZHiW1VShu3
MquxFe/EK16BMaQ5SWjEuTWkVh1WlKWuKEhKUKnFqkE3bXch1sDbmGSeIFf9MsmGEngdqf4oQK4w
m6oubd1h0l19LYgBqsFbLnnCl6NWVFS+rADylVFYY2VF82mZB78i9zGGZGh3jn2oTCuBWT8hyGM5
x7hn23G9LdExBnOUOFxBm9b/ncWBsJqwO9GH4W6DxLKU3TlQiEslHj4syHm6czxRBl9mtDxR1FIR
YEn+p2LLTEKUC1QzBEJlrJ7fWqqjiBqccN7ueOWfLOX24xVnQe66taSLyJFYkQc8Lq5f1ZYboxmI
XcijyQvJgW7lAggCy34yfFPf7uNpqZUaQaIql2+RTe8ZLtwgRXoNecHlgnVcb/hrNXLl+GyeZ9Tn
3GTE0OE/lXzUht2c/k9enuigd8GkL52d6HSR5E91Kyyl4igmoKMjCa6Z6H85hPolpPu7NIpyvnjC
U3M1U36UDpDcde/hBB0tEdoAq8YIxHljapU00m0mpQYvit/96s3pKwyiH7YCm9WMjMaOgWH66mX7
4P6RzMVk6x34Xh6Pq3/R0qAqp2FBe1kGgJsN1on/jQbdf0tO2FS/0isQRmWkTNdAuzORo1fKXpk+
6ZCzbzFyOejM7E7j+oRTconl7cgJ/IjPqUN/fCFnfFeOrzMsyjiWJkdQ3LilJBc816QRa8uM0SL3
ovQlHIvPqLRpIJ7ckj6P/G2XxPDNjPYOQaQQ1M/1dSgej9PeMZl0kWdnhtC8866qIuVzko8Y/w9g
3VNbEqxYsh3S1nqqS6DjXzR3HCn2FCQ7aFDO5CSMRfAV0NCdsfUrj40VWnjDrxgiy4PYLEQHjXg5
W/LBH1TWA3FjPzQFT91NvOLQZ5V59afHfaKUH6cykXXbEq2J+AIhu4nXnitIi4o7tjDRCmdxV4Ee
XZAltDXzokoujpnicZCPiAXW5YJ2WXax7BzxYpmmtQO8XLg0Pka0mRGUZgYc5tJ+XckVpIZmZToQ
apr0rrhRcdnvge0rcVQo/tINskHqGNw/0/SLK2t9IthxGppKxrg3tAKyQZjxqVMgAZWIPBqmx63h
uAjQuW3j1BAKqUTydRgOwLP1j7pQLV3ruKQxWL3QNmhR9N55A2/vpdK25SaxE91nd661XpVTHxQq
cIitna/oDvgh/8fcpiN8MIBIcRQ3eHWC9Sv8Vl7LTDgDaoMVWwPfmOONQ5pJuvMv07APg8jhNapJ
d5LWEu8Wb7c768bQXqwJvGFqLLWvHitW853zcv3ktl14J+p5vWW254EjSJ+lkqc5v2nSSy5j15+f
rRLuFLKWYDuyPCh///OGzYVYXF6cfp+BK5NER8jO1xk1iG96m+dZvEQZs8BoKRyCf12eO8tOHUVY
NrcVATN/IIk9Ux+GT2MiXRTtiHMln1Ngurhr0WB5a0e/p1BVmPOrGZ+oJpU+bhvcbUUbmnHXXjf/
B/6pi0mitoBl3mrGYnnWk8aGBDT5kHsrf4EEpX7JR1r8dajzQAeOpmGIBiCLVI6pQAdwcsaGeNhn
SHx/ewZbjDjG+YBlOwnFqEwtyrgHsxnpLJmROtQfBAzKaK84Px4zLHtaOhS+Ibe3zFROiP5Qskcz
ttSuuSrWJXBMyMjFODk5m0SSkREBjkMODqFL+8ZfEtQKtnrMrZAEwZNW3OFsa5KnF2of/znhweTg
+xqtZ9Y9GCJEOgjm5O7AV16PegzLc8u83AKbSod2+SvGlwjEp95eANNsQirqOtBXAtG3n+0033tX
sqiyJxyH2r94751gLqiWJwR/SisRNVS0BYg3W1G0H6SYYk2ca0TQ/UoXqw4fnYoQI6xKxffL9x7h
RVdVw724tPUGsiMR4o88E8dR6i+sHbu5CedOrXxY/03Nppg/SmA7ec2WZJe0USMsq1EWy2PTSTgb
ge4HZ5g7yhgGvqKlIVXfyQPFPe7dSd4QKVpcG+HRWMDRuL7qjJLKDcsG2Q7xyZO8oKyzXyR+KlyI
TkWBZ+HFQyOi3aP4SgpVTLynFDY9wnJNteHzw4ur1AcAVGl7mmhVqyb/Lg45jSm5XCqWww4lHHgy
iz+UBkbIF6/PL8SkcUMSFj6r7XEN13jNzSjZbpf63Ovb+ygqABN3aZQDNJatn4kKw8YY5o6s2B5V
lnOsVlxN8cIQAPG+zViiGq0/WRxdZ/H2K9kOf0qoEAGlbbqJRpqNDsG+cdq/wwySvBC4MtcY90hE
yn37433QR/6ZXqTYuUY007YEg7NpmRpqNMHrxPaQy/aqnaH75iR/CstOzPZOIh0xSYPYO7yCCY6v
eUfaqKjrFbhijRsXk/I3vGJVGz52sTcdTid052DQvB/ohPB5FWfIotgEpmQs5n0WA+YOqaHI/6hb
VW83rtABiPOX9wbnBcOaC0JjlmjgX0CheRHwKwAPvH3LWuL3jxNZgMUYBvwAsThKR2vX0KIsmee5
mjdtapAdb3WgqKgwGRmzoW6s3hIhG0+PFUTJJBSI0Fyh8i6EglVFIEMDJfmCPZxJdLLZAuJKbByG
+n+PPlpxUcjGyQw7/4W5ja8sLj9+mf2EL/jV5XuAAxJ4pmntxNXHR97GxW1dGzoJ3SzGnSxZNG6A
TQZB4cAtR5GUGd9UIg8g2t8LcASuL4pigOTU0/ayPq0UQDJmAKMX/O++wWXp/WOk5rQhBXtnjbj0
YnFu2cw7OZMjvW2y7fY+tm8OU2LPJYo2u4tGUBr4peR6kCf+pDM8SB2BXKUKxOHVFqtJj5HRWgw9
qLK8/z2+eDmWBrzpJfAYA+vQ96muQ/9xmdYcCyvpxhHMYEPynyw3xLo463y40acpbUyN8Jj2XsRE
hnl+ibPzWn4i6EMJocl3fw9lULJbAw1hr1PoFw71dhKYYTJBFISxGNnUJAPRimhrS45NGXn52ckn
r3gmuxY8o6SJVDRhwnAgGKBAKLZ2CEXbN+Qv+GPyZ8LZXEbrq0pURpnWg1DIiOrlXXrOULKYv2Ef
2/c3BZNp+izEcna/bv0Eal+b7lK5UYO4q5lAtV1gM/bxcmvYE2sJBqE97M9QuK1EjcDYuPPqj660
BHmQnotwcMEvmqzBOCvDge/MVnU/3u7Wk96A7TFwpdCU8U4QHrXaVO+OVWrx1WQ+2QPRoDLvzBRx
gQJeQjVv8AC3neOhmqm3FCDdEhKHZbVnUCn7rSbF37zxWTt4y/Z1HtgXedLtKH21YaHmqgqp4aQL
b6eJNnl1c7Rh4CZeLTqRTENwXvkul/6ySzNzwV8tnkMuSObOGk+Y/iqu6Trk5oOek7Sfvv+R0iz8
RKxS9lIICgBWl6wa1ZkDr0/o6KKlwWFKU/6TU9ZzeXDQ35ZPsur1UpqnrzT4vK3ax6JZcakpgMWb
8zyQBH0+BFoEJlcWkK79UnSE19lqRzpYhZIVzLJ36KMw1teO2nxBKrPZRUUCSL81HJZ+NUPym0Ie
1+FEFTBW3V7qYP3mRy3bG+Acimq0Zb24Ml7Sfb+1695G3ykfQQnuiJIT47Yyk4FsEIir4faIIW0M
KBrZ2HHIEmZzt23xvvqbyuzwCXpdUXGtAHPKfECAxnERHD1WxKYYNZTIc4wVdzWSGWbGjy8uj9pv
OswCDyWNNdATPS1Y3l8woGDzxlE1Q4cL+efgGwSf69S3uYHAsmmpGwhp+7C4cnbtd+EAxXwUzEPO
a00/MSwWsKIh52XkaIgTEjWyJPhH3B5VP7pbrdqOfiG73bRTJp8MoebeMY98J+S5rdPCrivDbM9x
OAL6foWlINmecl1kBsrmnYd+fnvQoQ/wo1nwXl76D1n8YkdDEJUBoHxcvLfTP6bzztWN0//UNSYL
dJp2kU586x10lhWzAJVFDa9aHxrlznsG7xdYPmYHCsq95FUJg2arppW0yBemVtqI6sunlAf2QqzL
NFqfZXlQXjDi9jNk8W0A0LpurKeccwsp2UW1HAGpEad1uEYtibnlpdcA/wUKRr9HNB0TtQ9Y4PTc
aXm42rdt03Ehge4eYLiPVKG+LlCvzgh22TtYtBqRzalJ3S/Fo/5mxmNCdJaQmR155h+nhaaLbr3p
GSWUU8DB8zkEv+ozelhHHMCybjlQn4T+Ki1b53OqcNLd3OMv1rR7lNJZCrIRQTOebZb2VnsVclJv
0Dyg4HM8no3euenATPq6CMbRRPbme3fUcIfAs3+YAmmn9SAuEjvbYs6kiOMle764OZw3iFsGbfOn
GlcKmkewvNNVG3OPz3FgqVHYXwnWTKFF8tpx7D034UbZ/Kfuv1rVLJkrvaDqjb4LZgMETQMHoM/Z
b8lHo8Fett5cX4u1b/rZSsF580nWR8LlBPd1LDO8hNyOu8c0Ldgl5LhVMbLI3DjESfphtZtPmezS
UAyGKedFJIjGEnNx+2jgWvOksq8mZDirF7NTMAHPa5irzYHw7gcJhumA8MLGNMGeU71Qli+PZJJm
XWPfTGQUQ1WWSXsVlb+YT7G2ndaDxMQAjAXSSTQqL8jEbsxYFCrPx7lHV9ngXTNtEZngCWyLR55X
gSq6tVrOUsCj1+9AM1uwnHJLeHSV/pBygqw+ny13+6uqqsOl//qlLe/zvOLKxpnrh6zjUCVj+efq
o2ACZB/TpllyrLUPLLzzSoTYOsqlPZg3gOeBrR9Sw0TDv5sPyWVvIe6pQvK1NVMw/ARozM2Gd46n
Kft4LxcMZmS3Ld7FqTiaiMCDZNs7Wm/coVHL0DVvxTCeIHKAiTn3K/+JuZN36mTiqAxZVhpl4AU/
x1oVhRur/TVs4Vi9otdsRHTgfjVuFIkzHx5TLNt00VhFDkygd2EJmQHbxRj3rMgtkwvnirQur3F3
kX1LeWvMqpjDoOadTPqzaonNkydLlI+C/xQuQnN7p571SCy6M7LHx96f0o5DdYW91kLWgWCNFADL
Hl0SdzWuNTGSC3ooSjcJna+V2Tzg3s2w2t6PD6W3ugfm1wo+8GNkr0FqtOTLkUqaUF1tfyRBMBND
B+NNWeRasP+v42OqczQFVTpQNxoac5HuEt/lG8JXQgwZCAGIrSNcm6Qm2uUtkf0hQCUe9xfVWtHT
P5Tgfg5xj4eKq1GvhHEdzxlXSnTTRT3zfKLBVUuqtewiDqykLHSoRReW00JZzCelL1lY8J6ps1eW
5kgHsq6c5nq5jyFIQ86k2evkdT5cAy+oPc+IkbKd3BWzOv2drjXF1fWRNI2tvJ2fThm1TfF8uMNu
2MBe5w9lzL3a0I3AAx+uCVNGiU0XtRTK1MYMPRfv3OUp+9OTY0gMm4Hlz2CJOLd3fF6nd7B5gg+r
IEwY8GfjNzPanmKPaXAByff59T1K4njsdvJnTnsp/U6PfdKIHIrSmVEgUkeg+Pm/pINEXwfFQnfP
Fe4py4VFiDwQ1ux2w6IK0ejpxpjoaFubUk+O5P9dx9aV5bXKfA8lrROf5epBshQDy2DLvTtGBp/A
bKEl89wNEQ27SRrHJRaoYIq0bPkVvM5+bHeXZ4Yo3ibnDVlHNcyKjvOanOnC+n5DUS7xme9RZfeW
GXAxYXVxlyfVezNyOD0ZIH1hl0OkqlGqJ27KJgzQ3mgMu/1K4qPvdXH0pW2j0bMRzjHW1XaKLQ0s
DY/LfoCaXz14PyjEJt/Uk8FUQRVP9eblLg1q4pv6TS2Cygn28gD6ftufzkwEzObBOjnS04Xqi2Bo
zEM2OxsSB4OxURNJqsoNwoZ1/UedwlK2tfp4b/j/olp/QTaVXEDxO6J/tq9oj6K6/cjFA0venNKg
NXNYJCCk8KvB1uuwj6aVQsG9e2ABjaNiQNCsys970GNKz0pbEAL7bWI7s1RhNFVDfR/udJDwBtZz
ASXwAO1nDJ751zPOgYJlPoQZ3GjImaCh2vAhRAoYFATfwAX5KU0wVHeVEhJzSa6pU0l00YvkDGR5
Sl9CvymyTWlxq0NCxwTbXZY8rkPJp0Rfdhfx/ngZeiyoImflUuIySuhMn1s5oZa/M/8J0Xv7eQE1
kh+i3BKCuZ0sNLDirt6T28tNgcqJs9rJFgK8/RWcEw8X6rno1yZiGmxWish4KGoGZV7ANxeXdWtA
w8l83FEvQUYl9Ef+o2X8SmbI+T3cnglPxs9DyDrHgc1r3rSlUlK/Yfp7Lna8VwerdW+o7sOKpPW5
464zKfisZ1ePECVae870TpokH5o5aIoJ+27QCHz6IlO+z/Cm0LqXfL2hYBnUoCK7cHUpNWiPRvaO
Dav5XVZ9nPnKwIA1maDHHOnKbzSEsAXIKvbT++fYRckCQdzbUX8c+BiwRw116SojnFs6Ns9TiIr1
1lbl29/9RSitxXHYpCUvYY59rHBETn8viS6yT/TxH+54d2omFNSbd9brkGBMOq9PfFvIynpROOh+
JSw7TiHPRyfev/JnV0AcosyZaGLhbglqIc0YmkQZAV5qXdJXxyyTZM476rOfJlhjOvJ4EmRkDHEj
CtRoCI5y2UErE5mqldB3fpYrmuB9mkVHl0/Il3jpvbx8yOiHUDW8Adyzb9v2x7TSrZJC7NgSbT5D
vYsuklIcEWmcf4+/LbJXDSsjFwj6wcEmSkaUBqtpoE8AIU7KIhvwMAgoY3invRhk0yTyV0LrDyLh
jnZWWPgJNkBmpO+d3RMDTAqeCml30BBt6bR9XLbuBFAq6Ez0ATvECsmXqKEcWivutQL2yCNcrnWq
gQGtRrGCWb5GR35qypjW0B6qv8FLOn8Gzi4ESIgZHTmEMygq59IrfrZYO8yrWpknDUqYmXOHV3Bp
fpYSacGBDauSe2sQD2zCsffGKEdQEKJv3YHa1gCqJBjWUnayYOLev4ynedbW50FBKAti7cU6mvIe
sa1sKqZl7QkPX6yL6cIjtCSdGegwX80VPGqBv52uEcEC5ixItp9wBEdhK9ZlXhnRPfW8NwCjrnqi
QOHgW47syLKpvmgkzG+c3qdlAnVd/1vnNCjmlUSENOjgnRuFG3/l7vfohMD8FwXT6GxGksrdEm2G
ohGa6KZ7v76otz6csGKzPlRNZXJlep+gQt5OsmC+HG38F2LLlvebnxJWUMiY8CNM/XLmBvmNmLRz
rYgOCJHmQPf9ZjrQ0Qwcs9yvGDyURH+Y5w5W4DqTKtgfWqUV6LCiw/l+r4cSDpDozRQvpFm3AuUV
qoOKu9Tsx0AkkdL81YQS/SlcCTvVPG7rk1oPwaQ+A1d3MGmrBI8wAMqFWp2RlvN8wIBjVtu++QCk
DMy9E2WD6uvEPn04hgBEe5/rtnkTSP3gE1epdbbHDMSef4qloEynu4O4g2iysl35lTZLRVhN6rDG
g7JTVKLvv7EGwo7H6q8GcbJw3JykxHSTkfVPJEDScVLRlkT9Y873O7nwrKCRylPa+1ZqW+HrqU15
M6Nba5evTpW/YJ2455NbNHcLj9AcRTHnRxR5uj5yMll5Sush+hBrkdlVeFWRmyFWav6L16uXA//U
O5KcOEGBahWe/7XtGZYaCrQNrZPFWiEAgGWXMMp3n0d2gOesRvV8FRfHjRrhk2DzzAnzkUTdIj/Q
W9QJM7fior7G/mN9yy801y9qyvKi88kbahTddu+yBDHStGQz8BEH07aRqWjfuInZbTrOA2m/ZP4m
vccjX9MSleMzt8vUdxKyVieVB8JOYIHKaSbPDbJrUsOqNW8J3WAuyI4leJp5BsQGPXDD8GdGop8a
jrOUKDiYpYiBKubwAQDqcDRk59fAMKcBQDSBbdXMSvRHrZWqaeO6ML+rRgrpicp+GxUxfSl7QZ9n
BZV+xS78XN3vtqU6yDwd88009ATo6at85Y6ImRPl2fURJ+ap0XInkzxdmmsfA4Dqh8B23OhnUUoH
bezxTtEGU0wjdJb5tMn6oa8E0b6mv9lkFWSqdcOR6J+Mt75GYjqAliryBAi7PhJRHVJ1G6hkK/bP
TujLwmyv/fVlGJbpFhSgoR3ab9MAs263wwjcH04rzmJXSBtR9U42dRwi7Ye0N6Fo8tUVBeYTxY9L
xq0sgKzSdHi7+5N0Tup0XSeYnca/RWT41YGIq4n3IQneBQHqbKxziV1G+KyoYDTCwWsr3OMW6doQ
EFRx4AvTFwBNvgpRgAforbqCO7f1+O9Ov9GhpbIb05uXDzCFRYqXJwXScvlU/oeL18pcOhQ8Na2J
r/eWj6gGjubXlazCIoFBfXnmPUNVZIfpnS2PgtvmDD1i5SpueEi+YQ6+hZaS+v6YQZObhh3s87+Y
33bC8iPdd+0Qh46O8DMpnNIIidvRqJegPLudEzkhDxMjhaOQiahsSpbSgj2oEmA2OjVFNDVmkHHQ
CRhl40QaBLVzGaXkK/09+TMCpjhWSowh7q9wS/J11+GHIM5e9eGhAdqpYQLa4ZFwSBT2wZ0A9OCP
jk3BC1q0OVoC0/hrfuha8zYl7klPOrLGilMzY1VXbaPQ+SpOJcaFcmn+ymBMN2DYQnIqSZV4pf3B
FR6ZjfYnAhFHKPfFFjitXZ2EA27OWWMGImyIyLaNiLs4QcHvH9jBaYgvX3bBj3kNvQtvNJXskHrZ
sAldYJvhTESg59inAvnWZ7ZrXMWALIoXb6W+vYA2IpjAa3ijagF+iqIcOX4DfmyEfclat6J7tC/P
lRRAgLu4VOU4F3+h7Cjf1AGETQXkIeu1m1RTRQgF3s1Lt7Fu6e3unV4OsmaYIYEqzBWwIibZZaGS
Xb/rQmRkiHyikiPzgvp9We+zxhydFttATvtyTVX97ko6C2EanA3fF/tk2XHhMmfLpY56sQlnJSiv
coJbAKflT0RrK5d9a6mjWNPeIDvb9B7XdCIcYEWYghruosmuqs1rtunewSYYn/JPe1Ghb+9AFrDN
ovkdx+5XHX5vd0dLB85NH+ohJgXIhPCewB1CtifDbvVMxgUDpv4M7ejyCkvhLp2Guy2a7RtZr20+
kyoxUcxk4xn6RzTWnW3BgaPUOSzBuk03WzLuo08TDN3MehadmHh8VtkZOeRFmI1p/DCJPJfaX6Uh
okAZVdE8nzCL62AG+ZvwE1qRIksJJafVUt7z0CHoepw9k5Xc9mrlG8Ssmao3hKw71aNHweqn0X4b
we9Vg8KuVQvSAEyWPHRtzktLMjZy/IikfGhb9CAthcL1j+ddn4zzdI/FC0mzEJIWye7cer+g7WTT
ZhaY8Jmza2M6+2nTvLYUpJmwzk6txunHg3KkoswezegDUwGFedQDCeaYQtdgc70gZ/m/FTsnjaRo
IxN1ThJH/ITj7jIszzNW6skWsb7MCj2/A9JwRwdUfio5Sf+c63y/3TEt1GR+WfJabUQp1tGIX88r
jfP++g8pavi+ABVnHQ4GZJ+rfxoE+ZRw3IBTmzctSeJKXk1OJEibBQrY3n3RTfRdnLHZkDRzjM59
dahKrmmZ2EXGyaUjhl1aEmBaOJgJtUDW4IG8RMPACZ5f+KEiBmgJ89oug7FvrjI02tay+usVLVIx
BCSTAGTGGL32X4ziF0KV15diuPgRvsFUndzw+MAMx09jeR04YxD2uwrt4YmheMp9ngT6IX1+Wypa
RvdYnwcm4PUsHvz13SALM75PiFIeSeIOhkS27+eF1lQfS3ezVOMUJNLVopPiad8q5pB2juCPb03r
nwpttNpytjaoXdO/KDdGEObO0li3Jca4wGXRv74eJ6otAN28nqxOgmRllmfPC+wGo2+OztJpvrfS
ryEmWhqNkwr7LG0wULWaNJqUGV59N8wSDmTBOv50yACeTADMNcC2kIzWAWt6HHaPaXfoYSNyj+yv
rKQFmcERjnOfNuPIkkG1CvL6yAhuHWHXxe6Z6WFwormNj7/tZEBAz4G9f+UepdmjpmionT7D+NXW
pxQwNbDOu7iGTp+cQ+12W1ozkcGQSWuiExLXgyKcP1TTf7hv9w0p5wb93dHke/0Sr8E+JXRZ/wT/
83I103vNBQK4Bx+Q+hHM3n3mAB0elJI48PfbO2Wq3xglicykbTnpuRlkhC/7LEFsGdJydx8icqIg
7VxDmKo7xSLmP4+hUWHxKs7FzWurt4A2N+5y93e1VJXy5RgF0Qk0AHUNYUVUraf0YL+qsl5n6Irb
DQ7vmXD8mZRHbisZiUcUKhwA+2YjbLjlIC2mE2UIvkeI0BskKPp0ZgN0w1fKdGvAW3T3GkAyZy41
KMfpX3CeQzVVOo5y26zGGlxH/4KJ1oHDs22OQnGrF++YcN1IfkQueyT6biMywGrLPPC+XzXde9Tr
nmuUyc7qolyLNiKouqLK5fniewtuV8G5HMxHpDB7vRH585jDPsW1Q3xeQPBFnSW96QuV6YB+vtd8
YukRrUgwfkSF4vgLr2yy4vb9aExGoLyyEckjTjAFMAn+U8jj15ymwr8KGior38xj93JBmHe6DQZq
83r440519oSOyI8DLGjklaMW4tDfDReD9pIQYUDNSfNeYNOG0LTgF42JH2zE/un+Q8tWSqcQPL4W
Nn+9Yt42WJ5PCzVf68GuwI9MhQm4uFMS7sFxomJ2aa2xEv0boZGW2igYAs5J/c+/EbiNT0MxFnQz
79tWlVYjBsiDh8D26krLHftk9BXNCqKnTBTnByhTElJM30OpvAYZVbPWCGUdV9ysmZTQPmmPwcLu
P56FetMK4BhIplf58tRVgqh35HVGvo+aF0x8p0Q/UGUu85fX+XrdBce5qsQwjArDkMUrm8oo+Vug
bks25e2QukMlWNC7+mW6fu0y7fXKW4hPoyo2yw7qzX5qcsP5Oin4dBYfAXTFO+Di9OuI+7J8TQBC
/gdLzHOc8tsN8aov+hn++iXcyHkPX2JoFYCiI4/g7yHaEdokNZC+raaF8X5fMfWv5VOAut30SVeC
uBQBJToZCjqYnlFGawlL35noKeexT8rw0v7gHIrSuhSZ3l/7VTCC3z5ISYuMPIAWX8SCArW4Gii/
ByX1bnKdHrlnaIRMmYPRfB5proOCo+sk4uWrq6gGHzrzMOpKCSwN2OJQ2+7fV3XgEOZhvR2NMYzs
3fsNEElkd3KPGXRXl774pIyiS0pehh6eFPfFN1fmUtjucixRcLsp4txQARe2OX4soeVzaM4OMc3S
p937yIDSiL4nTNv4LFvafURWVj5Ubt6habPzsZIeNrrGp3vvFQQGpAzVAE4ZJ4mPAjh0JjourM5n
O2muta2JXsVmYEOkNI51AFBusnRCqgXSzqfv4yiSO5UCdVI8AN9m+L8BOP11PTOaoic3LI+gKi7w
dQIFzC8bhKlJfNEjLlb4jEItL2sinXfdLLxHlp3udpW01eIkbq+rxiI2E3Y3HLviWB7F0hyeBO7q
XNgCEW5yF++tFrtsjUkcFoWzLneFt5OgbiWJYMr5oNA604pu50umhgUwEa1eeNJ29OFfQ9LYYbTt
WZx9kXgsNjnjhAphX8/sE2B69xewoEG7FzXglviVlXtF600iGgXLdQINKsHyyG5uCcKnLfWzpHA9
fLee5ryIURLr0WdM2DoEW3zxPZeFeW0y9SAvmFKE8DOYKd6zvgZnSo4wn9CjDr2WSS+ZgwxgiybX
FP30Dst6FgoDc65cApAdtbI0/2LK927ZBslVlhbc/IUx3O90SfiSwxXgcooIh8MsE3H4Hei8kSXw
of6uFmhL9qe0LSxn5T9dN8XcWhlzWa0a9U9iD9KFPgOXOxO3C1Yo1U3lbnlHalMw+c/m87CUwag8
mG0zpS6q5PaYmowQWYnmmbpPnocu1lcWfeRIxcqbW/vJVpxrNOXFRvIRlO9l2zS4/jv13YW56kop
F9qEV9tPYBeCkpUWWZBatX284PpFX+e4vtgvC6Lb8NCTUHHrynJvra/W42i62p5xw+1YGdQpucbK
bUT0zFzp3rYJx7Y+juNHDLXBAOpjkjsIFBVi2KL6MZngx0asFBa93LJv1pBZWq4geVl5O2dSUvZ8
reKtXDTl7UDNLP9ocl5TmlR/w2Aa0FxL6rgpCay+QenS+9JOdqUPB9JlrOA9gGy24UuQslHc7AvW
oH22n6Ymwmai+1/79s4klyekrHy8kh2IwadG0+oak/Trb+k1+xErODRLMzcRrWZKyqmRG8I6q79p
CiXBgdkAKVzC5FT0FbY7efSdiLvW/jV8zGvPKNbGdftIju/M4l4KPNarWaCUNKDmq/p+v5dKM193
5tJagYYWXPaPmoYZwqLTKtqYRTDju/x+8cFQbxCTTQXS2VOY5x7bcvte1epIBtxw4FXR1tlSHNOq
SYpdj68VQlGdnx5HLjIF/GO2sBAnjEfWFSCugOGyBGrIsWeCD6z2MiSun46AoVe7VQfDjxZmRahb
91L7nY7a75pkoGVy4B2yxCOeaXg6sZrd6seMjLd0r72xSm+N6hBIhBMLtEic3y2iNqtpZiLwYYLB
2yvrAn1KXlsuwKPqwYOyE0gXLchaZAhiltGKnTtXPHwiicZVWW8ZvZCOLWwteoTCe5LJWQp/dlI9
wIsKYA992MXIQtfquo8lITP4oVSKhs3VIyoOjBernHxVOTrKrgXIAZ95Y+qXFcTNYCdFGdEakdGS
WhQBnoJdrERdv/IUcOmiRXbf5iHGU0k37QBTyEsCM++YNmRVmJaI9Ap1Ng0izlZCMO8XfY68kjgp
avOMbOptBEhT1sy9E55xFN3j5lYI1GiTpLOCwufDGOVdI60JG4afMqmz4hlbQxvMIdiCUYFaU8sr
ImTDqGcI1LqI9zmk57XfS30WyNeIDBNvh2KWBSgVXa4duIl/aITJDXzwKuT/5YdjMdSmACRwlLn4
5uYslpzTeIv2cUPdTnVMILnNGrVGZ+W5YFzmGGa25TT5Ryensv8uMN3YTQgZrUtPxz7lAyb0r4OB
bQQK0YdxGeqkTz6tuOizWKcQK+ahPtgO0rHsnvdgEAGHrItFAuZ+B4zUcqG6/M0FX1ae9wdEj8Nc
bUZtKvx8Ohl6Z8hfFO6DkuIiBYMYYxV4aCh0HPxCCV7QK+BQX3WZ0htlyY8AHtoNlPZWHOTKmM80
mZxDvFIAVezvippoIXsCD/L+dh7Tsiymn1YYmykY9l3OQytA+qKyyxW9AawP0Bb77l6WjJKCBhdh
/JGoiikVJWrDf6PW0sElJXOYmNsIrKQ7+kRgOKnl/5chEPvZHikjt1hRDE1bNU1iAt1fE8fvVyEi
W9OmSA3xaYnvfgpEc9orq8B6IJDz8LsHg2yOh1Fpqs/ocDYWVeprT4B2dB8F2qRRbPU3mLB5UHnl
JROrJRCw2T1+mYbu6m0K1Pa6FvixjXnWcbg/2GESoB8Go94q2E2I/PcElhwwZ8906OOZ22fNFnKO
4ZiWSrfTruLZVfB54ptXD9lRinKR4BsFPP3eJvhI5hy81OXV+fXQwUA6Z76MpKmoe65NlaOKfyk4
ITEYx7CBKc6LCCZbIjByJs0OO9iUBslO4JlP7RlhTNCu3INRDa2hOSfJTOrx137DwHjbOKu3mt2a
/TMprlBDbv17vi0MENOtV0R/IQvdXgD/SYTZSWS1ymFd38pmi0HKqcto9sZhUnIymd/cK80Wo1JO
2+kjHJZvGasxB1Sh18J4cS0/sgU+MW7MB2WbQlewBdQCuy+0DvXfSY45FKViygY5cZTfWKl+fgZ2
nDJLqA+V/TkZumsCisTEopq+V9XO4JyD/Y+1oLxdS1AyYLa1aAunnlLohiel32ZJE+h5CkWBpida
Ax6wxsf7Qeh5rl2GCQ2kLhoVBWefd7Dip+CrnCWAefeApi843XHkPpKztiaOsu4ZEXAW1zgQesYO
vEQRRn/qB8M+2nHEYH+2Fr03CVnqIA80IHoNZGlXj1GjycJQfLOGf1sendisA1pGrJ3rlDNXJhET
4d7/tNa9NOfo6flPcdllP7dtifK0bWeoiBziFOAzOMp3K24NlI9D9rylFMTrvf0btWEEVgajgQKm
pI9EEUuiCvCkWB6Iz5fpxmdAS+gO+xn4LyobQggrPSI9ZW8TAxXpHKZaH0/F+cBCxvVkpfEbIwRx
9ka9Oyl2+yPLHgFK7pj+gIFYwOTR1rVVqmMwjACNHieBWJPF4NT8cvc0F1nWSZTltiMK+6CuRsbR
OFqIuOfXp+41hLdqWJ4haGeYBUnJ3t8cMJjgOR3Lg3lMnnpXm1klPiQYHeXh+0UIc5KnJ/OTXz+y
tvhoQKdQ+ZAi+WDOYPH+JK8609543TUjLDGsE52tk0BOi/fZBkDUXj0UI0RL3faqN3bzsBLaiHw8
j9OHqHQCGbnzv1i0deVZQKiut+8w1ETeccrvI1VJ+pJiqGuv3negCeVtU15o9nfluHVPnC1VGvEe
LkYjXF+iIgUzW9AvRck/KTWu+9fkHz3CCHnUQ4QsNu8dlfVugDCoDfj+lpv0Kze10VdeeLgo6W2o
OC+3t/EDbgts4DagApsfCfPnwE6xv5jXEB7EBv6UkWY5bC+1PBNB3IiC59w0R2R2PzgCOgi7EmcI
JpD31C2hLxK3MkPy+F7d+U3uKaYoXnqN9yTj/NxfgLLiiQx9iy2kSRNmZn7SLjpfA5pfhTENZFXT
AskBYn3c6aqQqCpAtDikWVJhJloGTqsZeglkcezRrPWSdqRlbkzhj+g3RIk3lgFMlvMr8rdiqrBa
vkJOlFebm5MboHKO5zGqLjUFBLEvcpyqVt8aTE4pb4AW2icmJmI47oYeyG6YIxouBMVuTnPskCjG
FKgzh9IGLmb9kfysaemOfTPlMzytEzTvDnduislhdsjn2q5hg1gtYhtRoDCRyQRQxoQShkosNRWn
oek4JcS0AvuWIK2XGLthJC06uUV4yIOSWkrDP2eD9TeNN7jDL96iDl1b4HyKb+MH3z9qisGNry4l
rJwyNB8kPyuj50Dyfay/ygOhlZcf050nezkTtcXLrieC/N+B3J3D+Jf12N4ui1LJi/+j7ZNitJ3q
N090nc77h31lKWgI4HQAuq95rYdkzAlyq8+Pe75HqoEOqO8zA/lKZCbNhFLFElh6sJ6ikRfE4Mjt
EKMcHkZ12uQMZENHIitFbob9GYT3HG0+jAoxG2+6fQG8hdNbQLy9a2s16vqw69AEUILK6Tbv6IvB
zAtYiVJq3p5lO2YXj1QplcG9X0orqds5SbxBGITa5KxfcA7dIKCGUwhnL5IuYkrB+PTRR+fy7chU
Xpx0sFqNfkFAfJpZ9jHQOWROi+DqC2J2s8uipIZyO1gxa5jEgFXiFDujBaTCSCtUYaVdS1DSlrEy
ROCJZo4jf/be0akrHgfkbDIZ2Y8E/Z2sL+0TKKnKarsIUT0hY31EeXKJETPstH0gBZQS55ktiHrA
Cw/7vQmBA721P8XMbb77+J9w11VlfD8RafN6QwgS7qM7u1haZnpRCRwf2E/FMjptrWCvS3f92uIL
EOoEoTz5sP9ZnZwCtwsXEW+X1GDWuvhJH3ERsvYXdk1GVbrAiGds90kvGewBlIxJNAxEDi78pWWD
DisIME0O1JBDNX94D7v+cunVLSqTzckKFK/I0WQb8kXHXy6+Y48zGhcgX4ziQg9weuRVxowwMrWh
PO76vMql1hhDo0jH04gtXL8eDWRrS1ARMVBN06Nacg04l1hMHjTr9Jje2IIMirXLBn8Zik5I09JZ
uqKoOPuN+7Km4M73d+Nm8mwN+/YUjBaMAckCZBQbU7vMzahMA5eZhiJCeYe63wUpKM+CImjg5wBX
jYf6Z96Ft5wWBu6GLwuYEc1+MDBN7btCi/FOI1hfqq1ySsTt/nBiIzfz4KIwEeD/0y3hZ1+B42pO
v6d6bpLI2gPRCT9iByGjfVB+ONV/aOcGidjOTJSYBDV9SlnVpBtUaGoLaXCXcT93lHuCvokN8oSU
QLH8EP7gRW9tnd6tW6koLAAfHMGF5ZAwF85j3mITFFKvwvsvoQ2vZyRuLqtXKSUny3BvZZlrs2w3
wzoCdpK3aL0ww9d74lJpJK9iWv/90XrZjHRrWK5Orji5GxpCDmkV7M9JmPYHVtlDyUXuKWuA8zBL
I6yX/SD7ucW6pmMX3XekySsheUG0mU/bRghT7oNkogRWdt+2/SFCcGFlEWsLgCFzDnYWhiULLya2
H/9t06t61ncbkuGB/5lH1mMfagURyeELIrX8m7aEnvvUsuKnb9AVpr7uFqyTFCP6cofLlv1Fe814
tzvHrYISvsvHZsLCPCuclJ5Cz1v/cPVmihWRKROA5fQhR6VRGL9lbH6BGMDQw0TL2Xr00P/3UGMJ
lk1EN4RKJX8m/+EQmQdHc7aC9yzfMVQoPXkbW1pqYO95zRlGuRdTu5iHVw/KdBjjMrC1PZl1nbcW
qriXPWPNzLUHod8OMSiRrUJcCOaD6I6txrX/0DqQxDT4J9UCXt4W9PGoc3GSP/6Cjz9udeJnO6vq
0gq4xwR1mxPcmpqYZR4Da7c7Pgt+MeGBtEVbfbbWt7kie6/tihEIfzOk9IvsajBt/NVyAsyIKrMO
sFTNfw7+ONyzdDt0BrxKzGD/p49uH7xANRStisi6IQZ5aLJ5LtvNttSF0Q+WaqNX3X93MjrFLaD4
CvzFIeZWNHMvWNKCoY0EyzG8VN1v2z8EBDHcLuJl94X3vh+b4wkr34JwDlK66aA49rnl3u7U4geQ
2MWu65X+uUaPzY6d1mcu8VgJS4l6VN9pXL+fTyb9wIkI6p6QOtCpqwEMc0ZnCge4TzPpbGp0DRI9
ngOemP8SmyeltNlY6ZEa/ff9dIheY5PCOxwd4yPobYlF2GkQxIxQZpcXbkPj6/V3p0nOsBi1IcRu
+P4sbJJ/0gC2xbESiaMFPEk849DH7TMt+kwgmJ6jz2VAjBjYWHws9FBHxy+b5BcExQGWq9y9h6LV
jmk3CH17SOYjo3jn9hvq9SmTJl9cjyl+3xhTxJNZ8zla3OmGUbHsQcCS4CTPTxRFXe+rmUNL2d4F
W56SVMfEDbLw/fY7RUWSaNHEGVuKnOMHicfzjf0pvyvM/rmR5AxCiqCVibAp2l2pE3hQhID0F4nX
Ttj14AIIP04R5d+5/31VfEeJemHAd+twQ/8QOHXOsLwY63t+A/r94R1Bs4kZEoSKYBBBbMFdb2fe
1AXSM2wRR68u4t3BlPr0GaSy6ou5t9l+mQrWluJE2wd8dWFPBB29UHah4IOB/qQJmVR0U3MNdPjL
H+29iJrMmBM2jP8fDZePM+nbme1F48Tz344piXRmtNEqHXBDNjDX67RjaXjG9wa8b6c3xvS4eLCt
bsQF6JEgZzwheCD8wgYUZhmgOMk0mDxLUKSGgnFzXhU+/dMNewc10N5z2gDz0znVZOwBq4IF+o2E
VCU5KVrwxCnmvuf1TxfNni561QsyALN5s6h3v5n/MgcGqmjt2/V41IxfaPFLHBGYOgblA+gIB1x6
FP+wRcIWlb39HdWbnDBm4YHjaM6Q60ykDtPJlsXRMYifM/F48DP35aXwy1EBqQ1KkWPXErrPmYcZ
LYm8W7kaLM1UwfgDOy0pHrVNK8x9cA5buVpiQ/BE9UJrPpnJOWgcAJgVk9BQRO0bjP+R6lfZeO6N
s+uqoRKwpKHZUXx1L3Sp7TWRePINYZVLNCQtp1OgnXlMkjDJOIeyfLt7cA81VBUi9F0xre3+fVw3
4iUYaxqnl4DIaYC5GRzavuvnLXwKe6j9jrk5FfuDFImsZ6YP9PdetEeHBOXHVeUVSITXTsNtHVjD
a+VNfukDLdFPUzPNHZxz5JDgNXWi9fknfAUKi1MK7FGTE3HcQ9ZAsoOeIcqViEzeqYlNkKR29NRB
z4BoyFu7fef9M50XbHLktPm5+Sja7kSAXmJV+mILIzyeJ/SBG/HhmYrMTVVpJZt4xrFPJ06mj/zA
RkiiR4x4kGGoysX/riQoW04DqHfV0edOwTPYKw11lYH4KHPwNDaH4QpZKp2omiqJ/TmvPdfz+p1g
MFRKv/WL4DnjXFXaFj3/zXf4xE0+PDNpcTMarmTixpV1KoW4EvstrwGzVN9ctknLaXRGXexsk9DJ
K92zcM+GB6MO2GGQJ8Yr4KzqsAwVy7xAPt8Q4iRIVbGVi39VkpEXoXYnwTjGxa89MJhn+HQg5rsI
4AqkHDU08BYA/KHB5EWl9B+jI/SYNo7gRP4Mx+nZfFxYwH6joGdod0QVQ8Yjw6SOx8t8N4XB4kaa
5WIJxOTFDC9Xsvj4mPi1gz8L8q96e+0B/Hahmti0KRa3x4a6SbcrHo7Wo0rMqlpfEaNuosLGJIA/
zUREDmWOfcQVpBMysZo08fhZzu/XLpp+nmVs7Sa+tsQ81X+gbzBtCXyVw/2hSFf8Gm7diMCoUMVM
w4cO/mdYjdGXdEcSJliyhTTFMv2tpe1qWUgk1QN4blKqMkKiIRb1nynbN5DYwkgO8H5Y7lxvoVrB
bESIYn86wDe/iO5Q8+OQe2fTjVx9KyszVOrHm7Oz/wd53+zn6vkjS8foWx0EILL5NgcLf4pdxsDc
KDT7J+AKGliENVjZV2UNQSU716cbu+KZ5bkbsngsTaeDpOegcFNMCzw49axXV8JBLWq4++bDii7m
1XfDfKSAk5xOspfU6VsVrAT0vWTT9iCKM10b+OTz1lsPnvIESpvWefMdXrXaAaV9L5SzunJO08vE
aaMQJuxfxgyT71uF5T+Sa6Lw51lUgi25P3ChPdTs4N7IPMnt3DS6HxNCBUaDSX1RAXezgv+2Ff8W
5paO42LkfaC13iu1FvakCNqQ7WQVdAceBA4ojwnWI00zJsgHbCJADMbDaleVr37z7ggMkNK5B9cX
6pryQyLlHGnO/RCz019eOKn+xIOFnMO8KgiO9DfeBDvWh35DdqosLDG1H3LiLJX7byO1Neszl8kr
AIRyizzyBQfJiovWPQqjBz4Pj47YOa00bNzCpqP48Dn9RMeL+shwgIZVlZ8bWnsxLM+ucSFuOdlr
zouWNGpRw5qkByActgnV7S3BeYzipcPccqYFlLtUvOEbcJI7uxLwrQjinvOQFJd4yikNqCpf9mN3
z0A2ZHrN76+pwYFH01TFzZyUP/U7C9Cuix8zhSrXigEdpDYGD6Q77mwoAm/n4DLHqITwOQcg/x2o
eaGKi0PXEevaMidqglq+by2ifYTLiojDd5M1Jr00MJ+e4YBSogouCRCull8wQLm/1oqudPaZXgDr
uZ2Z4DDIb0wnqmuec89JzlcK/nMHp6C1TJNkQpPoyU2VEku0oQBNDI0EHXl8jqOcg45gOC8Inmn3
E6KlxLYZrzZ1Y/YdfYAXu3xMrIVMW9MNcDukmv4dhIuoQtPRiefaM2oNt4sPIfYWyV+HnCLXM5wC
K532HgmrylKm1YwM0Wtxc8wAvy5gTqPK6WTWrR0ChY34r30LCmqSkpwh7Uw+PxlGLEQ2TnBsfEE3
tSYZ0YWlFeU+eOkPRlCm63jI+H3HYKk3UbWFUU6RI2Wk98wz7eJN1xC9HhsSpPq30Df6+x7EFRDa
UuOVFFpkUeDgBPdr6tv6KxAu2biQK5gsNJEidyyjBzFe6ZY8FJP+479QvUaUVFZVcTtJQJooQJ1Y
gX390kqsujeuXiQI7lBNHwGz8q+NI0JqQanOjFcOVJhTks7+7ue8v3EZkMocaxB3mt4HHvCIc6ZE
PQVjIuWxgreoIPBJvgqFOR9QGaKXsY/pJ4a6YMkUc9O9K8TIBps0xDhW5DhSwDyEldixc6RvZm91
16lSfX/ukZsG/RovZp60oz/ud7kV4cBzMjk+8bTBmbG7quScaVeq5v12F4gBnGbci7YO4Bud+8KN
7e4vOwnvhe5qwEgbxDIoR+UelrCJYgSXOpJmJEnjb4or96xCu4OExH16kh1MhMovzMZ84U6MO01K
H/iTfWdCYCl6dYtyqptzowO0RkB91N+QhVCKQFRxhXI+FJfdDGn8Hj10FLQxqACEN1fQqF6eZKZH
p5n+UtKUHFSIBjS4H5gJMIqC7I4Im/umY+6qiD9BMpdk2aEhAd3oLme9nhOprQgKkVHMTsFKja/b
eQGW8WQdwO32xQ1PGGod6LpjCGkZJnoOFkFeQ8A5VDCd3bvu1MSIuLN/ultSKJdpKlAcQQJV5T0b
LCF/KPk+uhNAF5vzB60xWiZx0VGBsfgp74oU71j2XkYUvev+4UTlmeCUsVcHxZ1pNjlvt6f/+kIh
Z9Nh32coIS7uWcbEVJ6zoLMOvxF49ZOcVQdaEUtoCKULcLOnvtGol9BNsmRKAIpqUdzcXkFPT44G
i1+Fv6TQV3F21EZnlpptF9qV7TFKqhFdbGjHmoUNPISYlC89kv4tUiKKI8A9oHRa0d0fQMmDJdg3
dYtgt90CrZMWLpEuE1UA1KUomOHIDn4V8yxCGv+pRGJeXiNyXjlGexcJL2EBDkRu1wFpkBCYACA7
QskLiBIq6+M1lmobzqnrTKxSIx1kmOs8z/OyGkBKXG7ZvKXQGigg181q2laZPPrER7vNs2glOP63
y8YwWjKvCFfJvRAMloaT1eiFDOqVhgGlhBK11nytM7Poxm0W2Rg8CtipooZKQobWqMi33W+mICnm
8O8cXATC6J1ruwMhQL7y9d0r9FOMLn6EQeJfDhJjio/gB18daav9iWEK7LQfD1wev0opr0HNGfyI
oASmoGZbkkpv8hfVYVwHBJuc93lNKWDepbsLJYO+hsiUadj5dcYpcIGNlgMpzXyCaLbka8k4e1CK
H1g3RpkRu3y2yIFNLNaze17PprZ+xTXbgZFRhvo8cQIzzZtlkXODw4KIOHsynrYSd1dleAssVLnS
1/EEiUsj31Fe3Dra4fW2AHjW0obRM5lqjaVpTKmGdyLkhg0dS/Pu2ZHgjc/i2hem1UgpWIua14qq
MlCzuB8/K4ffsMtwyc+FiNCJdAPaQC02PETpv7l9H94EyQDBFFayR12m2fJZQ2WSxH1+FO36YBcT
ich0m67t8hRVGyDRLKSS3prtKlErHvZipCAKYYaIia9f+3rOLo6tMrHrC9skDSVLKDdOxHb/aPyI
KUIqmUMl4iGqyvmB2vhJ73Qq6Vcy/ggJJBsxeWFdq9zybE76VE/FZlO4a+frcY86ITnGZOOxfOQu
E0zCn5JgqBRBatx4HVSNs7r3YycX/K1GmbK1RGQSz/VdWG50/jpWB+SvmADZd0i+HTeT8ddHxSo/
McV6yU8cWelViyum4of+32WlS3sWcaUeLyb74YtoOwitbWMuhGIsSXDUMcLqrrDLcbH7KKzRmGMC
+tXVLFYRXOFN/KOxxpsROlRg49tDfRp6hl/NfmMe5t1ztJeCvi/etSX4+cZjYI4M7ylCPKuSOpOG
+METItXECke+8LVtM7SxfeVEkauZEw0yF2LgpgndQ+zMDxUCQTAkpG1dJNuxXVFV7jTLJ3kUFYI/
ec/XFv+ySMSz8LfkBPrKPdpNixfeVNkYpLZOpxBRc14FuSNVndEs4VXZNGQ+f3esu24K3J8nbxRf
8Sie2QAnI5u3dj79Grra9S+18J44XMDgwnm4XRETm1kdc1vZiECCXSGX0/lYh2GnztSxzexAZf3V
r1rpmlWGiykBsKVnfIZMLDuEQJit+IeDrxqlXeHSQBD03sWggbbeZlJA2BfH5T2ut5QV9M3YWm6B
CXgsQ8A3KvPOmD+NEsUS4O1Cx9P9e+1hXFCZgqaE3Dg2sOSIuG8K91W0y4RNqhbNgJteMTlgzl3Z
80/m59h6bTNThssac8C6Y0EQMUrpXX/15m9Vu05q+9vrMxFaysFT6udZ5dqR2hOjYlELbTULXkfD
n0iVMql9lqjAmIKQP+nhxef0oB0lsNt62Axhb2nfqx9fRFpWZmG6YKo+eyiziwWd+oQ400OQw1D9
2HL3Wb5IZBNuclNmP4hWEegF3VlzFan53CWQOUJOJaQ4Wg64VxKVimlsq3HOwjESCmhu4MzSgfBx
zryCFYoTXFIdyT3bPI65UM8zjdtjBJcGvNvgBRpqudnJXovywPgXVwefxPyBtfQNYLN564pMDkqg
hKTbLXvjSBsfpvrgiX6jD9topDV3i6ijT38HI4onTF2wIyOW/bTSs9xYFlt1yB9cv/9+nAuON5it
5rvYBggBAgRC+Ej4sk0nkXxSH+gfVDG2QO/fyHQaF45s9uvEk5tfZxKVwbk57NEPIuhvqeezRdFX
pGYmopj0qi0EjVhvtI+2lQxeVgEul+t9n+anO4FUmB1sCBTQpPHoU4YD5qQmr/kIt+CaKSA29uuB
oJkc1sNDhxJN8XUJxkPF/fv4jiheJT/cMBI4ftoIjNBs0GxZ97N08bIfBNUqWzw3odg34zXu/x7a
X8hNH++UV/g64FQ39WuLq2GFRJtLjZR0Q6WJkhmBS7xEgsUJJE0WLRTY3xFj3KsRyhOsKeM2PedX
rhskdVTvbmNuqcWYGfKgD+WKyRBx1o3tv9PZHo6++2+hOLj8J7jlCgJGfJAYkjVfe8IuVJFn9Leq
gXmxMwZp1cF/TzgTSNL3zE5YOE3rfd6zNIF5wXHt3q14xhIFK5AJaDDmTKCVZe2jEbkVaE14NF/N
e3ghTwCW3VdZo+GDaoeMNVyxV6lb9Sat6NYds2G7FlNY9Drg6Pde8o8GTbNp9WkDgh7lgagoEOyt
y4snR9VOwm4CJLxX02x7GUj6VG7VxsQXq6E5TgP4rdSfEXw++vRa/JEp46Cok8siFnSwjRf+NLnV
qrEcfSuEiUR65D0wVeyOUtobrSzyZzQJ7Az4LWMnqDtSP6Eb+D689YTI/x/O1VOYHRq7YGkeRGyt
lGMNAQFU9nFBQUIY0y0hJAA/amMP6V8EPOAWJnfrniFJKW0PnMW9Ki5ED8CwKLJA+uzpJwsks7zj
m25iYE2o/ducdoNWNX/6L+VUXoI/kWt+AG1oTyU5sp81Z7K3OtTdyGiGSK65Ddnu6bW2TtN/dLqX
DawXdxVlTkcvLMqGi/zWBPimC9wXxEhM2hN+z16C93skAl4VO+uqqVLeaCFzbJBempkVJIlRj6SS
5zJHR8AvTlWiz8EkNpMs9PA8+hOyX+DjC0jcNCVTfZBRmPFc4CHRjZDEX1NtXmOTDa+v+cnX3OVv
xnbZMRWG2NHjN23ZRCGCNL6P1/Yc5kyw8l0Zal0KeIFjbnmSb8yLXgxsHhgR5LsOpgWIAXWPieGI
gdtqI8VkAkOSO/Lfuilpo/zSzC0HBAMBcvsG5qLdmfAEsta1CtVPM6s3i6KCt6oFzhHmrSR/NphJ
whSGt7Y1JdKPpLVVVRby9bjiPtFXBV/yGr8MoeYWKqS1JlC0mfNdYp3JTJjWN18y4QpX9isgoUxS
11/XOvYn7VFo0mEi1TBsxJWIEXAW/bKN/y+WpumJ9gqmH6IVELYl4uPBdwHUhPNLxhM3YgdDwBFq
LyA3PTyGSOxA8WLEIf2MOa8BB4BFVVNVANLRCdWuECy6jPZVbeLyHqPeKKD0fAaHn35PZhsl2Vv6
Uz9V6UqpV87z88Dq+WoSGjD7mgmv8eumbueXQFo7OztB3R6BE0E/d2AI8lCwP5zCXm0bWTfhRoFi
NQWWhIegp1LEfW6IE0cE+s4l4JITjilTpA7HK4BO1jhPEZjAs6/JEhttsI6tiO3FOPuWWfwF1YH4
MdNWW48BQ71r4I0KSvn9JTsH6xHST7AHfm7+oFoBCqcAuY0zsnbAK+MEhOAQsc6FX1NjDeFIGYeD
gvCynPoQYZmrAv4nPcKx//sOZpqXC5xmcJdA0IUOlANTIkePvVOJF1ZuqbGLNWzLhJY9v+4GDuqU
lXYS/lLyOwcN3fAgu2ABYcd8W9rnWMFgeLVJqE6VooODEcDXNY3VnXkRkqqmeIYTJrB0HY6xZ4al
NLK556LbvEVoAWVi4X0aQ8/zurqlhHoeI5XBkGLehS+GqNzlV81cJhprEu5R6hS3jQsOoSml4bZa
715OvkS8iX5ogEGXYIq5McVwxmFYqa44bNNwzGhbFSwNCKO61nx0Jln+B+EYkzo3qZIruiMgLRqt
roHxViWRnY6chtCH5nbeCjUeF+2YYzr036Bo2DUIg7WTNYYYZvty/ZQhPv/SDlrvMb/5gmL1nvdd
qpoTyV7GkBGix9Y50e3O4AE+hs2ztBelDi3mNhd58RC8OWjO3QUUOAgLmNIZwkj7E/lIQsbXZnAu
qOaCM8pVuf53xGtK7pucVMWyyk/sUW4lPB+V63VQJhxeGxuySLZY7AuNIHzhgKWIgIFvZkeQopHL
6eO+W4kxDRA+Pc4BodtjWFEQMnozTI6fuCgSoFMUF9TBAyC8L9lvEt82MBbdb2x372L086wiUkEF
Pe1qG/Jo4Jly+bgeLkDOYpPpvGA0R+yXYl4FHaS2giNXSLmCL420zUzId5Av1AhR6g+Ih7fcQSfj
9yCQ6Q+nX0ejmL0mnmcaQ8f/ETqPzTu1CKig8gk2YqSg+PRcVfqqY571pbeZCdQQkK5/a3whGvqj
sWfRUbId9NCJGyl/ydTcc0OWHME9IEK9PLcDWL89lnY+xJTwoziAKuHclI8qpU1Gr64uFZ0y2tDF
DUWFrE7ip9TcvOPhdb6yqGHNjiVmf8lC1KYk5iSRAcaVM6aGRqv+efkSYEOkCC0EFgNO73TtHJg3
7TGzNtA0IGZr1n6Boe88PDAoh37axbF+myB3zzaVZ08GtQVX2zMTg14dX2lWz9ztK3NNLIyLRYmn
mmQS+BRS2ceeqUQRcHBNrccRFfoJr87gV+ZTfedovlrfwh2cN0M9QP7y8avZw47J0X1nhgHw9Exu
159+nqAEdwrpI19imO/cQhJMU+WrRxFskAu5/gmQMLvdJjk6x1tVPJgTjwntKDfEnTGc1BQDsIOR
iujChBumAnnlEbD4TsU3MZzD4GmKugUeAHCtJINH8YCB2sX+W0l/ooN2Hig3y04HImjWoYCz0T4i
ZgEikFArSY15fP7u1NRBU/VO3Iv3+c3B67tLjIo/+iO1asRVKY20njjqs21Mgwcwj9qhI789fiO6
9vhmc6MwiVOe69mFGnZQb15bVevB4q+9kgR31RcvuwSXiYlbfZHk2VVe3pOfbQMRkMp+SqLwn2a4
CFTvWv42245AplINVJ30IDTbb69eAuI66fFQl7zY+GTMyfFO3JQledh1ayUWTfZSapAWlWnGc4oY
GpJckE6ovPPD6fhIMPTBsll6t/O77tD9HXwVs30h8jgs48o6n12Z3f3o5juXc39BXhwfPjTxSx+d
LzRF51YrfNP58m1IsirHvtZW8X9veUZ9zi7/YGdINV8h0XGUomSaCojPybwhEdGNDYUiFwMZBoW9
X2d41n5e6ueI1St0lvEf7cDb8CT8hGSaGdPmXdvUS8Djv5QxLs8yc7Ej0xfx9idHc0u9+jaQ6Td+
hL7FcBZU/Nva2slubwZM+K8ahjySUENjXmXY2icqIZmRuXV5JVON9e0LvFFCPuLUUEQdkxxMlsOP
g0D7AzWdWfifzqIHyjg0CFrAu8bIi5637VkX8whs1wsFDjzdNqhOu6pyrzNcO+seDxLsgvD81n2y
ZSv/TNLY4UA9YscNmXzG2qCjj+VA4LYve9qg1c9UnJ6PIF/MrfwaUsTyzhP1XzgfdwhAbO8yHTp6
r+4Os9e8j5+ICDuCvgQepEoZWYq5cijYO7kbwrz1/KB8AFKPkcuwmX37oki9pJikw8uSIDNjWT0u
TpkkDhfB/Gn1jVYDh7wiq2LOfJuFq7WRD7lDcAk/7JlbxWA3NKIy+cOQFdHU+hStA2cEyWna/doz
BzKKdUFTrrSvHXe17iLBnNgMEB39nTtBvnFJcPMP4+UvK3Y4kZ/r//Ez1VPNwlu9I1Lx9BaYOvEq
JB8yDkxSvnXRwC1MB3IoHd3gmrjg/xVZTNGIoLAQ03+1BjJuoz2ma5GkupBW/hp5kSNjKm9wbyXf
NMknpYlFB1hdSgF1GfVlABQDXP9Ih/hsQer5sYwSDVePKNhFXDZ8jzZ4HryIMJmfPa2/EPoQaXPK
VB6s1mqTEnEmxI0nB54opS0EK59Y25HlrATNHiCBTK1o49OCnGsFBoWCDRIqVWQLQWhWxcRs9WWA
syi8lOvn3NQs7JoBY8r5DxeQIOA8aMXottecF1R7HuXMm1Ig5zV7hDEe875hAoqEWAaAx7j0Ztps
s0DjZ0Y24rfKATga0cI39l+WmuMrybUl4mwqPJjHIB+SIPv/geXbUHsMRmyUXHAr4lVeSDxG1C0B
a3v3HfFa4qQkjtLkdk+WxBiCn4KdLBMdU6N/uIEjr6Jw793l26CXCETp/X5zpxB0IQ6ylKDBTeL1
OvH+5DAiUHmGODRs9oE3kAOuKXOkTVIItqvJTkXy07JIXXvXMuXuxjHoHumH+pVdquYMMjBEO/ks
0eX7+NgyK9t5Lrg7eqEngkhSqZp89vkAGac28CZ3tVKhqFG/tsByg/h39zer9vzZs2EcauQa0Xin
DDGnneZJ32q4zQtJ1+ohe3JbHzz7W9hFvr81Bv5lnWHdPX6I3k85op4sKFSUDK4ogudpTk5CB1+r
GgM/0J828vltT1VxGLeFWDOGNhmafanMgTB5qjZmzquch3MdNA6VhPS9DPLC30UJ3QwQkpxR8qXf
0LYbkxa1jnQcy9geXn2lXlE+Ztka7wU9B26bKv9CqlVkyCApaDGX5j5avlN7zD+pPL/1QpVZUd4J
0EA/d+ixv6Xx4pF+n/sHn+ZZMS5n3Vo2VE2PUyEZ8wm2Tku/xRTlWCDLoddEA+sEpOJ/cTAp3NuJ
zAtsD4yyBsj1ZlEgf2fmNXECp+hYGb+BiH83yW6FZfQkKKYS/Cp4FzBfQH0Go/sMPLvDdHcbZ53M
uHvFef0MrlMj5dvFMZo4BJG2j3gGJtMnfcI6Drhib5F+Yok27GIiYc6n9zIpIASsmTlo5KaYd103
CpB/MLX+xKztE8yj3E+w1GqU6rka3WTg6jiTyBZZ9VXQyVYUf/H5guovpte7O93Haic+0JoBPj63
PxFg2bpyKYqgtuZt63L8lVgj8zFwQtoZCD81uhT+qnu1OzpkukpTZy39zIxVfPIgGVL0K5R25Evh
bKQlLuqK5rJ+XTm2Etcxti9yY5ip3X11GPKoJ2Uxo0/Jub4+UwxKY06u2TLbD0MIMRDxSzRSgEgR
z6niebwbNAlJE4uF+7EJUY4ACgmW3jbR4P/NF7bbo7k82EuogNXAtDaHxYqwr+FoBND2SswIaKm8
kiQzuWvietRzyv9XCLAiCo6Ld8c5iLMTeUYWKT0rX1hQIzI8uH9U5dYcZ2gC7Yh1UhtJpsAntUIA
KGDlWFw9L3Vzr0G+Z9EQkInNFeY/NtP5k1QCVFNZWtOgWysx09zF6GrjA2VOQRBBd9EdpJx9fQmN
NiBakNsBJt8YxbKLmHDbBcIrIeO+ClOZFtUaVFhd4IxB88YqdDAZLd7clD9E6lBS69ofj+VwR4oI
SnxwSb2aRAKUnC0MJj9q5QZgvNGEAQpkW7SIQptpPP0/UFgMLtqbzd9O8UF7CzsTk4Z6/L/baIcr
1liMUm4jRPpqy36KBPjCSuR8E4NSJY7PNEWYGioclG485YTr3PwQ+5OUmWMiFTXr2Ey1Hq7SXjFx
2XIPIGOYLMDaKp1ngCqLd6F68vvCcI/HOMsjJc4SdurWx3egJLxGBKqPfkf9u7mzDjXPfa+RktGa
RowSIEt90KueJESzFMgIPuhvNcclf8T70AtO3e6CbEYDoORrlhe8MyMjGpI/zwvRD7XCifUmI0Ft
YOCH3dH2Z68v4/LhXXkIUdhSTkXtm3gDpsxaUItBBSiqDDF8dYgDfA5doregltuYPK1b6hcMair0
AHSjA6LriVrPBTQyqGq9NeRvfoiFt2rwCqLsKb7p1L/gSqQHTFj+rtpOxx36nQbyVBztgeP43Q/i
+XcCFERW9o7qglRBUj4B7yJWPD1U9MLkc8oxGe0zWoRNJM0r3Retn3pQdCxhHqgNWA4H8cnlK7pH
I3Czrw6IpvuNnsyMtY6E7j5tAQSxh+o/jM5IU10cyZoSwtuHlQuhUrRkWNl2HMRF28yq9PkgThWP
TQdM0G+4zFv1z+/rioaRH1hNqGMgcYurZT1Ku9bP/QU2nAlgjKjQ8aMKTxxi7NeJO/syxlapd5l0
0puYOdKv+yv0K9ZozkWaJlCzK9iWdct1uxtJT9D+I5uB+Z8uI/305O97IEvie5oD9TePiHdJdF22
UF3OHBXcW4YNDP86gBf2rDN0RJTfVsKeYSeWVE17Lc72+g3RRTPYJCfaA2bXlnzFpKeI5suFaU+u
FtgWyfDTe+F78MvqkDj1TcioHzvRCnl5KVLPxYSy27TzcIrUFLgzd+jBkajFRELPiXAsgUlRkkQg
vtFsA4k/mZ8LWZyFBqKt6NPlwuKMYGk6TQuZCiBkfnKPmebduQyxDUsU/qp0CdDpolbAgz2LEHUl
gFcmyxR76cpQsnQr9fnYw5e+P2xJq015MLkyRs+G+GfBNKcxs5CXkVVvtf1NYm2yhQ2itN3SUFaG
fRrqR+fmGB+T1z0ZxEynNOSte98ptverNVAn2mv4HpzHcMQ+SYMkwRsaV2FqUq0yVatqh5A1bBv2
feSne2FmMtadiG4jgaNuGxC7YyH1mYQlAjT/4YpRNHpgOvwy1C4F/5hiOLwIZMp4qQnsMeu2qlWL
dpE0aNsHH2E0MunSfFI+vzDi7xxuROrfmfYzOCOxUTUtjHSSYOChLOWalZKrwKO7VlTLgmcRABpf
oFvcq7ZStkAclOvRogNqeQkTheb4Osp+0P0xWf1+QjordnnWwL8hnymmrvGPcV0oFJi7zzHz6g8M
Qdk92jjrh8Wim2Pv2sugRMwOlDpaqIQz1nveNWX3FneA2fYBNQOi26HXbJGHgqNtLrb/fR9NiqTp
Rb8qO0BiKeJnkVwxuOHRH3GZ32oj92ewX5Bues6jw7Sp4I8ehXdofSH9nojW5c85bF8J6+RAJCdV
M+NzOCx7UR83413seq3kGfpNLNBwkQFbVPvwqwssExmAZLm14CB1k9l2L70LWes643j8AnUHueel
I1zine0EpDeJiy3HuLgGdT9YJM6j/gEDnHvp9wb5TOINUmNwhAw1n8DTnkZrMfWe75lO0uL4xC3W
oHuu06Sf7Qdzn3umkKYB0DKTbPUm3Z5NBgPQ0bFBM6nCJ5IkihRdGqScjhUMXT7jwPIZTZys4M45
TH7u9iW07K2bwIEM1wBJwJ6yzeQnEP84JaiMJzkzDfZlsevHpRsFJPvXXoGnuOryXbqYTXKA2Crl
ZeNoQ++p+rGdV/wxMWGwhlCCzSqaohEAMj9X4xkSLD6xOQrNmAM5we9SQdo1r/mfxlzexKJ/hHvk
ax7pxcYFjInqKozZCpjoBZilv19QzxNJuuUzD3kCImB1mX2lWFnehf+efDmxFjO/vgNt/jDmm4NE
trbV1orC3CvdhymAzg0S8PtKbp4jKVV7cPFBP4nSpvT8KqmTXHIhbv0CKMaerQwu8Wyssm7McjBJ
RVTpcZ8n4V3VkGW76xjWHSiaeZqjIvuZzmBtDD78NvhJpFovSpOmlYjXjNU3WZwp+DjeUqG5XO3j
qBdpGyLdFZSML6OdRiqbaSRufz3MBZoYbnWE+T1uYWgN3wt5362a81ehi/HmF8UyeR7+zJcBfOmd
xrLFvOvM2/NrN0ZJkQ++CkwyAXqhb3lKprBfvuTBQLL1y99JqNeEqImpKF4nyJiuhneyscQte+5k
C5wVNt76kxW5CyPuXDyejso+LOzsBPnkKL7mym3ATBuQNH2CrtveUux4jeVworW3rq74l1K/Cf3K
8AaFAdRPRlVNRa7kVTqU/pVIC3tWEGXPuEdbS1Ty5mRfLoZfp1RL4kulPViKQlLkyntOhe16K1lT
sLO+7yfIDxU8rhdM/yhwN2/xaUfq+Q0qkI7YXqYYokUQE0C+0INgrgegk80yf1YqHE/8GcQfkW4x
XW36/iXKXlMjTMt6IehJ/8XsoQa5DbyN9UJvFnAA6PMM+l2pXT/HGZ5ag5RSLFIpRNmYRmXlgiLu
/3qj+nu4KZ9X/7piHdC4m3tgPAgk8oJZXdhUQhBk13lJkdkzhauD2PEHA/thBXf2wL8ay5mMrd8X
f7j5fjdYFx9QiAxfn22jlN2IljB7b3VWx2DrRCAPqnb44WSGqd55VYLH0WeIcBkRGXm26LTCRsjw
Ulk8MrK5aNYv4n4fX0VJac5briFUvRwBnlf1DShlyb37Oh1swP6fsv64FSsMmT3H8+/7eeciyc53
AxKRl9PwkaDyHbMRk8s2aiUJ/1VGLgQcXwwlZzQAHNBYPR6hWytFdyn2fUsiO0uQNUsh94177xYX
QQAU5Fn5KN5vX/9NIv+srcDxlfZoLTuqRqo+vZAlWqW4z4AFYlLZnL6pzYXJC6M+tqMjcdzrFrdm
vYfshTHIIU96/V2DVVUYVRcsb0RFy/ZYukYQZfj+eb9K9SWJNiYNPc8Rn0cwQw5RTM0i8ghmZgCe
3I1rKijlXVrJwWDuvvSXd0F0D7FYpsOs1FSzjKhIcA2M+dLjxNkhpoWU4t67AgSeWsxs2Qs8vqjO
tfVdEcVpCGcDsCl4bv5buoQhys3bFBhHwi0L3UgUajkVHtUs0xMO8za6f/f6rTGH4DMDW2gZHWSZ
+fCwMH+yiOLDp1uAL1i786VV65ulyGZFOKV5JiQj5sjMWg/nFUSpdZv5mBBcBxjFquUTgRmgkK6Q
mT4c4AW+7MTZv1AkdVcyXeTcA52C/SfbX6bjuqnMPzhrXJS90PK2wZRZKiNhngGP3UVkqy1AThdw
bTosCv94VOb1mSiTdVLRiCAb84HGglIMpJck7/hCNx3e+BIeacU8LUuNVBfO3UrOqsVcvXaW9vC0
7khZTjLLqyEjLfmW4CIm05yJZL0RTw7iBjR56JsAFH5g7a5vATuu85K+n6HOM10RmjYLdgTl1M6Z
VGE5MH/0UKCAJJ2u6Yks9Hwjcm08jiZ1HEe2iLojp3ddMFf+1x9AFxV5FbHZveZEnUMzNmdbMd3W
fa3zrrBH/dabNAJYSFk9VCdv7XOMJCo9XhGVByEd2ie3HV96Md1zSeupG9oHv3cFYGaKrYlTJim0
WtjXIa19ZxDSi1ajfBKRWdRXiAbpcaNRu4J0hm2e+J1Zyi6B5b1ZKy81Khuw0+L5xmjhPeK7Yowf
up1LOnVJ5X53Ym9GStYltEcs+hrAl9SgetXaaHjrueuAOx1fJAytnoefDhI+DtL0IIQdioNR9Gnl
Y6Pl6k97FsWYfYBhHzWYD59wM9acHLdAGTIBx/tsvsxB0ITcgV8RD1sSC2tlci/cgTk5le+9V4kN
tgjKPp4Z8IOx5qExq312AfZ372U3UefHFMQW5jVJD6aSSW0FMXKjGY+sykpZhMEvAsSM5a62iz+/
CR10BiDKyMng6hgMsWdscFKJutrmrRKE3fQBO57PG9N0fpq2VU1m3Bsn7PtgGqbO1axhU8FyjNVA
e3aCn/85jNFk/9/fspakDeG9mngGTkNfdDNQ4W2QNgyffVe1elKsAZu0siz8gI0T/d+acbAOh5hw
S/burve5llfrV3+reiCqBkYPImes8eNQK0eensQHHVCy52NkVSY45FP+QQhThXSev2UjH/qQsX3n
RQ6yg64ewruUmNlioB+bcbNNnX4GaFAmJVeQ2jeAVCBWhRk67xL1YtOPovEbGv19KDaqT+0uh8sJ
Zkqgt/lb1Z+C+UP61OGtnbKI5uKndUrTwukrwJeG9K7LcfGPkYIo2fbZ5QPCwKyKm1X2VHNKeKdb
yxyjGneYe+fVnfNvHMe019Z7PnT/fQvqD+RmC0TuqCAtcAIt3y7MCsAt/SWBPj7FwnxmlcTAKHLx
euc2oXd06kGTlns7sSzRbpA0Ah2fX9p2+EGV1mwJdUztBkr9hGKP+FaDb9NDE3rGM6WVUSrT5s30
D1vtHFGbqbKEaiEmmB5XG39bYgj8oGzjEyK669ROAPIvfefoShjClKjC/qZ3zHgDKRYDBvi7gppV
eN9lOqupkKTytkTf2PARZe9YEmg4U4LgSCadrukiGuA5Mdn2HNvqI9ucq/DYbh4UtxlTaZCln1EX
Cz0rx4RYoLpMHKsuZcWGWqdWLFJQSD2kIqEO48BVmiiPE287t0AihimOcOC8mjrdTtCYg3eVwQTn
9pjVhVt+2/j4TCQlnHKED9NgDzXotqAvtkQDAqAaI77RlvaC7+VdsQAhXyWyEiLI1TWqA8ZG/uv3
KRNqyhC0DHWpcHJRpKflXpi42vMx5JEYx7W6xlqxceupowlTiPKzDV5rmER9ONhcoc6XQ2R5UQZ9
OoYcfOX+b5AwBmhYFtYd7jeogYf3nM05m9TPOk9vla+fCgZEu1K5OsY7IzM9a5eYZqtBgEi1gDhy
Kn+8TpB53tJxb5f2XW0Kc0owM4bMVsmVET7J3zmqMVN3mGKs5kbdt8K4wmW+/HC7QALJ46ZtGdvU
tNcxOnvvGiyQ9iY/LJIygUt8D4+jJsSudLNGAERV1uxwxgvAtwVH8oNKY+MVdrGrfLm9HR2uCcdw
MM8foq4xVIHBmrTeFIctHFDBQDlS/6osWF9keaWqxx/yCtPrujZ7pZB9mbSG+9mZJMLH0aiHp7t1
lofokllxXxPq36rnEM1aa5g9fWNbHsJ3TlArdPOKBztIgmDNcXcZOh8/F6Uuxs3Hu/+joiU5/Iap
ngpmY5mMVyNAK5NESA9HG5DriRJWFSHpkiVvav6L+VV3lW7of/rC0bIMMGM8gOupHQUrImbP/oaN
UEsPwdthwXwaLGPH5biRaxMsrjSu3ZcCwRa8LXcmp0sgsopSpr6F+USrzWHf4HmDlY0xIR1NCr5h
3oryQoXOOX13APjS8ms/eg3N44l65LhGEyfkyNoxtTZpzIw6f9/a7fgZZBGXCN85ivf103NWbJcN
o+pklpMrknPZ1gR4L2pyNuuF1S1Y0qrpJDo7fVMrHLo69MN4+BHK5wKgyQNqWKdDbW8U0X17l46t
u8J1iKgC7zUNmBrJJVEWisdRjbnFqqui+sKmLdsyFUc3pt3d5sZ8Z/9xS/lV0hu4w6Yoiv+N87Oz
tmqA16xnZgWimOPds0nmSlEwm6UteQjoL7+J2Svzify2YwzT6+9aOz7Xec7LjYPY8lQKV+qb8py2
9UnqEpW5+J50HVv82hc10Pm6kz1PsiS555WsEZS5n9XWzGf6jIlqwF9Jotei7wc7kXinZe58gIQE
mtqQEaSuM+L0D+cURUUjLS8CPK4CyOba39znW2rcLGw1SRmDdXeZG7BeAoyMqdlrb67lVVupngPX
R9Ij4LcNGQdR6FOyF8ujtCk+Pq8B5cdRYEDZeFx+/Kc7y0pCj9EAlzEIOF6cqXNOyh4Gyd3pEQDw
aDsuyg8hDp6kwx2PbHUAMx01lqdcCrOiJdQl9HwmRT3jqyBqHIDZePqfEQjJA7WeuA8egR9P/nXt
4E9Z95OiBMASERPXyu52yM1JkKzpSObFjh2UeRjtbDy9u/JnY7FgAe2UPybkZsfXBvX8GBUfnymM
EY/mQaYRAt9c3pQGheJg0Kd46yOTXp58k4RSGbzexwOvTiJjPeX7jTgbOlCZGxFDMUzU+cIbVFkl
Ia3juITYzc/5VAQWHDX1SsaeKIYT07fDBUSFqgHVA5+Y0EJHP1uKNtEKeUfVzLLCeIm6WyfoQkwX
zsSnAyXKcXNAputTBoPVoS2fR7usY/eJD0w6wktD3o2ahYzrGq22mJCoIeKlHKBVodUlyqXw1D7T
80fmBS1oPMD+eZBQJwvmlYZgdKnmlu8Yg7WX1RH6fXDz205AI/WED6ob8+CvFRQ5mRj+/16DUi1+
BqMZ2n+z7OV4lAy+IRZ8rJhzoEK2Y6NKesLVJknjhXNTukmchY2OVdiM/oStLaseDNA+ZW92YuVG
O2ieCDADeBhgmzez1iHCOK/ZJqoHn41rBaVGldX4vj4SFZ9rSuMDLF/scMS57ho/nY9h50iGYyRI
hV7xHZKWz4FdEAHlAMsvdAOKFMOatIaGXJULMroeMZSyQRh+5Tq1zS6+KfR2vsJZbx5/8H+tHIWA
j5OllFCrob9It6wunONaPT0Li6e0PLnVANXydfx/XvmuNxHJ9YV4eJPGeFp1rPTfgbAhMbxl7xRl
v8Vy4tk5qwgIN+dwvjg+ihN7hDe8kuN5erD5ImMKobfdiPb7Ty+HXVMy7LmZT41tQ00lIXRtBbvE
3lHiIlHEBJlInVq5T23uiML1+6hdJUWgfx1fRg4A7tmFCt7Bu+MNb9+PucWTQ3Vfj8K0ZYbs5CY4
U36O42kmipOOTAUlpgklcDVTKSEM7IHg1WMgdO5FCH7pLc33W68QGCjcD/QMHAPKpQnRUg3gKyfj
wb5eWCX4temGHaawcREIUJK54PUk1PeR427huqODJtzzT9TGsNLXuewFGcrP0a+f8fo+pyLbXeGM
LTW1dJBX7s14TCJxIrhcJGnZq+XcbLnx0oYcq2wcnKHM1g4jnr5HU+UQ/yYNf3OYyfxs7tVjFyFS
s024OiNWZPYr3V2AlR4mAvUEpjAkShm/oDE2ebpRAIaWKLqeZQtzCKam9x++aPnInWxsk/NjXWrU
7olMSOpc5uDUENP+62V80Ny6IWlD3/T+OtWJJlNUPEodcAfFm0RBdf9rB9FS2gg3OjI5vzSxV/+N
b+vC73ivVlCbCYyFd3dwPhqFNYzi3Umev0Mk6uyTw9xDIq4/dL0KCn0ZMBfY6URTrw+UMh+kU/Lf
xbFA+SwBnN44PKoWMUrV8gIR6oIUiDs07Mur3asFRhSdQ+5Byr6/AeprVIGYuYxWwOrhAObIli5r
uX368Dgs6GrMWdkO6eEr4B+5g99/dPRJ77gtAL2IyaoQWJSYcUnmfq0JCsGu+eM2HKRsiBXesbm2
yB+qxTNQ3AnwnA8Yme+7eUOj1Wg5RBFmfpD92ZOCBjRTbrkfhkDfqFrVbkWoBPRinUhMTR81l3nM
5bs29pyOLR8XRgrckUBwXCUPfhsK+MDH+sLcGWeTw9T2nETmudEn8wWBN4/M3tvdzyk79j+xicTR
MBim/9ff4wFlh5aCY7SOTuJZLnBG14uHTd2TvNXkohcUuQKYeqsk5sd/6wy58PcD+ZN5NznjJNJK
VjogmcOWCtpmEedNf6lv+Z18xQi8jyWQ20deRqj8wnzac5TX2eurTeWCONWmg+2gEaQyhSdHEQQv
oP51FpHkOquAMkqeHYZ/1Gn4/jTukba37ci0cBUhwb+xajjWnFHRO2udsXKNOExtYIiYPTa+ncoV
dkYnWcTo8sNMmiFySE3S9AX6JrOAUbh8G9yRbBEPsts6X2WR77n0ra177uHiYZCQb814e4qgAQYL
WKBA5U+3nLk5JolmyRq4gMLj4RniYLX5b5FVg8Bi0DfND2iNxFBrZXxaAIkfoCLTrvSaDE/BbDma
wVHMl/wUZdpt1PDQ1Q+wEItnkTNQpFl5qLkqECQIx94aQby4E7z+A+tn9t9jhuMJsY8NxEBKP5OS
t7ushc+POzZgORKW15TRRZw/aAccsfkXwJyYG1QBbcA2r0cXqrBASYaOGDG9SkHyynDcJHR+WF9y
jfFoPoz9InYq4x80M2HG3t7tqfHOoeoL3NErhhTFNJqRnjCZzrGcaGwIzMhhkg5+YSP2MRAUKcSd
9oLg0tyDTHqmvebTdN2cB6Ss19C8sSx8r6vqSSAl6p6BTUmH1m15/VlyZRyYMeMsY717HJTJk/3e
gJqAgDe+dRL/8QZCVQSUlzQpbyAJod/Eih8GsYkqu7BE5Pmbnsqii4Ho1Mdy+r244hlCpzXHztJ2
Z2SZFTRFGXVCyngxHbPAQV9WOJRN2LjceQ/NYILoy7L7xNIWKoe/6SPDiB7RLKO0zb7Atb7YXwYr
TB5OVx6TcMcY8NwsWu4A/SAXaUjFZy44/hKs/xR03MHVJMNYbacQHO13fZZ40u+VdarttSdTxXcu
Mwh+JUVrYTy0M8Rz1+ZVSeqPGGa7TXzC4eAUmwURoH4K4NhU4AlfUS2RuVOMhiKzJyee6NNw5Kdh
GIzuF+cxgvJPXj78JI9zwSb9ypokb67NYB9lQ4YmLIZJuHNGX+o3Cig/DZxKlwQiguBjEXrNRU9E
nE+OmiV7nuLbOxRvfp9ishCF+iHETnkma3LChdnqE+seOMCOXxIBhPqNmLpBuyucY0ZkY73l6DMG
ZPYEoSAujv4YlQqjpmqSBkhxOfuYrRcS7q3KfvcHBxBLWYdZ0Vh/qCEKt0q2DVJ1nvwnV0Y13X0n
ty33R4pqwqJElCTRvH9ShC+gPU2M/9lRGTbsVU1vgUd3FIzbjD3emLnmbx3C7u0uuRUd0Spzo22M
qMnZGtzIxKFKTJP8YKVK6oMASJUB6Ebz/XznQzaACpd7O+2ylN9qS6rRIqFdgS4x4eMEzlTkHGMn
Vc5Brr6EMWCc8TOZLbTCfuwMDODYbE6/olW7CgUQxni0kDBFJOSdXGwNLat4I79jc+mm3rX0BsD1
MNxpUmSoMECZoJMxFNcJ/nWahCxuej17oqeJlpkEGMYZkFViexYItuA28UCvnwR2XiNTtP2T4thI
9aHjBIbM587muPt/hsN+dlS7phaPmwjXMGwQARHIGDprnmhIrv1qH4aKrg4C/8jcGHq/Ffa16v1p
lGTfndQA1EBoCqje5PGDGboACdvsjAJYnXRcFkzb7TRUJlekn4Am/HbBh5udZT+PY9wmy115Dj/3
Z2w0RmjUZnm63X61x58Kg8XOU/y6I0Po97qoBp7336o8WwrcHJ7UyaO25MxxveAmTtrrYnNmUaIm
R64wpif9PMczuOUhu1VGeWydrdePDU6rp/4vSD+/4INSE9Cijex1or4Y/n1zuD5Q+NHvdnXckwsf
CiuGOLdqh0q2WS4VtbwQEhY5KhLa27TYeAbuHe+nDhIx3thbJ9UT5phHaC/O+wV+jr/mvN3Dur3U
VXZYxTNWhpY7kqZFvkzuBEAQPPgAL+w0GYaDiIl50vK4g9YCMjt/pAimd6vqxZvBzm2qmhOQUqHg
NYnu8KovOVDLbuBv3wKmZPEmzNwrMAQl0SXpkNyfroIa6fThhYIUS8DJchvzQxBZMO6PpCa4Ntwv
E7Bpywt92HPLOhzJkZsx+HBn3rE4cBm0ix+EfYeA0M0uUk/6/e88EcR5xGYX6iiG7I4dA/ps1In3
TgUx4oUvGESntOEJmhhGk5vlI7PYIdwmQrhq8F2E5qYOjTx0DHCVggC9VaXVmNOJy/SRlLUcuC+A
TeCTyagBZXXBsPRJS4IWSHTVeMMk6RIuOXOftm9qm3o4AjFWafiKBN0y0ktDdtZW+xD2JLd7Sqsx
L9cNR3bpu8jo3NR+76dIU9+2pusikOStqq9JwXQjEAaB6K+YhwqfVORjTevkWFMy1WRSYjZ9OOHs
oRn4XoQpQr4PyuEKUuuqdNhRwivKlv6iCmP1dUbO5BFQfRzv3tQaKnv9QKmJyivdX7SVvDa1S73j
fKC7q1mowO85pamiqHM34pob8RplH+7LFheEqMMipcxr/EcDOINTCgz3V1aUf0mvwW6XQ3RipFHy
C45txCNAZGTt/V+K2W8gvZfn2aWEPZg7OXtwvyyLakdmepwQ3ENQ9C7yfNxdvo7cpbuFm604lRM8
rccMT1EhkZzT0Ha+PWK1tW1hicb0T01zvHiB2jn5CJqfeV2kkk/ZPpJW2RTt2zvI15zHMRsEea/a
WkfZA1A77Bw1S2OEEUCBepPwyBJ9Q4rHGxAM+wvre62dvXeNtYQzcbLKyEdrQlv/FYKjKTHZxf62
ZX90RA0HlT3NC6Wpamq5cDnto+iBdTMNwEN9fGeHar0LIdAZJLcjLrOvCwx2gS6tK7bGhgo6DMs7
WmpJWRgU6vvuBtCOqKKLmpExczcs2107mH1rGALJjVoxHxFQ5Ya3PGUlyRGQjHdR2kn6EU3f1nj9
CWZi236q/6T/c9eKC1FpJRqFhtNPwdJkKmOhxY33fQfTF+yUgChdAcEStPKjuvXEIHkr+6McEGSQ
l4wiAYWGznBtke0tEgZyCTTH+/pIvGB4t5YEbNOJ7hGUmK0ynPSLAMi6XCYop63p2u8SLgU3iWP9
BMOt9YMpx30Nm3utnq3LNKh98uPoBYyxlAwAsm2dW6AHOLdzmbYvN7uM928xtI/z7jZT5UBCbTAf
qB5er2NC4nDLyC2cH9hVDwQpfc28XVMQ2QQP0voIVZ4ekiMw5TjE3NGbGLzm6wR3rcEyd/WFYBUK
kZd5cmmSti600ci+X4sxU7+omdcE54r6j+hiQBsOty7OENzE2kgF4cxXGDmH+KAxd70ugsMhUiBV
pWqjM7sjmdjPKuuv4t5MUYMjdzJz9ae0JcFmhBU0L6PBE+B+BYSkqXPUvhMeJWxt5Subo+kx3yZ7
j8iO0r3VymIUf8l2i4sWT0bZAPksT1HP3TNDYr/Jd7I2TijKvJSjR94c2qlrhzfgVG7W0quXRBaH
DkjQqs77oWzu0DMkG63o/a9RnKyd0EQDaGP7z0OUqUJerD3GzNGFDODFvKrUVbBsJsoqVeZUN9KA
PGMRn/BPZIuQeVNG9Jp2o90m1H8fFhwWMMFmWchLbZ7IDAI9gWTUTDNKHFDyIrG1vWdvOPEwZf0b
7SDg0Y9bGuFjy0mkTateL7iEV+LCMO+8uGC0xshtEqDZupZxUuSU0RDzIjhfVfx/l2wJ/XJUgXJu
UPS36K3tGQvcBqbHO3LIDitTcDWyjCPGpJWTQDcWP6KvZDT5wBqJvFdoi25vgg3KWukf3+4XfOgm
fjuM7OKn0OH9zgKTqea/8CzUr+EgLoLsTTWIrRjchbn+9e68EAXBhitQ37dZGUYzHWnLiDoVzgyz
JrFnZfxQz3JhSTEmvinHA9/Xi5YHuaizFDIT2IoHN74So6Ic4vGWje5uHzrX4P2fFDanwOtBCqqj
rhboJgDTla4cs/IAR3Ia9TeXCRcwxUSYv8s6C+GMaoMgYS0PHXrQB24aLKvZkz6e5vgqozd5i0q1
iBPtGyTI0Ep88rVkWfGXgm8gnLBjaEmiWfAy+turGtuuLCOz2KjFo7QRgEwxZCNjlDB0iMwXFDUB
qgelUXrIwTUKepMbKHr2OE0GEL4v8/H1AvyuLlNJ3py41iAppFa8DfRcCJS6l4JchIxRq3ZH17Zq
AI6Vho/U0RcF5i/5+23dSaSoxeMPl9XFN1Js/GaZM7G8tQycapgk+PHBiUS6ioHkIlhmgTBCK+Gl
cWZkOLQMw2c9BOmGRPFybRlFJniMsUMMWi9qeYJ7SSXrB7rrM7OQWWwpr2iVtDv1pHSUbUy87RBe
DfsG7icOCFs+GXyfljOs2rUOsxZ+GClUdXdoXytne2shjv8X/iCOe+Ncn3a/xHVmGLIEM6mEsUXP
RdbOA+BKav5oAk1erl27HJIUQ8KNM/7yyMlocJ00rpml2EjMrHFg5lFCjQEX4VyzdhLPiT0nh1WI
LPJY4FMcelNcQZCd5RrWVts6xDYZ8TU4CG27dy1k3cUbyc2KUjc4mLQtKQUUjWj106PSNWz0YYF5
kwOxTj8nUOGxELyZbRDuDh9CgLf54TDpNdH9CK5o1+C7ORoHwLw4eH0EmZ0pMTnNBLXT5nZM02qB
AYpHklgS17kFZ9geHP+XF5ZrTrRB2SqySlQhjPhwGHqDJRArSFQmMqiGhg8MqrpIGo7QXnUYPUzK
4sw/kYUCkxaeAO6EaJGm3poqNmxg8Rpsi5O77v4M0JiWBwZ2Z2QJxVWP5mPNlzeDeKDJJb2ssW6F
L20LtOqrlB1USPF+U56ubAspQ1ogaeYC9dSJnBcdCwKbwovU+25OibQftlE3Bb431eizXYZQbKq+
4/Kd6BAAenGlTi9BWX2MV8aNGJ1MKvxlR0Ln8pqyN1wjgPldSY9WpZgcb68Yjoxbj+yTyQlSv9rw
SvuTQUJv2GG6o/89ltFQq3VS/eYApywzo5Q5imWlLHLtjnwTAXAQ6lgoqszqKjuZkOkiY649Y0Yn
Yawp94/o0qj3f6jt8YeT87yb+aT1xgkD0h1XKnGcu122I/mJY+Tso4S9QH2GsUcXTm1w1em1LgZZ
wPE3Mg0oFOeq1/DAIxWLaqYaq3GaEbI9XUdqYWpp9S5hd93MdTbqYlZ3GR81mHkQ33fPir3gZAqa
lyMJioyFFkHhUhoUqgVhahtosGXmdqZqaKmO7ubg/OPh7ceVNRACMaD6ZUCVcrF49ekmZh3Oy++Y
0lhs2fyuVudmHVQLWS6EbT9naxZ1KYxzSxWhpkCvYQ46UCn9aSedS1SutV3Ga0kqsRwi6MWKLMnj
m8qRXDRnrlQZMTjPk62r0faVYV9iPcAOMuMelnMjLHVPWX0JcBlXJ/ovRzDcaN7dgnc2Ay4G+Zeh
1cdDjN3VAxWJ1+tji96YFcIn1i3m3e56UEYjKDFVySuqqmyaN0UU5bwt4HJz2MsSgFAsfCBN74NS
g0nY4K3Jw+I6eroDTTTOdEF/tB0NlGeGcmap9hRHXVgFOo54PvnEBkR32bqjD9/OLFHdcUU+TShS
eRjIiQPOPsKN2OkUhI+dai/2AL1UbkqN2KgFYnjRJ4WS2VYYoumdzRHgIX4HlUGfpEZQEaKIC+Oj
xsiqhK2GKUuL4gN2kY+G7CJblWrXYHl1x7zgMQKka+X6Vf6AZxNwjrTK7JqxgOi6tReFP8q7cynF
KYNUYoeGOuWjWUkA/C7NHdPh32PWcDVLyaBCEfw0IJtly0iJg2t8X7wCrY2K+bG8fohtPIu32bgW
lrl1e0eHPzJrQWnmVlV3+M/Z/kOrPhemnh8oiSKrYsKzx/z4QsAvktqSmdwcwLqjpCqx0JaNB6mw
vrvNyqur+zUP9BNBKj9/3Q8mLTAWLrd4Q0gLeXL9CQ6JhRy2lNihBrAqFqEgKN7hOjz6asuDpqsJ
IxaJszLxdZ18+IhrEA4MR8sD9a0E4yV0tgokpwDzZhqyiWSHVgSEvEI23tuZFT2ZnINPiSVXk9x6
QLN1ix4O8AwGUQkV+ESI35GBFKx1TB8gchyjkQM/nSC+bLl2ZBcPwP7QutfwFWi3qnGE9KMmaSi4
x3Ve/Z6SKIVa0lh5o3Hnfxu9ejB6dsP3L/MmLPQG7BKV2VaEbTd/yL9rZPLsctXbTyw2kLwE4Y6p
2z7lJLdI/II4uk/VO85kCf4N5+nYKwJRsfMkcohL8/r6boEE6gMhF+2Xnu4kN/NYRuPw++lZh5p1
FkZIM1UJ/sXPYKB0BZmEN9TS+mzdUcoPPYcMS0HUN6VWYCrxWtaVSqcxzDNR4wMfwvpUW0Ciaill
jDCGlREcotos/JQZqG4qMxVg8/e0hIxB+tMwvS9L0BxXbjqPtjMSRGc14oppcxxipRwt472zAYux
p+2fXWA603kx0wRK+BNUpieyDXNlaVm9yAC71IXF5S4yJ3ZXQtXVF3rvksqY0pTPTSvhDog6aeEU
XX57hx+PEqdJyfthSZv4jarm+eab6Ekfoq9XFyta1JJR6OeFd0PlO4xEDDtPno60+ITILBJrQpqn
2rihh8OT0+mohCjXuvKRTNJiisluHtwILMQ3OcHezf3MAw6Tzc50Z9/2xEmkVvjBEKQ8vx9VmzVj
6KrCyt7udzf7VyxhlKDWJPg46J4uqcQXEW26dlBUV5sBLUKisSLGDba2mDm7UQa2HeSr5PSieOuE
6urlS9+HXWxGKWTDyavm44EmOv99fXmocw8x3DIJhIi37nclf0FC15J+LWsF81mohJ8nereO81O6
k+7dgFyfarsG476xBLPQzMjZkO8STd7Ujbb7wJJMIi6KGJB0uid6S6lLioxltUNqdlvQRGcGPiV3
oYwVJPmjetzzYjL8rx3ZLTyYahr8IEP8/dQZIsFJxdR0BvfcZdPpQdRmASQZ1ojpSVht0HygH3R8
fUMVFKS1hnNl3o9y2/H7P5vyvsp2jGbayhEHcsr7Rc5ic81EA1KHslfWtIWn/yuCYDuJwAVKgi2+
1sUqHxUYtv6ZHXJ+TfU5iFXONZRkfBBFygV8ObqU2mYeWj6uJfNHWHPvzmIxBCEpMLwYwZkWrD/V
FoG+KoxJGX0Z6GBV8Mp7d2OzpfP6ECR7teIT5winrREpVGLNGEt5ulkSCz4OQrlqWj0IJpgCY8ZV
6xOixowE1ymNoX+qx+DWd+H7qLZiqCiLpzYuCa4BpBlSV0+MtXdM/t1CR9lKgYG2wDCyizG2srmY
kCBvXSOn9ddMAwskyyKy0piIFaz30D0t0zghUx9sWk3vehviWwy9w5s1DB/yfD1W0FKSq8ZsmYT+
hQFrOVuVwi9G5SsAfY/4Jxi9b+JIq7i3LdBjS2INr7kpzslYEFxsMaztMzwGpwxOjAd8LP+4/7yV
vYASuw7pv+M5rUuBqbyfEI7vULJJJuvM9PPyHGrtuf+bwsZXwgMFmWWCUo8D9c5S2eIpPtj+U5bu
LS487tjlqaCn5upvRJOl9IpHT0wB4pnCViFtrYFa94FNDa1SVz8lT7uIBO7BkdotvfikHVQEXzI1
k6OG6jGZLWGUq/PRlM1mb+5p+RP68TpwbPQG2X2jPn0+kB2xVrch08dt4mGWJMKOdUTkWZaVayen
Jt93fcqWxyFuIP1FTWy+NTqx7wtOPSyVV91YTxIwYQsdrr7ovk0sFn5e7r1mV/clkMnZqlbR+0YD
upRtqObppNRAYKWEywfSgKeH4BCwivVKENUrcdRORnl/MdBIHXauQzpI1kS462YRxmL2+7XWy1de
UXWBrwfncti0fr3CeOaabKVuuGdTk1inWMfpjoBLMFRrwgpiwPuvj79NyOsGFBQj/Nt+svpPQsxl
bfryPVV/EV+VBLfgs4uzzoX7cQxKFWLTAxgwt9BoF/q8CCskoepy3XPnEgkVAYlx5e+YD6sapsge
+L57CC540Vjss+xNwqln5x9kt3o66CF5nMlMn6CEpDwbjbBqEFgLeOtzzSztBg4SlGKj5sEfxrXO
gpbKiM/dVPpXt6/1PeLriXeXmidYqFBCanbbIuZvc0KuiYJEp0aVD/tsXe1H3r0szAfhbauSqleJ
I3bmLcHnRyCvSaBVXKboBznLMngTer2AoKcUJ8/BBnB8NpOZ7DWys9TLpq6n3+D9chb4OxtgrU0M
mHZMNUnXyCiXjJ9PQUq5S9BltMayo8mPCkL+wWGD0DiVR/MMm82UV9KTBVow/VccNSnMck+3Ik7O
9avAPTNYva3hb9jEwbCKTkrpSE1OhG9yBZdovmXiWPpiaCYB+0xYc11GJelJ6DYjQuAOrvW10RHX
R87wjwWtCtIe+9k1ct1Tl62fjea0Y2fhOzAQdpdqs9j6domyUEi+9p0km0Ii9aBc2YmYByGVkvA5
G3uDtyfqJjzNpj4uKDxzudoUifGsYiRG6C8wmLCBNQSo6DgqEpMSh5pUWqKj0q4lp611haXG7zla
E+42umklgBHBkbJHgoL5J7EFTMXRvml0iq8xZsPWafMf+FrBljSKQXmouKROok3NfM93jlXDKCpd
NNX0WjWW7f/lQhdt8uhjVPyIenFIcik1LaK6eF1YqYNDdSePYOP0lOOHcobf7nxk/VMU252YxizQ
JnLFAw3xp0p6iYstO/CULlSt1pOFLAgrBntt0i7XJp/+ye1BYUouFUykNLh3d5cQ9pLe+ClFYXuD
dxe51dv5cL4D2xt0gPbJlj0mdaf6wAXxi9mnU6MxUeWhIXPLSO4IimGpc9B87YOoZG+6kXiEYHXi
YcE7UJ3mVuA3lHALLBDk379RvZI9vC3W3/EDO05Cs+Upgh4MNhrwLakw4Piv68rhjPOEAMdG6png
tYC6HSVqL80E31D0NSvmmq911HlltsodutSLmbklNXFEChdVkWEn+YB/FPDX/HO+UFjxl90pdP2J
MSraAgQPh6dk1RfuKi8EnH8uLDt2xrx+7aj+lHrar3SqErnxaefTuTjfL3bhhES3kEU3mpnJJ0Cl
3fVo3qWJudck/8rl8WBxpln2en314nxDq+LMNJNN/xehO6YQ8eQXZ7BKWhf/QBenqRtkb45vjFKp
DQSmUW/dfdow9B6ROqsZxau392YJjJjepG3+xbQdqUGHsGk/k1bYq4rVos+apwO4oeUYRAHkqc3Y
jnmqumBpRAf/QHcTmnMt3D1/agZCPfALZ5OP31L8LUnLxi84P2MFsAgtkHDobbnyWfGDPiJeuPbp
DefGvsY4RZmBEx5vMPjrfqbgMttycGTbv2EuSaORrdrwByWNSPQVnzNwPDOtR9bGhVTTgNY+x9bG
WP5dEftvrU4mA5oIe4wggflA8XUDFVeMFdR1SqQIlfR+zp+mJhgm4gVmxtLK3qA5nohDx510cVBx
r0geFkCRLXiCmFbRvU6iYg7opOoUyo9MV6eDGeo2Ckkh+SdhDjD9AIwpjm2qfaiGp9N29j5ueaWJ
t6IdtahhORkzpUpnI9xyCGnPFcIjJSYh5xbRUST1eHIPPhIpobJc9OgkwgzQ+hfPhqoPildpopkz
aeE8vCw26j/gsof8nMIoCPGEpXL6omyLuRTSehhng+aLkvMqKFtQPaLZiUMC3wYmHDWQzVqJuYH4
qFMaSgLA2s8qQ4HZwMpKogcvxqtsKoDxxJTkoAWWXZEJCdUtYxSOEKWazABVK5x5bEkzAhXmSGqQ
HFcEw80OQEzht2GW1DqThtv8mngMi3bEk72Ow92BpaTtK1TeVabNwu/LllKdJeCivmmjh75WTYM5
YxbWCTUHIx8VoLd313zLYCV0oQpRiGy9AVt/64rupBLICAjiVvS9r6Rk4swA1cDVlfSiJCwt4q7z
mFzJPhUJzkBruy0k7XbUnpoxqVfOo02rl+V66zbYNDv4YZ5yJf98Hdq5BevXxtrev8JRh8tARUwD
U5NqchH8KVJEjdWOABOBJEagigdXGoqvxaBRRAnA/FyZAe7xAbXMXuW5+gqkyiTMexAWInyMs31t
bUhz+4psSdWagkRf/yiyz2sgSB9QVLe3H3+bwKP+fmE6epGg85zDHiZlN1996T7zQDOBLMWaqPY6
R5TnKq33ZpZADWDn6EVS1kq5R2WPf0mvzd9rrI3NLtYnhMAGx3mLDbpk+RaJ5K2mJ1KOVPFwdr9e
WN8LHx6orytzIGXYCLHCMaZlQAJS3mLfegkxvhia2Gj/qvQUtFYSfz7XI4Tqb5Gk1jef4Xi2+eV9
xgC0aIIOvodXMKMIwizZWScgcadBdnFF+tdyYmc0LHOJjRjWYJ6YGSWxQpRPSB9sKmYS7S94HXpB
3L18Cf81VrkFwXDxRjyVI2k5nx7dRyfAiW0X12fp1FCvppcNOVDlb+2PQJQK1p4sc1ZDILACgq6W
wDHTkWFnWswT8qF9hMZotfM460oTpNbvSscfOjYdwtMy/JNpKdAUwyKl46Kq5d0v7AiW0hh20fGG
IA7ey7oYIDpFp3dfqY2uJjkEvDkdg/qG649sGMm+TR24McAwLwqSIJyYUeaZplTZBr2++M6KF8AS
LnYEnJ6bPlV/pmjJRqxHyUi2LdPoHuMY2iljIx+dNYRAFGYMTX0TIc5grNcYKCQf5EeBh4vkaD5U
ml+t9s6DczWHfoiC/OXNhWiW2Lo40Nf+p4NjCbEqCqs5HKi/NV7bPayzBSsbmeHS1fEM99wTE/bS
BSdxeyHU40uHi5q3M4PiZDFbTDV+PhEN84DOF1dHTquBpZhyyfl2DzYplQ1xDTfBKFFMp1S5LSFl
h0lbxW+Cmi2FAziPF7qnjfOx8qKWFXywcElB4GGmn53a9ZpAp3s4G1jqygjaqKyxODSbD3+jwPtd
iK1etVaqeTCiC6X7U8+2u5CUnNHHob7ig0m0ZAPUS4ZG2btqlh1O8nxcHDlKc05xovkpCy2IfMst
p3cM+a6mI7rts0mwGyA5u8r+UWRad0a/+30/8nxvqncVoqNPZR9vRM4czGNS6o30fgA0CXGLpqvu
pu0ns7EsYDZfAhpxbN1/X6yN/8VTrsHuFhMiw4yf7JUX8C38jBKHuoDLd2Y3Wg47OImp365MRcs1
a41AIc3Hluq/54z507lBxEdnOswVoz8lqlxnscjKzwc8UBevkF5Qe7RiPxfTCZ38vAkOjoA2RSym
5/h7+GsH56jiMQ9MMfdWM7LyZ0+mfwlWQUCejKw/uf2CFFaOjR8M6EE6ysncGLXiJqauIr0DmYzn
rlQbvWElzijEeMHa/jK58VBbR27JnVYLL3FqQA2ztwiCsOSCfIwxRlpfaUsfN3ajUddpgOCmf8W2
PDIX4sqn2vPMh30v0U+Z5v2vhRylonPetU3qQzdU+wmIdzXYTphwKJQar1Dz18f1enLqsg9MaSvT
zLlIj5TzsTKUKhi1+aVfFw21+TSR+Fhqe6sGKtOsfQ5X8Xj4g3IzEc325uyCPkh5N9jQIkslJ2Tf
9+5ExGpKS2Z5uEn06UMAmpqQCYTWjSbNKNAX1ArXL7KYTLgGNMWI8bqzsBRSWtMcdmw/yGhMWkap
1bXisTp47LvqCtJwxOiwDV5EAO6cHc6UEhIAq+Wr4qzrnI/YyXvFMN+OjOcbqSPEvJwbIQ7TaV+Q
5Sz3/jPINpb5FFJT5eJnrpVaAV1NhNmxr6TWBGR5ffsa8NnUNAzeTvm6UJiAuDEpu1WB7wWFowRI
zcvx6fd23M3m4tDoh6J57am7Ccv1IpMDs1C/QKDEpge9Bxz4TSAbKt0/6j4rfGAOK/QlT3IDhdy/
p0Nz74wjRe2j65Cc73TQv+A81G6z2xDQcU5sgRK1mA9twHTlv7wh7kg4Z2GoI9EfZbbfQsBLtwPo
ivjt9vzrf0TSK1i5vfFslCw/oONzEPF2w5DGG3WWEKrnSPn3GxMuzDeYaWt+8zEoyBy7Spoar+Mn
Q4aoyg/wge1EjPpS99gILkrCdDu/P6WO6J4LG+rPM3DEQvIhKRt80MKOV+kug7kzgoE4dXeaCXz6
4ziGiPwJAPSqCjIKa3SLxDwX9QpTgL3PhOOHenDgE4iAZ6/vO1ehf+IqbNaClWpJsWtlF6OVGzWM
yu756XvrtrjNLZwxvjHz1sDYT+1EIJTAOMBNXiNnLjA9JJw0lpRktzdYxCDzSEPiOU6Uh/SN2xYP
PtgCTVa9HikhQeGNKg3aIOGF5zQroqpRfBa5FHCleM3AdLPen4uKEOGqIUrJt8mBji4/AkI3fK5i
PKMVMHsxGAbI/iGlb4/rw9vsS2v6zncqat7xH2kfIC8iCi0jj/LoCvrGVRa4E/M9ZYP3loP7oPZs
0XtPPeBHbs1CnCliWhZMjQz5KARo2+e7pH7Dwmi4Vng4HyxVeYAbufliVW5wywEKthOBgHiPIOsM
ZvoObaKPXTgwbpa/tJFkOndZQh4Dp3pWrEZJ1pQL9SIKpmwnqs9N4vKueCuwYtTcSG7GK6qKF2rs
fveRBhVHPU4mkg90SpQZ2cSDzCypR2Gj5mkAamyFmxPTKLRzONahqxQ+tVppQnrP7FZj10UeocVE
b28WNJhxTGATjBYQa/L27FAYXS8eFvEhNXnbUNFz7SDPE4XAzg4fvJu2J+RTtZNTOsDr1aZiUJqO
unQQedJqtvlrjNF/B2WtoESHh4DI8bfspnrSNve4lSF89SyDfbyJKQdKKglObozrHQXw8ivIHNGQ
aSV8kHk0bVg3zwrKPH2Sro4iBkgDSFsPw/V+Ut0RhPiIcedD07t1qAhTbGc+T5kVcBUdK824/ohM
vlaWP5COiffadeyn5/RZAdpafux256NPzTDTNaMe9tHZ141yJWOfK05EcT0b6SmU0/JTKBUHip5G
t3q5XRBLOIIt+d/ZMvSv2Ul0kPdVwwX+ElpzGkpAixrXiV5eEczufXcBEymRWvBRP2GMxX+dtciX
Hdl2icRWn5OV11Y2w/DS9Q5SNPPX5yS54W2N7oa1UQSlbc95UoD1AOaaSC9EOdishB+yW/Y48TCk
V/7J2JNbg0yb6QsplaBG7xCwxOXFoyqSW6nZqVW0cetUaLQCQxu4Y8KDXdCDzn8h1mACdm9aYrhj
56Ir0TEpd4DUYiOkC9G5iKsFkhBxYxrxAiif02hhDWlBaNrCeJDjirHxu9oaHqTHvuK07Efp0Tsg
yrKScHKOOyAZ02aQEc/W7+0mEXxnVi8Sr+N4TzSg3Aonrg0Os+Gol2QmgkAtZK1YSbdRkiwGjZ0T
/3c/OxCAxyXicVPoZKXtPq0s467qmFmVKX3qEKR/2kaeRIhy1PS59B+Dkxr4Es3ylbtZlAUuMG62
GPfu1SYLEKV+SH2OvpfLXn2kEwmQEwNgdxGRZWpdvGOS5kJl8pVZD8TIcph73rXW+KXa1Nt055e7
Ins+RHpZn2lFE/sVnxYwzX7tP2XeMOQ7b9fzJNH6fRBF3+kqw9FlCoH3pr238FRGLOPOaqppKcZu
Z85nwG0K4J2HfPaUqPCoR9cHSynxj5ZeDOsywVKzZ8Z201WzxnVBlV2zXp4IVmUDAdZp3ILXxDGa
WLVfr2uS3STQgi3i8Z6tYLnccFltTLZ5lkjiFmYSY3kU2fDdkjUJXl61YLf0eFxOLBF45x0SrlfH
FfvsXTzBmjgEJWBb/m40cejnJVV+DWzqvTNdat0NeYADAgzWNgKurfwLcTo7enONrVxWGzTmTpg8
IWXp47KpnvL33Hz4VrRh3HJsZbj187a4zoD2vx9MOjRUV8X0i9uLXkUaQPpaMhgMVERF8to8xGhi
b/u7OYcBEsSxZ+4/2px1scB6ufrHByT39TKaPj1+F5TUloW4tECR+BTbe/umvVkhYldtZCcqDpP0
yzu8yy4zCB4mRRvTuItS8m+B4b93Zv7KaoZyu4q2/u6AeZ6kcsuw8NAILew6Yb7639doRE7qwbnM
MY5DF3y85HMh65tZ4sH1cBZzyytoCZTd4W7Lr/C6X/BInvcMgaUSLJN/du0FYO9wyfFuR8HR2Bca
0IGT9P6aslKApCWbZDP697s6yya5vVnIJWvBXcQ2Vrx9OogdFNqYENd0TazzhRVXjp3R6yi9YB59
74eK32ZoSq7Juop9J9Q2o9u3grkRS/nLoZMvR/4pLtG+jlo2LDsvGSjbnn0KEe1pzbH5DYK8kRz9
DsAJkf8l6pvhPOQBc/Ol3GOuEgUSjJRuk6BKYfCH4Wn9rP6kLeFVMJtyKO3Kcu/qpfsqquXG1a6r
MVTHyks78l6twUFaWWHGttJM1ObwvGU0Bw4LXvHi7M91+h+SMGunzK0fxJCqFZ89y57rfz8U7+WK
e82xIuRdwxgMvdIFpQBNgmK6t6L0SoJI2eVMM6C7i3/77G0q+UgiZEWh373b4L5yuAxNuk1pVn0w
1Di/OM6VPZ7q2pupfw+dmND384G85qi/jAdjYL0roojPyhV8hY5R3/iWVd+DdrXWxi/Fpul0Z/xA
w4SWN8jSZz0GfniT66Q0IXyqrUyVrnp0AUCLPC4ILJjKY0PJQlX+55QLodOXTJGNisP2+Bju2Dsp
WgumQO4a60jJpJal7EJu9r2L+37TjqiWOiJTfU949xM3iB9XV1ovYhYwcd6NcTsZN/kRcV2ANHuk
r1Rc2QTDhoFRZT+E4hWQcKY35bLmjCQGSqBsW3Wim7mxuGtxzd8VxG+ltEz/aaxVxJZf2SeVjSUE
N0qwUb3QK+tot5YnJw2orw/9pWObHOhiBm50raeB0sIyMsbztRHeWwEYIcjPoVO/p2UcqCtI/B60
t5PUQKzEm+Hu+Xbopd9gR1oQb70Ear1YTfgTMiuN4Da17MPY5s7T/AxsttBxCe2pR4mtbI3hscLN
20U8dCUnK8kIbvxJy2LM7zBYpIM/CXmAgWROW1rjN4Dg2rKN/ZRxkng2EJPQOBzIOgCdtCFdMBhe
OPbVsmUnsqctObg9e+3VTIA7QSjtHDgCZiAcy+NBgxeYl06v2p3K/VNTNG5nOkCZ7ls1l9QNLwNu
7rqrH3eKzk5z0bkCV++PIAZXn558J4to/99HpHW+tBwUdg56eu1wh/3OO5zRtu1w8Xo0M6YjWCvv
8v5Lkyvk5I/un3CpnHh4qjn9B250fPboVC1SoGA0WQml7SyrRMkoaTTUEXW4+a81rewaLr1i0TfR
gXe8Ss6cSAVipmUxMar2iRrEZgDjclSRg9ij/50AYYhCBoSV5Amg3x2MIwZBLFJJ4lbA9cnUjQA8
dtilFQ4VYM9Hj5w9Bb6X6pBsxi+NOihtcgeKy+qiRh2O+A43klGOGGvxi5RhjaNd70sdmWpACG90
3rG8STeSl2I48eh+hRaNe2EOJ9c34F4oNbpP0WstM2hTvnPUXQ/gKajOullkKuuxL4z099tSXNDK
yzuda0a7tjQq5BDRv/1pRyGXDAHqw2OAvmp1hcjna4k8FDmRO1v3BNIz5CbK2JrNKFwJPq1rjNg4
nTTJnf3zI1vWLG6Pf21tWBlFufyr+PLN9Qcy+cv8kluX3QkwWdAoYlWjz7tI77rYwsDUxAOW5Sth
2TpaDQgipBJQnu3iIlCkli5LRvrOa8GjGBW/vdmPk8dnL4MS4VT91vzh0pa+GDZrBhsdvh7/nBm4
SnQdP46goxIuRboJzDKttjYGXGi9UmU2wr0tx3V9UW6q2gE5b599szMrVUtXgz8wKGh4zFf37lWx
9uE1SRDhuUWtBt5uodt2O8aWf+oWE4R1Hr2eW4etqgwk/trscy9mRxwiZoVs5VN6Af2rAvzqPwcw
o3eAAqTXvusdM0405GCRNYW05ooTdyz56B7v2XoMK4KBgL041+81KIei85VIKunNndPH0DNkL3rj
Hm97+P75EowEp8BGaUVmJ3u+XTQRIX9NVjEQV7Kbdp4xxZasPHNMRTBN6a0ABQoXfbPMIQ0Yeb3K
uFDTQoqnqxneEP6HBhsp89h6CsbqxqvaYpekwKyu8SuLfmY1WR78zK1nqk6isO03bKXVZKXb6xDV
7NuahNVwlZ169Whe1s9rOlEBCKMi92FU6etXuLVJbJY6HR8WlqXya2gqAfxF/dUc/SixV1ldEcL6
yOr3/ST3ks4QggbVG9m2a4Ki2f1C13Hn4fmgnLn4lubDfVeJuKcCfGCS2s1yG6orhiO0xbyGxO8u
HXkbUkAi/lAc2wv33Nk1xetyIxbKFdW+CI4q0CL1Wr8RrHB9AU0X3rX+bW9KvqCY9aW7RQEUBNGJ
Spdaolzqgv8qfWh2WzK/h9BYhH8r0YHh1nnHmYl7+ABQ2R3VQkMWcEWgBkBXwgKkQB0Pyfgyhc6n
8BQiMyJp/vqpgDXjtsAJU2jZ8jSZY0Xpg3EOYlnHG+bX3W7uBOtsaQeBrv7/V3Kx6Hi2oJ4G45kW
WyWrlLGXPB1Fq6Ni/Zfwo+H9m2MKYyAsPidkeMuMJeNFt8GL2hySjoQDvFofJGyE2faEES5is//a
itbkcZ/42IGKU2b0wyPFvhVRzeMLfYoeAWgZZDIefDu+CXlg0Jpqt4HKx3AAuSNkyfEwHdCv+J2I
zq9lkQeMNYpelgDv+PFNFS9i4x1f4Hf3eYkAGVBbsPNQSflWmBJu6ZJPW5AeWUDSoPkj2ABjqbXR
+kGZN+DWpniz+kBSo2CoNMOOcFUpoaj9ANmJBzVmz3HtifH1/9bVHYCJTUhx2hF6bjkJt5kF+HcO
xsVz+ADnttsXnzC8mfuXkE23F66Cdyn8MkV3pZrHkiEk2YpVaMCRfkw+ku/2CqrTMgnviy9gHQ+9
RzUvIM5B+9JyiSvmUzvl5DoVmTv5EEJJiPeW6/c0r+y3ri6p0eRg+IpU1JBG5iooSQMxdk1NQgUk
s4H+xi0jAOMPsr8NlvB6u3kqperTwcJkH649weKdafMKiqT05rS0c2VcYesUyYtg2QfljiQtVAel
sLJO13cSJRWhFMs9wydt90vR/8DTbgNZ/xMUcMK+ulawmF1HKv9CxQHinmd1Ad3Kt/brd8xQ9Bel
IXSQQcAb5EoGmwboOQvbD6roBXAt+Nh0Eq/QGOIv5NButbY5xNQ5op4GQyf6qLtJJ9hAJ4Bnunin
QWO5saGosfJWGXdP7AVcKe6RHcCueaF4iFlMRBqvBZRMX4rOkKOK1+FiWn7uqQZFG1/Zw7iLsgKD
EVzpCu9sOmRyrT8+AI5CvlH+H9biGnjjgY5cTLbhpYTyDy9AjnZXKRehzUiwC1tod8RRNB/YjVC1
ssd4lPazOzqicISjqiQaQKKM9ymaIWxZ9eSs0E0teYAhk9DPHsnoCKTXjECSozx9SNMZHsaQXGoB
WDi2G62iScz3Skv74gCDGjoEpRqv+2+6KmuiYpwOz5QGzcQqErASInHWc791eibZm90IOpzZy66X
D1U2i31zQ82oWKaobIB4lm466CKNh5JXd+tzF4ndJfSjcHxNQqs3gYhuJCpgkknNJ2BawShA+OPv
FCFtqL+hx6rj2gKV1DGNAZov18dk/+U/Ukr+onTn3vqjqYLa90nRnLhktSa8/9StctpbL2ItIqt6
RSkzI5Vtk0KNsGIMm9wDGNi1xyYwV8luDmsYOzPvT7zCZVwbZwDIx1o5VWR64aRECY0EiSn4/znH
o6C/QzjR/zFbZyeCdVXq8PCBvk5X+iLnxU6ZHanknvnrJFf/zf6hx8Urm3DkI1wxKk+n9uY8Bv6U
d4odzKVdFjkPLVsr8cCwxP8r5GzUVEa9vN1cvVj9X9KEZK9bDKZvjvA9/497zKGbrEqiH6YfCF+U
0qRVfUCk8a/k4JREW9Zx69AE8+hvT/OfzEYEACygogl5m0DFYWfauzOyCQWnMi0UtkSXNnAs5/gF
Ok1BhcYePDcMgnrKVseQagDl9pY3XZGb+G8QaI7/mUOp99f5R8JerqWVpb7mfgD2OCO8qaRp3DEB
GUfxCgRiH3vO6BTSf+kEmG59rVv+S8IWqgniBfjBx9Ngrpe7/3SuuwKr9wo8KCEvK8rEZZbGTu3n
+dOH6+oCHUYFe3Ehr2Ren0zNmhvWbV9eeyrl6QDIoDrcm1oKXi0xrcZ9C3mR8zGiMZGN1VZf2IQu
ITnQiqri7JoxxSVb0v9IxmJBMGNBmikbzISZvmfJkppYOG+h5GXwULWx7lWpZKx2UcUcee42zVog
0r99aCzOir/v5OfbDyaC5HrTXVwg0JnYxo98NdbudlL2piFd3VvqUd3DYFBOCeyVs5r2WdlwCQWX
2t+qQy8aZBzy5BwLIfFY6a/JRDNcJfnwQwotGGuqc5/SotKocekk2ejbkIIz5g8IF9qPI/Zzvote
TvXHfBc8GTadrgSJvv/X2CwbGwEgCR29xZ7FT488WUMhSs3B5T+ste9iYSMxBt5iimA7heQtkRjx
6lfZavJAxF7qTQibMSuy26/NjLUxM3O9OPYXO8HJ8hrT1/9TqtkZCdlu6nEQ6jd5o9qbj88ikPlI
3KI7gktGGn9dgWix0vT+B+5OlJCcN2wbyFxHmLYqcmsAhLaX5K9KmbrNxEFiJGdwE0zqRPz4w2mj
gZXI3nK8seIjv9pU6e3jeQHltkyG/38RLhuTt6Atz7QXaTU+onaps2u/UZM3D70H3W0FEzBpRh50
WTn0atvc938XtgK3JNFQfxViCAIXL/8wvwwMXc0/XGCN3/qv9hgOYWHdSfINEC/o4+Oz34052YVe
UoS3ch7zGzG+cLWyEtjS0qu2es/CkXGMmFZq3oSXenp8r7Kors6Ru3PK4VBOPO/VD4fRCNui2sII
fHemVmsc4ydVtVHym1PMe5faOZPWeQJZOxeaiUv60T0bYDpDv7cTIZnf5q2yXJ85XkdescSAoHje
L3ieyGQ9tgKsyimGTgHaNS96rxB2zDKqsDMNriZOSDpw9L4oOwBA7SNJ7ZUYf90w9V7N9/L7QjFv
u3b1a36bduu8jS4IyTjmDzmPlPekG++uzlnLyAC0WB4LVQsB93C09G+OdObAYSJFE2JYK4p+IbX0
XBaziFYJ2xUVvCP4txB6fHt63feQ0R9XNxZ9Macz4skEtw2lyZmk6U43GtDWtJu7nqiuP5SlrPmX
B7NUGzO9n3CdBpIQc4XbYQPLVDsD76ETMjzBXV8hi1fX99/GM6+q8YIVw+XUqbzD6BeTQfbPP3F7
STOMj1XPfHOtR+kR8+fyUnTGygfTHoe/xp4MgMomIKD+UfHSOGXJ6oOusL+QEkIEkUlKtk5Tru69
M6nqBdI7L68J5ZDfLR5owlenC2BUTOB4zb6p3yEa/zdSEKWA6F5VlYgYMT9pG+jdFoWdjzLsx2A6
belxgSDkMeTnvnsgohlVbCO7Qc3L4Gh6yIzHxyzi7RwAA7P9o4bS8Q7rcS0Ri+GFzyo4UJMd28j7
6yV7WJismOPzw2tQqyGILcCbsvq+1XCjgS4U2jgtjpA3gaL+7AibkrMiI2K9IKpn66LdJsm0bPu/
52nlCl06cq1utym/66/CpPVXfTN7LoNHv9u+fIlzAdxjG5viRS7UzSQbNywEmL8oxs23britulaE
uu4661uLbmxA0rEprErVoKDXrfo0sDm5DHQwxQZqkRIty65P3WC4ZeELMZK2kEkBnhYKZLxhc6MO
eqP+mfNxe4wjCnBw++GVMyevFfQWN4t3IgIb68kXJVe1XuLJfVp0ybK4CbAijR0bU8VKEsHkBu/T
SX3poZtXUhX9H+uKMpNd09J9RiUDuS/ChathTCSM555hvG85NVbcbdyIblCWQMyqdiG4ow5pQlGT
8vE8dPaN0tdle1+THx3la4UhffGSeX/7iFMEhEGp25SqYJ5fpANZkkQqhlV4EVXzYO351p+vGo+P
TOB5gQZuwMUsZSa+2JhT8fvrkxw3Go+DFk+4cah4obmfec6yYwJ25EhGr8SY4FEdDVUJKFCmKqhw
/ptc1DS0HU3YCTOZbMp9EKo44SrnshKClhI1Q5MqX5XnJ8zq/QoY2XvOTqMKMn4nqEGREZZfJ7G6
TayyLFHkGsf3kB+M2/UpQjIbZ7ON47Zs+KP16XQ8AS//svqI3tn0E1EH+zN1GjYLkcY+hopF+swc
Lh4pDWSsNx7SMC9Dln2EC3vyZTFjxDM/E9A6egCTljgRjcDgWQJQYy34JXnuekPIiGCuZyrkq0cp
V9RBiQzgIJvSIlnYgr1eybAzQYBHIkGljPHQ88rvgCr2UFqEKl+BcynNgudOQ+dsSBC51r+lFbxz
Xru3gVNKYH4i6mIRuUyUHL2KbjNJhUbEmc275zVqgiwQP1VdViqX5MoUiqCEx5zLb6Stbx3QQT7J
PslfCiFI0JlsCUS2dsnjEfxdOtlRHngM+dRVm1uTNGdV3GMuhUfN1fZx+75supxpB52HQuPWbutH
nBmFvEIf8r/OOILytdPIzAYDyawRJD01IWTlCSoFyJfTAGzA9VUWKPzSLk+59Iyv6JvyNJdUq0Ag
KApvD0WLIPpW0mrcfZn4NtZvmJHqUd4LnsqNtgFPITKF5xZNnqqNwRNxwBTq3sXWBeyz7RPJjvRt
pnVgiBW6Yk+v05OxdV+HO9Ec63x5d3nUuPQK7ibfs00tQ0eb6/aCZI9T/2RlUqD4lquFDMRGdZjq
hwjAjFwYpbL9kfm/LaUljOlPU9LF+ZoLmOcPVDIsWEeOHEKFAkjSEdIFHyI9nws1ai+5wqn8Dneh
bR2kccrsODAYlItWR/bG65hhwdSisKsAM8qSGOKhjMV0Cc0f2v/931FnlkB13sU2JfVzwk0ov4KX
kalNvwaGldRr/3jZYkKLmiJ2n9OnNDq6LFEc2Qi96ID9Q68+nXsUsrGFbt/hrA6LBOygBoccfb5Y
E9Xh3ybA5Yt8FU6jOAp2+sQukiM5vYVdVAdixjHoRP2qZzRzJLQ9yCcQ+HZ/5ZlfSp2+wvgmtrn8
AwhQG55lst1oT2MleAV1alV3DVSoztGOXv+RVr9BaRdhrR1O1LEccSie2FTEwUkq2Z+KZs7Kiq4c
TKrIoHCbOcKgMpU3aTSoLYH5rEfVwVKltfo/ak6o3wVgqZTpSV0+E9Cuv4V0wpUZmITX+Ny38u45
6g+VLzLC82uF49jQ/LjWegI8OVgADR7l3LjGCUsqAyWr/XzQBCGummxD1faH4+7Gx4FqN2kaYP6Z
MzHkc36NTa3uRO3CIXyKJ76TUuNKNozm/xRMJlYrMCBghqeXzsTWg5Wn22yijK2FV5u8SRb2VQzB
CzZKl2BlSpvlCd90U0W3desnKkayUwC1Nt6D+rMqaLRtE726GQNwmJtdKHGvKETfoNWhrFd7wQXf
N5QuEpcC/O1f1+AenvPEKHrfEbiXgxFjLnFY2ys7iCy1H9cGrIXVmrOV7ancaGvi6Ql7npX+4dy+
G20hBe/dMSADyhm7YHCnC8zGfhNZTb9NZgvLZWrhFogdcvXKUjtebK40zJpam+bxNaTacsEO9ECx
thAfLmPXlJj+6XddQViLR8v+A/WQr8WMJsbZ3Sj4jHmveUqfKL/nPRy74TDYsRyrVbVcjFQF4B0N
uh4RTSMuDQNuDTb4KJImW5/yMJQDANACljsS4WjX9F2siTXtgJna97UsT10FvaYxYtlfp/9M4A/2
ZDHqgFtHwMsx/fqsToODz7HVkUVHz7khfXg6c5mUObb55GGgEVaWNv1A4ISDz6nbsKxk7eqHnpfW
jKsRtsefqeQlrvCIJ7dI03A4ll3u+dAaYcmEY9OaMWkKVzQ4mzPmj+vaJE+ovAjTDGIA1qPP3MU1
FU+Fz7whkbIQ3b6Fe42iTymorpugC4Wp+FaNrUXlnR6FXnCCM6SyIHaFNo/WX/ZUp4Jjo7Q0k3YO
CkT14pkmrO/tZ9K/6atzCZop/Wzx2AS2VhA1yRNSCMmSDuDnEal6mbDNmZwNIs2MN/rrNx6apQ7V
vbLxpyl6r9i3tTXOhzaszbqTxWGvmFNdFxa8rGaWzCCT3bJHxi9ecbbSArXiuGeTe6kBltDRdEEw
qLbB6zWhR4prykFLaX2JhAfgf9+GnjDbARqIVjInZlR/ibEVdACZ1+ZN5bzySIWWNeD3O83AcVCu
0ITB6wV7xXRut2xXI4RAM7lqiDcYPUw1zzWBREABmchFNXT1L2H1kjb+KCC6DJQJ1eV3gJhjXt35
UE4nMEApMlsZW/0LCnx42/tMO5hi14s9l6iK0gz638dQu5Hx9LkjpzNoIE9ITTskhgg714JCPUTb
XQONwgEk+AVLzZ/uOKSJO1alEPb+kyAnitBjzOsleB8OI8jFiZZM+AYwiqyR9RkGMx/Mlr8hdvi6
XwCAhWxK8j+IEAkcl96mAncZ3YoN0xCLBRwEVm8JBctonsNUnE0YZsrlEgEMB05Q5rmSGZJpQEwx
rFQPpUKH/cOW0tRIW9E3v5q6KHUVKWIHcRnfv4vGGlsukX0GW01K+R5IXCclJNbMv0wLMYLXgtnM
bvfAJpR6spdJXDWqthx28BFnhM/EkBr9YIGuBJ++pmqBzw9AEuFyTROOc6xg7ylat2qv3KCEs2OZ
KR9AmtNSnx27VTeTmxmjtJU6uDyLY1TceYzPrGTeT8ILlm7Sm40k8j86B5c2EEcPGG5IwHn1ouQA
8E/DZw9sx4T5AuHjUgl2qMXYf7milnGjETweuDUKgFg43X2MShI+8CF/tmztKzQQ+RaG+uxyTqID
Gp6WkiBSN2oli6xsAxbtBv2P+5rCHmiSoj8xLvBRt8YbLAdq1FQ5VH0HslFtguWNI3BqFu/OJBya
6al7yWjiyeDHRwuv9SdMBiJ47ZoAy3lPeWVLcxMTR/qgFlFg23UHBb1i9JSWfY2Kw1UrC5lS5iVH
/1KkdI/60zIV3VdNZJO62DsX/YANlKiGGYwye1E5J19yfN7GXfL8lOY/LcvTgu/4yK8ZDwtTpxKY
EWyp+hRukBAtpAY2BejVVuI+Vl0fKXDoINcWMH2g7Jw7BwQbgb2a5phtSmsgxWjzm/ty8ckTfqR6
3aWLCWzmxjMBmr1nZD5cjpex2ww1BqhwjRr5tl/pNcFtH5C9USSZv3jkJnNj5vCaP7DvYsZZ6OCq
CRsgu2yoMUGHPip6xd+Xf0Kjyv8Czrl/ULRRoS9P1nrBKhvAPf5atruGh7z6m5GiWJ7/M/LxF1rE
NNa9Pew6A4rkwqSyQAyij8sbMa7Vud8KJPW0vowsvNX7EB4+aU7l8gAKGFCSY3NHiaZORuYjzkVz
MyDATosvK0NlgiVLLxEjpd30It6yLwWZhMpEhZ/boaKhr1T1UEmP3aGk4N+E1FmlicBzMwIsYHfS
yw1e5qJ6q15JYl9mmc9p7lXwW5PrGtFUZXpe9sw4pBgWAmM6xtcOfXttysDIyAkoHD+NPXeLwUnW
qq5aK80wx/JafZ6DZAornD0VHPtrF9WcmozIuM8QHDv6cRDNSHblv4684Jk/wa5OXa1lXW6O0/zA
7sEmjaIZixLYVuNGv8LgDT96Dv13+mGEmQs3YNmCxSGPBAtS4nYTGWA3IEWu7KpgGXWapkQ0DGJN
FXsX4nYr335fS0BhBD6gL90DRr/cWdk6wZI+kIyYXPd4W+eerBrLhkYCoHlSZAzX3QNWPM5IEJSF
nwqfecCdpuYuZ41cTrWSmXuLBpRm29xBwAQx0D0bD/L68dRlwmXK+pb5DoeQV23GVVTU3+O/sI7D
Zs0p+F60HwLVcxDKFEb4gDxZ64Y7U/XcWLIibvuYDF8LoOreX+4RNx4p2G57EUEchq4WqTDXXL10
Xa6WeO4F2Vb1JZV2gV23uT6+aoOjK78j6sLym19VW4OLKgVb4nDzyCdYZwFJEtIOFN77ANQ1kiPc
rCL+QgQZ+1tXYrYZdPAXqV0Feeyrn1vSuJSknyDOzr1UuXerJDFIJ3mk/ExdbiDXTOL8o9mqJrMi
vyKabviQt7B2kkhy9MCf6nA59+0ZOJoaUGK9ojbgnTMdkQhqW1W31U+z3avt01yGsbMQFtKttlPG
K+snsr/t6X1n6BHfbn51c5wr6A5ubcejDfQdAihB31uOnQ5mCoj5gXdhKb4Qlx8WahWVN3yzJ3TQ
6eepro4nJ5XCsMdZuPRN1VqVkq7VPMiajBQgVbR6RO/unVMdtU8MkmVDeoH+PAIxYxUfS/7+aIDO
NzVjmOdoQKW/ZHvAnqOpGh+EZPcMw8nmt4Q9Q+pWD0e0R0+h1oZdcoEs9bAhb3toNLQTEmRiRmJG
G+rprxsK7MQCzypF4a0bOUGtyA0rCRRMk+EOzBoK2FsptKaSxG3aaBx/CkmHvn0x/BOWjc6qCBQC
zOGYOqQv+PTdYaD1qffPzMOGOhxGZOq2tjTQPXO0EnQhgquvL+a8+B4KdZOQf/MLGwB44zMvqEF5
xyLGjZ927BtPkzk7FT+o9Ppz2vsQEEy2QBP6m8+XHWoNaPclf1ryKEm/SlY3SR4w6G/wyWClr5iQ
v8b+oXDS97R6HcYuhaCH401QQS7n0gb+oI//x8oWMDVWhCaskKTWVCya87pTHGmYmMjhVHMQRPaG
OORd20uCE6lwiP2bGdyoGa5kOnU6BYTbSsNk1eLTgotsNRpXg/+crbA3HgomUaafPjAGqgOt6zVG
kdi8hi7MKYgioE0kW1YOIiXN5sHcnINlS3oBDgQrP5gwfLUDP2JXAas5Rys1YpJSWiAIvqEQ2iot
K9iMoquScSp8zbrMywDrCYTd1n1MO8o7Zcs7G2i7BU1C5sl8u6rG4bQoRvAMNzohkeqtZ2Z/ZGgv
kFYrp+fAbqzAtZ/WcJQWjp2pCFD7OTjKbdHlrQ1HLrDDUmaDX3dIZS5hRuBitWp6KK3QMRipwYks
xBtsHCDyit3k/9q+v+8gYdjLPU8LZuopX+6tYhHrzakmcuIEtjsci7P3hdEWHiqdD5VRMYxrZAV5
nJT+CUznmDORIUWFVUG5Yjj4wyMaQDmSIUUJViAUD+tQ5vfBX6vSNBmrPVfL4uMUkLDtBlagdybq
Lzjx0msrx8jPPFspct22PQkEB+r0xcqB8E04kNPUvPvWBRtntqvO+VLgRpfxn0O/hKJX2apa3aUi
5pLI4MXYHshxFUCXlVJGy2woqxxy3/lbwlI2K3DahO/ulX+gXsjyDTO+yDDQDclHnjz5TVCG95YH
B6ZDNQDtAdeGy7Sj5sSuKecZNum1+u2OLcXvw3Bws6aHs2rjN17RMp8O1KTCVkocoCNeXCh+vFhN
gvlUZpLi2I3LGWZ0MYKCyIOVnp71hD9DVmIQXSN8hVCMzCrKpZpv2jz6PU0yxv1gg/pTiAaUxUGC
9s3kjMkCmTEVTaBhhbDNDuLAcmM1DYKlB33pUHd4G16FfEnpMB4HGY+++ONrvl+4Tu0EZ7FYn/Q5
68C3l0g/Tc5ZhLzxh+J/ONRST0pzzJ909v60yk7jCsAQ+lqpONqpOzX+UeVAFU8O6bQqknFooUWn
PVtCGBf3SvYLsj5w8BxzV+vltmuCY2HaiVr9O9arSgyZHfTMiKdokuIK4fO43TqJRaJpx9RFAki+
ZL30spoSQ+e7dbnhaUIAGylbgw781hLL/HzUnM6rela1VwMasW9+LcfbfZvHVBL1HgBWPjm/s63B
ocOEEwCmBl6MOAnFP8w5LCl06UR9V9mAVCBN5m6yH20Bzmqw2OANc8TbsHVSmogx6PVJ6JWN3vSW
ZkLPtU8EzD1tg67qC/10ZkhxWW9WSbFTixIeuK8erH3+aoenUGA2hcnY+FKNHL/bh4eFjN+N1WLz
qEIPzP8aLsowUaZ9H1wb7EamilX/JewIMNWKmNRIAD1++8wqbhTY24yqQD4pOdaSjGnWbJJbd5z9
lEhbvBoxLJX0vBOApBlQwKO8xRl6Fgk8VQfxCqrxOE9eohA4BGoajlTZXxggW7kuZX1eXO3cpQ3S
yW3zkyvLxtgjsPLeubZbBWwoZtHkYNttF1Hc3PGV4BT1qpuQ/GPibqrgDo/FT59I8AfFQD5Nvter
5EjGWNNmzPytFmq7YrdUmUsMV7ELVzi3AYIORXCGe6JOu8lCLoVPcNx4EAeVTTy1fJrDzt/Q1CyN
HJb7QzbkoZotpciVlpMdGw6IP8JDQ4xjL05V93A3v42GnMplScG++mlDGFnGw5gioEExpZnxcbVr
0EGKwhIKpXNKe5TsuIhmAkvFcWQMMVGrVf/p5iyk4AKx5+3Ei2yhlzkCGmsCTQrR86Jh3RMz6qnJ
W8mrOqH4GMP0jqbAhdSdYIf2v6pRsZI8RlljIvvNKg0L4THQp0zv2LqTlk3J4cNaZUpvtaFN8o3+
RlGJcsah4Rm5pk7bRIu9EZDKv682EjelLYMq88pKxv4LTDxFP4C8I4Zf4xcL2X4Ra/28lM65/XAW
fZABWHuMmgb0zM6gBRWv6rQiSKtQn1fku62NxPBav7QsWo2zI45sGg46v5tA+BuhDKYJIQfG6Sio
T6cJ6OcUNv9G/W+255HW76391yrYYT+7dwJnNm1280pz661rUQEbH2oQ/tT1xWjv15EyhhbcfjzW
JZXe3qpjsQfVvCJyZrHTG3w+8/WJ1uUb57HaBT9n6SiD2DRaT4ziiMRfpUcyvmaGaQ6w51vFz0Ei
RvG4DAnkjtxAFLkNFYQmCsTQKeau7q+oZD4/VzF1nSOUEBpOPO+ZQtI+vOUepfa+Grnhm1JUt8Ir
+5nih9UkP1bLmlZUHBOCAx37bn1LwjcMvaEQLYVYRph46X2PRG3SaSHNkrPzCqkBPlYTE4lfUT+l
vCf3Bi+CGF7SSubtWsjkfdXdcBTWj+lQxcMT7CRvHS1dTybC3XY8ASsfHMlKbveoeb3vhQeIQcOr
Vw71ZQUxuKugZN1pUX+rP7itFLn/67bIGHx7zONJTa7ij1lgy1f4zEVOdeY7Jk2V3ak7ZEOAzR5Y
d9zGk/KVcrEk+Hk5Gz4eLXHONPZV034gcenJkvVfTpjb9rkTR6DnOwjWrbk4Xz7Wioy65iMz3AU/
HU5/6Ga484XkI+zalp7XSV63fCcJ62t4lTTvQhGsaPhnrHSa6syMJKUnq3iLZYmWrqmgIXJXqKzn
RnEEnyjrvUD+cD8FE/RWdHQAd4bxopKiINh29hjNFVmrSvsJIR10irL6tUCmaTpgdVGmd0zbCapG
TEvf3RbfstDen7nb0UZg6YkeuRefhs8T5sFqWtoyF+7+y1oxeLc794LTiF/GJRQJpxpZfySLVXQq
xzNBEeg/pyE+y0cUF4Mu3ZIidDBHehv8IdyLHN2ANfKaAkd/alvMxcA/OFiwg18USNKuBXRaSCZE
Yv6opfGEYnl8ktCsvVxxvgMf7TAn+q9Za3UKifSSJnLt6Sk3Yvp3bw+sBGIdsaCdUFrBa24R+4fU
9svuLKFHK7eU8NW02HrSNSTonJHNrtO3jm2oJEvRd6XPEN3ALM/OCffnjXp7I5w8zz0Ql2vgb/VZ
kX/x1Hqmi0GIa/ZQkmeZJjk3OjgkwTCwB5QJjtWsxj6+iJZMCs+DlqktRIXLS0MM+Zzg9McSxxIR
Kq65Phf3LcdXPUMFU+pTTL2UYkGwjQ8aaxFvopGo8+kTD3EmuMjFQgWfxXeQ8dSoO4fK2HjwWsAY
5yzRYlamNDAQjKIAs9c4lLMYL1xn1UCIxcqESvf4u+vFV0b4mTfeyzCTOu5m10hU5LvwfeOaXqZ3
ZOGjg9RC94YMY0jO5itufKUI29Px3KzUv2MFIvuO59S9B1ouKsGdz5So55v5qsOuglS0qY5+1pvg
BNl4S1girov58Z5iagfjauCrikFHxMRnVOdRSKJReLcxVIhnpHCD3UJT4VnPEvAtyuwkFTGEnbe8
ipfABxsOTCA/eDnrrvCGjnVhXfC+t8tyni1kBkA0J6gUJZUPiehrTBsPJaMbbnb5kMjbwQcdsDT0
hrqu+cN3574kHL+wj62RwKUiuDW0XiISMo1LGYkT8OJPujSPHrKHpDfEAusIsXvANfffG2QGjcsn
7yFJI0v8G2WkUJhZgNyV3GFyDKS9ayuCe1ICJqhEQahuEAWPu4A281FdA8tTdUgpIlTXb466LeQ7
onx6MB5f7G+CXl+seAeuEcuuaqyYMmQPTsCDDcvo56E8h1EgnFaYqtP5NO+Bu90d/cPGFGUcRwSa
c9QvzkPAKj8du5Eg5glB9JwdknGRvPdCZZzX2AjPullLMumHroBue9u2csKW7GGsOWZ2EvmN0cnN
nrwdskh4OsNQmL+8vtRBKZwswjOohOg1oMuk2O0SkrHCeERfmqqVXxZkkOHolsgjLKcW88xSRdyr
Q6mFRzSLYpekxQ03URwUqspQcv5qhZCt58jd1IGHAfbEPerzqSpMJyi7ZoYbcVI2k1a/PGaLXYDt
b4fTzT56CFf6QvrwsfNu9eVtU7bReVv5yrFHHUJSd/cmVZYWZAJ27dgaPgv6mH0i3UZQXpXhKx38
5dxxIncxGI03m9FZFWkmcAhV48DNDeedOtifT2LRuJeuES5FBFc62LnXwGgeOP4T9UK8OYWmtQkb
bHySrGXYbaKO1pPBWPwo5IU19qsvaxYZZN3wBe3mQ9sDdOQXbocorw4Wa3NcNN/t/TEQQvoxzRuH
gQWiI/YszI7AmIL4lN3M37GGBqMZu/iY8u/HDkDMHD6doMU2a3VxrJGy1FErn6MYrvBcDR5pW/S2
EH60qGpp/gkiUQKbbEkNBDZYvhgw1j9Gh0jEqz8Tsai6E8Yw2U33LUo8nqvJRPH4HxObsQB6Swc5
qumizNgN6LFripZeodR0Hj2XPXMYf4XW4ouqQub71LCFxXBRPZvmyp7bs6POo2PA95cGb9ctNcR5
LPdL3rzISQzMspbk6A/+WEZXyFLpH7KIqtRL8XPLpB3UA23liSDX8i+CfGCEtwbzkW1PmaoEs2b7
1i24I7TWooG/sBuf81lAXope2O1JHYHEbsWttnT6iRQvpVnq4HgGxNkoF5cs7IGI+3N7G+kJ1Mk1
4n5RtaQwVDgSyE0mzMi9/MaE41OmlEv6R81GLXkMCw3Ptv1pNW3oirCgGCsqRMgjGPGwwebwO8JV
aj5/1EsSCv1zVkm16DZE2j1YXUtb26441rC0LrF1IT59D801xFSZU82eK7OpuiqkT1gu8Svxlx3n
Yn6Bh7ifxBM1KqxkBAFfNmycrJ4dX+xhi+wQIdmZGYMYcuwgLQVZ23jAAo6+Mnn0Bpz9hqMVWS/M
M4LWQSIpirJHYLZnRLeCkefcWc4O6sS+0oK597q4QP3D+8sOYXu+m6t8nN2EY9ENKrDtZ/HyAW/o
DMa6E2DTVsI9W7IXhuDqYXQL0Pyd6znKU1SoA2qyH8uf1PqpCREEakZ7q1NKH8OcTyO788ul0Jxs
BgTuoSJ2bLocmKg1RqqraRRDecJ8afRdpdbecs+MQJZOYtvcQkZ5PudEYbxyfX3uqfSRTRWzidrn
Rnv0U78SpIgwgkVyXEe3qTup3JUMBxBhTp99LpZcMWjCNzUcq2a4F7rZ6WIwmZtkSiwW8x5EYTDO
FQb1fzEPReQD0Z2skj36cSlkSb4SWYeVBJbBbijV+m/KxlmRm7hySaA7+lnEw5iPyqqDU9fWItD1
35iP7oE8qGqYT6/29xkOTknyGWDAT4Ci3QqJItnS+J+KfZSO3MUOQOPV70ug/ffGmN7WmPESm3gv
h5QDBBEb8njXNoUTfvXt+AazIkzJKCTMmFv513fGYDu8aBJU1ogSZqanMvSJmrC4emHayGCjPyfP
E3UmXh6LRISJfGKVF3YaCWCPFTdCu777Xrfv0flg2OTfMSgwZzSwZW3BYwjfQzTlQHnefwlhmyXW
JdWJJaDQYhcdeYaK+geFQV53EXIEOt3SGDa8kdrPqXDFQnrkG2ZYf92QMCdQ+gjpdDoY2rTytKeY
W1L5AQMFK64cUf0447wJLqNlenhO1hfci5DILjCaMgYQF6i3mnpZKVptDH8CPrQFX5acHIznX5ix
mAdHpeHzQ1PX1LVk6bG4/2KeYkB+ZDXPVla40YWHV6Gi/ExgY0LvL01Y1VGB3cD0e0w9YmxkPYqX
JUzwLiMYV1cQJSSwUN6W+UVsU/YztVHcfmTBhXpCuRoBepoGT6jmAId9qPA2TFn3QJGSCfdEdR2t
FIkUdaS9H8amoIzjMTigZZZeP9raXHeAHLk3GPDcdnyXp67up5FUYcvJKbvo6HhibHq2PKfop/uc
P2r6YrkrMjRUpTKZFrLs1Cs6/UuCNwKMG1hB1woO+PBatVuEHZfWPlp3Q/noeYJYn6W0gL9LP1Nm
zzGIQ16f1Iz0v7FepADwoi3hqX4wiNexO1NKSFpYGzmru0EpegnhSJ/MayvMeSppJEKotA945KvB
7lXKSnYp5Q1FHsd7NNFvu/LmbYt/TAPwkLXPKlCAWij3GHk53ISiPtu8ug0Xtt4RA4jD4Cavf0sy
sedvI7v4olQ4oXonHLWirkSqMR3A2mcjR9V5OF/HYrHT7mA1ZCpjeXcDaZshZRR1tYn3vFKHN7K3
25PYAK5zVH6OwtW38/glmoue+DcyzKHGvW9k4yqialIjTew0OtiwREE1e3OVI/wUqlfuD5CkiuPV
HEYk2m5PhZAdEbHinLlV4gbXfAeEtK8YQJbnL4mOgUtzujDvVCR34em4eWrlIxWTKKyyEU5YEPFo
sk3i+bDiHuFyAt0OOBaT5fi/6EZ4Qh7BXGyp70OWfaoT7DzrFg9t6gGPdz5HrqyD4tdKGK89iq7I
Fw9kl6SiPz/ZtFXGZ+Sd1aF0fJAehTiPvUjRafj2fxyG5QUsZVMcVnobXBXDwl7Q/3HXg2WUmRlB
4POCbU/soyRHievXnxKEIdS3GW1yNYKanWhTaRm4rLqWjdKrESCZK3SwCqXY0V5tSlz6R87RxRBV
oFvFC62t0mCmW3MV+hXn5ESFjxTZAzeJlx3eBd1K3XNOAIlhUlVO19Gb11pZMot9Cm5UQ/+x0f9R
7SbNXlRTwkiCsH7p+MELXW9VTxTQEWw5O5dd7BNJysEPHjA3/3NFNjoTd1aAbbUjjKqxzzjO9A97
SbelchN9cI2EbJgTu4OC2usHaIe32x4+KSh303FkSQMxroABq0Xe+jYfp76L0svGyDV0Xm9hGjKS
qh+1a8SRJnEMAFEXJ8zAVA/jt/++eCjkFe1UCnHLeY+yvjw0oY2eAPyfRnlf9Vgt8n7Et36tg4FU
FGKN/KdFQz2LZ25eV2/WipjY8LsXdhB1Y2opJ2jC3KH3pRLpMwEZG/t0imBvC+HOnRVc3TsDcKhw
4nJeJ6lXCp+CwIUlwNlolHA8pGc6MUoWEcYYICiOoUb+Ehmv1qsiHx6ZSBDxToG3NjUMmmFBLhRI
FcugLZufGxy4Fp8OS7AB8YBJDXtf+eie3qSE+qn4zll1aJL6naETL0J0Gyg55SYoW68NfXOn64YZ
qJ7BQYFbm5TO+yCgmik8sa0QXG3JE7Uh+MXgwYXjN27jgmzleNTp5ryq6LBEPfS25iGzh79ovyET
n+DpC1n391i7Rnh8erYh2UNZNfbQIpX43gdPH9ml0UbtcdFxc5sTIHw6Q9X5/nrhAXA1ltY4tV14
T7PlctXEvCehizl3PagRh68F7WpxvRWC9pAciFqY6WF+h36RnPmK4jkcW58Bkn80AMkuHGDae/ZJ
Xtjk4mRNYwWpbbciZChKR5sxFl4lKNDlKljh0oO+DxEsUwQSdqllF0l/EZru1fKIv4IFy+MyoBia
AsTFB5Nh0DT29tsY/MQkk0SyUHqswPR65a45RBMmN+KLh8skZwfu3DBIINHf0aqe2iy4hVHz/VMF
azZxQUSAMFxJUUrw17EZ96dWWycEFGMVi6qcTJj1dYYdN1gkQrqGg9hg99Dw4czLl42fn8mHCb7L
unMA/jRxY9ekRt+GlbgeEGgy2cml2H0JqD8wCxs3SEdN81YWWZLEJPMGzsm1g0Ww7wZwu30X/Ik8
OFPPGItCQFGp0KIRT5K4UFFEsT6xRt+HJbtKyu91gc3novWWnzwcHGl1UiL44ZPy9KI14y2FGVpz
DemQzcNewplVMsHzBA1vhtJM9gOQycwAtMJ0NEkqbpPXY3nxFRkEk5M/2vLmNfQJaAE0LmIXsncQ
5mjl+v9VYNAZxlPFv2nIVEYTSwecvLcyobJzsoaiYHrpBd0mtAVu9GGC5HIe9ORq44U4Bn/LwxRU
6Qsh/VDsEW1HnjXuRxHTkYSbq0GMlWUwsPOhmFclwGSVtoa1d8+fIoWgITrpqdE8pnv4l5utT9p3
H2Hr4g8eZqdjLU9QzwFQJcCMNO2W6QHNbqoeQh4i6gH6l1fOG5Xg33iKoy1qTtkRdrF/i0667hIP
Wb1z8TSP8UBOwxkX2W1HObeZDuoiqL5C1Ga6b+Im26+p1cJuU2QnpWYpIc1Av0By02ucoYwDvv3T
Cw8NVOoJ3iwGZhCRPklGi8Wc+QcpkimcxhprC7rSaOsrBuRDJoe9qDAF0YdKBB2R09mWjWK+yoA3
lzOA7u/N7iVeqiA4TEW0qNc+SU9JExYvtD0LQuNGyh57s/qDUfDFIsoz+v1y/DLpI29TZtsK880L
KpyzHQjlTwzsgiiWOwxfZCn6PW65YWLNd66RDaFtDEtGT7arbPKy9onDXlsPm1GE/z++5Jljrd2y
mWNGCKDdR0k0hU8BeVMDIIt3Bxob57V6ryOuVUIecWQbyOrdnHgCG3O4Ye3qUKahO2OsP4r3SYKE
u3UWMtErBl3npPVzobYFBBeHxts78oHM9lk5rfKaSKemCuUqPxY/NsoglTwA5jw4dBB1qbium0N2
7GRSwI7c0bdBjslqOlI0NvMahk9UsVkDbapWOBkeY7wOL60+jn0ULj2DjIQFa1Z/p0qIixW8TCOQ
m34TNtCWnX/vbWLiH/esLE7CX4abg43skcexPQT/GIj1Ss+Djptcx5XtyuyxjQjZuh3vYlQtaqaS
s5FzErXeNx6xLJR6DUTFoUSUfAlGuNSTtgOI4ybebkPcb9OaW3TvUIwvtxZR6j33cpQSJm/PqRTb
nieJkCr8bi5mcyavoI7PbcCapTC8tX3YMIOCTGC18alS0eSxWwi0eK1UdUBLjFrJPeLiFGn9QAnu
m1ksiT/5BmhHCsVb8H7HkgpQcoD6rEOUHRpN58fC66B1aNXLR6revxhvIJDiGvjSfFN4UtwpwLOk
NLh8Svd/1RtKIr65vq8bGBTa06BE3CM/5Vbmxol0tEWk7Et+4o+SJEVKVUVRBRiUQL834TeLN0VF
wEirD9jPrsSVGC/eczsF9iysBPYY280nyxXYiXntRNIcv1tTe5ZKI2P4GpTt2MIIB8aThYyIRYlT
LNCitAOr24IbGY54TR9i17lNwphZM7c5//mwx/8zTAmCYn74uotlkdLwzq6gBkvy1G4qRt/qDXis
roeT3G95PwwhQZQUDnW6pEUi6zUEt3GX5geF1QSCQL8ZyTqN+rfEdZfzKExfYGajeT1SHepHCG3K
lczBSUnSXCTvhcpe6Zc2+QIFwEIyngUp/t/osYQE6Zrd3dwz9W1q7OdmWCddGgJvlK1QzOt6INg6
TU0tlDfwVh4jIuDGvgXdfmggTblZRcXpLh7sxDxIwvOdkBy/Ad9PME8MVhiOYNvfzGm56Pr6Iqj4
ZBGao0Y6b+U5I3hIhzzLkWYcnh18MtH8C8Rv6sCCAxm19l7fQxicoANG29eVX0Y6sPCdhrKnUJuE
FLDw+sZJ3PZKEGOFWlgrljcDaiMiOCfTfPe0VClaTMTA3lz2odvQxlCRhV9MTWf+/b4mnx+gi+tj
gC3akr0tqh3ISKZx6L6fVMlAheE7yWYk8RjLPfe4sRDl57otai4Cp8svyIfEJRhcfVR5JhFa0AVe
4M6lJ6rAlwfe5kKJ28qawZszuBS9pvPaIiQvm63WTbpPCFBJgQLz4VkgemOmuzj9FZIF95c0hfLh
lRrGfrKWIh1TxJrrrlK50ALRmw+yFTLVXzyPlXPgouzBl3F4FCi151hRnp8yAzqTokd/8qgyPeWu
iFUGuBQkKieXdt7C51YzIh60YBw5UZfW95msWAY6gnseJuqkWpuc3Jynz21HFswMDYnyFFTxw4TZ
LH0GmKMA9qPD5EjKYv77TV21MVh718LJGVG8Gaeo/rmVhd9d3T3ET43QRlwJ4LyILtZj91APmQ+k
0sKAwAs821cmztLUVcqq8gyV58r2QGKJEiQwcpoXLQa584skpSsm9QdbpYH1jUyN/4dAkbyQwc1A
RKFFzO08Eou6PDa+1VUyG3s3ZT1iSScSQpVxOg5xQnSV/pI493VYaPqBijYzJWWmg7KQedqvSslf
MLxwHmSgrr3G/RUmoXv0iL8Q90Y9JtfG+6DXpT+eM1H3Gt28ZfzL+m/HhCMNlOEnzMKzJE7qdtiT
NP0T8FyQBKCwqlValrqbaPbMlrTBafBJa80Zo3QzyA/jmhaQqE3/BQFebrLcxQxFNqFIXCJfjxP5
DQDpOKvsIZCZlxIxlruyIDehGIR6rQf4o9ikcxpq8nExx+oBvH1gb6rUsf1lJTu3rZTbFD5gEmhe
D0vAvJW3mskDGM2oL/ll0waibx9tTn8OWVx5whRMEBcYgWeDvHO2KhghjUUkhHAuY68bfA2aex+j
KQNHeuNymChFhkcFSuKas4JMxS6jfCEbBhCqIIoX4imwAQC6J6hTa2QzAjAH9r3YQVC8J/pMZr/E
Qq8xGkcKmU0PTvh3V1Szfo0ysDSrOg5+N9xqfqfRdwY3MT/ud7VJ+UsaK6e3qO7n6ey1y3XQZ9Bz
JbF0bmEjKZJbLMsX6zmS+jCRBAv1i0Cv9VkoIEng07YN/G2KQnK9Hj8jncqz28Ytf8X+DeDpRMbD
2ElXJ1o4/WZ5aFvCaHa3MIDwf3XWoikV35ctidlYMm3xZKF9F/p8ACVVPJUF8WhFhcx2L/70TCCp
rpVxWBwc8nwvYFm6IBSyZV//ZA+67G6g92Cp8pYXCA/N4tpJT2ztU55Hlphs2LGlbgwdXbiwnk/y
7NhoEejvyKYpxuS0lsGAucToKWc4JhXuSOr4aHMBZDhcsN0Dlt7LDjJRv0FOP2N21NhqwzXmHmw9
tSGVYuayRt+XKPuIlFhCEHZwXOz0futuUBr0rqGcCT0PslVBzsV35e7Qq+Qj38TWZCB/DzpzpB1B
R2/R1WpjuMcOeCiRAcjCVb5xpKBch3qrVrlhnPv5icAn7ZdLOf4t5vddGCKiwJd7AlkFuA0v5sTr
rSExQluRQBT3Ugkp3w7p5Mr8rQ1OitDrsQRqV4MYsoOXcCao+ZpOj+6mLGfzlA9n8JHwQzVm5/3s
EAlgsAl5FoHxImSf8cWY50dG09HZZQLUt3lp+994I29XwoJ1DHO77WN5fQeDv+aH5cfCQRz//LeO
E5TCsqOEQhl+mPZrc09ORoV5Vx0iZcoeserDHo2Sd3Xo60CB6E0qadfS8Ybp6D77VjFTzYyQzzfL
zSJPpMxePidf/KLT0x4tjNA5NdqFAFkCpNrAZ5Hj+XBRO54lZVyoEuw3vlTGcYPNyTJCmf6cejkx
kOIAjEgWak+DoFSzOYUg4K7jtZMh7SGQwYDdxdY4r/Tfbe777TzXBOUj74kRqQo452ku2XrbIfd7
r2P6kRIpm0x49b7/S0ZgIELfBz9omeQMy7KdYO/81mhhWYQID2g7UnxjzzJIqzDki5rnzNluzv2b
CV+O8YUxgPI54kUr5vAk38IhF4slRagG2c3KDLpdpwifAcVFUOappqWfepS6RqgywgPgh/Owv89X
Nu2yx9a98aG7ubGLwdIUrpn2nhySnOGzs9aqf281sQHQN8AkvzxKU4wOzIkFj5Ky4/tziMvPfwOo
67DuNI3LbFq6Iah200u6U2sWZVf3MBZfPKv6vOiMSrxebGJZB/jM0HZqEV68es9nArpR/942ap+8
Oz+s7BnZdlvyprkxuyi0VeDVjOIRuE/J9hsWd7sk03+RNEdCe4hrowjWCa5Fi6wYOqBKAUWZ9ZgL
3h9b8xgT4WArioBDu6y4rYrvIp+D0F3cCzMmLHum0D57jTVYpV9EDCoVP82o9xXqgEEvdbZDS1jN
WUesSrfcWevyPnozifzigaXBZ9mMsU73IeSAyBOxW9Zcn5kPa8LedfoP2AvhNxBTFQhp9an2K1kP
XJuMmje9U4LZ6/szPKP6neHbZ7skYxiVQ4yK0f0+g25n0knm6SAtwjRHKc2A/ibkL3lUBOcV/APG
rwSM5D5auK151N0YOe4QSLb1Qt7NmJffEmIO4B3HWKlq0JZ6DHCxr24qvBtELJU5irceXkLFOb1x
B87v1Pyxssl7W60n9KkU4N4IVQTbJXjGIhfhabyYPLnlavDnRZUzROz/Jid3lcJlS6l6aIiebGBm
eQnja9nEyg4CGZd3WHT1BuZN3vlQhbQToGd6wNl86ALumhg1ku/68KtCpw3YUBApjTLVjbhsvrJ1
k9RC6l2JgMOfHPC/EqJWYnuHIvnfrGsmSBrFWDDwcGu+7F8LKICheUR4qBtBLzm7dcpYRDcCmlF+
PYRgpOgej7+reBKqh6k6RjV7AGgNW5Web/k8lDRbHSsepCkdNC+URadvv5U4ExeVT9wx81a5wawj
P0hNH7b0MXS1UW5cPEOj3MLKLB/xP4Ty2W0MPV3s/5s8tdD52H1YO/fjCsjqoGcH9sGLrh8UIp9F
WS/qO+6E4owO90b8/Ncdyrwn2GwKDJziDqwUt6kBKwS41J7YldMVJT4uqtH5F4JV4wIJzrXpSUN7
pYn94XL01H9x+l0kaDEmXKkrF1pDHNcSdaX7zgAU+QXmzfPXO12EfiU9ijDbO5pYKFi7YhEFifkm
mciEAHiiGFXR5WxcdbHmUYZaz+ISbU1TXEtMhSlKxMb+yy9BhyJBTDcamAvqjpy6Qbh11CXivgTm
7+/68krpjys2YFY8fUFZNDsU4MPxOoY4K7UMFDCbltDQTotwiow726doXQVdGjzSvU5vZDEq7CFT
U9KlOUVPYOfi0ecBiYZZGm2ZeNrzJ35ZTfW22dbUhhlzvT9LKiRm5HP3DPQyE8A/uZ53YfC0Q2X/
2xvBJktOhAFpvqJFwfH7CV+v3Z8q36n7AAbXfQzqTq03htMmIwyc5QpqA2H+Fgu76MlFF5DXciJX
mL4DnJO/mzTrqM750BxIH8z2ysc7k2nrY7C+rTvGBi2PHnNUF0Tl9yrTqecuKeTWhLQbTHNfWac8
RWMSzaikcRoeESXzVEkzrqEBZUatQ2DU5m1knU2C1iZhapb/xefQDRtxxo4i1rRSq7twFUngGdxr
9dfa60+iSSyi1pFQn6vyJmHe8vkINhh9ogWvxFjIMPD4kzbvlwiZfTiHLMteqT+BEz+tqBiMivIL
81N60W6ft++R/3PpX6Cc32vnve0/aNm8r7FYTbDnCwmNo13WRxIUPy/HZeUhvIjcC/rD/UWLnDw2
+fesnTKejyH2P/MZH8DCFLUMJKY3B1OJgywB6nnus1eLZkDZ1VpzB8Xu2N4BqEx8iTT4AhlAthZp
YY64qJDezuvQwdg1tGmsLY0XzyZFGmLZieeJqVcImX0hCFocvwfKa57KRNdbJxu0GanaqSpVcD9F
GY4v+aIMNc7jnV/1j0QmlhQ7myMsPvRt5SDjEl2QYEWMFsMa0WrDKNRJ2i3K8Lpw8/ZyzdSlscY6
bTR8+8zRDvwZTMafCIWLjWbZ7HxYtAn4X8u3edrbjxmp5CvWh7CoQBYfUeDmyY9hspaeOPqHmBBj
ZWyrwZOoKlV+32moU09Xo3AYV4YIaciHNTRTHQQ4VGXjOw/34pZe6aLVKhaZuSSYDqvoiwNSXixY
iC7OUV2iiDer3ZovcoTw72uNvr2G6Jsu8h2yeCMVBictspgz4mp+Da4soU26DyKtKvsqz1CtiXlQ
h+hCZcTHTLpG+e5/b+GYi1Mu8Nm9u9MnnyBhWP72LR4R/A0u09mGnDGQ1DrgzJLRdUXgVW/1IaZE
hPL14eArcyXw3Pg/QMjI4LbzPxxI3UUUR0bgZjmcxhtCCn99aYqy0q0eLVV8lCUZS2gaT7EMXsWi
VolPm8G1bzsae34dWARa6ErQrp+J08kuiYWApXdlgDdU8rC+eoRdfzQWl3CreX6/+9rUuH5br25B
7KLNHsVGjPIkvLw3syM9lOSa26h76RcGjiVDH24iL6HiRo+bP6M+j/2Rp9jiSrtUBlT+d7oJB6yG
P4b1LfCEc1XP8KHofWcQSOquoaLoHdDI7/gmV5Tp3b4oxRBk5KpuUipBq6/H9OkKO7da+SZZyBno
cjaiQ0I8vW/6CogTRo5G72IUwzd8pwYWvv2g76thz+hTekeFhzSI4mXS/3iGeq1UCS73W0YavgCK
tz3OeR6xRC1TASErxHpsfcgxlesDcm0Qimqsod7tW/5ppxn/0jZyUO3Ew+zdChwFVLnI3euSzwPZ
S5Ett9eTuxK9uKLJiBfAQuwsmuQezK1ZMA90lYi8I5TfFUA8nAlHRIASXgEbDX3rzIpvdAbpk+85
gJ7xm6W6PW0NGin7XBB5dJoFh5IOSy0n8RL5kMDrqdpfiBqnjd+tOM6qDDKv2sjnuJpkAPyJXhkI
67q0ixjvWwJh2EeIQ/dXLTSaSkJZbXq6a0hxIv1N3W7HKL8Vz4mQQ38XqgTKOf4CFlX5tm3G01KH
VKG/VIAdNc7Nuv5PSqSC/5X89A62gpaGx9YOFKYBEZjLoIxxrGd0SV755HA28ngK3AxuRoji++Op
tWIuEhN1JBOJku4yeGjtvwJaJxrYWFv4p5Q2DWS4ZEOrfia3RRIcvlF1kWDrzHjmUtMuHLn2U3Tl
L4CCNU10MVhfe3b6xc4bahxo3w/A4J/6XsUp/0fX4Egk8Uh4OKc0F+3Pb9O8HAJ3sSYMiXcBv5eW
XJPEXZQhC6YJASJvzJd3SbyExxE+4lEdqxmEqwtWwnumhuxx6xvVcR6zWcI/MZ9RW7rGS7ugYYw9
+6ypQHVr2LG0a+OHBdgVV/V1BvzROd3cfddXzP89t3hO5A6YbOM7JT1BBtCKf+onZHN5Tluk7ml0
L7RAlkdai+6NQTLHOLu7KFI3PyJS9xgaAtd4sPugkVr7NPoA7pr4nPIkSBlt7V79X/+deR7HFkS+
V4KOkIjuyC8wjyg3UeaueAdbKqE+7JMzyd+V4isZgBSj0LRkqMFRQuYlF9QI7Cddd4ZnpOHQv/T5
0PLXTvi70m7q1fa2OQz7X+kBNgnpyJ4+3Ly4xwkYW8zGUQV6MlpfZ8Z3HAaJK3ozWVTAy5PgbuOD
G/REqBnznzHCMz1oSWRget36RYhIOkbGxfiXFqf2Hsj/XoKd87El2UcfMfAd/TjFoKqZbo4RCbN2
ilnavOSdl+VdkDqLgpz39cXjTrmrcBEyIWQvsuEXEZLy/uOBpU3eHFjolA7jkZGy4L21PH6Jj1lL
mjYGvsoZqeOQy6MsGJ1snNYUOr1r4P6rSuxhSeZpVdzWLM2eoBcYsPkD+zrOz96hQYhpLB60+8BS
mpZihXdoQcevsHwgSfVq+I+pQD37wr0Iw9rXHnqnWAtlTh3K4J5ApzRJdoJLU32L8OlUM7WMnBUK
zvmVEafdw+4RNjcKoB6ITqyjBnCQqYbGp3HCFubU6x+Yffb9hnoUA8Ane8zhkX2UJabkUwIkPf95
dINOK0ujY6H8A2X4faDhv8qaBrF9HOyYGc5/1km5uVAbt5DvCAIJ4uZ148Ewi5vxIpEKy1nHnIEO
X0PcCph4KhRJaJkZaWfNQebm6VJ56d5MR+GK3ooG1vqxTohi/SbC2AeIoS+qdM5F288HshDMN/dL
HsJI5p4sBsWg+GX+MUNZlP1uAhoBLmNiG1NaQ3X+PDjajg1Nzp7BeoAMxG29Jge/8sWwSmdpt9R4
cssd4Q/whI7hIO+TUYKIMLVCeAS2HqVpKIi20dyVFj0gx4qRaEGOdtSLfO7uzabNyxNf+sdQz3Tf
DXpU1OGHksEIOusRiEd75SjMfdNI/gHuu1ENdu+e9e7IdAtCQAaQtVzMSIlSc8MV67bggllJSpkW
r6uX2Wnfbdflp9DdQ95qGIyv+IPI+WExMnBEGAotF+wuGVxnWCdEocl0xAC/R/bqrZUag9mUQ09n
Tw7kPkMqZZBQfgljjHoBoxCjPg1lV6+XPtFUllskn0bnn9vl/MizElqRvP/XHu9tLKLtXwq+qoKd
glB+WKzfwCBUqMln51upp1yFIMIrdYUtz2xD2whbTo2BQ8ttLGRoMoQnb3go9xUrWMcOIWmgAV3/
EeYaV8WpAKIA4V2S8PLjhhH/r2Isk8xZa0wQeVdJjwLo9IAs1cwmLCg4Sy8Lvl1tBvBSamZSmHqS
1VT8n2xWLh36A6Vm4gB7fWEEuK2Zu9pJmS6BJU1vEEK2CKXA62FJS5G7rlrbdgJj9y9q2PKZRpoS
VyArPHq7l3AAyePFfjA0MP4w0GalxmIdq0WYmwlceocrxu9B1l/P+u11tTL+V+9tuvIVW/qGNzjz
97bxmCvs/YdIkFXsiIjvn9l3dnxhMGR0I0F10RZJxfeYGsLIWWKVvVOJJ5WTGwk2tqMzaI6gmcDz
C4Le48gHzybdDyh3z36lwjTrCSFQ/QeO9/56/8W9JhcKYsZbDGJ9XlV4n0HKle/07/5tR9WmK1Mo
y4eQKznyXpefVvMnJlZWU/4kOb2PDb1IQEAGM/3La2cdwPW/+txfwhW8y2303j445FWz8FR9sXs5
3Oh70m102CfTHFv4Gj9LBdvH/vJCwiylLfdedwleeMAlwCWMtZnb7rcjDsW90B4rEh6V/dEdwDq+
sYK7bHdKThgL3GGc+hC06AHUr2zRbiaKH6eSuGv7j04fF97HqnfM9eYQOCvp6ibUMqoiq0JYK+LD
UviqO5wvyuxH5yeV3ZkK0toLZxpVmIsrJkisKZZf4CWNXxkbF7gZInljXB+M8GpSgSYIBTPlM79a
N6OnWnXUeVVlHbu2ZG+/0m0kUf4ZxP7vvBqtioUmg6INuwHkgpuebLdS+F6ruCvtrf7BsoPkA6gA
kzdHMWuUvRY5zyZbK5G8647Ias+pXOb0lwJ13OPjDr9Vpm08hsSz+FYos6n3Axe+2KJQso9hn7ei
k7PWQNvXMq8EE2XP4uIqa76rCvm9fEVcaPHBvdO8TFmK67TpBP8f4haqwoXN75xFi+howzve88W8
DNiX/xeycvz5UwEhqgRpgx6A+ihP+hCe1Of+zymGQwrLzYvjIrGGp4CAbMMc75zFOvgyfgxgmyrl
PbJ4XzKR5fDGT8BzB8H9xIU7iyqmrxptV9lYSBlH3ZaIKM7snDKwCe5F7WZk+t4S3ELYraH6Bbh8
gOK2wS90J+iVkRqTR7Flfh3hmNxwsXDrODbLwQWCjJAdKiosUKAjZsartI2bhUPLXhN3nu5NnEaH
Oi1VSFDoGqcloDZfjQzchgF/7VnsmXSb1eNUQoOfhd/Q0XRK5TtJdQbkZiLKdH2iOEsdTWYlB1uf
JQJ0m7dZg4cl92RZKiTy82tEl6JSLzokZjUrVUBhqZyRtYRt8wyu/Gj9a37fRr8nQYZk3+bTzIEF
Ny0VDnanpfOf7Ua7Ih9DyliSYUzCIsEfSLCVQ3asl0+N3S0umuvMm7T6um27iXUeUrQZBy41h3vP
JRM36WXlds0UfjBJSpyc9o9S4r+FvCgN3CV2yqCdaGulvdw7LhFZMz12s8WTPk6mUXkaWh4Ja5VD
srtQ1gQqk8AWSBkuKVj3NIgNeIR6YQknsTst/hj5IwGkH4bxvb3qyjLatBaH2FXqhOR6RvgTVdYp
sKcEy8nLf3i6nmm+JA/uadGjFBD9MXRUjIygy2cYnxUBr6IZ6QqPDwP6Ccn02nUuWUIe3RCb76uw
uPh+482v8CYNlIjVCDdiDSYmm+qXgLf+rJy7gqhRYNG5FOGde8TGQqLmbpwWoiOz9DeOX1to1Roa
xXWlH8HHBop+/PlFF05pEs+VP6+u92OyhQ1oMiZQ0azNYytZnJOl+2sV59soyydhiaDO2XFK8220
JEPUT9HXRMKHaNEh1hqyj+5z42vfkdKCxetA5ZqgrHMqTa/tWBTXlk88bnszI4ofIjmxM2gxWNpe
vIMvbrKnob884OTIGcobmxl/Xr9ndS3OuSUalucaztCNdDeWuivM85omKga9XAfiZ15VetfbZD7B
Hq7/6koRmUQqL8d2XTdSjndfgRYSslb3CjiFStZwP/xpxClr5aHvrIrnPyvigbKZvdwfA37XIzh5
da5M8Js5CGdjwWejsmsEvy3T1zcn6wTMN2sRRJwrjkoeXkTWENxHa3LGFk+miINMlAYWGmHehg0R
N4pufSKIuF2Qvp6/jGTlpm3WpbIgXqx4ukiDe1vqfgcF38hPXtt/MYYRvEZCL1O//QdMAzoP2JQc
3mCJJDezivz1PnUPS9BNRAdAAXKioTtUz4RNyzE/RiE5m7ffl66YUc7E7bAlDOIneOZdD6JUJiGD
5sQCNZ3auu4CmokvR3mX/W61C1wbUXkW+DfIsnplK9g1Jn4llBz1Jxg29PjE/9HVno3dGgdx1TwN
QtSsbZ3hnMFOcw7dn+I3nTzfKcQX3WY1fZ/sKUiB9quW41SxwIAY48ecINWuSRVEYsIU0giaYQo2
Vdp6D2UOOYL7lnoPmYXfjgDkPGTVnNqLPpPXmVn8vF+ptyztUpYIkZ4I0KXWaa5qKXFuB1fIzfE+
Tx9Few+lVHY39O9r6KzwIibdTf5y2A5jMXox+JTc7rE6qwaVTp75g3DVbKjXaAMS9lra61rC9HRM
KbbWu+E8As46TZQZvkW6XA92Xf5gxEyzApwxmOew5hemd+R+bXDNKeEZs0PiQz4gC3vAN3+IpQg9
aw22uO+m6ykAP+mk7kAOADZohA7ob/+QgDGkcPVmo/apC50j62OQW9eoB0dCTEQ7W+msAdObe8Xa
cojMC93QLWqnO01EPl8KU/hQ3vT4sUFOTq2v/4NsvsPdwLse0F1BzTsVzLC+qABAEaWcLeZ7YFXk
Ev5AfPOImXE1cdOVHaKw2SQ2EFb/yQXiisqDNnzYqwIDeRivQM6aw9OtAjP3jsVaBDCHvn0ipuLC
2nVFIEv6mnJlu3Np+pXz+r9FzV4NUTAFkyfOJDwXBzYuByz0PvAsf4Ic4chD7qEpBiYtNOy1LFzL
DO2juJ/rXKVSrkGGzj5Y45xFRL+cS1VOmIIEBHHL9lt4vBA9fzBMiiLI4eF0krpBeat0PO2LbxaH
cAgQwPowMjf0xmWHVOIsOTO9FZsPWwWlUmAV/gIzug+HC5lNw8YpX8arlsITj1NVptwfQOwjpmbC
qgDNufaXfwgNwn8xK9Cq9qzqx4tbGSYcA4wf7pnYcl6Dhsy0I5ssDXhBjl5EQafn2SXLMrijIsl2
jY1SCobJteeYk6uzB3G9HxjurnCF5G1eF2bzFWReSSqWS3EI/kk5pipNb9H0cW6jvWZkL7BiS+bw
EOBomLZMjyRcYRcPcB2ea6jHDnMnCpyi3QTw0RmG6I4ObJwVKCLDV+c9C2zNSmrqzXR+OyBYUunK
yPyQlD+eqbk+UiMmpW9ON6rWwTr2K8FWd2EFSXy/P8yQlij8F9Y9emVHphas87993RuxA2jyy6de
mPgS9ezLis/dMXl4x6BXmcc7GhAWmU8rckcOPNIiS8F8aJ23HHbjONxGqPREsYQXoRNfaAaDKMmt
OMx6ddtJBm5WiFnWiMgp7111GSoS/lZrgDFabFthB8ljX0a/xuZAKIUXTLxG4+pvF2P0g/lpzRpt
zfbltkD/mZcLPeICStnjmMfGjinTMK2oQpNOKLC2QqNJSCqjjeIxckLrHDN59/QlyjHlpuNEbq6f
aI8cdqoemzViw75s2JLugBWC3XYEn/UjVrJcvHQyR61o117K/dW0/QYEXwWSD5YOqU91DrlgK4jU
hF7McSS2xPNbj5/8q50tobRzvc8p0GtLoFp9KWMJWgiczWHrhsK614cER2K7xrwD6au8IKywElGF
93gdZX9ruWEPpiFcjYLsQA6nmd87BuJ+U5ROSaiHMlk0dvgTynsstmLiFp3SMABf0752fMUecGuk
OdVm7PBlPHQAqoJzj+ILVceD7sdagOJoOIfqUCDc1qg4qU9cjivRLU16ApWJ04qba+9dYPK7HcA+
ZJA1KBmKY2b/LglXO6Kv8Ixiy55UhXOBHlotLTah3u4qSSUYjkG41gYrcrHFsAR9Dc9+YqZIyTKM
4WEb1VCA/YwG2tgdC0TGELOfAA2mBSuai3o2Bh2Ip3XhQ1/XtW3VIY97V9xEdBiQ9JSoo8LQkHkJ
iTYNsd42woQN5L7qiUPgdwbQaOm74cBN2PlQjUGsqxY11WKFTq41j+uYWRb+wBY13bdxG19wnI6e
I7gbq1x77Uv8LnR95H9Lgj/lSLY/Qqm/3b7riQKd/Fyze9RBf+F9jDSlQA5fF/ohnKgdewuxFdYt
l+4hDDsM4vOc09g89hzQb67Nd6Y9ueMfRHXV08GGeVosX25nBCF0AR7BqAqC49tlwLug5RmLJV1T
SGsNN+TZ+VF6JQvqmro2SJqCe3IGyMZM1TfRg3WJSxR2tA3SYcRpSeieO+2YTzoZqE5tGhG+10/5
vfuOzxfs/Im6l3YevzA51r8OiDiE0woQNmXU0m9hl9bZtk6whddYksqaZyHD5sOqGlRyy0qIiS2J
efmYgf55NP5TopsP4Q1nDczxsFiclnq+LI4VVLUKAQo8JozpcpaFLrNmDFvVP4+v5ISIQEaQZAkb
HYXGVplB1HLVQM/o4jx1qiZxYB4rn1WTFwt1o3UWsmZo57sNhU1IbOx8mGejklvAQbOAiaOrpsB9
opuW98S6JqzKErUr3NgbR/SY9c+byj4WHXRWjgM2FbQ/hya+Mr59Ey5TBJoaIYvwECohCXm4MsFX
h7EvtHS2Z1Zh78PyoTU4z9lZzv5Y8O62ldqom6GzmE6Ej/B8D0Gd1WlaOYLrXdombMTUwITcVd+S
6WXvgO3rWmcD2bZgjzXEn6c2bCkzG8NQOWwGnkWbf4zn79O7qpzOoP9f0mi3pDUA2mtBnR7Kf0F9
Xnx+QaHSd/6/j3h+yATo7yUbCIcM6zM8Jq2z5iMFCP5kyOrX+aE15E9RrfIFaTADj6udVTSEXV5i
lFPFk4uMCTsE3h6r7nD/9OA38y54XelflQ5D010GALyuttOcJsmaYCS5PLH6tXl329qxI0Q88IYQ
2x7oDpLEl7wIxRB0RTmcqpPUs02+Dhk7i791HL7X9//P1gftrFuKOGwTMEEgC2nhqTOkV7i7EPMr
UMruiNcH5W1dSGULSJSpCEbOVj56eOtYVeOyDOtBzhDgozdZbwa51T04NNuE8aN8IRdQHqcjDWvA
WNG0HTXXg0WmrkVQ9nvSoU96KLp/Nx1ZscWOda9NJqEJ2FdWuJFtyCDAuL7Ief2rD2WxXEtAduc9
PhPv9romsGAFfcHxfcRBBaPMJqpHfslVbZf/b+i8MNTTKPhq9kpfUftnakQx6H/dncy22Zto7q1h
2G/wk9RRVIOViCJ5dfW7bu4lMJb4B/oYfvJY55wP/avuJ3xxaw36g1BtKFY6IsQ6IF2qXG4h+NDG
x631TRbpH7nYls0xBzlkp8f1kZnlhLMKPkyYclR6mRztLz9Kdvs7aC+j59/MNJv5c6druPmtrEVK
YYdF9mAc/GkxxVlo6tVU2a2N3pUzxJqHCVuxBtPzatrzxILj2V1xqzJq2FFz7LIHrI0chOjrxDa/
TqXAffZ3066SLvrnY/MNJ4r8oc8LjHoWmba4iVJl9kngeg0U5wtwkFCbB9QxHyvx1SKh18reNRe+
NpamtiqQKRfTFf8x4kEDsW//RS/fMj424bnIBgDS+4uIucGA/bnwgSdAeEtQ7fE0pHmsP7vxDXvQ
WGWBrVTZwFdahp6E5Pj9xrJdMWMOp4N2m8bTm3UaXMePS4bs/dgJEOCpioCDrMUak1GGXkgnXiOV
+ZBxHbg4EojFzWZ0++Ut36/iLbCEoNFgtsD1hHTXkxfWq7ORfUj/gkDnKiFIjCHpa0sLAW9uTFAf
pVxGGkEozARCcA7Y8BSyzHvJZOBXNXCKZbMF4fSPFOEbzFsNmuCdNejq2hswnEI39DqIC54uxD0f
VCpyNxGJTEMpTXPyqlCwyG9O2KmsgoqQKo5CPywWrxWHb0o2KoTzYIhXVkPYz7l3ygZffA4U5iiE
2R704Q5IzWOlJlGsvlMBfUVvl1EhUDRqAFSLIVoI5CqWRubBb60/dM6z9dYCLhZ2Neen4uicp2rJ
pyRk8LBgTKK1aGmOMQlrGNm7o9o7OwWIGXroAJMaPoti5Wc3OK8hEF+5PreP2XnQmyEabitlVUch
7Wt6jfFHAzuGbSWGMJajyhg8fMIbyBdueGeOJC0p04HFF1sV3i8/kiyK38KDEF71pQOiTWxTqA/c
ui/ZF7h70DV7UJ8Unt6neEvc3/TY/KM5dFDFticcENdt7+rWtTd0hrnNPVn+fWRxrHc+wHr3aPZC
NJ7syBIyx7VS2XyPGxYwv0MX2UGZNvprfbtw+amkCJE9ccqWEDa7+1x3J3u+UXf50E2oaxlpLtBb
wh6aPbHhtf6Og6Hr9cvyGQm98p9Br9TnGqlllm5wMKiWt0zR0xa9esUFsH63B70xsMtvPM5gpwMx
V32vVhDq5IUJKAdjiFSTJRzm8QAYCqVrovReaorqJ2VCeafOQ+I7LTkkyqYbcr+FATCFbaH9rdyw
QvXsjHy9QFe4Pmf3AWmpuqGAvkM6XXOjPBY2EbKagadg1Dv73E3KZCSJQcBt+JeR429q7KV3cG4+
yIHTHLF05O0Y8R/cjxKr6dV6CiBuAKRc9XXExjQ/Xfa6tAA0bRqKDatEVzBfhGcYjKtqUNMJAP8x
NpQVHrDbiRqSKcdXeAboQfa17egXB0D/1wOf4PAkuckZ1Pvu8PHgqo+uB8ZZiMYd6IgH+eGtC0IA
9jWFa7+IK7UseejDSElI3Yajf5IVQKhUyJrRm4IttNz7drSX39wfDQyJfSKB6eYuwWMnc4UXgokn
MIzB6cO5Z1Q/U6PC18NH5oUnkuIDj6KfRIIVWlSdHeVpq8DCORyrkkAksVFvG9TPfI1K4FfZ0p+l
HfMDGKN5JYUxyB8EbwaG0GOaE3LSxow9EO2F7kduxFSAQbUZVDcA78Y3lYME7qQ1+5FlYxg2Lm2o
NLmWk+uA5eBPaZQXMQ7UAjLkBbc4xLVYu+y9g4bL8f3MQyHzdeObEt0wOYDweG9wLXgjJzw2MjE+
BwyhqihPItpbYMBgbdvWoezg/4pDybslMe6YTWPFfsDeSC1L3M8HhFooS/AuJm/eAeQsQSjy34Ha
geRBWSb0swOejAjKmj2R2I3kYHwS32p8VmO53ZrXcEKiWwVOhepCM7av/GGuCmKRWA0IL6XXpN/K
AeDMxzaetl2apwPAUUbsy7pYZouJHwi/uu0AcHHzi6txW44CoMXcFHSCOAXLaBTzopNjdJp4m8nU
adBLOCngsy7xdKVz1vB6475Ut+Kq67b0jZ4KxBTfn6OELm0poJW8O0VIw/mFVco1W4OgGQHp1zfj
umcqLRpebQPMciKOwi2UxV8BkIIO2VZ3ewpzYoZZnhirGzTRt8P2dZ4itYujZ2139qj4080j11Qq
uqT2zp8RwML0kzXwa6v3+CbhNyPkEg/r9hvaDE00trHVfrIsa/FQLDNueGvhqrEdIgZeztMUXr/B
l8MhmvEE+2HniI1tDtT8ib2nUybqJHESxSap7ErNHAlORYJsetTqs/99lZMBu8orLgN+0TMmxCYl
qRInhCl6an+FXyLJEtZe121tcHHm/Zw763cf5ndqVLx2mCWZg5DV7t44dA3RK5VMeS0ks62svOXS
O2ojchTvtJgMJhouWNGDFC2NiFfrHkqFI2qIZUreSlRVPn3PBPbaAl6T+HPW8CGc5+wIC2QnmjXS
S5GARFZMFVow1IFaqQWQ2Nel8EvhA9L5FM1mjwxhRutJTQNxLoNcybKy/lzNQJukeECycYeW6Y1s
8h4hgn58KaxAq1V3fJcUSbtb+7gzVCk+/YaFP52+q5+dFWvsC0yoIbZxxDfHGTjkr548C0SqZv/A
V/lMFi5SqpLCpSw8Eo8ntr5Uam+QaBoOOo4Zk5/2ixJDEl5lCrhjacthk/MEDMeAYnYt2YT0AExz
nibUumClq2iLijJyPDuZf3KwQc0zUHOvXQDlugKl1fk/ZuE/dwQGUCmlKTcpBO9CRN/xDWKU7fq4
ZLyJTUcALzuDkADgllBBRhd6xSNO9mxFsZR/0AeM67o9DA7FTnuPYsVMQW/OeG1+YloEGkqM5Kl6
q+kL4Q/kANTX18UPJCVaDPc5aqPxVUkiNQ6PRP3+F+yCIW6r1d8IcTarI8eh5n5/QdTI3Gz/Tm58
7caj3W6cMo5nqsxCPnniww7hHY746FX9NYNpUGbEWw2Ii1MFsAMxjZso3qeiD6h6NlGIxLBH+mno
ati+s/yqlq5wWUP3FoX0HAZuEF9i30yWX2HH0ZnxFKF8JnrJTLSa5EABherFJ2fUKD62Tf37j1fn
ppYk58olWyKb3uMYDQyYDq+GWlhI0onV4U8C9UbiMHQv9PZa1i0YL+Fi/zMFOTc0uvdkUi6ZDLBo
MBMEok3rgwRUPNVic0hikFa890qxhV4XkGW4+bKc+x4vi+9GyDR8zHvWFpZYVf++0xS+1Flkd2hy
lWlSPutUe2qICGkcx9EJXIATAx78HIJxvTr3H4WAUPDc1hXdpbIUAqSW+rLJOWDy9hyfVWArmi6c
xTwlvOPyU7jOL55liT1cz0g8ZYg9nPofA4KepWO6ynIsM5IUzFX0zPdRseaRM9aN7OK+x6HdQVWD
i/M0iS+ww9cCmhsRDrLO7hXmI/wHrttIwy36Lmdij6qHM4sEwp5Gln4Mv0GZ6P3D883f2+K/fOn4
Fnzsua+MQaQLf6x7r1FE0Oo3TLgJMIy+UWZJxSlANlTsTBkBHojoXiM4ALzXTdPxcGmHIFmRdeGP
t1+Pb3HKDw33o6VddXUtfAahQ2Wbgo2mZYmLUuoQCdwkFFVNhbOB4hOuOMg+VpbaPy/utrniXEQ+
hRlqc98lSzxCZfh8O3vrQTtEGIDP40HM8tThWJQDKwYx94dmepysNn0Fj004a+ppm1I5+uH5ePWV
YHNyW10dT/wA9W3p6ww4Wrb9y5AUBi8+yPsvZ/aqvvtOcqNHB9nOJh40Mn7+HibYetgAlRv1puPj
JDxPiaT+e3EUxfuzkpFE/ClzJFtPkxcPDcSR/IbZWVfbCMgbOqbLHyjCZY4G6vnZsFHpRg0kFGjk
R43CJW5/5iodiuaM5OiBLNrjLOs14jK1Z1vhMNt29JNThR2eBrQ1R5FsbuzOteyoGYvMonNeqTkI
bls8pZz2KkPDfaycCsibOnVMCA7ii7UkzwcqaHbXau7gnyuXVnxRJiLkxdygtJpHC69TzKtn3ts0
8dczHjR3swb0AZVkVOeme+eoLCRppgGrqnCOcmLTobJZTunyZoxauXjdOwG0uI8s37hhCSbGmtS7
/rkjFMfiEZCvOovFvMHdpSRmsE4sM5bzGryEWBtfUIN7oqN2F5ByRdVsc3EIcYUPsvGl5Fx85LdA
NRevE7SOeGNLPZpax8LoAxdUBv7ZbCWQXjZDDpp+qORVHCIDFbJ8iJUH+pqK8IjsJD2a/nLjhkxq
eIRGwpVnyYQSeDCIQry0RFesSN1VbJ6WNFH6+WqBdWty8aByWzYRiEGE/U4gjWNMcUMdsA1hQZyn
vS4N9v+nATjtDVO3AzWxdVcpMi70+VRh8GtoniP1wsX18P52aiJIphYmGZT3uKeGYz4I9XpVhVu/
KY/GsHzqTBtJzPCx/bdD29Eq1ByOyacwrZtPDo/IHFnRfXVfdB6TWjebCazhw3cEAQzVFy44OLpw
hyYaiELp0YPHwqBtRlG4Ib2n689W3ic3BIjO+gnScTgBPvDMxsZ/0xDpw0VSFJSkfQeCZvpxNWtM
L2EvQsp1ME5XvyxbF6J2flO9w3rxsotlaeOzQntT3mB9aSHrHTC2mCF4QVl9kMDLOE9WcRCCBQpk
8e3RBNIuTUlSb094pnHjFtE7UYIhYrtkSsKo5yFIToN5xdM6mcuj1ixW0h6H/tNlQu+pC2LiT1iv
UB/YBpDQRSHQFgPN6VYxB6hRrtH9t/Mo8lawOC/+hShep6V/YnHiEDtLZN9irWu0a1xs0OS+8QAg
W1tNlWN0XZ0LHziBfiGG0jXSFDjubzEI0ohCIRv0iNEMZ2jFQrCdvOi+2d8IuEjg4E/iWa/RByvz
hS9VaZ4hD6JJHMcFKnoh1Tqu0pNeJYBgAwGKRiMTDdiGRah8gTuhshEfjZQUrvqzFmZBYT/EOhxn
nPj2j2FTIKIqtzp2TANWZqBc0E/dWKOjKxbUDGhD4z+Mmp4D/PRM+CfLq3qw6lEJlU3SP9xOvIBk
vTm6fJa18GHW8kmmFYo6y95QUYiFRVMwYjd5VC+WZ4YvCFZ1qfqaTNpefrxac0tbY3jZYEKqv/YW
cOpBfbyUh59Z+ceoxtxcQgbX8c5QrJvG/QdXMq2Xd9kISrwdXpX95oaxWbyqehfk1dEQ9BTytWsM
JxXyHD/Xrsyws34DmdZ4ggd6Ovr8wjo3HcEWMf8hxRtXHoyYXaHXeP+HI9KN9Aq0JVHSy8qFUB//
DJkB6nBo8UyJfoCiqDObnnRoW6qWHMDYVcgsemjKtfvReZiz7jFqe1VQx579mj4Qn/7dacwlBAD1
XdVgn2c/0bC0MK/GA9HaWVTl6VR04BaZdmyXjinlDNzjFMBkXi1FC71UsOidHBloiTHSo4CTHeuC
JwR6XARMZE4QWhVclBHdHAajiKqfB002Z/gUF+tHPV4/IZR0n9hIrklta/VktaZO70m7UQG9pmCa
4Q+ytK7pCk/QZZ7i3aK5YMlE+l/9OUhzPd+AZGwld6GUEWvgLBObbQ1jKIfeKk+/aDguVYq7/WmC
UBbQfn+rxoWnBgQEHPJiSHdvGmjCxClfuc4gub9BARp6tbh6BnDHstUupmUASXYo78yNMIvltlzd
KEAzR70/8QdDdJXjIza07uwABtyL/Is6pKjY4b+1VJbL2+rOMuk1yRsgrFlws5WKUWcE2twPTpAV
sXUqzassdXesP2xFtXL9tEIFigVU2U5O1WNfHRopUqw+tp99eeZPvFWEZ3wmRk+eQkHVCjPuYyd4
EJNWDxU2phA4f/GuffH72Z32fJcHtkanCv60KvvY+PPHbeRDVhWzVBK5GBAClrh44gBgk4JqcvIj
DH5FOg9uf0h48o9mocxGTfaTEICyX/1AXtfDYK9/eUKtBZJ4vdC9Z09Iq3P83YsMIZN9+jdoQO6k
im42iJosW1uUgYMsrTlrIlfgI7NFKguiFnMo4SE/SETNlHdwq+vxOGN6arZ0WmuEHXTIzq/l4zFo
1TM3VzfgNGSR2S5vHQakIMGWRR5n1SrOQMN7eor1nbbuvypMAyLBtZdg0Us/BwqOgjgVILObEibD
66zK8SUyBuaB9PG8nY4LXCpYoX/jfsa9B4Z5/5iK+EV5hS6vXuW7SsDz3aE41OGI0N7SVpz+WlTu
eb8UAy9Kj+bEy9pSYljAFuTRe/cbb1QcB1PdusCPsgRFgIaTbe2T8zUDq0h5P5DDZ8xhAiEMyeKV
mh/Prl1mYgEG81OI31XIiJN8Z3nXGftDF1Z4QL1+LvUXDbmJTEYxYA0GOGQPXCKhblumrKLMZlGS
M5NUXWj6+NCNEW0U8s+UMbfwgvM74VkR87K7sGKNa2m379Sgqopahv3EDohBVJE9TrZXY2J/rZNa
tYRIzJW5xEm0QeLVyYzwmIuK1RgAPP7ncjBK1UjlJ0Oi4GoWVoPJjkWXJfiGyI/Ier4ReYA34WFA
ozfseQSNtrE9lFR4wg0vaPCsm+FFRVFjgff0h8juVBidILkMaOvhr6KcR7t2u8882AfNol/aNU4D
3qi7eWAkwj81j4ZVByDB3cNtKu3tiHVsCtwJuRNSz13oOBEHfaUKBBL+zEwzHpISWIDOMk5CvfXz
hMkPnua7/nJMPwuJVWkdmOICbwK2JsOkhaSXX56zFDH5qRFLAGBOv+/57zUxtZP9VSQ9k44WXOR7
WRX20pudut2p69k2ZXfD4RIvZ+PtS57kZ0yshRlaTbCz2HwklZrPSszkay6lAcxtH6Gr2SHv3lZA
iAvkBBtGIICNWNj48wcqKxNGH0apoZBzTMGwpqYET9uKebL6APeiOxFyHjKEJ/9hwhpJjIXl/IG1
Pikn18pnoEt/PgsL41HdVX70KZI5DgDaTyHh+lUCwW8i1/YPVzAZjGGlUUQe6cXM00IRYszCqTGe
UtROhE6VYrGQx7MAl3KYE2wGmZ8NnO5BR8OXY/Sl3m6NezntyP5UffzjDSvHbYf3xE+4ctEAxBZg
RlML7da7lHOCtZA+6ImdJtz6u2N0bDMQVUcQ6VBHbTIn9FQi1nbXqvvTow55iobktCUAMyYopFi8
Thn0cF/c35A20UJmQRQaWd4dmES2gvcfaQQE8wma5vrDhbdO2RyqmTRGi7Jz+SFb/owuy4yGlwse
5pr0b0v154Ci7AyVYqLO3Ol2zhSOrHmjZ+pVhhgeDcbzAUsRKQWmvnm/X79yqn/2e+w+4J8SWZO6
BynBELIwQvhJ8EtY1Y+EoqWEVp+SRZSyzw7M3tNVmBpDIOVbEDnd9tDoIE5Hb5J9zmXoMgUudBh0
ho/g5YGwmyT1/ElLLfNXF0PpSzTIj6JiqUgSUSfOqpjDUYCB7sdydjkniJfQ/tfZMa7Q5S04SmKh
RpytYEnWXKSMNxi6JZWrK5nv52lMJ08DLCC44D4H5bs4ayuNJLS6WesDn1B+1siXS26Dw5mH3Gum
wg8LpCOt5vYAh2iT9jB1dTKg5ZXw2zRzPnFR6Vr1A+pDNmVj/pSOY1JwnRVL7GZfi84Sqr+ng0Zj
TOnyjg5w61g7qaTkHPkEaA0pC3/RQS82MIJ1kyntJ0wxU5kJsTAFAfbQNhF2tpfBjnJCEuz0Sfq+
y7ftr5x+TElwQZQBxqjHKnyR0VBrrr4NSFX6gqyzz124s7fff4QU4A/WF0iiusVyfYXX6XH/jeAR
dz7gNxymsN3E+d1+whtOEjooRl1SXoxVZrVXPk8Ihe28/8YXIK4IBSFq2ti3erzKyVnsSyKYd0BN
ctNJuYM7+oDV0TM0++tE56jRLySlZwj+rQE5EGY2EugbCWNn6kdMFdff6H+ioao6hOE5VNuKjrPp
LTmQFOpNqiNolz4UDC9oT3o+3eLg737g+hJYlchALnyvMPQP7n/A+WNhsePhxRYZiGgV0zzc6A73
JgeRYa6umXX7Kz3p9BNjeDFhVN2Gzv6X8OdlW33SdA7bVT5m9ZYEB8L0FoyRVGknR8U23a2ROOe9
4G3i3zjJyEJihfMPUW95Su+gPIOHnwME9UypTv2t21Dq6r7cAElttYFfZSzeu6v7pTG6axRD0FlO
3nOmfny4JJwBTpO1SeGyN65u3U3GicNda0VGnxHKHhujz8CDcXIzWl/DLtL2dWqX50xRjKMeNSFV
0A4kyRH7mgAi7+5/uBgwhGDBHw+C6IUsC+AtOXKHADglcQz3DKOdtFl+OdMQmSJjNk/Ia2ouV2Dj
hQgrgxpzg7yDf0KG3wkHHouPlchkYNLiJK6vkOP/tbmlVCVZFdZEuEcEoBlCAh2ySmyMt07U08vi
qwI+QDeOPSEtPh4QLxvTlfsCB7DJSblRdJvQhrej6Jyh/8IVzj6J6UIS/Hg4hj/4DYvI+l/Q5WJo
jx/MXaEZ+TnpUIdi8qZiX1KXb3ZInyEgynBGgXEj+FKHhLwESPns/rOheaSHHxHNzJfcCt115f/T
4TlR/79WY2oEar86tYbih7s82N/Wp93iLTAnXIrGgntuqdka+mNGYJu+PANpD/LTYKaol5OV5Nrr
4B5VNMeMugtnpCV6LQwwGXYdCuFw4BjgPl5c6y7Xl7AQAlLrXqnwzFac6AMJ7XIEVIAwTVD6IKH1
JJFggZ4U363tCTanVyc18H+ZCUEHjYaKQ9n3qPKOXExynRZ0e+wLL25/30fUe1M37v0wvRhCb+/V
jZa3ZHYAhNzXy408XIx2xZ7w6XGwFQuRro1nCGbHG65JU88OSotWNDyWckS9m7pLnSmiXYjenaCs
MFoELbCQKLot+76nPt8didMf9KaaFzsSMXroIzWZJ6QBNPzzh9fXGacgQqJ0DWxlyqYoEQIcXDs7
beqh0A0BpmiJhLTeuQJk4GnEXoeQCfhOnfMMtANm2tF6NXXDEftD0Shg/TPUeYTvHKmtL/FwJ2Kh
6JRFnFNfk2ZbRix800kRudNMj+rF/zFHWOMk2Tng4FbBYDNyUVO8da5Gk5d3zd7RcHmwbXn3yvdS
G+oTZYvxU/WMGzYtU6+2YrZVfsO+kOKVMHLkq/UTSTipRxObGO7yOEQgRvZfvzLkEbaXHO4mqvpM
lud++A9rBIqdj27mtGIrkHfpys7jpCYQZzEw5Tqehdc5ayoo+wDPR94fr65kIdKGOoJcOw2xVZXO
7SdDmqvxQDy4y28POG/hKddkIg3KHjHlkn7pgxyI+yKQoRQO8pS7HmDe6oumOaM6S9DEo20WD5yU
SQEUvBc5EU5nnaGoXa7Ct0vedV/5rEKFsLzLe4mzq+l/veymkN5VmdflAsLxPcNVC3HjLpQcUmGx
d87bkqQLPfV0YIg0+fsAdUp0PtnBlaTj1bhblkJ1RTR8MZT5rElz88fANDWjoR1GzWXX9aYRbReR
sLIwAUAgGB1C+BQHipgm9uLQTqvJui+qka5fuTbSLyJwP7BSEOhnjUFmEsoeWK5ZNJqS4uy0sYdC
7lKDAaTQTCAQi0xkalrlPsoLekSQI4d7+PrOE/55MnWTezF9i37JgsGQpnl0LruN8xUo15B60LUT
NqLOsOvuO+4hySg3wptYbGDSRXoOVPVxtyu54+h+uGwdIjgJiphADDeBIZSxm7xPHHJPSuFVkbtR
egbAIKNB6YH6MbClYq16+SUdZynRs1Ku8q+WgskF/+y54uz7hqiaDP2E5e8NygMKali0Sb/y9+Ds
/09SAFeJwLb6/OH4E6CYDVTFRslujO3g8Kq5fToGhM6ztdOAXufjq3I2DiKMC4w52lmVATIUTXk+
V1K1XZfmK8OjACAjCci1XbDDDZFDSmt7jYSV5dFK+mgnQBgzQhah1tY/OulV75NnM0bNfpUEDuR8
1ExP10SOCg6yPIxV1BqMiEReo7gX0SG0J8lT45M8jYXnmN2xYUnYVj/zlSwu4/GVav8BuUALJQZF
wZxr5CzMqLQAdyhCsqwJoJCeXFBQqO1//wjbtyukU17jyVNVXtJ31jLG9VVc0dXQ1oBYPulUmEnY
C9h/4rgKZhCJ++Ld9WAGukhO7z0g1/6bO0uv9alJBMqEQJUyBCZ/qfpsBtXExDckHwt4TW8owVIY
EBPc4xAayH2BpXy0DN5vGi6N8nFe9UlaR87CNF0jrNY48fTZJACqxNMdOXwIHq+xrA+P9xJoyajt
UN4jp4WrW6pVd9ceIay0RwbnTUJSQ42g4AUFXdAOtO2vWJTOyZVnfZ+efQhYb6uR6tSUWrrlSVJX
uAgo7Hf9AW5dr1ax0M/gUerOW1rqj1HSMnfyCZ0QKKn/I9d8BBWdVEn/y5ic6dsUWXJJ8+KaWS28
jj9ZJ4/XrtSs07I+Aa0CAXqqBfiEQOmiwMI5+UnBonevNOcv8KtvoH9+C+pclujLqpH+6N8VS3F1
+lOBbascBGeCfokx5writYjklGmTOsjG5TCqXAveKDFAT7672dcBTVBbAAVA/LX6IBwYiWLVG69O
6BhY8weS16eRAQuND7a9CdPE/wAHdCarw0vSElRliKbUZRCqBSlNorRO1wFccLTPx2RQpPz9ih//
7Maef5YGV3yQKHzFPdeKq0I2u0KseP/ik7rMWYzfbaWzhYahkUAt42YVD7CX2s0KdjxmzyAVa977
LvMVHCKpWcwNZCqggbbY+7arxnNGR2+D49bhiJtMYMlOLqfD7PfyKW0yyUHt4AUJ34a/U1+NOlcc
uRCuuIQ6FeuCRMXYjAZywmZ/iojRJqakWIcCUq3PWXU9EB0Le46zTXwPWyAn7PUapRp/onccdEaL
8tkkKh19uSXrqojdE7TnsrNVNI853z9cmix6uG5b5nQ+hMP3cSCH8h3LA2/y5myTD680kEZwaayV
PaEPK4Rc4lCN0CNP1zhidmctCh9B8WVCro7rMNAp8+ZkQnkCSPZT/G5KRPM/duoNo4w+I7slDg6w
1NMusvUIu3A0MMQiNpC7KkujKZF50iwsu8zm6ZKQN1KE4iVXpMPRkE7wA+Yz9wZmvUpMFZ9lepFZ
bSerK+a/PW2nKVZC+2tQTa2XnRk5Ic2ITLAllvABWXOLeNNqmm4gI92RxlHdoZ0mrGFyQ2xTxgKN
9GHOr4PY17eauAkEGLXLLxDMW9n3IbydzeW6mrRdc6xYSwBxQFrYKHxI8//MS4qmyUwLt4uHFaoo
+HkBR5+SYQNTjB9C7W+TKAeG7ZIeeqcaXeUOPM52lqVUcN7kCQvbJXTLaqqLX0Z6w10k/as9JtDG
XwVlXV6+ozELNWpOK6pi2UhVXWpWb3Ha2ohsptWMIQMn23cuhcXS4SLb5coT3MB7sMc+vLZxPFVm
K7FJp/QSPrQfVsD0J+h3SEL8fTWdHEjDfnlIiYG0CaiW+T/KY+F29jHh+/6bXUFRg5ZZTl8HhlCA
d605Lv6hYjd0J//K93xsQ5mB5jRMnNBhnbnT1IqOXlDFgaFgeKeesy+hhwaot15eEQLdU4wpBNS7
4rE4/hfFV9ZgyAx0FK7NQlr9yS2ZXfEuDfNIz8mcY/a6MpfFY9tVpaFKRJIoAIbRCnb9IQcOlsRY
4lt9+k+kF6kVFWLzUQno8+ekMwNk8ChtXpktr0zXKFa2EQOMWcZNfLefQu7ZCjB0EF8+RDTUkPR9
++8p6bZpyDVa8GQtzoH6M6TTzwyc9O46hlnJc43R+Npa2Ni6i9J0DNsIPeY+ZNhYZWVwkO+Nn28r
73KuW3c7qQLdHvbmTAejgeAZyxFJ05K20Z/uFkaas3qHDGD+MZ/AqUzo8fCvzWxEbZLkh03wcRab
L8JwAyFybSDjijdku1SkkbqL9B6zi1/y6ADIZGA6Rh+LF3K1SheTwG2IsnAhNwQV83654HaKPaUA
GiuJ+jzNsv9Y1gY2gwPDUmXOYjQUmGYr4CAzGCvMroj45dotOxOZEOAuSm4tMI1FXbjdJKh9OnPv
dLhVDr+xTNbhOgndNVSa+pOWEkzEp+SSxOyaiaj1OvQGTdRlQFn2YgH6towlk5Rm3YGjNTkAxNZU
kMeWmYFA1WIYYfdqSeTH1Kdqq6hW0d3kiEGgrW2goPOQrRgTKX1JgNxgR5aBjNo7brzStiOHfiAz
FrBpZ9NMT6LMPxo/56FvTwqgOvjeI4gE3hxY4X1z3nBFGS2lVs02DcP6nHkS0OdnM/AA0dbfvp5J
CmVkpKrfvjg1dO/1B0ICA69x+TwoljtBBpSROgLW6ZhvIAdH45h6TWWkRFwDDlq2m5fNmXUCtscu
BkLV5nFcsKpfq79iTstkw5cBhRNph0v4eoaVhMt2m7X7Z+nVozhP7MaIb09oTyQFISspN4+JSqS1
tvZ/CyCU8Z1wRVTD2svuDY9s+AEjf19/KbAy1OOoAfefEXgNlk912ef0O68YWo6lHr7JIA1G5WMf
6GyLaGPyRM3a2EuYECsBgkMfQ9VRcmU5V5b2Fm83UYCK3L8xmfVLeKl8TwS4Qt6h6Z6jr6sgKKZ0
vkCLy1JqrcMZtQptnoSkSP+S+Mfj0xHBGVtrkXqjdWKH5P/nqIX5JUt4k04SMwTrfGkAExZAKut8
Vnscca1buU+i6dSkVAcB5gjqTuSECdhMgB8iuAAHz1OnYJV566RXQXh7hmFYAjaGfiAmUuZIB7GL
xocIMIjrR+Rx0GB9XHfuVFfLFCLAhajTCtFx6RjbdXqJZcndInF4C0nRcUjnP9/grqTr7QJdk21v
vjSO4+i/ELT+wlUVAULKO71YKPzFKzsP7a7asihXzLRBTNEI1VCYKIxF7CqQZje1bLJRO/YqA4Bm
iFb0f7HdNfR1MXf/3cqniLn1lO6bubNH02+ioaIe27jOrQlcjaPHJlSfp24nkp+7Or+Nson7JtX3
zxd8XJLJZZxhy7ZrjtLVb9d3BzG3JTWpi/A5ri8ycKWJDNEx9s/9PVeT9p0DbdhfVQ9xRn3Nar10
QNzml88U8/ipcnJ44bi3qXH+2uyyWFt52LevXdWMRolrsD7hlGxki0/y8tI84uqoKIGltuWR90GI
MOA1VIkn+4vkLr/6I/TpVcLpPxIiODiRFxMMshR6bjXax7K7hFqdE8rOKx5faOUM++2kqlISz7bi
jMUgetc51dg5BoyPjOJ1hCPrhvF6B6VjTV0QtE3klc/4GEHzWvHAblDOAFxz/rtURgL9lyFhiG8k
a7MwIKrr1hf6XKdXKwMmpU01c55w8+mFmHmcqRrMfnop3klLQkug/0lz+eveXo8c0XKUeY9fRDL3
5JU/fotNLinYfFH06qKKKJW/CUwnskY88HQXUsH5t1HIseFxmOqhBl8zf3Ju3ZfHJJA0fuigAeSz
fAaMdSGIzBVzv/kqUGg6TfisZgPDNY+nq6OhDGZJ4BgTaZpY6UnGeQTP1RCeDZX41aUlhFmhtANo
WBKItDEBYfWsphQEGLHu5pBI2rnAzLBK7oIa0CYkuydwnvMnrOivl/WrCIbAxTVCU5pkBk5Tu8TO
ktYQJn+xQE/IioQdj889uVk54GOrrEWYHdOIqLC3MlvUTw1vvmYe9aWh/a7RnXTAJwTKIAq20i/2
tzZtGvRlsxlT/yrKQ7+OQAMtmhEiiBc5T6vVNoKGQH3SGBPayrRv2g4vCq1D3EC/f2Fz45EOv7G6
7yClbCH8+/RSIjXZ1nTw48boF4JzXP1/TeITuJlOmZdzoGnR65mi5HtUG3fuKs6fXda+wq73cbOB
GG+IYegdE5tSVjeic6X8bWRR41muwfM3GfqtkdP8e6hG+Up+FWxD09Jo5oBTez66411ADsR+71Ip
RTVCSr75+aVonMReDSdqJXa39+MHM6WOHR1YUgMPuP6+YSjDOH+7gfUfgx/VKXZPmrQ+sFR3XKBu
yFu7wFQY9JAqTl21Mmp25W26UPjWXpNCpXQkEgMWLkciymxiEdxEf2I5ywSReFk0fUmGd7zhO9vp
iZelSZx/eyxk0cCcIMQ70ILK/kIGBGgTczp42TfT6io5/apbTn0LddEF5q+w8xlWI4pAwrLtALxX
jiME0vuZ3tbFJoaLSvxrB8Fx/xuiQV0PKXLnaRIFB+Bk/AqKlSUGB5hbh2dqQnqQUfhvihKwvLi4
N0k0oxnRXXk883+e8PcDCTQtWoeFcmaADAw9OsAB8vjoTW1qQmChB9X9DxAF9vqFSeDcr+wLN7J+
fouO/W8sMYy+mC4mRbagFe3ZjdIte3BDP4bEiGbF4je5ButZF8+5D3L3zm+MnXNXTLWD0LE9bWyn
Y8QzelMwV2jYxlGKjBSlhSFOlREaOzO4ezteotGnpp2VKvGCpGZaKR8o3hk8zQy0ijA/RftBAtbb
8NhngjDf2HhjScXFWM2vgAUF1Y3Uraq4kdQlNUnWsPqqqDyelj6zoG+m9v4WRHgos46j7Y9qf3gR
o8KhPZAep3Iz/1pp8XOTV9C+OmInuNnJ6jDF0p+4eL5L8GtEYOWPjcAu+Kb7wBoCfDihi2fN8oh3
Sda7jX43r4HNlqDMwM+qCDee2QviP+yib8fwNlLj1+mzLkUiCTRJ5cBC8qsNtcqJAm7bbY6AOsT4
N234W53EJpN5F8jFAYNTaxH2+YhrM7QCji7wzU05WtjiNHAWntrSMXs2uja7MOFpMXIoTZ30/Haq
KvPGjbyMxQut9K2T/joLhzcfb/xotqQublRaWhk5Ww8QZGOn7957TsFmxl/OzCmRLL7GkYf0fDiR
ioVUMtTexwZOGr7/Ky44WmF9xvY/w4AT577JBr8gAmBtCBnx587+CFg6yxJeCwSfCF/OkIsZ9fpo
EgPQ7lnQrkFZ/UVahb3waa9bWr1s/Gk4ELOpIW1r7KSORL4nTj9Ka2EJFDH/Gg/vrd5nW8xoMCmp
BzISDNLT4/dTgOkLwwlgVxFOLrqX98rm4z9AZXy4N6yn/LuKYMs8sZBmFEC2GBykz8rAFqU8mAWc
AFHQIRc2WS/WbMyM90zBk4f9q7umKBPQZimk3aZRtHMjE8CjF7fSSIcYM+lMyGEcocwyOktriHHD
AqAeNpNTf2ixKFyviTlVr9nl+VnkKs4g0RPnhaZYPa/twhf8rrft/r8Vf3e8I3o/TE2YA9O1GXyZ
59swwYJWWZE3fCLZr3uQHmkKpAnnobM9+gDJFwEj/zcjweAPnucyA4YSHJm1RwB/TZ6KNtXcdHbR
1nHbOqjBXjC6VtZp2gLZ/PQlbWxqaR1xfPPk1TMgBJKC5bFXfgvSwGbDv53JjCFyV6qk9gVbOKxA
CAF0D9fZ4K+Y5tFjQasQjJKiIonqQeaDPcm5WTB0VBZGtlFkiA0SZgsdcQZd+3G+paiYb/ijEB3+
lny4KzRuoAy9fZGa8AhVBy988/JoB8AkYNTXNCIp/JC+P4nN06KYA7jAjF5rA8Y+U+tyxZ4fQ/a5
VOEWkuX8c6oamc5Wz3a1xWQNrm1duJCnRX0TeyL8MLyGlLcSakm+nF8ZO0SfIx+0MHv9k5TIwpam
mLh65Ud2XMMho555xFKTWkePiIkAKKiaDTHcsA4PLfa6e67/FpnTK6JcD2VKOjDFCehmywRLETVs
TIxgZF/6hvqoaqaJxrNEHDDF+1HDj6BxJqXkAPM3vXWioDANkUDK8UyM459iCorkzL2+1/TsWkWF
VewnVrhXCRu2D98LF+kahv1llVin3hUUNzNXE8OTG1e52AVm3u+U1+okeibGiQQVp0K49v0WdMe6
vSlw3IRAxif63xM8vngcFo71NXxXi4dRdBvMUCHMe56ZEnkgCJ9X02fhUVB4+fiGi5b1Lq22ju5W
lbAHggYxx81bvP667c5AydqthT7AjNgOm/5jN+ELwUV+xFovtiO/GYw9IRFsEDgEW45WaUW5l4JZ
3T1dG/7SljeeTTtd1xlQMgbs49KMCOb5OP1uCl4IggMd4JEXNgcX0eRXlkRXq1+Mxz8zYhsfvUzk
gR8oskE+J3AjnDT/PfmhFQzy1fw6FupLdYJ1YGQalKegfDu6uZsl+CWSmMqF2Sti3na9Y+8VsGvI
QW1N11WyETFVoeWrFaNXke34EyJ6OrKEYaKxxj/ynDcAtclWP1UGGoB/JjnDAztP2w0Ljh5MDQRi
IdrZD7USsUxhCLPyoeTZ2QrLo1N9Tc+KEY+Tzj9aE9EIgSAXo8p/NWG1nxc96EREx9pkphKINy2Q
O2jn20Q2dpfKbP7fg8LQ6tHiB435h8EpCsS4j3IYdiWkRzW63rD0SzwRhbTxm1LIqfy+EhdMaOn1
Dn8AzXOtSKsyS6UugWzaQy0gpWgBFyok4TSdxE9yWUTQWejs17/Q5PKIjkx6YGBp+4GiVu1RdT9T
UfD0Nrkz8kCChD1xWXms7Pq0vFJ5oH7Xn73dP8jI0HZnJ1qVXYAwSdpXQa9mN1FFpi5lK7ZFh58r
Y2DPfni0biLAPQdy3a2bTzymMRC3aE7iJXRwOAWkGpUXDrNpilWR1Hgdr1n7U2OYODlSFeK1j55z
Feql+uH9dBcL6og/7SSBunAFmB7Q2dQjPx/XBaAivrHWqkwmxg0BoQDCIKocvgn4amUzy1GwUhH0
JjqloB93dfeOOy5kCKGl4qS9AqQmSrdM4DhhBFNelWZBGlqAa2U1hF7QSigyOf+gbu3kN2qONGTx
+TimM96jtv4EyDTfMwLT2cFglhZQTYpJ4BJKz5MO5w3ULZ6/pfH9MohFKj4e6kWiuYymLaTI3OWy
Z8fEOlxDMzzXR4obaIvod9yG7b+mS9tzcHsN8SKdTLffcVdB7ZpnA7mDozV4bNPMW2SLSF5XoQrG
BCzKNw0T7JOSW0EqVe34iwXF/Lf+UlZx3JayXfiQ/+u0AfSghFmPIzExZDyjbbKta8hxgJDPqpF3
HDyzVKvqCTgrv8YgA25b/BgCpz84DqGLAXPJoXI+qxeDHrCh3BexuiRzEzx/Qa4VootOSPlYqoUX
bRZJnm7GsbgiPTZMv/tvUjmp4bD0EA3SbZuqq2nFD4u2GlGNOb8da+R3NpEWriK2z5UUII38/DP5
gTlNDazEg76LUFZ4XfTROiLSOrBLsUjcwOqQHjh4c0ATZ41yyOGKgEwGpdXnw8t9tLNM/mmTdK/u
Ud3YpDkb+l5Qg7Kq2G6M4drX+AV9wN0dNG0uO5uR3e6vMkPn5FfhaG3LNJRNxM5l1jNCr9gK2jMr
u0lTrgWxKeuigkG4AnrdVaCpLrdXEXpht2WRhYoBlixT7YJ2RATu8OFpZIqVRp92spDFuM71gxH0
3wU/cMcyhEofLojrPLQcFg1+61Be0+evyHIbfKe2u6QI98mkwgXxH0dUE9Pl8TqCncHqgM1c4bJr
GVcBZRwdLQavUCp5ynAxqHefXHxzz92j3a5AxPoruKZBXzK2ZbS0qYQRpTxJvLp5C8sO0fjgcWwK
JE6SX8YKnqmhTSSyn3lYowY3f/1fS7mnoJAp6iVMz2xINJRpujUV0kLdI1cjaYh88JkdLOl98fQj
blku1HKBNy81cmlCuNtD1I/QsEP2PoD7USK9NT7ySESbTCvxqNj0B6iqnuyhawhfWDKZ381M1fXd
4FKyWyzMmykfoCjF/LcnOOOgovmgeHWpUsmFRZJ9J2+XE+RTw1vZjUFdYW3+0pFgVcGZLqjprBPK
3uOSv3hBzzYVyhYcKe35VuIPYY5ZvRuJsh6e5m0VYdSN47UoylEr1JM7CMF2tVFMOa1zEAefZiB7
KUMUQQimHyevEA6j7ZgGSZDTLPS6oWUoIgYO6FUDtqEE6szI6aV9XKsIK0FjJaxk8965Cg8obhxB
HOobqoNOCLY31TMPHdWTwftKXsPOcaJ1ljbvyqQ+FXma832kiGpQkhPLWztCgW+n1y+Ib2yzi5Ve
Ru4B4YrgQkXj6xdK7mdey0dV5ygmDdlIUXuvrQ1lsyKA/+vE20r2scrKqHxKY3kftTygi4Jsb4oz
UIBVcMOJwmI+zQ40NtSHyi7l7p1+r+ytchzK65MGKIgmg+HsYMxIZ0nrbuvxoMtnBDjqDpVJnjy3
p1ajxcl2jMlLryWsT1cprJ4okWqsNgQJHbNtQbfb7ujxC1sxBekpTEoMNpOK/XccR8sKJOyud1cq
owKy1v155HxaHDRXRJqq+I/5UyPnBXWVECPqRLvGkrx1wQSMUgP9hnn81AaH4AcpU5RvGM0hvCLM
xvPBH0UQxdOZkg8m2GenRCrWZ2vL9uCJ6t8SzZDe0fn3Ov8P+66nArxDHZAwivxqLb2qbk3/gqPB
+H1iPFkSJ+xfDR2FYhxuwJOq5995kMif1YnCr98Bs3qQbNoUjgaqoWwJGYZXWgn3fNlOJ6y6MqcN
T/UY9gRNoeT0sON6aWamaFnSI8yfXWaJPoSZfeAAIBEBaT9qAFpSUZY505spkvf4koSi7tOGFuAj
BL/rzfJQdBbWpqMUgxgcZxtymBq/nfPmBAYZPYNvMz2xXl9KHGQaLcxPBN/SnpqWooSaJ246Pat0
ReQjXAeFAqOekeyt2qGkm7qTG6uMV+lStEWQqtJORJVXqKXgEceICiW3GgmlIiGyuU5E3wvyh7Rj
kV9UQ22UNcTKmTnXxdkcE5/P7oSaBns6lq5cxpYCAhIM5FaZQt9zD3/JjxJx/KxbhDiMcFQIj9Fi
lLU1OWwJ6o5dMtbNhkHbinSy8mkMNvaC3+PtM7qrUEIPJdZa9OB9naPTBMDPWu0hFAzzRc1Y6LBj
+HYWqNYlJfV1MpbsCW4FXj9ZP5PeKy3Ks5S6XKAiCqZhtGJTdHJRTXhcbUZE//DJHDSoLUBapAkn
QQoRI/ICJIgByVBZyquQFpBTJnFAxl8U3fH6LPVVTLjRwkxYIISu3gJzjOTe6LajF7NcJ1RXu/QS
T2PAaYX7gKqH+PFU6QXcj1YZuqAQ5+C0Xu+Et16FqbBVzACXnDHLPHVWzdWLXpb8VwZH+IiIES4j
2QNgdO0mpvRsdol7/e3Dn+L1Oi1npoRE5iPvl2bc9IsGWBi1BaSp3P7Up7RsVSqVIQpze0Kg8kdU
eA0llEVgS7HhIJaoFaLISJh4AD7GKnCZMeiwXHRseRV1NjyS8gv4XgULNNlDIoKynxGYZAM9AbqX
BR0iQZUyiMlsxZCuEIIrFcItzr2Hh1MCttD+gobpevLWkkfgWhio8/b5L53UJ7s5MmQGFj+/KZwb
tOsVWnMJoaHUnFNoSJrlDayC3OfI7chQrDfv0mcPfKDdNGeg2ZNAmuAqQrp51MDb5JoVaLUjT00i
hbxo2NnNmnrDP0s37Ek2i33YIWC13N9l98EVrlb/Q2HkpuxPV1608cSBfCTMpZOoMwaIkeClBGSm
l2anZ41YyzJ00KjUUEy1ME842skB1KSXJgr+6JrW6vJ3U8SRkaavqDyQE2Bbfi3Lk8BaeS8wz3io
oBpewoyJ7R5FKI8ywQ/KXaTiOfNdUYopqfrrz/3i0VRqYFXfpEX6WHQ68t8QntvH8u+WdUAb3CWY
LTTQa7gztvXuVa+QzvsbIDb4qObKlddirthKCctt9wnop4HKN7p+1Va6vnU6ea0fKO1FzwsOkxO0
0cQU01zC8hMPSPSznv438zp5T0zsv1pO70vskgLCX9Kpkfvb9b9/wdjszvoY0N3JteEB9HpljqIi
QPaJ2OtT1dt1lanEjL3+zaRaH7CDie+uknYc/Kni8TX8qcFaZStSAw+t+xP0D15K9obrE+D4CaUF
Y5PWPYzEk9MD/SioI00RbZMBt0f7nGF4ih0Fx0fQwTjsxw/gKICX7OmGAX2Mo+GDXCcP2n+pBSf4
qjIwCX979ipskcBF+x4GTAqlQNYoOSojWK8b5d+/M5GdP9IyuFIXM6gnhek7V9GNExCa57GPCy3v
lisBtcufaslFIKyhI3EkHA9Bc2VG0zxP27o4kvi3w/7JDs4jbHKSWwgoTRCs8GLYYxZXEym1oZam
3dshwC2JZFUhSCKNxufhmmpx3BSCZZTWV6Lm0s2zYayEpX3Nu9tHEmLbVbJrCL7Cj8xnurnGbHRv
eVZlXdK5sGh/C1QlhKIGR/gUTZNInFkdNT07XXX1N4C2g+Vs+dOEEEKOcLPHf96Nl5nv8ezjIu05
iUF32CE7X5YlO7jK0wKt0YFElyVaodbPl0+ynlMAcI30JYFzvNpzUgQlhhCQYfiTS/qixqvj++IN
etmu6DXoKIclcXpLoXwbnP62QyDKkVD8K02mdXC0LgFe7jDZt+5PEdFiOnUThWNScuR/2/Q7kFBi
TLrRgBQxBgGxRDxvsNxsv0bEsXLVkXc88NkHrCc2Jqflay0tdED5d+HshxGbP2D4+GhKXSuAbOaC
MYKid7ClhO1f0pG2mQJuQx4GYrVXhUGBcycDoQnLXwCUXFnNUqt5wz7fNPujqkc2VlvjNMsmLIC3
N5ovqAWiVqhXnV52wD/JvXbvfsHOoEPy3ZCjfQNndOEiyqfKtkVZIgqAxzVuso/NrQ8UFNr348Ib
gvyoTSusm9feqmlcz0O4YE6YgvHcgFKGX9fY7hF95m76kacETUOeetmh7FFiunC4o1770sK8g7nl
N2KS7LLsaO+Ru9mPEaZXVjl7lleqTYnfOLXeVmY8A2EMRSLkt3fXygTykN/KUbjMdYLcJBLwqukI
Z5e5eeGMiw5uMPR6Cycoke4lKuW9m/VWgSsx3J8250wgl/8cY0oRBkTaAuAt+Ahe2pqGotAIxmvB
vhY6CYGz9ouCgX0Wd1hAw3KV8G8dRuBOmjLBPikzoL6tzmDGKLc4azl0VGYIleWZ6OR2DqI2etEB
io9xY41FcoURcwp0OgXJOPQljuee3DC39sI/R/Qn8SjlXAs/6rxomdo00slDcyH0ewEgiIfNt9WI
db7DZDV7/pLfYNUfx/WcZLlFd3wDGsStZtva9LPdOCo+GO7fFCmjqbSy4txXtsmVMkg2qltkJ7TK
voqANnxrFeJBZooKkaJmntb9OfeWosQa/oZ0evUUdBWSiMF6AahHX6rw9XBK2cWKWkdxxE2sRdEz
+5K6BUpivyYtzL6xsBvn0MKzWvk9YLw84INzVnV4z1pRHbCQMphxzDwN9QnhDq62vO0gH7A7ePR8
98qltIJx42Ao9TYrzaO+Md7vHUKnr+1j53of6C97TaMC4UHgkUCJpwp9cBO3lJOdfXTx4qXRvbJ0
BHe7r1Bxxue5UqgqxHSzafMa9g58SBnVdk1TXMVBDDURLpnK/qfjvmqpfhrmPXRBKMT5QiiQZeNV
7YzlNuBlolWi7DgwKkOd0UUJTRnQjD006/MjidWbAar58vLWAtxfUoyKZWgWAcz/z5WuwjzemyAn
M38RPYxpBOcztE6hGk5bGhUy3hQqwElCO5XFlO6y/KXtUrFcvF/yt5FCY/YWp+mVkbAFoGE+UVuY
Ozi7kgNWJXTorQawp/xho/FveD2DrVgGyVFfvvSrrXdJ8PociquJYsF4LjJYf4lDWLKg+bBtyNgb
J+qGd3s0OivmME2M+0OoqYkwxcThZ+wIMEHcOcQgWshMfF2GPUhPRm6Bbxe2pSZHcw/42Dudl7ou
mupeCB9VUyIln+7x43KUiqnIkgz+32OpW0qGbETxOSEpRUQDo3SG7wQdGXVCZlJE+Xy0QD47gZp6
IEUPsqJRgYRpBh//u6An70ou4V7j+Fjrpq1rqE3dsKiIIHMN6J2uZuSt8XJUEUG1eyF52uDNchPm
ASoCKe7tIiIIskifeaFNF1RChdisojiGVPCmLwPG/l5/qIygINABpIYLj8ryVYyEQrpTIgGuUxJ/
4ATD7n8cRlNQMk0c+6CP/lyz26a/Svulax2nsqemSpLq6SnrzLuRVlmtjqxv4DQ8HQswZU4XCZjF
C9cNEqIEdzlV6tC3RGS2jQwqmOjvnJDDV9nauueGkggsg1bkLTxhefhVayYoR9jO4vJjF7PwiJ+n
c7GhTvKGFDpzmtGdHppnP0rLsyA+kFBbokLfoN5N2wuCPJ4T6P6fBX8qpcsHtMsDvQcnVqzKzW6A
txci0IErENAQZkvERpCp8IwH9P/1OJ/bVyjT88P8P/5L41SRuuodxEd9Pux5z3O2v/bE0r4IE2j+
mkHYFCJM4KykiwLmnbeMQ4O9YGV1I3N3U8rhNoUmQbazEwVLJi2IKhX8nY5DUisVhQluG3vNHDlI
J7RS442v2FsXZ7U9/4TBpugPbQ14LUcdHN6itlP/FDRgtp0U8pjwcjMKbbPVAuvzJhr0a04hWMUm
LTBPyhGyE38poVayV9wAhmMuNYzZeiUy3qt9qjR8HluQnFRfuk8ClriGpXFxsfrX7TL8slMwQOFT
4Q2PJNfJ/M3fqG0fBGEjtBQUcaYZMtMKHfBm5ghAhr/tqpEVHf6ABVE8fxgZsHL1ELdOiXowfjN5
mDJltn04ToP8L3luVOp73gJPRSZ4PB8hfXnN2pQY3X2434Hh1YWFZMtuyMnBc1csjio7fhRboWGA
RS2cf9e8UaNFvpU/EeGDDIfxMEhRknLtqGGzKVTy2Kcp7cc+yWGoc8zJv/xxuI5xlWirAd7d/s9o
NgkIr6Xdu4/4rsLLP56kM/Xh7NUY5Dm5U+e4OpP5LPhB3+ufeo1GtqTl5Z+DXYGXm7x76/xUf33n
jWG6S8PkpedbXGBxDczjCpztQgkztUlcJSHjWmrTkzIVCeC664JPh7Ya3Iepf1mtrh2Jfxg6i3y2
ctGLFne9jHpLpUIUXiiiVnTWpaRdN92kA1VoWXXykw+SGxXxwcSGYeMNntHRYrs4/GeQLRCclay6
lh3VQIC5n3NoJyKOmK1jD7e5IzljqFP/eL5HVGG7X6LTXKkHOsYXzgqjhlAVe6MWuL1fEvrwPjQv
Pe0TkaYpwJA/CvXHzgTeWmeChNXLQkyo2SV3/0BQ24J8l4TowXhJAI//HfPVz+tTaoK+cWjemrtc
HWi44446fVgttad5NN8VppmIsPrTrQ47h/Kad642VKnMx4G1zas6ou4UXeMb0YdEP+E9Ewp9AUDz
0vqKZzhEcjzXz0Pg06S7VeFpo+2RMtRigwebg2+Gm3MPBa4r/S/EYUvSeSOtfh6TL6OKbHnzbRZ2
mVYMTvzbdN2i9OmHwJ6RiZXR24LsUW7xK+GcnYPnoNtqTII0GgIiVslx0D+ijxll5OJVHLjQ0uV9
Lb+m85rEP5Mun4HO2evJDAbgwKM7CRLNTDSJmHXIihDA60DYWJM5kWxS3gs7Fcyabto7OVY5VTkF
iV/biv7suWZIgohFufB2XLOnMeIgTnATuJskQMnkwipitwtdHc2y8u+p1dQyfJg3U21CyqTC0f1x
Ei/TGBw+44g9VtwJW1X7r8IhgzLW+8vzRe+Xc9fqcI1v8W5TKu5Ak2g2+1f1JCXEHcUVOc9cO0S/
D37vdw1+HFkzm+kIvma84+gyOje4LV9xThTQQSI+TmU/T3CTJDv9e/AFWHqsA/rgHwKCO0LwuBwB
J8NmtMRhkTYJdxI8Aiz2vulWwAt+d6kYmyckqzVCvPyyTqg1hIwQoHXvXnSLG0LKZiubvVKkFPUQ
BpkrC2Qr7K+feBV4FuTWzIk7aSSZkEx5Jv509vU3yhbuabtQrpQc/x8qRETlSexga+Y6Lq6GIsED
xu+KYK7mO6fP2u/fYrDCV73VtBxOBc+tCTKMeF7zcAC/VJGaOFdFHDLu2d2NWd8SDoIVovhN9Ht3
kPJeYCHWxnta2YIsyEdtcnnRdbxk5blUUn6VJhu4WHxhnOACc3tpGls6ZFZV7g8CVtlfdRHkrNVN
OsEPCZ6Sp4OUJrYL5hB+iwj9DJWNfI3swp8c2kngrYiIneffshOVQedg6Mh03S1WXQU2riCCEplJ
AlEg+Wwdiw4E/tFXwj41Y85lXe0l1fwH9TMk5Wwry2RBlDhOi6Nxj9MFhmlAnLfxWDc47h92Ho0L
aRbMAodqIoPgcDicvFyDdc+N4bkm7h0uslywA3C9PRvfg0hC8fWjrKiYD89k2Ds2sUDvC4y/35xy
WjFLfFWNVmuGUXSx/U+pJyurstjOnd10vCAHydI9AAtD3vM8OtvmIr5MHaoADluH2/dIxjGJHI8i
D4VbtFNrJUGTVFpipgzF3pCptYBQrkdZbBHliPO6EPaneTd0EqNd5KcR8W75dThJxhrUhX4ZolzL
Q6Iaz7u5FIOTD+Wm3GpDtmII6EVdn2KUv3VOopk6Rn1FKBkHAFFGwQL7NIRZSMXexAZlxtkC04hZ
19dpNPEh0+dtYR6XR06sD2Q005qLmzxaLN9T+amdP/7ua4DUgtElBgO0SEKg+BXMcR0KVX6xCREf
Sg+KuAwfhEkfwn6PNFNwi9lwC8WWRYf0LQehuHqz4yyDm6ouXIUgfxUgoPsY8/REaJ4a8W0bncW+
lr4tLVy2CjloQmVKFeCUdfX7h0TCEa9zGUI0mSnf1XIZUgPsodmY+ivzJKD1rPo29liLfvEB8CA0
gTrofLa8IG0JuJ9qIaDOh+RW7MOfQFfhiyUeA+7RCQobwLR7g6IET6Y4BHU3zMFtg7Ys4kK6UQZ8
5FShEZCzwdFcn+yCcPndv+G6uFuvuzJ2dpDwp/ByLVIc9IUQeirYdJXfEn/BKs42GP3PrTC/92YA
HH22YujrKyjTJh93W9Q3EO86ggkpeYw+1Nycq5xEUOREiIPgoZGCj/lX0HYbLbIWFssMw4JztZkh
6fxkbryBrWVcpnQ2XSxqxTd6fLYgS34w9XGozldrf0J5nHk98TmpXAZnopsUT3EyT31RMIL+WbZM
H7gs2Bh/ZdYklbkWzlKXefIifTkIXMrUrhSNpM+ym9e+msbtvzeW3kTnXZPUrfSxILQWenFyT1rg
7jwZaz02HSoSnKTebMm+JsVCr9TPQ37fenIwhtn+Lwi6G739IHyCttK1Zv2KtF9ydYPLKABfaLmp
y3CAPoevDwcoxGLzcTjkUZX/kDBUQM50GDNFBSxDNaW4y0af802lXvBeXDBU97o8dWngylhtzMMX
yDLXV4fmwamkxsihiKkmMOsl0EEF99inroBFMyuqwrRZqqAIf6sqhAbirf7wIJyFHDolBj91jg8R
4dxQEuWHfOFy1jpSkALp7Sg/diMM94wXH2TQ+JNVz1e/S2c1zayngnvGgx0jQvpCO50tX3A/ST3A
JGqn5xM1Zrfe9nuNfJi6kkCSwmcPvNzUUv2nUWWSmsdeccUnuP9hBWTbL6v970zU+vZAQm9Kbhku
LmKdKK4p5D5HMlMvurAyHMhwN39c6Fvva8B8hkr9q+CVW7P3WuH9SwTDLc9HgDtDH/b7krSsp7Sh
WQdKjEGAgeicis/7uKnk5SemMjJ0TRA8EHW2QOQ4Od5fFYSPgZjqrcf/EkDPe8kiB4Wykn0uVIPN
JZuYBXEphOAiFswpxWFLifPW8vkWLOoVbJQNuRgMCz0FiAfB0gEFFqggnCHwsrphBkwPJ0ZRFIHS
TKCoaOzTR7gdZra0uNoFJ2XT/yuFuyMHVuZHh80g8+UJ5JdGLiuS/ZBFfD3msuX63rNzm3o380g+
kyJlg+cHU/1YTt6YV+ObWrjkblvL1D7dxodDjG6ld2FcQsrqveFhEbA8arJ5s3mT1o0iu3l8V1lh
jh7x4GJMsWNvzTrLgv7enNXPakzt+09xwFhbvYLVDY6MS5RCEEyheW9VARDdL0h6oandzWS31KAV
XlmZW2pPLXph+YfDhs5vI9K669C+vFM4ZTgxLkFY6E1GNodzM/hlTkiJh4b8XbXjOTZ9dwFakK/E
5dB1fssZY0/eTAI6WRoe0IKRFd0XeB80sDm+0qkfR1leKODqIXU4zkjREmnPtAqynbEwfUehtVdE
SlZOAJytN5TCoCrAr2j2FKkg/AXcZuSFn3JgKpUpUXjc2q9WPErarRRoz2ude3TJPlJG0KVu/KDY
ytUxKsbMUi3JgDKlAuOLzQKfiCsK/MIiAVbmaQz/eEtZjN9tozZxDshSvw6zZGT3SfqyYcj/2bLa
Imi3ZoBeiyTeSodbhaaNIZm9SQhBMrgPPihNZX+eeXSjf2FsdFThQbJfDwt4fa1ISJ4SJ2UYMPIU
HvOw6ruLKjdIZr9DqN4F9HFqxMJv/DlwYfYGYqyQgnajMdB75JQyJzLtp0wCFWikriu+nt/YlhGN
+J/yjk9QLz09el05UentoOvxHQOYnJk1dosQ0Xnu6tM/PeefB8T8summY9gdtqMbDafcGvFcx+A0
owlZ5XVEY4iGZ9uSQmqmFvx8KZZmj6/IUuAAWeYc7C/8RGMehT3CcFcrOeZWk/AvbXd/cI0iC4dK
3aOIcnX8xzeT4UEMO9tne8CPIeVu3qqQKCq9TsWGItKxQLQF/RMmcCWnd6FcEpqmwX+sLfYfWjlO
bpq2ZucvnrHy7RMw2dTAbnfjZ13ojGwCDnPfB3LA6f0aAiMCDzMS2ivolgHw70UHDIrKNvyVhUwn
p9tdxtdXJtzQ5O2WqMf4XTflLh06koUrPmGiF6xWSoPl/R/H756VJcf2ImR4CovZGciJVre02kM8
qHorbysW0kGYJWwamd3WM4ZBaRd5WgLaHFuSn8T4XGBrVEAzvL7OM/UQOusPrhGDIP8ZyrfLgX6u
GmtWyVAPYTCFCqQ1iP4DnqrgInbQV0MCrgnazeW7zEMjxR+8Hg3GOmoAYQQ6ip88xpUkI3PWeH6+
K+VdlBZorvK1xg4f7zxTVVcoBkk6QWIjK5pSrxpGKMfWWcpRkBuQAD7kPJxgQrcZ1MBCe8ZjtzXE
tkcSXIJHsw6F3SI73mtdgb9qccj1m8RxFNzBaZ0s/XGOVVQ12Gk+5NRiaAr+IHhCjhT014JL+O3O
K5asjRi1mxfnd74WJHeLYwyuany0UkSe41CW0gGgwnwLk6OHBIjITrZ1IUexzwg6NegLxWWcOrJh
ZgdGOvkqWWt3ValGHg94wumL0hWLYGQ/78fMJi+YTCmcYy/pTeCJMzFkakJQzaig5cImW8mLv337
i+9Fb9hPFRjJXkLLeldvzgbk4KrIwnJyO3HNS3EWhIfFtQHbLzROvUimfl+bWnJ6QhYZnYPa3/vp
/fglzvloLknVZG/zE0u6sFgMD/Kcf6R6truM1kE3NQ0kQN7XJ3NcJoN59QnK1917hlRIkYM3j8lR
zqLplHNq+7PU81ByojhuKVZ8Y3Fx16ADrKpHPM8SB1+j6fmlLNC5oaJFnI7T3XAFDmrq7YlD6gLq
UoprT2c4GwC8T6e08CmIFoojHsRkByCu8OUiDjjuSaPJzT+g2P232XctNHkBOqh+8KXW0eOys48g
48u2CzBj5QdpEu3VQlIJ15hy47Iqx0cQlrD5gMxnuncfmkJI4U9JwuzyInhECKaNmwQe7E0XniAy
tcJ5TDvy05LY3cSGUyIXA8QD3Y+HTDg7ApJzeWbtECbxOCOXAqe1/WjQVv5sPyJGuqjAbHBs4KWG
YffMgXwpov+e6NzAMk8PLq2zCgRS4IXotMZgfYLdpSPdAmXQcin7gPrmEGkYYFAp4dLIUMkcclKK
40+/eNOAnCxTQG4ifXl8DuQDs2tnADv9o/JjHZPO3CtY1LrcgbUhX6IYGnod7caiLjTJhxTS3USN
RAWangLdiscgUmiiMFgKMdu6DE5tzG3IWZ8kqcfg+uivD2ge7YmVdjY8ejVezvHd8sqa0wxZDvpk
Jo5fCfnh92t6CxcQIiAb22KX6PpAh/CG5oCDjFvPUuF6GG6oxfX379W/M9zMjI+q4djA/gbFcDDb
EmY/j6r97vyxqGUwNc2oeYDSDnfODdaGFOnrPtSxdxvm8ypVY8iOJxqenLIBXheNtSrc7Rr9o+Cz
t37a2Q/xUTW3VTDD/HwjFD2heLZtOKV2RHf5ac2q8xpPQho1YLZPFNGmyJ8cun0wb8RU6zJly5Uw
MMOMv+VSqAzzMKBtc4vlkGdnrkOj5hKkikR4XRsj6+T3S3gCh6swX23BXKuY5gFnNV1hj5tv5uM0
E6RS8FUvjrdHVSSyhFilqfr/2ceiR/4+ZPIBCkMRDEfIOMWdzO/WmMrWuvgI/8UE233sxyqhJ/X7
DP0F2tXvf/kG4hGaVPX88JuBBzj0HkZ0v213yAxGHFGj8pzcAfCwMHebxMwQE79EHDXx4ocU6+Yy
oQhAJmI+03ioXXDUEhg4Dmigr+z5v/d+5F5Qi5YgVNWPMlxlCkZaz8Vs2zQtw1YjO/hHFLDV8uqC
CJqvNlEMwU8O02LWs/S5VpJHiH6oZuJCHczTyjivTsWaWhtj8Z6LGnj6kHsCVBp8ZQKiHHc+9w4N
T2ZDn6jZlIRL3ktP1dqORVmvfXlUYZCARxKW+VEo+GKt7sFx5TZHIMScErQf9op8zq7bHZVDkDP7
9vpqhVnB8JqXQ5f3cMLv227Itr+9og3TeC/iZqvxsWEXOgWo0d/gYR8LkcmAmTBm5jo9gqWF/s4A
3jXSCNgGNMnhvb6qjiwDIlC3fZADlv+4WUDhFvDwefZiLCnUw/SuFuVVHD4I3MYYYG7612Vww0YZ
cHYlxz6hFbwuIj4FpBfqptb3Ptv3bdqYd9sF9z2GBfLmZT9NqbbFm1lm8F6yRTYPpWGpvUBOWzy+
ozKs/0XdUUi1rbVocYtQc+DsrwEcwlif+xz2LRZ+v/6KYaW35QJ8o80p51w3gFUZ2bnG23b+vJEA
LJL3YIf1A2iq/MUgfx7tBD+0KMX6Pa4rIoJ4emkwx7xX2R/cig726YhyeDnGbaZRrTv97Pk6wLQO
hQNl9s+mpBuJP+szPAcWNcqRKdNnf2OJ91R2hiPgG/G6Q0iDDjD/nrAdjTRLibQDSrfjjFrRcFRM
eALD+f+4Wxo3ScsijwbHU/IHDDMC9FSMM31CS5W+fK2MPAm8qkI4eA+OwoVnCv3nXT42fAY5tq1R
hPIIALKlyfG43jowu0UEOtpmblJRwllatckzvXCH8DeU7KoRTtDZHFIbXCUdLi7/L23yboxLi1Dw
A4RAjaYP1SRiuIVLXY4heWM7vtN3QCno0zBSocOdYkOjjWzooOxVIDeowteCto1GSt4vRVfs4vPn
/b05RA3+9YnHfU6Rbb+E8WM4gAgSkbIAf8tHYPlzqlw8MAssfquU5yZA/xt3u5EYGFWv+6aC6qkL
BxPEuw5iS3tEdtsl1zjWQnYXj3cAivNkuTvXe8zO+Rtmrfm0/IcfsBl6+7s2WpGXpvcKfveZodVM
5oa+IPdxBOWrYFoKvMcOnqINfDvxbAB8rR6ZRCekp3QWzUUwjN07St1VWfjzRdd6LXAjLmNEKzxJ
COiJM6lL9tcyykjvLl5MUPzOOSKJnNeHtackv5kqYhmukINuUpipHc+kZvvx1ylOjfO4WjvZ/Jc4
oei71TGLGoSAb1ld05QYssG0t//qSGcqEuTMryBU8WHi2YIwIf3GPS31oTQp9qR8ZgOJ5MWqfBiI
eQHkl+0gUQFMFDPx3frRSA7RYB8nicRa9OKVV6onj7+wWj4/bLpsec/BxkEAMOFeLtgRs3PXOGQV
YNG2lCG6dtd5ex62tVt+QCj2/XYDIqVHEDMWKjNJyB28npebnFfcXFk6brg89dZzR3Zr88tp1QW9
312RR+Nq9L0ygF1dQ6azx6tm7vVRTx51Sj6qF3IWYUdcJCrNUpmfQHcm0GJNvESIRfh0sx4TrUud
fgo0UBiy7pPBPkN8eG7GawVBAcaTtCeI+FnEbBZUlWAQBxcVdoIrYqOsC4tkFd15a7b8H/Vx/kbP
FReya+7GvuVRppYOXbvFqhDAuSgkttPzjd+IowD+I4yiyVXRnTcUrZ15yVnwENf/aMVGY7LEkKX0
Nbq0lfmIRDVTpacTWK2v4pywfEXSjw/+Tmqh7osM+c2XnwEYGz8eekQdRtixCRn93iYxVivNL8Hg
6rj0POabbMBwrbRY65W2mVNDj0ohNUdgC5R7LA8hkUUClUu51PEVpYzqC82IbwhCD3eeeQ7e6tXw
qGxVFtHoQX9MP11u4DmYlRZvi6h8Wm8+S2v0zYnTxvLIWKZSyEO4DyfvtIuSZ3Ivp+am+ILMTyMs
TyREdASuzGggR4AfsGg8qjCArFfR69rxmJZOtoeZh4LTAy8CHicvdoffz40fZ7wEcfaq/CYYAm+d
I6KoXhV5sP8e1y5w3DfAa4+JhGmm9QDR7X2W67z+zlp+OeIOYxsGZ16W/80XmOcVTkTDHlpknla1
6RB/mDcbahugwIZYNm3FDX4eQwhNBXiStKX09GyA6MKYzwS5DD0oco28KABFSfjtQNSiYlP+yp9+
x4TbpISuEGfeDR1p4jgOT0e603ME7lxj8IGnXHfcEPA+QeU45pE59/Wr8E/LEB2mXWmqlSmR69Pw
xg/PR42rzaV0BPPqA5oiaQYyMIb5I9kaPkPD/bfC5qmtrdlu1kHWXceJkheCcCo7K2ZgbUNT/P9f
IL6vCGhhQWS0pS34zn+FBJx/wshbpfLfk8jOW8wfpI86YTPjM0BM2tLgAY1rLJUplVolX3cEX11a
xk3kjjlOmJd3QrRadR1gBwepMlFvRS1RYA+0ukT9No1eQdaE+bwKeRu1relzeQ0dD4f6oLP3qe8T
EawB1NNogYGgf52munN4Z0GruTee5ul9X9PhaIxHW5c/RaHHLsfWNkWwUow+eeeV9vZcvVK/blHT
HqrNx5thnlH67eJkpYoY/ZCsTwtII8FKFrm1JrRJpeX5HRT/+P/qDXU42OVgBl5FANf56HCzvxeS
O/cKygmzgckoYKxyRR6BmLSWwZumMKh25mnPYFAjavrO0NmPrrGQYak8JiknSfaRMnE7cJIMG1YL
CeCXb4TnKFxaY5zMWm66q3sgBo26zbAPGb5l88VD7rEGOsosQLgiYx85RW/5gwRanquPs1lCe+wZ
BvK+FTywVpEearV6H5oLix0NuzmJaGYkX2g6KMSohYbR/cD8rnihDmOLKZnoqKhrW74sgb8kKM9V
zxJbkE8p+H+ev9PdqHLCCTqKiIXT5nrzVYgXP6hl3fWBy0MpDn6F9JESBeNMjTwDBB/ov023ERI8
uYRwTMNCRdguI3dXBh1l5lGimO0EbtwDbJb2Sf/WVBrXF3Q3Qfd0R9JkqNVS0LUoJFEcMkaI65WK
lEdI7tW325EP2qpfIRVSciit4tCKppDdp8B3IwMWqLo0YuCmkFk6kJjc5Ck5GLhx1SNnuAE3Z15R
Y3inCGsm5N+DY49ReuEEbP6RAW9KI5PTWZ3RzoXb3pxHebMgSIP4ykDh73B4gN4lzgppWiRrwioO
LUGjc1cMAvvQPt5JknA0njOVtrQMYPnf1gyY2+zNU0Ttc0uBDJc1ur+OFwn2QE1WYXWm5e9BlPvg
ZVLGe0KCmg945dOz1uerLJD2GaEZiSAq95ZaLoxlNjmiNXPrrOXPncmki9PkI0hqMWjxjjaUP3VH
Izy5Oirjrh0JhmiQmWuixxjmLmpHWJ4JY15m1z9WyBzUL7+drfYloFUcpAJyb90bSAfEEHey2Dgd
TzhpGHxZiijujUoAnTE42dpI8hrZ7eclMfDYDFVh1Hml+JGf0glIl+JZ9YDTl8+lYaPcPfGXo+tA
FfXVdh0y3WUGg0Rox78pyvnQpSrkNJgAz2z9BEPzO6eSpT7fHQVZhe7FQSsFKJSVYS/SgOB/XDGQ
4E8obMc0hobwUZQR/Xfwn5JMwA83YLLf3G+ssGcGBdGET47m9Y5VOLVWqIO4Yud9LdgSr1C3vfAC
KgxHTzON/mjGU50RqqhzDkJlJzu8yMy6ccqvo+ZxO1IubZf9GOHR02evZI6NOIMn70d1P+e2M3fa
ASGD5rKHXf707DxJHFbovOW4qQJYucr+9GRsrez5quCN+hBow2ikTX5ula11Fi7sDjrRP1sh/ddd
APqeN2eL48K1rz8xgG6J+ngzbxS0LtzDWDiBjk3XEK1sJPOZ+9vmaDSPxZxtxgxGNSfCjQiN3gz0
JjKIRlF2WePeY0A23nMyl2sZrlQUbTI80Ocp+Sf4gMAgAOqDd5HZ9yAzBrmCa7FOvMuCqkCjZVyt
Vin3YiPHrK1246EWQ5kcWHU+7NVCOPAY7o52AXNPZ7GggUgBx51WdFF3QFaWzppzRmLx0xeTu3Jg
0QPBUSg8Nihb3vT3ggaWIAnAwRAbuhfV3lGhwx7o4b2Kusus9KsP1zVvr6L4X7onX/wFRcaO1/t0
L14WikxiDQgfHspWaXMdsIV1zFAXaj8QQ7W1nOUs/yrkWVDBd7hQHbGe4KqJbXu99kccr3Kn71KU
+vshpmroHN2hDhpdjUpzFXGx2eOTS/7OzN9aiPf/UMuTWGPBkOwzFzt9NUc9SkVGAirbeNQPxq3y
QirH3vPWxTEE49MTUp6dZHjEmZLdnS9FGD2IMgLvtyhdS9iYgRLWJ7N+a1Io2hDo9fAc28YR7/iY
74Miv5Q0A2XARtXc5l0YVghgxX1U4QoHhB66/jnIqcoCHtldkrQi4DH4yO2CxSPbw96sfh5a4uLW
SOJlbXPgkGivfzsEcGeabVgV8+8sAl05UlXs0h7tWfmQIJDBYxSbHd5+/QbDvPvaHEvVBrDFz4j5
Ov/Gthl7C9afZ9eRiCCrtzEMGWlTbjrCUoIUQrSuecakj3Q68IW1JyT2uznIIEv2ES8cDCFPJOQN
L70yS3c923H/zPet4qpKwYX2n/+nDr1yWa4vQGb3mVzFoGhGuvqxHnQO9vJOTwMoZj/XQgn7f429
PAdk9pFZ0lWf09hkitIpmrlRViMHlOGgxgoFkHjIabUEsNnNURDVMFI5gRNUGb4fZXO5uJMotvC1
/goVjQ6y2dJi9gZW1OM2KiVY9p0/WVlEIuv4VfTV8OT1Xfwc2HhoMPrK83SuAgTNsmtiHrvc/lQz
TW+4McTB4y5udMpu9xHseOfoEpjAzSHGRwlAbre6RYnJujbB/pSys/0pzmYWOlBMa3a411LbXmhm
/bJdREbpk05Gou5K6+Y+4dEaUL+5X4Gaw9ltPNyR6zYpXay2DZMF19ZRqF2+whK8oCLPLN2yuIs/
ikTAbGUfhmlk5v4XPvigUbYEMEi/Tjg51uvm/L4APXPumDd1G6rnSh0eYKfaU024omKyBCGVAyWS
zVjJ1B6Mw9fsVYj4grzVFvRAUlh/z+17KGuAToefBvUHJBEAE99rNoBDvryIgGw2bpmNkuvyJPhk
FSkCOm0DrkAGho0ToAz0io9zUyX1NiXN5bxzJe/+Vbaj10vUauc++YFqejxfN1RnjGsvr+x9cJRt
y8JGLSM9KrQ20v0sIHP3ygNLkmZSuo5rrfS/ZWPijFcwu3kyL4idnGqkJu+RIScZSBryCvC+Vv9p
o/FYiVP7WxigqDeKd2XuRYN2xrCdElD4tP5NHKty7/f+tR54gkaYxbdfIGXuE5YkaIdfoOdS1p6L
+8TL4j0aofaScjWeO94T5UaIrGu/h3/MpJheR0JerQTo4kW+432n4dWKZzhjf41WqhatXum64/gk
ZH3qQQCWzgb8589uP1QnESAXu6me7iuJoF2L1449uRZPE/P25/K0BweMFH5lhUTNWilZPpcs0puD
FF2Vkk4y880QavB2p/v8n+YTulQRlvxvc2dnBe0sgzB6tdpiuYt1cEkC8T6sOmN/z3abXa3xOYqH
Hcthp7NJJxm/ZhJWvjWG7GUgM5Aff6VWkodjzwTaW3nltC1CKiMAV23eligbPuxjPrwDqqGKtHLc
0cKg4EIDP3Xm5XPaeyaKi9enTLQVIBq39m5tRFtlBtZHNKHIrWCaDO+MqZ/ucZCJ7vFvcN8Tjc89
mXlZIfUuAO29VAQb3Aod+FcHtlg0IJJDazDcpqJOXHe4M3TABSqrOniAvfwFRI/gLdUXslFPV8ix
mt4Q6+jB5f4trtZzGFFQX0nYlVLsj4hHaEIXqw1LabIpdJgZVYOHeNVzNVm4w+xrHQ6x5xBjQv+b
Ih9jHxEFwiBsMqaA2SrOvVv3NENAj2AJWEGWXXneImqXWRYgUwkSAmBO/a3d+LcCGbimF+gIOn3R
hMKdpShaik2HyKMmISksNPFcfgPM8Y4CdRDrLywM28Ww6e6oBswEfqxbANcy2JrEM3Emi/0aHDRm
G+0GJDOyb7Qs+QzuMMnaID7hvRsF8k/q872jQW8PpkBcFJZ90qXcl5tPtt1hqmOmdpI3XvUs63tR
j/wMuv71i+8kkWQlFcAKoN5G0H03awdfLCAEfR7DKPpPMps8rKGdOyGoceT4XuvrfyzkvgORDxkX
Waw9+RhwQR01p0i91YrXMCXGjvrtlB1XME7dTuNNQczKKDlhz85NYmX7z3SDHNwuQrBX9MAQwOz5
5BJJYaSggB6963z8DPelIan5zAfkcD6HyyDLCMibFG+GIHxwndiXwM9lx4M7zvnn9MG6EViObXf6
7apqfy3YeITDvwranK2JpVDg2ZQUrmtbGh6x6Ar4s8zCV71qiU6QtBcVifDu/hs+UJUr+nSlIw+3
vYM+kPw8CPvPlNKKcC29FKcZX5wlF8y32gv9NhXVxgyUqw6/UvQG6idACCBY8E8VLpTMZzfr2p/k
deeFhV/zQRfl9HPPqVblmcONNQvwgggF8kfzTYUon4kE7VtKJYs5Ai1IDcNNRWwv6dTVGaeAtzd4
FtjkYtuXg8nzsz8eAjuNSXgE90X14+kX3tWG/C823J9MUgLHQ1bmTU+CjUtgABWLTmmkvc0w6lno
Bd1KE60rsEsn4/7TFHRFIMsqFYuX9HAwvn5jkjnAYLgPac9WoWIvEJkSDS9uCBHT2nUwcpF+pafq
Q3NT1WNtXNNtK9PizUv6gyxZGrZfztkua1G9kV4N39Def65qAJ2lvnExsOOnx7gibaPzTYJGCaUP
TeGQegdPLwvY5WeA06fy70cnMytVmgEfhDG+iY48V3fcIK3e3M9yKO/aqNm4Si0ReSxMANxDZc9n
H2eW0d7qoDWa0NtR3nSp7ESKdL1YFhvHW6r8tspf1Bgk2PEAQyUsuvVpifeE/zfOrZHoq+GtlcBF
OHGhtzEHoRX565N8jdio9ZOvT/qrNGDBnJUipm5u6ASO9QIZJpekdwmBYDY37E3E+Fz53Nq/pIpO
sGCI5HJMbiLA70QgsubPbuZP959IfpYgigH/WCL+PU5K35N44Q9NJxPV1zWyrf9SwK40+8IGDTx1
pZ0B9T96VNf4RDy8WrJVV1Sdp09Jz0ZeFTguMp37vlbUEQj1C9hNIegjAtA0nr+/c6PEhV28Ppwa
JJvF9dcu0Gt4Oc6DVSVAggBB/Cfu0rOBBBtFA2zjPejv+SPm2V0OaE430+3tEC6md2eyPtEJRYPT
jYLgyuO6Ixp7CvcI+WAQuzkp4qlfZylgt+RGtI/zAYBHTMGpsCHSTX2zU6fDYuKJfAtMjGnFwXmD
75icc5LcMksi1WdFfGcgASMpDaeyaEBpgLfy3b5FKxWCbQPZMwuApEnELPBg9lCc50R/mUTnZEGN
/HvQ+ZOqHTlftZzt+9i+JQiwX1L5hxnsSVySQJMQLzXLlsbLH1z5XsQPF2bEF5hsTGVdjgjMjTRD
/lnfQ87DQzBJAPstbqFDzVHDkq6SYVT7hFMVk4zDAz+X3hZ4cYtOuN0GBKWcypadjUK03TI14NuD
NN+g6Sw5OXs/M06FGmxJ4PUh5dk756iMyu/YGFlh7fYLEdVzJZ8LrdgnsZiECFFGTXSu+Rwjb9qU
cxMQx0Ck7TCujwFbkjUDq+LLhgEnS/2MJh/A/UsvQs9V+9Hlk8C/nvnM1Wspu4ac+5HUcxvpHQI4
H7Q/TNEWoyXTSGjtCzKgcIbZbciZZwrLC3VuiL7l/1SoXGiFVTZ0eEJP05/Gsyhk9KZnKC3pr514
38XkQaun83fxaioBv8cJ6lh+37fQxIwWI3qA4QuBypUOMtPpAZDtdHDO3azJVuqXzH72oK6olAHo
J1HQCXug1isO9FVQsUYWUsO8XZUDwoWG/FmRcykpMaMce2fWfqQWbBsnNeGTXdFseUoXG5AZPHcA
n61BED6cfNx/0paZm+tocH2vhg8aApUlaULTr1+j4jcDuAFruYkTQFQzBB6Hah0VjMidDJNoWu9y
lUDqrHYPhWNuLgSJHltJ8PqL+VKN6r8ZXd6bw7NMr+24E8PrCtiihvf44qGIPRHDYK9i6C1zaddm
S45goQz+PWziF86N27pUgtdhgoByEegUlZsD43dbfLng8kla0mA7qS1U8K/ivOw9nVEz1LDc5JB/
xm15jcW+B1dYeMh1LOnuH/CMgbNiz/m121kM8JVfqXmrnK09hXwFWb3XY+Z+O2qEiIDEN7p//mnq
pVAAJlSBJUMDmLN4s5u9tWNkJ2AVp9653shfedM/8YjQOhuk68RqeX/prLG60erF3DLQ+4OZrPND
dIX1QOvX6RGZ2YunMfW7aDI7/LSAn/d8gX2gnccY8HDSDu3zXgLYDGOf9DSLrJk/I5js8Xghlf9a
IrXe8B+S2QHlydqhjWinawP4YXHsii+ODNdw/l8evsMU5BwyfvW363Ma9UdV9gUsWa6u0TSHR1T3
s4ysu+A4gAdqWyJP47o6ku0pAgCfGqyQCauHkHg8+bqT4dEDath8Z6MTaJvO5wJ3BCwsu22BqbcG
uSJQ1X2ghE39jTrVRY05KbUT1PVW57RKYzw+yBNRtZhiEjb7RhS1tVIzPipvc/fyMwJy4FaiRGgZ
0OyUKc2NgSi1Gpr1c9jzPoKiJcSpPyX0UXnmqeULjDgBIiEp44XQhOCWNAD9nH+sLjuA8oeH5uyL
xc88y1P5NlozasQgJ4rxsk52Fq/BGwLFyaHALvVhRDG+UbDO8G7GyVm01KYcpp3kvLmaQFQ6W6Mn
nV1sZ9FDBWwsdTnUqdGU3kX9aytNrCB+lEC6oCC1ifyEjnTuaLGjFY9UBKKbnmflEidrWi2k4Vm5
CD0yt+QsCqapvp+by5d6Ya4Hy9Ixx+1pcF4eP0OO9vU90IcL0MaGhKGepzcl8iWx0rVI/1V7zM+X
2t7oG1qbMO6Nkz5Qs+IVjjAsBxixsVUeDMzUxleSXYcDLN+KH1ECVnlYSAYs803oZgAc0+8unGhX
QF8us9MrzSaezNnbPZL/GdA5nBGd61yWVVh0LnA6fdxHcUsL/WaCbyQQDJ1xwv1c1laux1/MtZDn
bizVOmlmJL63BXxIdghEI4SSaqdy2U+Fx73Vj4pGrCFNbLAlNZECTnekKMBfxXKWppqq00bSQ+fv
fwJXZklwmsi/h7+ZI0fIEMCnyV0BRYB1GRlw2dVAlXmGoUuc4wWO8+H5bu2d4xgqh+3bDe1ayy/r
SwHiiD+dUVrnH1Pdm5fjUO3GwvzcOXA9cMarshI8vIWv1EJWXlTzRKv8i3PWCfv/WS3pNNNlhbxF
vMyskappiNsu9+QSRV3iZKWZrdZApttDvfgKSlcNxhKW1qxNhzlWWKN1s++cbEEg0d9XxNclxAR0
i77EC4E/EuJHR0gLBv3q66r0pdNK5el9HB1FSUwQDwDdui3x/pYN8HIi1a9pOIocs0DGk9NmTTwl
xGWmfEqxZ7rbLWDA105gH9XpysGZL0NALXodJ6G7uJJ2un7hFxItvuijSSak/9Pml01mLrICL5oM
KWNP2y92fJbwKmU6yvbh1MG5q8uLDZV5Ujaxt+5rLTDkrV5QF5MFTZQY/PZIDco0FzJVS/lEupVs
OsL2ROSqtMn1Xk80Ob8YTO8wgn3MGk7iXoqMwt9wut+4Fyx7n9n47lwXxGZm6HBs450fC1Ph9qc8
0FfgXcUKcqBT6m6bhSdf7S1h/f3hWmhGQ2CI2AyD62SbAyS/ichKPbRIZAEUlUijx3xB1kIj6giR
bkXAHj80qlryAeNE8m0KKc+LTUa6P6PBQtivrSFs2YcjEQJqjPWgMN7AUhlJfRQz0INIGOCigdET
xFkxheF9kBHhWCJpkRE5jJR111KUmrQKcVhPcBEilJqCXK8tYWJ7OVNyehd8nGY90Ku6ltJfWmfd
PNHgTfnAYiffzSQCQKeOz/KuTXcjgh9KvbY0a5rBIqfRq8u95iR3mTFS4cfE2fug87XHjS17jQDt
F4NgaFIfqUEKK2/gM5rVquLFD7AF8CLProFfLOerFdriurkePT6Oiw6m9vLPW/f7jxrOcg3BmtmE
x9CkFM+ynEvY20Z8oGdXuaPe3OPvr/B3i0aGZ/YoBEQYd8ymeG1xgvLf4ej5ERaS/ogwGVvbf4Oi
vwpgFCsoS5BylUxWWID1E8ILBnAakUa7ZnKJZTQKVjKdAN4Gpempgrkahsf6LYlxaItJELBdowxp
TxyFOvCYyw6ZcFfy39x4S9Sko29548TOq17sGdp6khLMnFkdvvHlx50zsw/6IkqdSl/eOLmL+ZKI
Dd89sRwUsLOzSDI/7RAa9oBCqiDkNpR8d0wMDGTz1ObBkU78YvTxLhog/srDqwJwkvkWdoWhJosK
Mhnkz5O8EuzWxOHSxbhdbBupNBEomWFoz8KxZIJUHAnt8xZ6HQrLAi1uPQShYg+4hHzRHMu3iX6j
QU8hKbzrWoePnHc1vT9+2DE7CeuBkyYhNbwJq/kKraDUj+jZIxBF6c2+PciYCuW6rrHtHDUo6tDw
HEoN5h8wKzCgerpK00h2DMv5GApw+t28C28q3QIg7/aN0YnK74lWD1+O4tnuU8kH70N0/3R4Vy7a
tYcWSc7eaG5tfaIcX3uC93LzvW2GW+4ZamM8dYaKvD5Jyvo7QpVQskBLPMn9a167yT6OzzLaKwg6
XLnH4zZE/fIbb+wJDhX9HwLUslEFBl1tDIk59YjQUcHE+QZsRyYDENx0apIrNKhgPTwC/5ub94fn
L9GG4GCd794dwd2vB8hVBzGiuLhTnyO23zg002OqM0hN3GC0ya6gtUcA9UhL/bT08uefw7g5Ujv5
cDzpe/WA0Gw6NIB2xlSXowSQaBxNeLZR9qKxVqGdvL+kHN4VDkswP4d9TbVtm/KGq3qe75l2DPY0
u5zQT6ky6xbH5MdprouEsjfUr6Ib2YRNvqfAoxchmpMi7MPVIbaN8MpD7YkVSDv5PvQwnzy8OfmC
mlpWiiUflDJZWjgd66Dhmg5H82X5LIq5h7ATjnkquukM9evOUeDSqI4lPdyNQ6jgKWMDUoaaXAk3
yVIuAsLylREWJUNY6KlE3n/XgYRfzCsVICmSsx/cf+1H/WQh3ZAF+yZtB1KKVxH1s7mK1lxI21QG
XFvVe+KyvCm5JFUnSuLRA4hDEkNTinyriVqiuBGgEEErcrqfqGlcaLFXkJ3BoINjsbITH+cvSPci
1waq0QlISTlPEQ8GQUTj7xdCVLPZ9nSGhaMBkyiKOkq1OkN3O/qO/+exg7mzZJAw/5+/duf8wnPv
s8np9NTcKjymU3o8yxQMlBR4ELec/Jd4gdLTPKTLijTNEbRp4SiHTGaBKH6a9bg6x1kljkefmtXR
2kEbEaCSEwzUZHOTfUd7WPs1xvw4W5qYBF+6zfXOvlyXDUU+AWwRGKwaezifcc9tOISD5sH6Qy+u
DOO2eJlBeuYAJRRWS0yqbiwhszx7TPhBmVjTsv6/4bganeHIeouOtmjkem8Ic9cD1cJXhAvnJENM
O3ZASlqT/LmnteiFSckKLWJlX2v5PPC+gfAHnE2/X97GJT8YufJ3CUH5W6HWmEKbfeuxAPDUkuCO
VJPcEx7Pqq+87dy4PY2II34RZuGopY+xp9yHlzQECDd9Ki8we/kNlte6L6sfJtLL1OP4wt9ZlkOD
g/K1+pZRrHPnBaurK19ZEX0H2t7cQ/TSfk0aGNFf954zHNoBIG+YABf44iKBGmUZNpnnMYPg5HUk
L0uBna7nNkuPJC8VRo4wbFHabf7JDCiSfIUYtjpy+leJNy+3btoB8F6rpa6IoTepQtZgv/CkXRRT
6a0E6h7tXxohJJpMvw3z9D32v9sCqEXHgp+8ibqHOxOm54Nbr72RQnnrVfRqQerXI2AT6MMt1rg1
fpxaKTU7q7eFuLMQvFgF8+N7lxJ/0W8U9vObuE3GQSVOAnZlNkS57uRvSuRoPfe0u6F/yumaEgKS
d895TltdW/TQDddcW6vNmwUvFX8HaYyENRe3oVHrtoB4cQesIDoO6S2KskfnDMPmlAz4YfSB+5OC
lJYC929XbSEh2WF6OqAowdvFUiRlZAFCN68FITT7nYPvU99yLrLOgB8/yVpFcPYmaNr7+EQSwW37
nV5NgOjdErVFCgGy5CnB3BvTPKdxBrU+uozi7dGps76wd6L+Tv+4AAetmFEP6cFtnO//Sttikft+
C0/LDVUfpM1vkS0L46NR2DHC9DXAFo7vAbE+shiIqBqmX6Xly2wTcFikyWXnvOnpkcOTnhfCOYSi
Yjq8K5EsQkokAi5kh5vKVpOkvGPKov82lDHs/2HAJ6eCTzhU0yXT5UBn2kdYg9djP4i3z5pDD4tS
Z5nrkIBdlA1dy7U9zt9JuhrY/ZzNdjoU769y363+VpHSsaqX6RYn0JG+K+4XByZLltrKZd66LI3t
P7tOtUlR8TnIqyoJZwmgW/PGlvPNoQtWKUleu3sIckjpJ8UyIyNgqjrMyUGusVau57mTG51I0fZB
VotShKHj4QCR3lopgGeci4y5t38ylo+2Du6ElpKT2yJkKYPwTCjJSU/Zuqqkh6/pRQFwvYb3yh4p
g3/aMZKMUY1F4TKwDtoeZH/jGVBp1MqwfvlUiusDFHi3zPdqFNNncnebDlneisszC29rkB3PJ5Mc
ujua5FWQ6zVd5DbYanIr0rS4greE1AybU/o9kllmbZQwk/nhnFWTbOUjmJPYmNzkQk1dVoHTwhWk
XkXc9rVpwRtwzf1kIhZuaEDOg/b3NZypOz5Em9uciI55wTK+j/eCarTjQXRrRyH1GRqnH828BltR
+1tB/8YV23VuCfjpQQgP2CFx/sqxz6n2jllKAbOwyjQrtb6M3kPcwmI3elX7dDz0rDcyebNwgVeO
yW1s6VxcojrcSZV/NMBpBd5tmme8VMQdOuxpaG0u/UqLOWM+NSJPxd+bSm7ButhWobJvuvpLJfGr
/gU6PN3QyaiQWhtV9G47f4FUtzOVHJT+NmKY4lCkDI/8ZyD1ndyCsuM7Xgi0nW6QQK5Gu10EuvMV
oyW1qp/urauJZ8n7Qez1Kn8AD8I607/2mY+s+WqRuXfQFoMcmq1B+pQfYpeItW2t8ssbVQSk21l4
nBq0UpCCWFNAC7m8jx6poR3jrd/14/R6zkw6jbHjUXPim8xNQHc39Wwkolmu4DuG0Xhps+D2fWwR
3CwnlKlW+RBH18AmjkPU3FU4I5IagLenmfrgJoTeUssKOwMbRTV0fausp2SifACm0QUjJztPX53I
rcRaKFuTr5rAXDaNuaxoZns+88gmSGeu/IlRWW0VzDY0dc9N2+E+XlIaxUrbblC6WN0OwkEFh285
sVnsuwC1kDuCU267NdF1oRhHQT20z/lPZGPTZUZbY36yPb9FdZHiQuptsszzEPe29lnfWp0vuIoA
BLbwlkrjRjWnWoU1Hq3eC486oeffFo05X/NHimLGn2kP6m1QCtkeX6uELgRxuHNx949xCyZaHc1P
82SgHOoCplsmU4xjAlUJ6v0gIHw5IuRCa39SrOlBVaBuarv49Yn8gFGG6MhbQe066ZMY/o/0jeSt
OBe9ejA6zklGHSeT1dVJUSWldLI9r6rx4t1NDnSkPP09gCTyQv1MsanvrZoVaFj0eG4RM2zpfCuk
UtPNHzrz6Ou1q3KKJAunqPs6txS7zr7HhUG1XAStPyeJzqvJEU4NBURuDZns0u19/Z0wJ+bg5TNQ
KzpcyYEDXL6XcDc1c3usiPAk7SBfbKYv/LKApA6jAQ5SPQf+t6meYYRpY2Am3esppKzRfuuovYUr
ZqaKLte78FJ9fIdCFWUf6Zp/sVC81TZ80qDP0txX7zKLjpCKCXdZG3QBFClbK+TlhUfm/T5Gmvps
DSqGFVTfSzsNLQ6V6BLx2TtJet332R86LgDL1ebOpySK+vXswY4rFOlNLAsKKir4PGaQmzryrjN0
Eeq1bCnD4dhemhBs++ifHynY+3lMQ8Vv1IrFBJJIq8uNNw4njyjwXmFcBrwsCvUVRPfq7ogiQ09h
4zyyu2GHKkSAJzxTWufaapxFrCsLwfcJeXrMNDap9rZoT5mZT4sWVLvfvNfvUsQS+CQxZoAwhfP9
m/qojh9O5vCu7ort6HFD7huWNFBFJL9PVAO+ANEN770KJjni8lkvk8Mi9vmGgB+ExFt1mXGuWynf
KsTNwgCIdnAtodrwZkARIwpgGLm08b9kFjm8+3L3IDFWC/90Id1lRRBJdJ/3sB2OTh2Ixqxiw5vh
O5b3/iqbsAbuSRcng2qcWien/fRXjI6gAyG6YIo5fbCqceNsV5lu4e8jsDmurqeCE6DLIFcp4dbP
PQmyK4KSdptC7a7qyfBM1URvpNjOeL+jnDZgiirEXssKvzWzJ/rKmTI3YUvd/H+D250Dde6kmP6x
YUObvNg/5iUUb9H9naoadwlQ2Ps2xo6xAxagPNd9DNGLANycmGO8qRerF69ADvXWXTr1DDyz+YKD
Fd19Thoi01XNQF6sypF17G8DYf1kGx4kwFciF5Y1g2/cJ9uG4k8haYunkrP9Q/kkMVau1nDjl4xW
A7O1GE1c2LFQFnvAlsTvrKeD/ubjg5Lu4as5qrgjtUA0VxMeMUSmFL1DzxzP7su8Pnu+y9QuWImW
+v+oDjEdCF8b2PYjBtdqBCJoi7UL3m5Uu/x0KxaBbEM7rygnoRCdhluKBBx8ObPSmTNJD07TdZL+
4PzNXALn9VljweitwrB2fJUkMwgpUqflMCXTLKGCVEye2V03D/KumyMGQlm1eaQRSU9U4r4+Ne0C
1Oaa0js6DNJHOletnSutDSLu4LKvoc+EJoBCnD7d/AMJax1xBFeqaNDelBc5LkSF6o4T4qfoIIYY
/5zCBYQCDPVo97l54oAMAuozexvlxEqIR5WpCay33qrPZRphU19CDWft/D12gmOJfgDXkmdFzAf6
bjn7B44D0zBOSJS/5dQ4Hpm1xjRiUICCCoYfrBTsp2EoBxUDPBFYcY36MKAN0OWx//Wbbe0z4Afr
zG2jmHulteXsNO4EvWWi9SGEgNoYFiuL2zj0KXxfZKUCCiqEYwlh5N6uXSIvBOZOniajecvAh5d+
WEJVVYCLBHyPyVWTg9R2TZW6GIMBEYefg9hIUmIgnJMjFmILdoAQQGe1UyXyJbllax7yIpT46fVg
muxUuui/ganB/4nHyxYTt9wKjw+1y7k0/Jgr0QilGEFq57IaRuQVoiRsJhQX2g77BvTsWCgFt1Jf
9zHygV9l6dPmHoYEaEU1sVrNyWkBl4dAiNnrtCUx1K/qEDxgcRICpgzrvgb8LoW//nyB/K9E6DqY
aA6YZVa4q7hwz6oKwuUh5pgxHGG2kU+acW6Oy/aQUAdpn5SeV4UG+T0Wrty0sIXLMy96dHVYd92m
cXbvCiuNI71eN/365pM2iO2b/TxOEALu5qPFydqCqRa7FBN3SN/DgVm+ufkqP7CMZYh+obmBDBKz
pe/QkCuK/3tNRQfS+l6sw9LHy67fGBK21Wxgyu9Thx3NBUmRCgEpXgXQncl4gnesBl/foG3qqst+
KErv55FbtfsCzDtyh1+cvo2tcsAzkzoxpiOXzIUTopToGGGkNM/740A7+nSQ3PwRMtT/aQrI+rTn
aHDDqK3JsYKPI4bLh5/qlDcoonwMAGyrwClyT4Mw/Uj00pq/TvBDhQQqWdudIHdrjM3KVn8XoCeZ
6/urqx9GO7iFE3/l+4zSHYSu01Xou+jhj6ObfV/lIWE1ejvUyI/0+6wmd+G2WjLogUpt6uSV8dqS
wcyWBFu7qzGQkPsD/yxtTE6qmBUh6xVzRZM3OA5UvEimNpP2T75ANbHIOHJWqVrC09t5ZVyiy4Nx
EC1LNYlF5t6FxeBh2nRp959vOJOxOXsVG+fLAZoEc35ZK98NvZ5HPonCVzbK3LluqXW0vnZv+WKa
IJvCFthDTkploclS2MpuerUMxflyxIjT4di1/pPy5th03ohgdNLmOcfvG9i3SYWMjetPMAnytrp2
c2xmL47I1gRc+WeETAh0245NMMixnFKYj53dq4vqlts6juKE5D+X8sgp60a2t1asnkxvtFDDtu1Z
kHSylJx4eeJiAkenQj3C2WlDKRg47sETQ9odO2TrGqJ995osuideeaTdLaL0uOi6c/cAYO9Sy9Nq
/H8IeTzfgNDfVyTp7n60dAZLGN9a3K7CvCUSNWCLm473hCq2hRO7c0CAWRKDCBBpgvRXlz2NY5Z7
ilbU7I0S/sd0mrxmCVTOi53xtLbg/MFFoBMyC0m4SsPgeTtHLO4l1pKz3Jmpoefq/HYGq0tAHVb0
5MxlQD5QH6ULGAmO+Z3WP/Hzo2xSh1d0RMWcMvxo5Nj2knniMI4rCRvlnvG+AWyEfMCMytclFtw+
gStVsfPBsFv4U8NaEkWUkweuiUWAfrR6RkeXrdRhJRM1AawzfuIO7yRQ+VQsRYBfU64kZVLNFqpB
CrsgCjjzhanOT3bQlA701j6tCbeYjjKIix72Tbh4zisKYqELRSFRCJ4q7RTKxsW3TgVvjnLDjrU4
ext81IGrRVQSEyflihiyvs07UwowAC+jhmf7QIPejZBu7V5/dUJ8VsXurrmQkWj6qe6DZOZv17nw
UQPZoTIzPz/pC3ha87/sOnFymMRNn9uB7kvsBa6JoUYzvepXp8grfvrwcNRvWYimVR8SuoFn1pRY
2Dq/S2UPuCSI06IAvVtDShW/0xNcoGhUadR/dUImiP5O0hMCjtVjurWjsUT2ZM1Z7thG116Y9lZC
DnYK7PZtCeTexwAXbrlH+2CsVmgu0Kxs47vPjfSksayc5HNHfLk9yzAIfgcwrdZfKYCVOQOyKbD3
B5bSV8EUR8cMrm9Y2Dc1caXKtAtEynNGbyDe457pgyboTVY1nDjm2mqti3HaRzP0GogBo7Pvf9eU
tApeePzgkJsrSH/LnDJyrI8TJMOgt9rCTAXDv2egZdkPgLnmXASjtK7CJe/nJGClAfj7myUgTjHL
viwl44w/4vfIN4tShhUZCh992lyZPnkBOqlfwD0oQdL+wCIXPfxy4/1YeSBKpZwRELysdXq6DafG
eKcOaEtek+7zt2W44d1HyFJDdJ9LKqoWtRR3t9X87E6f7teWghVWitJtRhb8X+S42NKfA4K0OXaL
HsIUOCPkSyomXgFafTfZuUGpAZlCxdb1QYPaD2HckWMeleCO6dKvpECrT4oosU6qfUEb6Xfq2JSc
eZ5V6oosc9UK3IdLGAUUUY9aFq+rnLGdM6M4iiKJ9OyKYBldR4AADOZqtQaqKmzT2OAa9K3FcLHK
bpB06MfsrHar+BUyFARs7zJzl2BHY+o9BK5iuV5AA2cOEGMBamikfpFPJJcL
`protect end_protected




`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
oYYUZ0MeKqJUJoI7DJiuvSB+q5Ix+Iwj9N3EwG3d9aznfrZuw1+Fc2PVy4cVNiksbh9EhD023m7N
/1rZI7UBsA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BmgMGlUziZwp4Aeom40PM0gFb+Lk4HIg7NJ8Ke6/iR/nzJgqwxvBOYZHlsOO/Hp8XOgAeNb9Zd4o
mPFcvStSgKrLqxBJrTC4jOtTOOUVOGECik9X7RElVDiKeZuCTuuYfKks1rnTANMNKsXOPeJj6Svr
YyXA9D2NRP6YkUNuPRY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1jtnTjcMZBAylJ3gewlkrSdkM4rrC/SF7w+2Gpl8C9SK/D8Tzq+D0qrZVMnmX2MWMKbqqYu6bkIj
sy7Xox+kttnLUyhBRsrBNs6gr3T0xsxsJ7Gnyco/P3Bde80gstdJ+PNfjg9uJOXa0R4ym9WtfNGf
swawtPDRNO3XB4oPqX/YBORxc12Z2+Xzlc5kJQDf1WM1UoKUm0j7+JBzjmig2WrmokL853BM29jT
4Ht91JL1B2bOy9A+fEpZnVLxL5NzuQ9svrSJluHfL94vaMxePXlPq6InH4B+XQp0TAFlIitjElNz
4mBAF7U6zb9GPz8ite7f9+Ofg2sCbTc7qhRaHA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gQeqr96ZiBT2MmGHCpbhB9Ma/ONapmaS0FJH16GFlg7E/VRDUjqbqiiC9oovpVsOBnNDQZNmXNgv
dI/YoLxA/mPd3NXizDTj33SvvwJdHC+sPFJrC6pT5rNUHqY3WkLW4EktYj3xtwACazlM0R3H+N1W
ZL2jtTv4hCIZZw83DISHIwGMevxP0unAXWFpAlJTyOmzC5wsjnlwvjA6I18++KC1ECVIFCC+grSL
XEAA1xdZCU131f12m2UaGi1yGaQH3scoEe37TXsoGUkWCMAn3jD7PddNt1X5zhoSRxPsOfUDmtSO
kCNVtrnPznMY8kVS/SdMToJlnwH2sKbHJZ6YoQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aYbz66wynlNa4RYsWnE11uoqAUkMOGD1rK3oC0qHnHAmOdMhPdz4cV/CAQENwbN3ryQY7/k4qEBR
2l3bOqYxA0+CBRl+jt8CXXxWU8WE2qwf32lPVes4/pVAbKANmE02/Ysj4IR7MGLvUvtr934XOsBK
cCc/KqvEbWgnnzkEdl16nzyz9Je6iY7Ni836+/z9BA/OYPszoNI5lKgO/06ni9esrcL9aCuvKXjM
Vplsu70i86fjOGURYjM2YFmCk8Xng1M6ROF+0KD+TufNMvK1W5if6MPJr/BsB83OF/hzcDKyULpB
p2+Eliq8StuhC0n7jUXEo6ZGATEY2a8DWEYVhQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
B8e2xR5DNyjb6SEEOPCOnfB9/yUC8O8izWpzVz5s4/hfcHkvr1SHS13gqMQDj1DN3uSpaoGxcSIv
a3uLHDL4nIDztAAEPOvl5rp/eCLKhGUauWJKGzgIaInIPCBXw0hsptiyzlIicQEO3rsxoS+LR4e9
ltN4asLfvR5i5+Aru5E=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o08P3wLx4KXr1Q02DiaLH2vPxf0H1jXIwF3rbwsiMxYgYGWIJGF4/mxUFC7J/WeIjcsQFoTUns3o
ZlNZWWRR36HJ1r2GmZoMunV8HAWjNjCUrk6RBWvB/4dYllizQVzRhb+3YUjmiSEMr4rkGsWsR9/t
W+i6luLQskwMDbMnn7puINFUehSDaOzDytgvFigNs9cj7haJi7XjPeMPUBa/JbbTJGFnxz8xzl03
55+BSHF5m9JHUn2eN7uDkExSgYolpcYI1EQnoCH8U6Zfcweg7A+n5SfklkTKUeWInYHoz9tHbIHA
y9aJwNoT7f6uxEt4GVf7oKjEfFlxUe/yajXHuw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 132672)
`protect data_block
rvmvtIUYJGgsJuXvSwzCskoYqheZhuUdadvYWJRjo3wwSEV475aeGau/5GdEhAki224BmMZO84qr
yW39LtmFODfPaA/pfxVq2MNlJk8Z8Uge9MMCDDWipLrc2//jysQzSt849mMKf1YJ6SKVFPRIltZ3
9CCXRMtrodg2tfHcuIxA3VX4MefAdlNfqjqAII315trU/dSWfFPVLsbxYAigpgBkMgxWaasv/Z3W
p8QPdV0r8ql8jtbWafzQTteWU0fxCPF3KyN4QUkOgU07BK1Wi+7iLwxgRtVvSL3ZsM24Dm7zB5mz
fBxqovjMflpQE4ufmTqG3jDuCNOcIbuy3TgIMRybgt756qH+pXC+6AMH6DY0uAa7EE7qAhNkmqxj
MKjRDQtmeTADOxO0oYInY13+tmxPBCx0Pvym+JNltHYfG5ddmr7QaXBEw02xyyQxxVI9JoHMLg+/
6uB5XkC3cD/9TUNJjNU+Fz7iqi4igBwL0/e4eicBD2rh77KNHxdMZkI2WNryY9WuniZ+m6uW6NaN
AyalqXgmzUSHX8nAMFS1dEWkagDEhXAHeEsNADlSINupKCoVgFUwSTd5TVl9kqALzD1OqXVdW2Df
uGMwPjVuGigpHMe8DegtQ/TOToviU1ubK33OVkl/1wS93EEX3Vq+v6vVvrKbenswXP9otAqu/Tbn
mEeMQUNwW/gMUG4vwvcd8KrGozCqFRAmAq6z/iZQk72mI6flwmLzneZjSDoUwEa/kRFSKwle1oO4
haELh9Vwc61stjPcPh1j0qe0B2tIHIeV5zZlWf2O63WuwJeL9AOmqOgmnAqRKk9bha/bjBBZR9u9
3VyPNbS7xwpi+qe6n4ceUxkMlz/W6KdYWGKYw2Grvp/snJ7iV8q6OabHP0bLGV9p7FDyle93PI6P
xS9H7UQUyR2rgQY58ZTrnvUpLXr652l4TGABmP8AfFCktD1LocZTF/1ZHXckEJfKtoOgorpVwgl6
BHwHalooUB2XspITJHLAA7qHyfo6p1Ijd8gu+X1y3BTAhrwmcVcevJN9TYt3UytkEYa1w9isBU7r
zwy06TzcmVDcsTsbPDOWq6+xos+W3qgKEYj/01kaZDiOT4vZPkQXInep1RQLn1uoO9G7YS/WapYy
zpYmqO/sx/dfdVDFkiB9R/mrBYq7WH4VGb614oZRXmpL4SH+/f1kLSpPDpYESXIEBsn1/dROHLDm
Xgm3/MaZDSjkCsbczUe7MSCHAIqsJGjeBx4mjx7v59df6kQp8gU7zfL8dNFG6MZb8ve2pSPuxfkl
KceWCt6UN4WuirSv1Euen1PlyoS7qXuwGfIxkSnEB3fYsVwVmrEiyO47E2vv+eMPwUp9z1pD/AZd
xz+pL9quNRvztyLOTvCbCAepOxkHRN+kYjNKjQPH3cvIOCQxFupIy1BLdxhyVVj9Cg5bZEtVJG0g
t83WFSRcIF9WVSFfIx0XGEGDzBa4alKn6BmwVc4UUMmf7PcUfb9IA1DRuuDzodlPJJqfjHCpzb/B
ghK3F6snKBg/67lw2tWiTkqJYAPkw3manXPTZt7Zc9NukXMj9spA67QAev2TTaThqHu4Ri80u2dw
zP5ihBQf26vi7wWukwnIWfHQHSR4u6NsAeKg5bTLn6FL8p7n3dILIkxuIeP35/93f4Q0YUHRNHIH
Cs0feSAD/Yicfop0oEYirLkpV1oLsrMhnh/P0MuyyeGMCxKPygj4ra69Ymo5YEPDB1k4Mt1a1k07
Fc00OgWSPkHMsu5kEFl1yWvv+R48dBS6MsJb1MOIenC/kMwQJvuuIXUl5H1E8I2S7UySqlP/Mf7P
C2E2BNPUY+xQWlQ4d/wGgS+uSRPlwYK62sc9icRj8toX2FOaWzHxuYTYh1SfrF6tObHYRCT709pV
OfFYXzSB7BPfwYXP4a+t5uE203rtOODzTyilaA/klwRulfFjkC89QsW4uCYbcS1DxsvCTRtbIm1x
aWGdwqGCGAleYldkuhcAiLiXPxSc9/Kl/BOG7DWOWa+46cZv+FQGOi4v2UvfWOo5Q9jRlihlPXYh
kKkShQzj393zURHiFS2iZMOiysbP7+Ohpg9QPzVH3VorNUCKks0Nnqff5c0ckWF2ESuoP14QEmVk
qva3SIPgqyAXlYzfFGPhGWKKa/qODDXh6QEIYY77ZGyHf9oj9IcTRZf91QvzoMZXwrds2o335Kiu
UhMKzTnTKdo0TDuZRMTH3LRu4iUJJGu/CoNQrEZgdEQH3PrIyQ8bilPicfXtnyvM0BhLmPZTUSQd
+kpK8tBMC0EDyRmZokZnaS3bJg+CD9VcZaWatIOalI9Pn5wJLpjcs9arzNCKfQGWTxK0e3yfF1w3
jZZsIjshaJ09Q1wcbkzBzPlwUpFXVC9N3GAOXSS3mT67023eb5qAVc4ScCxF0XmelBmPfDs/Mma2
FkO06hdBERRglaw9G77WhHiOmz0N1jBoEChCnmvx534iBVQl0onJ/F8iGQmoCA2rOnl+PbE8Dg+G
veCJO8gzNyCCmc9kuRHzCxfMu9ZUBu+Te9XeXjAVbvZC5VNVuiY0fmLHXfU16muISZBgNGhor/Q0
fBim4t6wPPi6020zA4rT3TA4jHWujdimzrF+3wfD5Q/+LbKpaiM3pUF4E7tm6FkwBtZlB6bKo1JK
KwhJCRyW/FlrM2fl6pvcMvcoV2yUo01Pa4iX+XZtmBOzKfKQANCxYJdyqQFAQj52CcX+iFOLeKWR
FzgrqZsAL0RwaeK1j6C+rYYX81ltsxbY3pLeKT8aJ9n19isLcaTYxDjPgVQXx6YUjN3/PjizMe2Q
xtHoHygZLm40cj4uwu4DBdyIJksNliLmq+faDmMzKr1X1GPQNlhbhS/iajQ9VRbeEb2mjh2U4aiC
zgkf+gKWg/4/LdxWRPxL5Vj7UWoNKc0LgIVYz3QdMansE5yNvjjlZotE0YJVlrz3jrQq0eZg78hk
5M3A0rjY4EATPqfhU1BuRO7n2TJQ3y3ZRYYjlEvO59eGj3o1kP0VjQbKm4e1yDeKRPAQywmZXNuZ
zUzKUGmVpu1KiUOkd+xh/JVjeXepASTloas6S8AHN+p9GMg2QN+UCogaGITAluBmIH7G4WdLXUH2
lezRdQRuu7szWNTUmOdrZcGru/HKuqfzZDaVrVO6IV3Qjd4Aa5Hffg8oSF670Oy0RibteiHvautb
kOVxRV0Jbvb/eHNyNLDhWmpiNHRY4a/EadadKguOcddtYeybg1ajKo2Y1Fy1vRTfb7BaSn1AnE0Z
RLAfAtn1fkif/W17SF1NZDC3xWB/GfO4V0IroWSjiV7vgc3Q7SC1FemstTezw1LQovCzocFbkMsL
8qtTH4raGhv8+iJhHOlwZz/YY7WVJ1AAWde5+nDkokjUH2bEyGu1EkdbmuDVM1Og0uUF/GC9H/Dq
kFZxQRBzonE6tDzhcOqGgDkZpD+sYY+IZ7xIloNJboUCrxvUrXyDBjqhX36wxw/aEzHT4tDH6B8J
iQz0EpnRB+kVWgTb8F1D+etygXE3t0TIL+ouHiYeozPkhVzM7RvWXujNv9dPewCdvOmGjfXqDDvq
Q+xM0qsYF5EQXpEpl2rMIe5MpZH19d6jslzEGNm1lTeA/1erpAFOL3z+5tw6/6D6HgUlPeTKz0my
Kz9daO4DUTgxmK/Oxc/h16H0UXm0ebwVpPeaUpinr63tihMRPso5SPO25T6j7cZT3oLCkQxT+bvB
FXgZuhwyP6wui5mpf/w8buu1EOKoQJWOC6jjlVTwKjhc4ShCGYeDKDrK0ZXum4nqGYWUj7gSmkTp
hUm1mNKqh5Y7c3xTkHKh5M7lWDJiZT811LsmNiS+ckjqqKnboc6L/QsXMshd+vGFzKcmK2nP7gNm
vu6pxzK8B8INPGJKnlamPrZwy/+0jW2XUlsJPAACrjh5MjmT6jihGCKArQXKaWfDNr6wHauA/vfL
l5QDhbuwrDqtzww0TT/l9uTwWoQpzoqHZciEp7WBjY2gBh93zwSJckGHs+M15y/9dlHrPZzbFe38
/pnqmMkPfH04IhGkiaRCoDjaKAUZ6Tqc6gzqkafSu/jT2bNsmesaS0Ae+iHgoOLhbYdaz9t+DQoa
Z6dsA81Kb7RQIdtwfAmipGzMfl+4de7DqEPFY33rYJ0WtsedC/zpsIzUm+w/UqO0iZbNAiYcWlpj
idz+4MBNcLYmkL62hwuXL0j66RGp1f+rZo3KlfpyVT/kyo+NRTTAaBBn2Or40ELEOP2rrDIo+nyY
3dWJIwPyfO2HgHCOb96bR3w+nGAG25gFtMRaeGGLwJhSTIqPIqevOlOSKH00dUuxgUfrAy+1lU1T
nlRBmQNjbPFPmGiz8E3VDX70fPpRvw/utfBVTsHzaylhXe9JqBKVci0VuuPOiBcJCQnC7OIaphKw
zTD0JCovbMba8F9Yo/dBX0PmAoyEsttTvC5kzFwv/uCoyaxbL3V6dHA2bKBnefXfJYld4LVWf66y
cjjjCLXC1JqasimgcUBaeh32oTbEyeLn3y0BohSSr7k6c65s0zUzgeWm7qNrQu3vNvG7WPX9s2JV
G/X32mNkSsR99xrO6UgNBmb+nT/htE7oiqdsgFvydRWQDqHi8dd9C8JPu82/veBkcWwwwYkuAtJS
56SKrh/W1MgCojY5rUR4L6OZ8FYpHMJ0rRaB9sQxzr0n6l2dgnh5ypf0aasSmSUZwVpErYduQ8k7
VKEvY3iMFUI3+H9v6sncrXVniOKcvMrfI5ln0gMFOerW4Gv4IVFqU5jcdDLxwLTFJtuINOeukk1w
hdxJ35lxrf3Q8paCGFVD0D1phq9DZL69EWekDbuDTo82AWh+HXzJZpRSzr73YjLWvRGctRQFU13Y
ynKS67LXQLK1CkQUFDSjpaH3lFOpBBpbeFHWcO4nygZ68XUzLdhRLn1ty/0TSmWzJNi3lO82SERI
vMdjCB941REImWBKID2J04bbtkOWuAE5qi3SedjHAD7i49GRCGS3lLPkuoDnOXziYNVX8miX46pr
MMaUZTMk02m9qZDWDPReVnvsE3sy8ySO5nHdZt2I1dU/g1gLJ5djv2GBYiE5X/uNDi95BkCnJ7aH
ywBJgg2R844mMgteDDY2aETthPQaFwmxguutjN+f5c5CKCBj8AheOoIRwG+kPo6hFgLGBYziZzqn
okFS9PziCEdzDgaRgrEqxXEnWWgZiceqCVcHSZHkX67phwiPDG0pc/EdJg7uTMNmXw7IsBZr38+6
AxhOAGSjQ0lkziFkv3/Dz/cDnuMCPnXscpOr8fX43rGV7hD5F6WwD9ZM4KFyyEmya4jcf9AbTNa7
KMjb4Lm9Outcd3m1XA+pyINBBjlhzLQY5B7EnrwTFo0ExZxTEuhipoC1gxbp78SaGA+4hLaaT7LD
tpYn5GOAOEFOUU1d+VJJ3Rn6JgPN03F7/1XeP8Ls1j0BjJprYosHhRedYj2i7097D/D36fq9Pu7p
fepGc/t1LGqh9sH133oGbOCRQpxfHPrLnn43ybzIBkc/fBHUIlo7U6+li+o3Knp+OIILaOtxxJ7Q
zF8dla2Bu4hVyyQBGjajCK8G7DmBvUvF3GUWwHEuQFOJ19K8mW+PQszFMyCuTCHg81P3kx2wF1q1
qiCBrK+wCMh54FmH5LEfN8JVqajTSsVbZ0JqAne8bcLg9a6x/JxGvHgs+bjtWRCWKrg33YdNreRp
dkHsrZdQodT9ibUmf7PkoA/F8dWOSJIrI589Sb41fdjt/rztx5OLXA+ELN8f4iJjrDwKxcj1R0WP
EUpg/YhJKlH0NZTryRmUP58Gyul/60hVrJmmmXlh6mjmaqjmyaAEeJf0T1FSszKZhdzqqZGzyK3p
hqST/dYiRnbbeOOCzJBhFz2wn5menXyAq5rXNfBc+gPaMh7lQ7TXqiw1ct/9QwurzbpSntwU36vb
0JVkbJjOUH8tZnXPt2zTs1HGixkX8MfBF0qZt92uC8DbtvBqU4zviHZCqpTpKoDUGkbWv1fJoM4X
p7k8m9qFTEQYwiEqAtPP3SE8GO6OzNh8gWmCVi6ikuqAlNmcIUV/Pl6e683GFPqa+cvuGGwMKUMq
cTogmnm2F8EeJrPA4eJu1GHpPIsOMEfsg5ZnrfRn+fSTdUyIFMo6BKebpbjxcs/kxYYaZ7D7fEvV
TuKixA+y2WhKMXxfAu8bryqi70niTPJelAd2DkmV7kOEz3o06hAgcQC93aWQYZ2zoPpf0EelWP7a
q2JeyYyalDRAoSZuH0A7dSHaeobxtqPRxm3ORD5QiqE2Cg7yUwv+GzA8m5TyOLtxxdJh6zrX2qGf
hYew0i7uNMJLjaxJfkWV7fbdVROpipSXfjvV2kfffjIUvBWOEgY/AtzZewvCYPICqfPpayO99UeB
WywJGBYy5pH3Lc9VHpnrqvrCTqk8Gevl9Sy9DPmz+W2mjxX9Q2FfO3bA8Msqus/9cLXiKT2/IwTW
MHl8hkvka8SqP4r72CFzBaC7dO75NDOChctDY0yXZXo4sqXGQ/q+NsD46KNHvPYUls5tZhW7Ur4g
x1JI156oULReJkO5zDZZXn6OafCsbeRUNeRHZP+txoOKUu1YkisAAfhwkcSnIGRiWY94RutyPgbl
BVO3VLIW7eGH047KkotPH0ya0SGTvvch/LOrK8/t0xYzURy1XnOuPbgLA36WoCpGDIblQxDKVBrl
JLdzoy1EKBxnJC+VVckmXj2nKGMKxQkPZMybbhtLMhj9LMXuPpf4kwsEiTy/JtNjF2c+qT6b7hrj
SnGkIJP1mH2IvdO8XNGh0jzS7BhrVaepa68Z5jXiXHTVoHWDlN39WbrZZhZ/1hsnc61X0ApZeJJG
8qc3hV64hsOoan8uO+mPzWm1XxxewL3W0jx8zzU091PRmBNnTq+wCZOGpBtj864nHMuI17+hUpop
R9YHi0DhHsS1FBf+c1EO2Lvsz06DGl3UgY8A/Bf7rJ9VVWsDmxcAYKY0qJTMdgLz/RMWgtEjZiZP
Kn37iURmqUP/jCVId09qdVzI5jN2hJf2vnEzW/h1WyZzUGYZbtKXh9oql81p57DvnZxndVSKEdjF
runk2XPcMhyToiFGgN/NIBCZEzBxyezoXRFPVItp+6YXGLHvnLGCXlG6B6zAc6IxuDyoicXAbTLb
las/PkerEfcyo5hu7VtFGIjt7fNJgJKe1MVLR1B8lwP05x1tLPEkfM0sJyHXVgk0QXU+2Ym49wmg
6aSyilfkuluewp3aq9ZoSRMGiZUh0p1O60UwK6rCMMBWN2D49HGNwIF15EBYyn6FnYHnH67k+7Dl
MzgnTdl/ForpoWbPikTGOioGEutnkO+ZzS5j7f829QFsSJ93flZQPQ34M5Vvqasn+KYfP+XUlzIr
4Pt0amRl9h3CUrbzLP78XsLgIJqmMHpX0ilojDJf05Dm96NVcp9vNG67IqjEMfa8Uwc/9tvYnhY4
jE0jRmq95ItnwcjyALpNNsxLPPH6EmNDi8+wz/RWlIpKJBAjt2hSPhItW9Mj0BL599KokyVW9pLs
fy/YRbwQ+lZemK74l2S3cP9qMBUe/xDpo9b9mmLK1N7NDmYE5X2E5mClZLOs4PO5AuH+Xat9ukpN
jK08KszThKoaAjT3nRJBZrk7w7Mq7FtpaHrd+hL5MR7G85sBOm441JrrPsbEEODCnvzqP4t20/wb
P0/p4CTZJuPTzdBjwUdYMhKTAyhoyCVsRQxCC6ArhDSJP485Osr65yzHZqH25Z4cv/QgH05S+/9G
68yBmtzw5hPv66lU2hvr7/yJ/YEU+NT3RDNZMGLMDzXZApRJgvdu/BBUtOdYg2rsGkql86Y4K9ez
zFhBI3PtIcyNcmyzEtXat+vuzLLjUJ6D2mvzRFvs8cfnOo8mRXY4PEVYaIeRHnTB5LYHG2lMDlIJ
Qso/wvtLM/embfgrVOfPco5f6AQkqmlnZ/3fXgfhBwhhBZQX+TcypKvysTv/IWj/nWzwwvCi7lWE
O+JtgluEqTqE5tcv3LhGJO44BTqefL8/KrnKAl6lokrb5YPyROPiViNkuZ8jCJJoN1InBrXeIJ3G
78Sm8SkCyKr1w9srn/9+DHTNp8zM7N7ACzukgr9P8Axlifx/Nwo0kAwseznWxmeTQmFQiqLO9sdF
RG4wM8nxPnELSYShROOX+7GC73SYKtp0QtO+Bk9U1/8i9VrY3GImR/Q+C/ydL47NLO0H8309ehDl
tSMhcRO9i67tOHH4S7X4UabUH+1u8AgwpKpSY2VR0old80C7qTmA4UfU12h3Cmobp18MHYtsG1Wk
1aGjoZzafbr3qkxaXsdRl4L0Cei87QkhExgK/RrlkQD2BphNSMwLbpTQeq8lGYwLS467RNhqjbY7
o0jlzdd4x3D7mn8Dmt4ukRbE0rC6ftIXMAEnMdJze2ba0GfK/6DGfqafjukFo9DhCl6NXIN34qOR
GSPXfynXL9Ig9uj++Mm+OGubrnafyG8u9VKBrmsL53fLeBrbt9Y0/5fURALsTUWnaL/92gecskbj
B7WkjZcweB5tTDo94/rZLDQ6tNfElf5oWOnLyGaNMvory7YiK8L/FdSqJ2bvi0ENmVAteqk3bfPv
3daAGuHW1b1fyGIvhgVmM+OhHq+ooyNgzZYRcxxrJGwB3DkNS/q5BQaqs5TTtHXgZHlNeSt5Xmkd
tav23TSoQerJCn6r8HqImxb+7ZbZrCcnU83BwObcoX+jJKjLko8zq2iE7CbpWWw0NkXuT//zoOIP
bu34xVQN+R/PPHdYbjGBilR5LqSAO8+GYunULLgHyrSdZ/dttfiHD5+zxwki7QjHW6IHRzMWT3vX
G+GmWhVDXMLMzZlNQUIwWNFKuhalqRG6Jw9/DPfwU/hepes7lvL+62mEHXXdpzH/ejkZ107jbkMc
bnfy8lOv2U7DtUjHUIqFb6UxmEn5mimVYmFKu7lXEBqBclM9lf4y8Z6VJO4VHNUBk7KjiZekNmY/
Lp57Lco4bOVyXVfoK8+Mv9ucirB8WrwPPeTnO6OxdSVKvd/uOXzsFR+L4N4XZv0PErsBLSf0Qhsv
GqXWpqa/ou05+9UHod2kOh3C7FHmHieP7hhJgfREzjrCJRrpg1KDMhV6AeAY9GcyUHMvAIV/P4Or
/HBjRp9DXBVVdOkU4G00y2ZlTqOZeml66MbPe+pXZE1QjS13O5W1oWEzFqty1OBlGQrrCu0PExfo
P/M3KTPtUEYkrLep6MV7HQaOzQ6YGLPH1tQrc7ILHayZUINPlyg3BDIz1z2FCrWoB/3QBcazKodQ
HybIEbEFjlU+sO5rsFR+Gu+klgL26RUzsYq22DXmAy93MW7rnorfQ4gZduMdnw5q+TKE3sGHz5Oc
Bk/zBG/zHJNGe/Pe1i+RFV2YWZ6DzmOE4QyImZJCimgfzz7qMzNvv20Hg0kYungUo+J1TFGP0qbg
Wn8cY/QqnMtKBudJXEPs5yHyQM/b224+61DH7RU6qUUyxboda9O1Q3FYQvVeRYMLFa43MmZBVWif
1N5waUaWw3HuqaXBMHSIUHzxco12DkHRzOeB7zjDbfhawMRUiHi38d2Mi9DMw3WDJZsvni1/HM+y
WA8y4V7ZmL0P96rFsd8pQe1oVOGTincfq9p1FwoHrPskyaNMM4n8HdbdpL9y5GFd6jd8/qzI5Dir
slkRFDGlF+fDDEBz+OXxpCnJaEQPD59sdz7S1z6QU83j1mQqrlTkSZpYEpSV9FWNpfMvlICHenI9
/yDDrsvIhzmcb7MWH8T4h9groLUUxN7WgqQEKrO4JBc11rU+jDw70WFc1hhehu0kmwwkGLmbCUoE
etSVzBnn8hS5TAmdTYSCQuZyXV3gEIpTuYN6oz+dHZnql2TSpp2Vxj9EXJVh5sqWxDVSacor+KL/
3V1oUBaBqLPWqW5cCAYBiwyr/bmiESxBCpfdF3TNMwGybZflINThj3WsMVojlj5daQQMtiFZ9zJq
h2kU8YbRmSTKamYW3A4WhrMW1EZC2+nRWCrImcNQB/j53vPeEr0xmHcsauhZ7p9AMrJ2Tj4TwFvK
ji/rk85X8OVHqgCQjQus3i7hlnUuz91FjRcFUxlr4SncBVbzbUNPDPzAXKlOaXd9WW+jExn/5wwn
wBD9jzjokjPCkB7d+SB3VFpP0nRxg6InIHpqVlbUx8Kukj3+b9Mfk2ciZuo7CySaIwGQoSJecb4z
KXgUL8h27eynepZJKgD9ihQLZVZO67MhWNGKECsy60EmgPa9/2/LbdpADQeWzgIn06lGywzv3bTV
/PrZ/9aI/fLGvFrdoI8CEd8/KuGHTT3XsH7ZLDE6rW1DGC18szb0OVdeqdhomBRTcejytEHwJGhL
JAlSpo0ko8Y4QzRVSDdhCGWGwuqz9sBP7cJYZTUYnuBONROifIzgrcBbtIVlYt5jqq83YMKzlNmW
A+3aVNq5Is4K5I08k3KUF1+qwLG90mDhl+Ak7lZRzHjpbZoDByjRSQOSYz200peFyf3ftFZOt3Wk
qukOBPmxAem8Fw7q/LRCgTtfz7YQiI+QSSzKxq4d7zzKQ5N9kYUoManfQNcPvipj53B/V+0p+7Wc
OK4sQ8bi3m5US0DKKX8Y2GVclB13NS03Ck9IcVAh1WOG/Rf/gBl/tpkwBIVqbBbjx+4ZyjpiOdGL
l3aovgq+KritqoQZ0A7YoRCsXiyRw19+OhtJ2SwT5Q4NYhxzBR/WgSQNwNMoM3Hs2nSHy4v97347
EI+Rp4Nechihiru/s4uI2g7/gPsd36nUOOLVss5pUrkNvw9vCobazMNXuTW2JWjWCJ3fFd28E9jz
PW7AyLAnH38VsfAvzlfliHYfRJ+79k9mhpEsC5YHOYjy0BIJBvuftViLP3h926mRQa62Z589qvrp
pdGQ5k9rie3SZhtOqrsYi14rt1E6A6gkBT8HriEl8Gk3tbPDN8HPN4goEDt99NEKnYQt7EsLst7o
dfWHqn8HSz739xRhUct5EWfOtkqoXMSPaMXoKmGwkA5riRSETqDwDPG22gAAU0PI40e2+DR6krCc
llMNhHXM3c+uDYNDdH/VlMgvbmO05DVef9+ldrra90p8BGUTiwaUqxlEM6TZuCfYt47fgTVeonFO
gxzFiYQ4h2UMMryFJMgi2X2eKnRE5rJTAVqOI3RzUcIRWWK823nbaK2MV5+FapoSDdZp9Z8+UYA/
aQizeAkimpjDVqIQlfqcj+g3z32YnWeyciiT9+hCx+vRiYlaL9PkUQz/c01g1W2+Yuow3R09WZgf
WbobP+4Hrku+wpPocuhVJ7CdTel+UfGeVlIxeGfDE0UGTqGWYjumS7DE/PseXmPizr84oQ+l3xS8
twP9G0/YCqJMbT3yjFIH3CPJqHkTzz+Vjtiobr+fEBWSEZgBFPh1G2I4PbohVCOU/Sk/UPjcuKch
qnTqyd8AzghxiEnOE7bF+FAihe1ZtIybhZ2WXmXSlzYnzHVYaX5iSLzmINf+CvYtqIKVGcaYlvP/
uJtWosKdYiaMrFyZvCVPjReLBxuEdgF0N1f5pkHToEaqMk5sQShwrNr1fGrOQ8ruYK5/O+ENHDJj
ykGBTduZoLgG6RdLXryonoePvdWWxWujgDBO4v1E+Qgf+VVTNzNDDlDRIbTeyqZ28hxhkVUsFmg9
tUX0PPZpEhJ9m1DnQn7hLosJap1zX+tg/qdwAH0vVKxA7CCivKZcl9X0oAja7NZdQbkWRoCLQHDr
ac+M5QCzv58EU5U7otit7a8gsBKk6+amUZJCodvBe547o3PFppDKflFazWgxgZR1eDru9mDvfHsJ
bhVbQIlg0XxVnCxzuaCb2PyZap9Q774SdPafOzEUdINqCQYea4osr2Z6mhUT/qWENXtE8xWlWpSt
m0Ol/J7hOWstf9uzVatDaMTzfdMfRUXyWOLBTk1mVtYnegGENuuvHQJQlJ+qj0a8QKGer+4VynkX
X+IeHo9DOWEOW/z/t2DUZt/904j1QsqbdmvWqq6FYIMuZOPE7nhHHY2tgakQ3wvEBZdf34CjXrSt
gUDpZON2QSNi1y6xs1Cs+vEzxYNC9r1t53txewFZs4WYWg9mEWYxU9YkpiJsdU4O2XDYzE9Af5a0
fPmX7PPKnJhJR9FeuLklkuaoQL4RDaOUhP07+wIzYe1yJpomrPGyXdtM3JfX99t2k3FwsnZp0pXo
2tHNTht+dYaiyJSuBQ0olSzmUkDnT6uyMOe1eU2/QvmhwkRjOhJxBar9XMy1PhnqwpbO4fC1rcHB
REVR6XhKgAtCV7hSnudQ5MSpuci3HOXcrXXXhzmfUT3e9tQVW0rTYe8ByEc5dEnv+FraUpZi0hSy
qT4f5XDZRoIzmVWv/tOmJsRwGKdeeoxwGFAkRs8JRzC++MtN6/CpnxOXKN6XpHI9AeZ0uWzQaGyR
Z9VwbaRVx9o5dA9PEhOqg9dmm6gNPQxG1dopWxG8zMApQOhv7gP2SWy/Cw/UQi8O5bUwA66t+TFG
PdJzX9ZM1Ct1ycKmc2vmCKVPmPGX0trqbKKRsLxb3dCkyGhgpurs4a5+GNL+WaCLXGYGLCYenoRs
Cag2Edf4aEVA+s3vzPGej4GIbKf/q4ms9HonkSVxfsZ1pEUgg6XVDHHJxbD6oPMUfilZHnECvcO+
9ZRI9ecsSvUmBtgXgqw0gKmJY2vaw6uhG7LPLTmGDqKJEEq7flB8BqAj+5ErnYzF52Sb+N0CDtlN
HWQFRGwAy/RfRMEta00v9qVXZRm8szjq1BVlrty8I0MyDhLaWXwtFvAg0P3dEXnE3TISX8s/iyjI
4E0ASiBhKU+H0w4aCoerumvHcGXpLOBuHOafgA8zcQrLM7+fK6/xKYT1k//eQ23Bo5LjInaw54CS
g8K+FrWDljG8da4KDoD6meN30VDfwKDA5xJuKb7+miykabgo6zayLGDAd/acKlujPq+yvmfZBkyB
R0T/7EcDWgFrimSL3I6sAEL6IeUAUv0IQDvWjn6+CFOqrmPo7mraL/EtaI27p1Xpyao6VbTpSQdb
NxEZp9owc8E12OTmbsxp11cY75RYghb6Ph15AIRttHmh0q4PypmH6yfKvknLvZHwemu7xvz2gIfI
JSaIVsR+YFHUAMR3d0Zjs6LqRzKT5hhlH9qnLIt0ty+2Gewqun3xz1IQyLrbPX7pxFybdrA2ORN0
cHylk9tLJO22z4VncGxLPJvtHR+kwbD5DnnmLhPyeYlbe5T3jnuWHL4QPDM8chpN+yfiQLodwCx4
03hx4vBwiPjcA9J6wacgoNfKs9Xvcb8jSe0fUco4xDF1P2nmOU2b4Q58wFQyLzWLNuPyCE4zS1jK
r78l2oauJTaQfZg4xB8aPqCUnkCbTosXc2QiDswu48IukYoO0dReA02+ZI0378JA2FjqdGhqnMDN
MLhCyjVA6XF9WyTkmLGFSNRrSEE69FOBXfCB90buZkgld2cjqWQBhHDo62fuESockPBUSVmt0TQn
C3JNpak9e96bke20equ6Q+jqhmKvoq4D2FCUed8ZEjVVXnyVBZolfpYi97kDxP4wDQQhWbOFlvFF
6SCCOqXMkXe9CTamIuksNiTo6hBn7CvOcnuhmO5IWASSnZvP2kyDYO4YXmbRMKdiEklgfHjbgaII
jTvHk3OutsaLVhkqWZI66MMSSIZnbJtP6/AcvWF9NOkmWTYFwvl1FAkcpiIjykx7rnuIROqoBpf4
T7gBJECnBbjWt/btMU87fLTAJu90U77ubkuyoB3W9c/VeNYXqvgZlA66LOmXyzDDA8/2tZ2dLPE+
8QsycnS0+vQpDpif9hOJqmTfk9uwJos/qqR0BxrJS7oDyp97iM/WF2YHOA2EPSqJVwzHj5VP7EFz
cN3Nsx1a6JJyrdXEuhFQWH9G70Bv0xJnS9XqORm8heyFmUZ3gMNL40DjBM4fPTbGSwSgmzhvRrYH
c6sIOIIqyx4bYZaRjiDKrV/qShyXpwJl2NZ+hMHtcMejdySVYKNugUzXSTMZxqOLyjVzxv6FAVQR
zqyoqf9HSAyc13m2nlzU5CE+281Hw8DgUZrmcvj1lwSAtSgO1U76iXDPoXWPSwReNLLMsKrhB01v
5E+OzFL8923d49eLMF7Ox4CDbftA3qf6Y4sC1h+RUmfWJCoAdimQcdOp+/4HMyUe7VkzVJfl4qoZ
7BpOoISu1XX0r8GiEyvkRf57wxBbWgPzFPUpGHhZ4W/1I+s/51gcdk4YULWHJivm/jpiFUT796l8
tBNsGxH7xcgAEm8hw4sZB7/xVfutMGz8+K2hxjS5fd5fPZNQVEY+3hptU9MOkqNuUUXeTq7720Lx
VpkKM2IFJhxCnIHAR0GPNLPtGPjKL2x+h1ETzAvLIF0AzYhlyBWOq4wsJTc8v+OOfi5RUPRhJVsv
9xUfExbQhW2cthmpdFkuCGx/C907HXUQ+2HIvgK9SfB8b1tki29oBR16xivoQsdcjfwAwp4QFMPL
N9oC8kTfpvCq8fx2AXU3gfg2Ru5BSq1s8wI2cS4Aijcx91HQLarfMHgihTENGnCyTfpji54IeBfm
NIKHP2COFmjV3Dus+DOiB/UJ8+g7cfqeY9heOjBZbS9aKXiKAf9k9J/HqpDnwqCZXfStJYdgdKVu
cKx5CjW7z1HU0WxHjcXoXTUR/ACRsukvE/9aByIbbvlMYvGyFrnHBYDsN1dtL5oHA3We8Hnhpw0d
j34CAfkK1GtjuHd864G1vfI8CqFWtZO1e8mxDIs7mc0hjkAvlsGsAtaHlXIpwLWOJSaUZuB1tGma
2+hsroukt21zQm7foxfcCQgquPCiCpwkjkONZ0ORRsG5imRj3peSO530ZaAsmZdXxAndFD3PRSYN
3lP6nvwUp/tO+s3iX88I7sdobwQkj1a30OTcz42L3xfeestbCw4bBQHaJL1Zb3Q2l65y9XWMDld0
gGO2+jMtaN3h6gmTAWN/vbSxnyi1ZK7Fnsg2B1CgzynZWyhwBAofhZa3UH7v4/eUuWnQKEUOJAao
dBMfE8v2k2rN1RyQtuiuOKfApfd1blA7/jdSM4oITLe0ah+vjqUxu6n4tlbvTBi7sPLpZQ/4jcJO
a5FjZSzzbgA7FgxldwSVX5/WphdQsuP7pCRzZ7f5KhUkkbouwsZaBuxd4EMAXRKj71IWYGam8SB1
8vLWh3P6F0hl1JdqLNKCaAuNS2H1Un2adbRorOEYT7QciJGBObWEPRCjHfaLgHYKASy7TEgQRsGv
MAjB6eMQRawjG8h8BaIw24pdJexCiWkeRX72IbUuIY7/+tcF86LJdpyeGCQp7QJRULO8hO11ZbYQ
KjrL/n3i9A17UjS6JHT7BN8akmyDH/71jIBNaqR5DY94zxxm8BgurZ7qH0FjKTota1ZgYi1Lq85L
t5kIBHlvk7SO8n/k4d9Wg3g0WmBq22n1Dd94fgALPzFd/x/HIMvSEQTqUb1az3y/NBlE2YeoxTih
tn19hfdsC5TIW719W1vPSWwgbg6C4/J9UGnPmvD1MoFk8ZFD4NFS2ujr7bWXwRFH2vN8duSuyVgw
d9pyP4RDy3EGpFL4WBvhQxfiVr1KsN6bGHghNfRHGUnXNlluCIziqMgdTMFDIydzlycXgj4ne2c9
gffoPYY7NEdGVidMWrW9e3T7TDnRlnE735Rr/hWcHW53X2lvjU1FxT7yn1MsYu/nwtgL3pZF9utR
h/vlcPmQB/4mTMFmb00mjY9oTcVXMiNgqLWEcWyCkrcltIFiAHLgEodjcZYclX/GEz0+D1t43PAz
QQrhefMrTGZbdIoB5Koo7/8N406sEHSGAsl+vg8aPbVVB/i+/x4nmEnwSskacu/VwI/v720yi0dj
szThRVh9D5kzQLA3kK8K8ITTpZByUjD7K6lpV+xnrOwpgsBb946OA0VEcjAuL72akMC8Y/SPKdIB
D8rDaOTb2RmfIgATgJdlxeaiQ7Hb/PWrmH3CN+e87k3O2DQ5TqcLaa3T3Q0r6NunnYiG4TP9ngd8
V9h3zu4wXsgcHhgOj/Svmww9CdkmWuEcW1Op/di4C09rBOl3FLeb7OwWEZGWWZ8LR17ERhI1cEgm
awL6YCgzfvXomzZ4fc/4zKqp8x/r7Vf2CIGrWruGXVORWdZlY3VK7mwZ+gKG2ZmgR6ZWdz/GzdHg
U3lVWtPzANyIE0RQBkYqxO/8vErQVgmEdjOUsmI/tHO+mNnNlgB5GOuRZB1sWVRtRtZbjVGybV1z
J+x63o+pMz0o7zcPnmgnyzL2yQDFBxVynPsOiqil8W38kkT3A8zf1l8S6FuHZucE0wR14m4EAFy4
rzzlqWKoNj6F25q6PvwcmxNEc1bUvWEF5UB9kENOrkQgW/29ecTdil5bKjD2PLpOFd8bbjCQXlwM
ykJX4qrs3vuuRw2S+2Dc3v2das/4D050uKEWUexT2nTP2covzcA2kHv+gtPx3pdayuridx1nO2zB
hBlfWMFAepJFfLiqxUQm1PkkZbDckppCQ44XZmaVyFRTLbaKLxod/R4zCAvkr4VisOKe0YfKNzvO
3q+DBy+y4uSXX14L4lvIktpV26RMRvzQ8M7WxihoHocpVZMhfDtZwtqDepfTyhaWK5oEKDbEDsi3
hAU4GDMx3/nuKh3R3E51r28SrxlZq9ZaEx/OKM50VUKulnLroWlx5AZdfh4Gc3twOxlocIiQDcO2
FGYHXaszVIs+RQIiugq3rbO4/fnTKevzLuZ7JrepPEGpD0TUKebVRyTX6dhjQES+Vxwf9CzScAlD
GdAIg31JWgr9fi2xnWbXOFIjpTAYjiFCw7zmRI4kg96bz3O7YT4wZKrDSIfT90HEc3ikMoQwqKn+
54dAiLmj3XdB5KqTvKZiUaLu43TjWwi32VbOLpatsJ2jpbMYy262Qpgqh66ubizN2Dj2bHC5h3v0
pFyk/FqXrvgVHyZZ9XicvI3dVkcbONcmU20pT44lW7OWmijjKUyjw3VfCe5fUUgxuAnHhLvjlBwa
BVmq7SOvRMaIv5Q5dMMhe+l1d5SXV/u0JnzxFOOtcqsJzRPBzd9JNgznvxgK0jxckQE6WpQuNV5/
3NCAnYIXsbAnsaItQ53r4IC+kzKv4fR/NZeVyArxy1PrmGePcSAGoQjbjtDyLiXX0oV9NuuuI8fm
XhhnesRFWEL+8VaD1ZuOZta8mjUbWuUP8uqmZTdi+k2f2aw/YOieqFp0vvQV6ODpdmsZt76q9sR1
3OxOTyqbFQOCdqh5LLUGVkIKdMmtGZVuu1PpR0UEO185lTRXjRoG5m2dOK4kc4zNnS3OwzipOWqh
jlZMgOI1VbAEDOaOwowSdeOR51QGep56MY6zVBcHxoB3+tKMKfpeYS2Q2q66/kIBu/4+XXnvD1U/
UsMBsw2RgDAb8kBryzt0h8L9dKfjYEJcSuaCNPEC+g+zo0OuZhDs3/pYTBeOdERC2Tiu7s5bdy/N
Pp6BkJLH7qq69osyZlL33LNY2eEy8zv4aHTlyOo9BuTp+D7+y277pV2N1eUWnPhv6GxSHDpSOFXd
CpZ8L0ujB4Sm20xb/5anlg9XCVqu9MXitpUuypZ1E8OhsLBHx4U4dueaPSgvfzuzNOZKDI0r+DxQ
D54K7SGxctukIQBXEp/M0gt1rHEDy7mMhcSj5YpTtru7mgzZL5xyPUKqOQGji7ImrRQcrWbK7ES/
SQVcfEmYJT7Dn40R9HQZXpfdWmB8qv6soTH2he1JIX1EIPApquVoafBygfA7oHEu+J1UIuvIBfVw
Txy3rP7wbzyV6WAyuM61gAKgOckcwW23tGu5CUBjd2rk5+lUhDKbuR4dm8dHWELt0DgI4zYNOwTj
HSzhRr+wzf7JqEgYzy7Vu21koonCZzvHqQfXwAovsHAYLcdVbqM6L54DrJIeMAxcBTMqcTImFLOz
O2POwNF+ISxAmjANNcmd+/WdtBmL9bk9M99S4UJUBT+04P380mgekZv8ych3ZmpNmzZcYZwGwkqG
g/d0F8JDhnrrhxpyEIMFqrELB8jlsGiJX5gFUGcAxcrOclu06NsMQJ8+jLSla3PfE6VnzA3kmu6E
ZKJ/DOzcLYfNznufoCtlsb+BKAd3inoPOEKCmzGy9kfhu0GBg4h5cOp5otSpxXZmv2NVbH74Le6I
22xA5GwsPkNmJPy7KEnZn5/QQvP4DsbDx0wMrHcbJuc/zm+WeZsV6Ps+nDUHesMN7tuJVSvCy0ia
GrCIWm+qMWabDSznDQWq8jzkGvPFc6ar3wzHktxf5wHmSmiWZI4gn0jkwCCzVbmY/s5Q1xPt7yFT
Z1KTnwhhjVC2/isOfjLDv/08UHcsuUY1jhMhbL10OQKg5wphR+/N+gM2TUzxrcSDlBOED3yARlkc
qmD+9QQ19vR2DfrqIHcuiH4xFulTaMfedbrTUERDOguBeReOfp7W23epiY4+aH5YokfOlpBXwY3O
HMDMdZqz6jlEuxsvgskyAf3xXS82pC9KTMBlXd9dHwxvlSpN5o1EAbspM20r2hbCkV4OQLltVZaT
rTgPFlOlixc1CidjdQVLX8+czstUY3R0Y/OOMam+8OzNDo6GTRBDMI23i30GVUyk961rr6Jk53zW
PjDE+7fyimGDgVmPcE1608nc/8jYnOtEDjqJRudDQuswxQTBrL/NOOUF1SIVrefnb8bTsjdlZJKe
FPJL3ENfc34geKQZJ3hJVZoTVJrD2eNzTGmYYf2Uz64S2z5l12iJs9rEZjvD6muiv7B75r3tNxAv
wu2AWd2cHixeYvkgMN3Ut1K75+3SiTJ87UTJDr4FP4R2CpMlzuDU8wTO21zxXJ2XbVNJZkpe99Uo
jGRn5Tt3BA4soELu7NMebU+LvEqISr58FD7lUOFBn90VKaUDUG2GmN9RiY/9rmIj1fTRLxqFHY58
PIQEL2fRsrVKwLyv26cs1HMhM+3MSqG6AuNDHfJGjs4IgUDsd9jjGkMpKix822Pu45aUdv74PW8K
GdiMrQK4mfCEsgXd9++0uENr01377vkkAY/aiSO5xRlPgJj9WIbldYVdLIgtsz+saS8CbIzdOgLR
4Er31VOmTBhTCp6zhM/E3M6TMBs4aB4bxzF3AKkIBqqerWEL3ENqTV5tacxOZHNtg6u64uXmIiII
v1hgo+C7yYTZ/1nplUuNkRr4cJ3r4gHMixB4IQ+pqcriF60wTd9jFsNszZNEc8hDG4URQjOgWQb1
t1KoY/YsDCby/zZ1HQgPXRmlV2SpogX5AB67AyiEOy7CQ7gbMw/zTcHJGqQH6+NSjAgcKtdgfTJo
cUED/paCZYxzQIPKJDlejTnDRlQmONRHUkM+RAMyeBsfqaHe7jdNLpAWc32SE1FI2wajV5ysrsR5
MYjEu/owzVSYq737+XtylNEwmrtUK1yFsnfxx/W5OIdcIFO9AdJzVy1cggU9lffZ2GJQrayMBkjM
s+WRvtkB0iq/s8s0G3uDeEH77+wQnvJ1QB2zzcLWdFSgSvKtcwKKA4XJD1ltAgNS5/29rQTiXIV4
h/mrZkMItqi8czvzRCak2ACRcxRjAtWCZkvSsFN1flnDeC0pET/wlJ47yS/KCOeXn7JL0UAmISd9
bGE+CLh45bUZeYkS2FgnOgl+N2wS2Wunu+FMXLM6daiwn35U2LNs9L5LEGGRc/PaeCbj2EALwaJ9
h/z5a9hiprxpayZ8HtwhHpp0CNFUnPzlwKVhiqfoTFq+Fq+Z9yqaSLv7piZmV5+m6HDSuKqnssJp
LtlrXAXfZnRDCQacaN89ydpk7/tksBFtcgwj/OhCrLjRpbY7OilHel6bOoqLJrykEcjfWp84g6YO
ZcgKDKFoAPmfvy7MkjlplnioI9IsBtiW4MDmjVVm14Y7lV2wv0yBP7+5pitPDeCa2JUbyMVO6rwP
HHy0oLAPUQPpz3+D0snBC9sWU0e6qDjNyLQvBg77PvmQcm6TDWPNeUC5AtS3//a91i5/a09M38Px
uDNlYEpRL6XVtgyttJb+UYbW97xYtEyQRlNw2kXbGAEu9ph/iPaORBYwAl5c8zSa1YoVjqlqkLty
b2hSn3KgsU1Lr/Dz2aL9YQEYrBHUr5vgK1ZRMFhCyDYFusMzJFkao3IifxV+F/RrAKtyys7MuRI+
ajv8FljLDvp4FnRqL3QNPZ9wD9LTCO2WvwShs4WOwb3VdYF/mOv0PJ2B/wtERvLrmOS5v9ItPJI6
iohRXnK5m8eTddcc4lchfjOFlH4+Ka4KNkXcdXhCmOpKc/tSvzWduaDbV9xoBgbvSlP7T7Zs3n2M
pp5aOA2T0J720caCa4vA5CZQEyME6GvH+vli40n8iKqR4CinCPW8dxHTqL20MngFRf61mE+cLDDr
JSOnhCYiSLNDDkJoR1BG9N4b8z2Oxo5Rv0ocjLBmJlhAxnwEMpuG1/AwdpdNyZftR4yVIjqf+MYT
6DWJnRsd/xRXnvFs8KTrZJ+dZ0a9BPDnR/v3VFwR2EX/dMf1OJ/teYcZYDpm4yTz0EnvcL4Gtyg8
5os8hPfSnbE+VWlgBzIiAA6EUJYLH3mZmxuLcoMGagCqkxf1szWdVNfrTLlHBXsSIoexgbaEy/nb
vaMdXDfRWPNYTRBBXcHzzbFcd2WYzc3z4jZtliAgRoy4yZfG3/tYnXWNDyz44exhpOqK7OGpQIlA
YCbuDbed+jMNHLMLOaVmM5izOFRcxGFyfxbGt8QAlhyvitwTKIIdENTzv5uUT6jLpAHfC/qdF5Dz
N+RAQCHhi0n2JWfmcryvfNH1SgX1xMcHq4yo3jPkv0L4y4YkuNZ6I0Mf7SutafxAIVgAPRguhk1h
ftD04MhnGP+ORpW/9OXktn048vcBmBugALEegzG9j8xtN0+s5aBIk2ON4CK3gFOYymCjtSA7zV1b
wUW8OnzRL4rsQ5V6ppjUV7tXGVD0rzPUDGQNWgq8Cy75qi79iCN8OVpXKhyojIx7oQqP6TNVxBK2
Gr67S8haavJSl/1hiv7FtPSvszhdbXfgi8foJzAEVTtSbBcHdRgrqVj7o2f7lVGdH21oA5tawpvm
/03ifI7wkS0KggCGIs75xqf1NGcomSgj2FMJo0m4NS73kSALoYCF1v7RHd/0C2eOiMs1qzofrGhW
FUBZuY1jaGCFQrHbQN8aPJYYXo2vEsoFWZoP3Z9cib6cgvmmFyzCQqTNnmopaHVxlkiilRWbVoTq
nVRjCm9wVDg7usGtV7MvxS69hLG55Jl9t0dMirGnC+JoiJ51xZ29+pz5VCJAYCjKG+2aaVOESBmZ
oXxhhBZByruOKACSaP8VadnQkCP4QPai0j0qOP6FBOCjXS4j1doeiIBW6JowgQdTvPGsUu1JRSZM
SXW4uytBo5/bjoFwHy9L+GlhXS3PoVwrMx6jNUu9IraejyF2QyxkNKUWlfCmt9jKa7U1efEiTWVN
siTxgZji53pL+66Ta4CdOOkkEizI+n6WIvcQH0O2GAUtnhA/XvghKVTqpMX+FrK3c6qQ2X1dgId7
KbAJAli+edtpMjfhTlFL/bsTZosgaJHptrUuUhN7cRIHI2V6vrvjpMt6w5vI6TUYE+vHbl4/RUes
y5ii82781Y0o3vO+hd3YKyAMCOo400NpY66VqPJD0eWaJ3JnDZU/cwGWqNgIGJTkqwFXdUi++3s2
sdoJiVQ5/nu1iYiQoYngJPF6csuFR+o0sxAgppupKNrisuXpe/miynZfL0xFcKULpT1zQA17vHFD
n8AHkZtpo8expfqtWjE7wa/weE80BHaQFTgfJMnkt9JBdK2CMbYLC7LTKXGvKFW0ScoQkK8+PIjT
VOhlK7y0QzUY9B9BT2x9+SqSuec1N+oeSLIiYNzH3uHF8RGtD0WDIbLxSVC/z4jD3YYl/zwrCOjy
RdTUBk8XFp000U1ZKgKw8W7i1ulx8gFJPmQ+zOsfN1CLAGU8MYqIAmdQufjb44BwAu79F7R29fAj
gzP/mba+zmS+ON0gWxlPoS46p0vOu6gZJED/DUe9e97Y5gUj5jH/LSVTJXwM7eK5tNYR+EpAMS3x
u8iVlzZsiiMIFuxDCZKzmT3Inmu188BSuo5gtaoBxn/RqKEq94s8dAlFSrrW4vUJxhezWwTKnSdT
8XRPOwFugIGKhSweNMPVyHPolpE91+i+c8qs3XxYJyVjPrsqHs8SQGI1J9R93W59kxSmxDe+xp2F
X1laZTc6UQpF2Yw1LQCKbuIqKNT5QlCh7BZIaktM+dkjArkPxJ+4IwMdHYbA8raiyCX/QljPGl/0
rk20SnMRcaMBAjCkM80n4xZ1gaOtd4plK/NtzoRSbgY7rFWKtlvI2CpM1TdvjrJo4DDGJ+mgXArf
YMLUrpsmzBhE+EZQA0fS0XqoZ61U0sivwV6UzfM6rcYj7vmEUChWF0qVikdmQCRiL1IC+dT/zvrD
OLQQXopK/n1f+GDKjqF7Wz5H9MjAgsvEr8cLL4MqofkN8LFiGib5Cy0AOKfBUMjc/7KXPteuvmnQ
xMAQzLAUCJoXdUfdQR/WFWGHK1ZfZbrXK3r/UYgpnAUN31FPhlx1rpKE9eEr8x3JNI0z6JQ3tvNl
aNbFLaLD+yiftVJsqTJSjDTl2ZUdMkGFnohIE5XDJQPCz7BXjrXn6hoqHCq0PKlA/K3iOO3ESiVK
Zi0CeYJCAjA1mI/0Q38NjACYT6nDvecreuxKnPIdYjEsjAJS2dZm2MVnEWX65yUnYH66+HN0HJpJ
qj/OPOLcPWlu12WvVY68TaSgSdPhhQZlfa2OcLtdx4Ib2J0b/yhvZN1P3FYVmrtjGvr/SZNTVhdV
IrNial9F6WLEAEZtRArlL8iDa9ZU43qcjXldnKuLymJQU57VMK/P8bn8y+suzwK03JZFE1umrxZl
8A8gjm7/GVpJSnWXj1VztUgYQC7X3Bd5jSXZrhTIFhLb3npY8XaceGLdGyWLta5VIBjJCJsup6JZ
rOWewtWQfvjhz6/3LF+ambWA9RFXUBrekdAd+qF6eUTeULfqnzHn87CwbjR1P1hMKZWhJtJq5Z+S
MoWEh2OTkpKaEd6yCAbuQiKXzcF5w6EgMv0ZJvDiDnd2g87inzcgsEwj6Pz4KB8riZQij9SRjiCv
Iok8pxDJaCLvcvzqG5RfXcP0H+orCJqEvyX1IC6q3jyLEjE8KWC/7zz4E80d1dWVy0mf90Hgwn0c
Q5lK1RbbM/z+kp9ljZUMe/JUz61k80ium9DxZyUlrsKMV1+Na46JXj8MWVFssFUmPigLEhZbHowi
tJSZgUw+J23Y+dT7+A9e9vcdL0O+/WGrpgUif9gPWbos6g0eLToelJezhrEED+zdXpioPNdk/TTN
9E2Yr1OZgYzz1oQhS2CbWQGEP+VpjEmbqsIXWqndXYYGoV2nx82M6mI/+AKYyDr0kW+4BqM0YJtS
2imgfkDdhjBS0JMsdzEK9z3c2wJiP7gAlkyZ8rsNNCduOGFL2CWh6zBolTooYTTAsVTcfeFwJtXL
+UaMRk//MFbSAXMY+KGlned0A/CBPVw5H0ApxFOX4yLWcZU2Jx25M7fQjuAL2FhLszL6D7rKclPN
NqdXZElqxqZzsKH2u5LJ3X+lM/IX7gQTLiYXqS0KjpsVit5DLR5J/BLJBEVTqOf5eZ2Le2I8PUUZ
/usGt1JfGoxPNRfPdgCLztb8QJf8X3xCHrEaXUqhbLqcDVFWYRt07uzB+jpbPGrZ1FJGysb67Alq
tNtF0xpp04vX1mYF7Hced6xZGlCLSkq3lPxY3y/33/C9tWEkr5DF2q7n5tHmvfVJerqPGrTXAivk
P9mjPQi4FTJCC26OVqyN5dcd2DtuUdoTEAka9sN75DQbZal8fl5beQ3uxqTwT2SMcDKE5r2JGwXZ
/yf3Q4xBbH4X38rILu7BgjMU9HvGkTYS5L0yl6RtB3pLYIkZO//wjdr1EfWHVLro+NA0jL8Ij8fG
XuENBiAz5t939PGo7CktQw7OjJoHvuHcLJw3bEoX86HE6bufE1mHACgVdU9R67NPM4bjh6FC+1WX
G1mTfw7SLlQFr8SbnNbWsS1Ha3L+bRbYsJa4BgO16rdbK0Z//Qchbqkd9Apzg6nsZ0zK2LZAKE0y
mpceAnb3/VwhO4LTePC1qfJ3sk+n4gDAsLIL0UbLb2h18bzTCBEhtYgRKwr25fBV94H8OUvXezx8
cvCKJYmnd9e5Sd0fpQlEemypAt/PI6mYuEnCrZBsOHEC27rLfARkVdMt3WuakCGUU23bN70tLMeJ
IDoISk/JC+by48r6jX8SWBFV5I5aGOWvHXvZiWgpCSbjllxtbfKMm/Qopkzz+76Y0jtLgYiZGn7w
Suk0X821ffnfuQezb1y6c1F1v/12dWztJhf6RXv36lgCBBx0IOAYMUDPIK/TOp9NVKE/2dZSHPiF
mGMrRiL8bOH2+7qe3zNX92v29WipumWU3Th5pmBovtNBIEtFDwLMSqjX+jRg1NL6BRrbGr/5yRaX
DfdxF0KTZlu7H9glox3Gn/yPv5YyGwo2NCEUseyGdIfciByHMiFIuPJpqA1llysSRgHp1bFQpehG
fy4MHM8OmoFFxQ940Di0jlXBP1GLNq5shLO7EvWjuMgdlMOv9vg9yWctKjv6Fp3Js+VPe4t5wNSi
NJJlzhuIgzre+/fYr03MFflGnhF+cMFUrJ4kkViq1aA6GBVex2nHuENBDLxm4ne99DS0vRea8K7k
AjaYj3riNj/sFtypuibC2NrFkk6xr342zk062NQuHFkEgSltoshmXUSFXCVFah9aned6g/+WuqoT
sM+GoveusF4mzu+d1gKi7qLygkMsRApxy0P13Ns9wgCVmC420dQ9A2K6yAlhwHpdGq2L7921DeoO
dhnFnujxyylL2xCbKGluJ/pHiagQmt1Cg5NkQ3oP7UdR1/gEFEx9bqzAXQxpYO7mvsZyd12PSpZ2
t1rCiSK37gLYViqzkfpB4lxjkTKbAPg3PW2IgUGUdt8R7XMDWpTqAvn1GJ8hYPWAh2i6AuvKiO8Z
EEUrnHv0u9ub1ZuxNFaNfjz3Z5s9c0OSz1mzqe1wzfz8w3aulwn0gAJaHI57Xe3J24cmKX9liwG/
NP+CDDlQxSMlF7igrg2jktvTeoL85fI54UL8KOT+tRPG8nj/fvXivgVWS/7i52TjHIZyGpsPzRYc
E+3FO3/DW4RN7/8WNc8gyBJBEl37qgjFpKM2sQMuvBbI2o7hRjTMr0rTx8DBxgXjnxMk7r+6ostZ
iCjUYfoOEi4y4Wf68vO/XUBVgvMONb9QPrLJRWeoI8p9rL8wo90QBKKgExV1wrkyWbaxoOUXW/3N
3kjjjYnR2rKOnbP4/s2ZawJvdnZONhC11w33Qelh/JVY+iE+yHRC9TImr80iaDg9EfEzNVpcAg+o
xi5pJmVA9r2m4zIhjJbzhRsegB7WJoT49+fjkP5kcO2YQ+sO8lykGGwiWkWJL/KWe08cYuVL53db
rCWEJ4TQ1oRyZp85QE7AhQ3PP4Dgr8lIAaQVXb0LBQfYR1crAeDDER44K3UX/7kzf2++V1NDFk68
jNAwR1Q/WAWrO18JWM/Nanb2A2hXCof5YJn058UrhnZIskWUX3c+rCmbvUfMTvlXICsvwcqwqVv4
mrbvzIcirUFXHPMVg0bk136tHh0xKVBrsyQuDPrF20qLpmFpe3F3adTK8V7oN10d+I7sUQUIXeU7
Ul2fm6z8ZF56AF2/lrI6BZ5CEtclTkS0jx4XvB4P/a6sagXNsToPOAq0Pz5Hwb7htqMaDJEDTNvw
Dh41OsQmXNiiJKG9PYbT5ad8nFjM3VVAbSi+uKJZvSMkvCPanHg+jstZqsvtEu5MjWiii42TT4iS
cgJG1b77uZwSsXgiHyNG3YEQ0GOxZoQ+2aHBDA6FidI3mCQ8VaBKT0FUPBKFC/icvScczcISjIaD
7iYkVu/tA/h3EA7ls9ZZj7Iqm4KyTROOyYFpbGMeI+tb5Z4jbNeK8qb4aYt0kcFlZrd2tqe/xZJb
FJKjSR3o8mlEHCIiSIPdiL1a+sf8+wnZ1/MjJNEFCCkrjqF9SVVT/Utfyf6JtqLZmhCn4DuHeWfK
F/STd6jAJWAIEKf/sDZoLdUgRKdSWEB4RZ9Uzd0cvaxI0SVy0M/mMhLA6bWV7vk6F31kpZmpwjng
DaUdg3sqSmBGYR2RerNWe4oNxmXbLZBjXabUYQuE2WU1zw8ml1bmtloyTVPoe0xE2k6p1uQBpjTm
OH8I2Xa2SJx4h68TDN7xWTkAlH8/r9Kgn7lyfb4KesVvOUn0ml1w0vqbiyG0ja83rmM8d93UWQu1
dc6ZJfShx8iiUMcV15xcYb0UgS/kiPz/KqBLXf87l/MyzsVl6wcxPsvjcg/3Beiqkne7PXgzZR0r
lOnReQj3wtoVq1CWOAnCKAUwkAvL37GzZ5TVd2ECvTeYHEWOapjuxwhzhvinOI34qh7YMJB6iVUI
OX2IP1bkgXvRljd/xxX0Bhci1ausn+Z4ZG+Ue2FJ5QtDS9tx1CbtAVdey25BhqkqyFfwAl00SOT1
0UZb3NWZACuPvHTstLm1ziOEEUTTtWIra7FDnHCGVkMebSZAixbiyenJRfoTFj0GYMGkNXuO2t+E
NKaMY/DQ0/mBi5ezXzXSWvxvvUzow6pkWB1exYjYnM5HWQTNcd52tVsTFuOAKVPiU8b+2hVgA9HB
PNWeaYmhlRrTmrCu+QD16MfghBKS+4D9hRwFEom/ZtVaEx7/Uo3RsB+zRCX+wvQc7YrCDXaPXAZN
P7CzdX311pyuOMUsam8VOgDlzSFJj05Qb73sn+RTvJ84hdbSLvzmO1C5hBcWLpSsTQsng+tCh1/m
Y9THE6mKMoryxeS6ZfqdcfmBsTycuUAGlKd9VxVCKsV/FCjVp2djlkQQ9GgolW50g3oEuXtPIs3Y
gyeJvBy9l2UEAMS33xVLqVzVy3DVsM135ZwesfNcog3mtl7BYIiGdxj1w/lEz7PaBI4bC4zZqW9Y
R9XzloBw+mfC99OXyrUnvEYva2J0z4A0H+kzHMpUyzTQ+/oNSYf8if2R+p/l/qvYRQMnIvNgojPm
THndcpZyFTKEbDvXA48XmCGOHP2lEsoSOhsnKJdNdTcE10XtP4KANZduKuFpN4HVwrvyiTqeSygb
31lfYMKvWzpDp2tIhXTz6lxiZUZG+HgKS46LmC9PiEtUWlXGpGs1Ldg35jgsLyfUslYRB7Zhg+zO
dqOMWbU6il85osZL01ex+DQJZRlO5dsQyYAscqYNG9j02EfaXjPovwIlVYaBe2p2byXx+8GLZOTQ
iOJ67RCWiCsgCq1acZ8WaNIOUjLFwbV+rlXlZGwuFQZbc44Pk2JwlVabH9wW2zbQycMmjdkHo2UX
fEGSTJ8LlqwmmEGB0ilIBIA5MUJxa4zlll7f+Rk1wZCyg/gwksuhiVkb7/Mj8OajPNJo9JGlAXJS
80zcNR9TZtxv7fP3NEQUXflcmZNE29bjlB2J9LZRCKgLtr3b43hv3cnS4rvrVLuKgegmaHwprFVp
7zhKVq/2CdU4mwHq0zb2TqdNveUuabV9G6K7myuoresKMjtrwzMs9BCGXyJF0BKhscpmPJfzcC4/
AYMHM/20tHd6g3fplHSzArpYLxQVDzJ1ZmKGoGvpOTysMZ8Iv4sJzeY3v8pohtGQsQdUjogE2eBv
9NxLHkMihG+2mZUZd9YUqHWjDBaBuPzOqNrO/OaF+/qY5x6jU5PZJQj1oX9ppo0gP1yuoaTEMEPl
8W7tcw1XUeDTy8owmnKSc2SlxdiR5eHQpTEPGz6EBp+sdDvQdo56seqXQ0/iddMgvdmvDb0xnQc+
Sem15QVE3SiJ+3u0d1VZSpaIkHq/XxxB7ztNn3oDt4z/BVitfzuDYROU+2RagdUe3LdIH6T4MpZm
GOXiQ2vy8ivVb4mKvSVs55+q7a1uCJxo6FyooXI/FzFqs77AwOZR4Td9jj9Ru+njicGXgYYjuT8n
iP2fVTxZv6x7ZS7+HJmUZFdxWylUn2sBSi5W9ncErTl8323QewYUVWWbynbT3UwmlZPLz55OD13U
Bj6IlM6jZFvvLS15HZdxLBX5nCPE6ieZRM8PGqXWLCHkhtt9bP7XVKtqW1+wece6kahMs14syE+m
dUrpWd7z+iueD65JCOy48/YgsY6egRYffA9fQ7Cg6FRv6pslAFZXHGRMqpk53Zu3675ln39Obx8A
bcDVMR2e5hu9zwyoaWp7nhTB8yXLC2UjX4FPTWQ8utBcgDcob++yM+m2vZCRb5J0N6jb/8iXyMWO
7lMk5itKk9i26uXs8AwJ05r1DdLtIlHjzYYCk7HFqX0kUFZjb9b75/nlC1nwjK1nttFqz2/dN02c
cXCoYlHbvC+VkbxkD2HfdOnWNg0kmWmtFg20jHt/KeDvSRvvXpUxiMRaB/X5By3/GcPSY6QQMiR/
j0dQhghuonMMsF1paVXE9Moc2SrwNvyxLfrLFVKbqOGNNCwxeIg0Yq/ec9X02mGoloMZT+1JFmBv
B08o4TYJXzBuITyzv6ifVPXFcoMG3+sb9B9/gisOxdY6HDneMQxy8g5AGKW+HIR36croSsmbu61y
L3/XaWLbE7n4SPeN9fpu1G3xZMpTP+hwgc/iqSQGbXstAXvt8zEH6kwxkRWURPHRUe/Cld7CpmE/
AyyjWvjjF9vn6cwJmgHMlMGkw/zCvCM4VQe9S/ED2aFSH66J2SDOxRtY9e8MLgIm2AEB/ObVEJkH
urDrjnrri5X1BZ3sZnfju8DrKXVTMUUjPy2JTlLsO20uTjDEBJGQnTO+qpZvgId8cv8rrxUeApe8
1VE5qiD6JU983gBra5gEpYSZ3lyoiJrIirGqSRRP9YSiPya0G56WwyHtc34S1c+gusxI7oIcFtuK
I/rEGCuD/f/A0ikAJaDWFkpy9/sjhfUByhpAQIHDFoLXBb+v4TkQIdpYs3pH1zB0EmnO4io3WhE2
+8D9EgfGR5ONpU0RebGODkvPXdDb/UQM1/r7oSf66OIxetdTqv79m86UyfqKAJJ8CUE4A8Qbfg8n
9ND/7OmtH6pDdmS4A2E8pdZil+xvUZlc9XqPv1QetJWKn7s5u4qJnY8TO+0jW7yWKy2xZhwNZ2oy
RAxUirdqRtqjrWOX+i1JFk3n8bzYd4HT6gXzrv07N8yqzAMsGOagtU/3uRVT4gKLo1hlo7sjIldl
VS88Vd29g6afij8DRnmkg5R/Jm1icjp/U6bc/H9z26iixnb47qjbux71LVmgKOKHdX+7x1hujjmK
Y9xj3dNu0fllRzIdK92iG//BTvvqKztbH1VRebgjCsTnr66/8RpxnbpctSAWQ7gVS1S86QTFt1ON
jM2M7pOykQgFL83vwAiMqTgS7NThbmLQ0W53NuXQmaopCUBDUexsPp3BzXaLLj7qKWteqvUYDv/B
2IvzuCqwLeKza2ihWt5Wylu2+wQZUII8lTt/0NeFHg8MqwcdJEMwHhqQUqDO2u4qZMIQiVhahWF8
ePFk/NKnhPnOn3d90np3Y2EJITe6w7fIIJsiiNU3YuvjXGrHX04wWulY0V7fv7L7FfCaIp7ZEKG/
txFjRDMqrLuRMyufzXIc6D//vyuf1mzTbLm8pnX4kowiESipIFzWbM64HJtOFEa6D9JoDFVOhPMx
GWLVwNm0Hsv/NIK0s3Z8n0DgMpNWA2AqQfNr0TQJWJBGSwjJxtk97HcR6dS9Ghob4VBS8oU+3mVv
+rg6/tzVST55JEd3wY+tGNA3x9MuSRVT0cYqcHKLBQH701hrFz3pk1vhudg0IK720xTRSgtGom3B
KTiFB/1/UemsJmpESGSdCNOI8fEDt/VtJadNGbH/+xN/2/u7WFfLaOaN+g7m6UqSELSKkljEbo/c
Qn04lmxw5Zpa8brc+tIqH939H/MdOl+BI0VEM5W5Do0Ab6b0wx+6VSRyzZH2eNUdf8ZwYdDiJiT9
Ua/5powNzINmUCRvc1UEoqFzFrbhoFAbZLaDxfREHGcZnKMtFdbRT4oWucUhL9Dd90ac6u4VH6Z1
nfu5Ua4ro+G5Dk6A7Cub/HaSPHc0zPIXUMRsj/gpm1zNBswWtpFD+X9Kr7OuCzOF0+gsK0y38AaX
cwLEJP3qnoHu4MjDW8sbOyNSVvLnXMWfByiuJ7bO0wXAQPBx4UgtEsBtRNnnxQDsaoodi93JDEQF
PInjybKo/J/AOcAfv3BhPjmT/hx7vTwznPTE9/taNv4QXs8E7/hyQrudbZukXi4fqfdzwYtVyCSy
DZfXWzXINImY9+GGhuBysIzVqTnxwAWOKgp85eAOEcXqTc/pANT7mjTP1EFnVrH9CcsidHJnuV3E
hz3E0G3ZaUfskMxWZ4ZGJlk2Pqh+r2jmMWTBGQxF9B2dV86WAIq4hD0RWeojF1yWhzHEC9ffzEzQ
Xc7AT2wOfF1IPJULESIYkYiVnq4WMsbGjMr6CkzFVwcw/FgAarg5PDDlrGiN7mZeD2IdOFMbl9hH
/z8nXqJouExUcEMY1lfP2yQQ48hBEnQf9m5MdsItD2NQdTG8zURVh/5IMqixxV7wWOQZJCFK874Q
rRla0Uoc2ExV/SCbxX0YKEVK8TTYpJ1XfUGkfnuyFsfXFE+nrwQ1TPE9qbpSXHkRNpTnbsDhI476
RmBpNuGu0S+v31PO4SpJvz+KPqngvAIwat5O7I9t6yY1QbBu6InW8T0VG9N6Gfnoo3TEwdWUpp0O
+wgk1vPTsbLcvJ+/pNaotJPDBCy1eGdm8ME7lOsJNeq32y9sMvpCe5PuIiqdH4WMc7N0VlT6GtEU
DxE4DB39HbSg9MXP43fr/vrxAARJnbyu3MeRIDpXLqBJs5DYtn4gtPJfMGRvO8MRMqr7vl/p7HCt
5KyrM0jVNRq/QliXJlyxlcz+Ppn6RAkqxMwdMl9UkWjc08/Ql81cC6gMEgq5Y6kF9jBVy8kthKsA
Ft4zUcD1nKrOsa4aPTDT375sL1nly9+7xz+EtYELggEK+C65R2gfg8kF0HXJE+1kMmc9v0YaeVow
01ARJYJqYrcxPQKTXD4beS4hwuzDFGEu67O3GENft8M+NzBIzUMJ+Nr21vtQFT9qUafxRBXF0+3S
PJvm2koJYBWEKm8vHxmDx0ULmXOtMVtp7tCXOCSIGMkwyrN0nODH2N71Eheql3Lo+01n/R0cTWJH
EiNmeR6TI0o+zI0sk73aJdly8Ddf+L3aqchMh6uLKF0uUfLr2+UJyzCQcg4tmJL2V2x7uyIKUYPr
CKa2ad8vWmm2G/3X6AYXy/0nXAQHk2bT5yTJbNGSeExGaj78A/vPHitecu25PHN1Mjgx20rzqRHZ
lzSL9hec/67BgMoO2JtGJFwLE11ndZ0pVo7gMasFphTVeh6QjM99pFehFzhISgFkfJcx7qFEeHIX
R2/xNuvI9c6vum2jqaFGB0wdn+SEgEGBqExzMWjaz5uPuyZq7BH6Y7Z3USPgn170SKaUjfBY2uMc
8t7rEAXi6TKhkos24oN7gxP43EXJlzH8aY4SoSqnEUMuFf+DFgliARQan496q6ieKKD9FIRoMEav
fo2UkwFiay+DSjAkVzf7kp5bQXV+kSYsUwe4Fo8lrsAUKd9JHa9dekLcPql0LQLmXYYTNeXRT/z9
yGtVlfw0QxvGl+CMzvyHPe5X5gLHA2D+kenf9svd9juI/5WyX5LkscVRg0fNuGnYKxR+BUVWjJE3
MnRqHC5HxaHpkOdqeflnNONVLO26u+pidBlAWoSYEqmKFgecluY9BZljmxduG2ix7ZzMJw966KZJ
uUdkWJfFHJDhhtimeEQHT6XKSbC3nnxG6O9TMk8hQETcSXMKReoJE3pLgFDsY88GVklYhNqF7JDG
zEoOnCBjl9oTliizrRx0DYPEvU37doiRDb7k/StB//pJeW3yO6HF1nxi3cjjjXsHs0F5+YqGe/+E
oLcsBvYKkgk7X4Wn2Yzi0Mn+lLLZ52r/ytga2+AEYQXoanculnTpsrAVeiMyCqaA6SisFKKwvaCt
2PUk1zHf1ahK0maqvQ6xqcdA8zi6rAuApDhaNBs6Gbj1As048jxwa1K9MMhhHgiOQHryJfxOx+9B
OuO6sMrtdQ200/tGy5cKs4grGF0kThg4qcoxPbPBNINzyuO0UYmcGMpoTy18NRS7kf/ikpikk7at
tANJtfQ6gTelh1oWMHTz8z9dEWyaYS49s3eOKFyDe1dtglhG0rQyC1ymaw+U05s50McMnO2JpLrE
Sgpk79RX+WJ2zGqfDLwJho4U3/YgspOyHd6K/4B6h2tP22SNCsZF1R1OSYN9Z7WyoWGaUw6AHRvL
66iILNOJXobqG75c2heMUA/oyLWQ49gaXqRawh9PE14E2aobo9lTdxb6a2QWBg9I4YvorLhebVGJ
nIWF5+4e9wJrlBp9nzIgUHrMFcthGU8M+r/thOvaG6GTOWRTzxrQ5IOn0lSNteipmh2NUC134nGa
7J6PmEzva+BNnyXc5zXOb4yJK7cgWLH39LJas2IueDhKyNYBxT9/FEbLeioowkfRz29Kqv2djVPt
8nhz28940+HEldMKTATggs8kFefVA8WTmuZFexM4MbxDAxjy/Ppxgy1jTTjxqL4aQ35NKVpDc4Z0
XaxSnlpqqLNIYCqg43/1JfKsRBV9YZ8H4A4G17BycNgMwP6gnCVttGxhcXQZW41L20CRxv7WK2Qm
VnDSE9GfLI7jT/Uqxgm8TUpaD+37CGUKpgbC7LYhLLZk0FPqZm+NKn03ZvO5hMRnpIwmTnXm4ANK
M6GcYX+T1qAIbuxb2V9IG4xn4l7ry6iRqiBbhbJvn72cASxpHVxseFvGm62MWskrRUiwIpKZ/c7G
jQbkexXs5jjnThZeWmmWpQa+ozrqtV9nvwRSMhbGEt6wqknZoLuUozfmhBOYRcf61PfObB9z9moI
kpwfZ+pYM0Lg63RAlp3f5G5mA7TykA6C7BAv6Wd0A/u/nxXevbulLSBIfKy0vZ5PvTkT2OtTETQe
1erNeSwIH1KRUyRJlRwKwxA9JHhUBcKxmMFmz242mUzhdp5bbSYkq4IUZoukxo/96CrmeKrRIh9N
3FGnoDKenuKK/jD8KWKyj4HHaQSeL+0xLFD+Ei9FmCn81yc5Wi43Wn2Zh6N6yYaG3GpubGhOFJv3
xBCrSdZQfSwNbD8PZvFpvAsKhY361t0zJCJvtKUyRQ6nmA849WHdxqDWZiLVS/hBtw1CTZxNQ0sr
3xFown+1YHAEFA++BqVPxdCvPJTw3M3ZIzMFf1HD/0T+QrkUXAqcO5jbNdLKPSj6b2LQWPI+zzDv
p/oyTPcvvNc7SOXCqjIMDSedgQdgSHxTX6EKJghtUNMBP41HoYohz9mhbdDDHO57oIxB9NjyoEPY
vDnxTT8YG+6MpZ6+0CzN3LR/5s1vSbTo1aWs4o+ZSngCThcStTbRpuCB4IpJGXzD/b9KQ9xCTEXn
9zPLvX48BtNHZEeZjvhj79VH+wWjcYV+JmsOuFod6EqU1SaIqx1gD4zkusWMXVFvPtLwjCD2V4N+
U/tY4U2s/fyqMxS91fHEjlQccYCoZNQtAWrWCNsXcK02iz2CecwJBN/26DOKCi0WesHfsvUxgqfb
3EADmkOv3tn/1VXbX1KFqxOtc7tUGJQ1u0oZOjG4K2vPUd5QqEwUyMD3miybgJbSLuxX1OQdElgv
rvGcTzqGtrGc475ClJjeTDLKJgnTyBz2G6ya1Li9pL8NmHjkJtOoohfXzcJy18Aplyuy1Om9yFkk
gsQoVkDWWg/V3GS2JZl9FxlNOJYqolO7/bigH94p6nLLV4ByAMiz8lUND3gK6zMCZB7IwL/f0RG+
S4rQEkFGrC/z3imDo0IEaz380+anDe3vZHH3yeJxdTzAMYJJFkRTDV78mL8b00rd27GdFiCVpRVG
/vt9/rl9+/lPVhX/mf5NlvXTw2jWcKmhDmGbVngASslE4uaNlLhjbAXHENyjJYKM4mJfzf1ku6LJ
7PyPPJtTzxIJqiaHC5YTNoQZch9iKki7Skbh9yOXw630lwrRCDm/ZvlZ9eKAeh+1a/GB0YKQOlpI
sSLM2yUEtCTJN5i8aU9qdXAAAOx1O4QjtV9E5LQoViUM2RI4Ihsj62UXgfekNyuEwf04cysWGO4G
64SNLAmZS4xXgEzgLLYrMHskW+cmboOtB1OuYIuuRdwS7Z9uncREXeuNofR26JN031lzEZnRI14h
Gflpe0zAYp3uqpHJkQnK91w+HxHIphrGroiX+KzwJxy2qbnWYIzC7UqmqMyLIV+YdNryWP0BJXxo
9tG2cz3sz9n7y191kT/C2d9YYSFQrU3DycEb/fwikoxUC1d883D50dAGmGOmkw+UHpj3pJ4MUM7x
RKoVZkOITN1tLAU54O+9eLuFr785YIeWzUveBIFvbc1niSc6oF+2qXNA8diByvx5Xg06Fpxl2r2A
Qia+x+GKTUbpfmf3MnCK3MHnnUOJs/EPG/HOkjwMHCTreuIy3G31rCL+/E9nOBe3VCiUIQ4iENdH
N0XjLkJyX4Z/2521tNQYA/6cl9qKDqVsN7vDNtdvW4rijGNsCw63ChYMlxUVl327NjwYmrTVQuyE
pfTua+0FnyeUamn5wepxMtugqSwVtXXLvJYn5H0fLDYxsObwMEPCTQkVjCnklIHuhveKEw/3kqKO
cn5qEHY2mg94kqHJtesdfoK4tMDQK2nqhclFHlif7U9VnoR6ghu1DHbJlUqXU5JKMAtKcWCu9T7u
OWnWeQNZHIB5U7KVFkE4MFJaVSTDE6myIYhGx2oOuWZbDrZ2ZDC++K48pJa4zzrouA8i5qkQ2rCD
g/1NAg/h8MkTfvSnfLZ89w5E4XM5zA5jG9F5O66CAaTfW5FrBmhj9OV+BNZX1EYSnCh0YAlg6UNK
XLok6IPCsb9dTUtl80EJR6bZyVYJnkfOv9xfE8H6jmfkQ2BD6RQhbjjzQr8pgfnYu22csxAevRMv
6nIxxa4A0ljDOacRV/YcwblOEbmiasqtWrRVifb91FvQJB0EOCChAZUyiAcfKWn8ooaI/91A20BM
ZNTi/iHK+XjV7exVQ+94MjPuNWzekHkTSsqdE9Qqs6GdNX/xZle5LOpvJVkNq11//nD7cjwpQV3V
Wlsna7/S513WC83VEezWIC/J9Z4Eo+36aDbKymT/fzChPWF2HHHIXIvZ2xrrhnvniamxk5rU0pbK
Y7nV5oIQLNyS+WZy/LxGif70wd3R1ledTvi3BzBnMQdthv6f6mBQOdKcMry4mt9L0ioVSK7hcwPw
myrK0C6jcFCFV1f85gqAuNKS2seuIq+5WO0Ics0IM5fH3MQZ+MgUL1JWkZN1COh+EP2uqKvBpZlz
ZZiwSraSE0IQnfpSJMoebZ+sjCigLFxrhEGUGz3x0n/JWrHYcMve4iiAzgd3xNgAgkTtiZzF2HYj
neuWKLRh4lbz7YkJoXz7+OW67+UHB4WeH6es7gXQm/wB+0cwUXakNtpJkL1th1kmcTM30os9SZhW
Z1KKjkzbhvCFm7xnl7RonBTCiqLtTHPHVHxL9L+xG32ELtjJtViFxkqPswCw3Lrzzu50zP61zuSe
CTMskhIlIS3Oz5KhdS+h0q5xALXJY53TgKLuHhrCXYWC8x34eV2Pw4KdD+r0iO14gzcNegS3l2+L
eFza0o3oXKR6zuBbhyWb+h5m44ExKW0YVWbjsAuipQDCbMR6hcFdzmt24s1Lbc8yYUv8zeFxdbnN
avaHkpvXWrpRVoEGabWULqOnaBNMHMj1YbcHAxKL1H2RzGgwRD7xMEJqjJjkqkCOukU0PpwMHfxa
Q+BZSl2XIdyPV+ZEp+Y7pvSV5W01EwYdbvTK85UG4BZ8V3nJCJeECWa8vWBYi3+aoYTiKiD83Hlh
ub0IvSWfVL1w99Eb7tfLX8KekwgGxQx75abzNARhnJ5qmCK50PlEvY9C82os0ZtsBGhWYv4InWcr
KntuxNQEWAt3UzgwUKDcvju0dMIJOnSpi/fD+mKL+mFJtlUsEL2SbcCSXRFesT1V7AGUUOVXjfZq
fbU/NJV/kneacHY2wqQYU6dj15bj3/Mf3oQHrqqTiqeM6FGzjRPePQuaBem6cpj7GU6u+0KA711S
RUJb05T7jVWuqfiSqf6HTQsqQkEE3KVjhfX6dVL2NhEiSfEOi4pfgP0JK2dyHXvv+YKIUiLgj/+y
Lefw7o4qUYo4A0JMx/F8BQERavDN8UmP/Eo7ZzwCijXXr+3l2Q6fmGSfSqWzu5LTl5aV2VNdWWSg
beihpyS6xVAOcOlleQoYakWoQhsIa8byl0EBPK33ZUDAbWB80DrEHYy/RNv0zGYEd9AKkyGfCsL2
MvRSpl+p73w8xu4BipRCU0dixHpD0q7TXBkHoIToBkDRAhu03LnH0qHfcU5eDeEaV49uaOLHbyzn
XT/ev6NRLHZNcOJ9m7zCVrFrcqlI3e9/5l0dLdZmm/JkSyxt7SOTnpuJwAiQ54fbg3oHRfhq5Li5
ceGzGLyDFVnc6Vj4DchHcT8IZo/Z51I+ovlgPT3qD8UkY7qpNPvMotKaqhYvbmfbfHPpqXJwITkx
T8S6drrXXl/PW80beo0uFo0yMEPkiK/Z55rzGfNzFaVZH63U8o5Rdk7e9rCWJ+x+O4xNbuScNeor
cMiRkS2plNHzm+PAVlMX59ip51zorzFjabS7AKa6TvsQ6Xht9JujhxBK52ciOdjmJmkZktj00uyD
wBXo+eMmrhRMXp4Tg9KjP3biksRAJFwjeJcucY8P6ZZfLBE4wlLQVnPIvVugNir5uWLHNymYJsZ8
+Pu8CYnxws4nZ//EhmgTOeuR8uZpBQsvRskxf2wTJxSh/dnbzAJmTnEzwD3gpMEgRnMrebhTqM71
jfEzUpFO+SGxtz5TwO/WEN0WtipsoUT3uQh5ZeOCErzobqZ8gd3e2PkvU2imbd0AIyBiudeHQ6O4
SaK82HJF4Bux0VslJm+1LHR8TZKt4F4QbFNRYnY1a5Ip84GFWzzdlr3W9IHMZ6QgYc7u4350wVWF
N6RdPI8YzFDRCLN2QDuFv17oXi3L7lTkn2NUgCSB7ErU+lrIf3PRFK8uAuYK6jAMxlc/Sl3+9ZAQ
tVPHYNIsHL6uUNWUEK8gl9gtYf/eATKpVZ0FkvkBkp4BUdaM9Slyx/GwdmkP8ssrMeHkaPeIuoqf
rOSFSTKmsCLZdE18iWnB425goESiwD3+7NLdUi6vYnnfP4mKi/ek3IHhLQDM3/e+QtfXwPr3hhem
zDLFx2jSFY9/50pQwmIw2Q1z1U7rgpAcoEUSTiSgH4Qkvf28ix8J/3KeYYCH3rFC7E8trs0jwCL0
sW14aAuNt1lrPt879HVdzNUsQ8e3YHOTjDQ6QjSLQ4vXoUHo1zfs7ipDAou6kXdK8oqBaljMIEOh
f/F331A78hV7rX1Itwnh/l8gr+alHwOFxSf/qssxmlMrjBRJCMY9AevuSZs1yiswObZGnGb9l3rg
yA08aaDRBk5nzWeT/e2C2fQE7IsZLVDyOYlGpFtjxdMIQChtYVp05uTKptwQ6cOhwb7NoMbIrbTr
GBkZFcjRHKdaTjXsrDkqllBXnYVDoALL/1J0JSU/cu0lOnF5WPiOPTYU9AL7Wim+RDvFIOED4Chi
qoGOcwj752QEeCMt0FNIeU6f3tgybNzbcFMa5flF+tkOGNsii9GfOQhWIHqD/z1ptQRSZIoDVTNK
aNz9Rm6VrMRhAwGWpilgn/RruAteO5lXudEYMf+tvFrygmnSu6MshMLbmXcCgkP1y9g9eIPuFzZL
E/ydBJVKVBC4TctVP06BQHjLMsg8T+LhqaP/vX2VgwvSXyu5KpR9v7g/zgep7ZfODezOewEhdAdi
CbsWpf7LDXgR3Luc5uTP4GSYa2pTSBDCbEZvN4Ixz6SPeJWre2V4jtsI+5hVfJBjfjk+1zvZmKPV
ZyVhl0+Q4PmwBBtl7NYLlubsOq2KnImUNB2uSSTDnWegSceAQopWsC30+++EGFjDg7r9S3LyxYvI
6Ma5KZj7ZmF5HfmhuCjFpwWpzXoB9mbt0ZzuAFy/FphUMBo4bvHTdMLeGgDndW8x614UQzQR+F4s
ROO3N1pEaWK9xqTBT2umX47X/x8zWu6hIP86cK0GtBtwiB8lQXqD/lgQ//qS4rC2D+kJ1XFFLxYD
9Y83vhuXHNpKYT8iqkAeNnL2Lf56yVQpgxRj5IZsD3kgNcEGthHxWyy4csrYdtedONgJnnLeynif
3ZiiA1M/91yU1kf+IAkTLwO94U2AUxNbogxVv0lc/dqkUMHUG+UuyXu5u/dWUEd0kWksIJspSpWz
0FucmmvxH/rbbMAEAjRzTclRZ3/prNbS1zwtiwweLpiWZl8QFfUncM61fsw6oitUGe0xegXaook4
tIK2QpXqvbfjSDgaV/cwuclf4BcWSBs1RmPKMN/gvETvbr5/plvPG9iouus6E11bsJy/pNWBt/si
qeYQgE8yoYalVUXgbbaTH2WHZm8VHlEZ4CqAf1VBayJntFrHNGSSzzZKutBZV71ouwFlRllXvKpH
zr14RkfLGFsH6B9hNf1+6XU+O9Et8XCubbu9mxKT6CTuKTp50/mdsI0PpRXxptIzQ3+m+88shRLL
5VI4wim+ooVFZRUYjYOZDF3wf9EwC/4ceIdn7ZaXIuMWk9FYdbjdr7yxGhazuMuJ9W0puTEf8A2e
dEceWgNBnOh7H4c9kb3egy2kJ56GHBOo2NkSKf3h5wmrbqwjyP5B95GZEW9gOleio0TnrAoQCN7e
2Tqg4ZcyeKRXxE8gx1CrenAg4FtfaEVrFpNYTUDHy12gzjjMsqh+YZGjpiKNjDmZAMYZOkOJqyxm
XkUoNM373X3W1wmCmnQ2TJQPwRk45M3cFW38GYRdcWNCV46MSzx72Zg7txO9NOmh/jXRtrM3xSuK
m1xxKFUNz5Oj4puO48H4YUTD3n/dVndlTNRV/VMTbRwr3KDzW2CT3e2fBNOmnzRgOdysjDnlPmx3
wbzVfDBrePM9Cn0qqH1RIkY7JVEgXoM/GduPZ/MxnqRV6WrgKBlXNGa8MsmfXnuFyl32Ajgq6Jll
q0FP1Td/pa+YvlfiB+KxxyJ36eJ2ce//9/iOknEh6htaADllCDK53uCvWgXaUvFfIu+0e745CJ/3
uGK/qvoDuVG1ygswcCcRJvrr2Tru5RFd+KWYEcRVH1x0N5zjlpxWpKmXuLn3BPLHlZ2h0L/Nq+oC
Nxqcu2Ugx+Swl1qdRi2I1IyM8KtZNbWRQetfk+DgipAZGT+q/5Uc76ffuTAAR1vTGjCcY2RZtq6S
XWqlN51vXW3wdj/K/heAKiS7RJrOPrPMy5RhHBPDYF5oobJeqouM87Vwp9aOj6R1PjCPcRlEFcNi
DaCFMGIpFylV/xC2RSfYYIEfamOwy704HT/G2/g/9SNjPvE6D/z0xzCg1UzD4mSayI7jhkTtK+K4
YJhYAcSqAWyL0QgwQ/pLH2cnUFeW8JlBqGvah19qtV8sdGEPc+FoYM2BnPt1OCD6VZuLsZ7Nd3FP
5bKG+Dl+kiuBgpeQ2eln5sT4QjU/7KkvdAqaySjlIcmTE+ANxN4Ehk4RKl0GQ+DpWEw+jLUCwK8g
8op9gmklq9CcFKdyoRZxKy1E+79kycrB0LuDVI/H4pyryJMTVY2SrhvD5WoqXHXuBOiS1cVK1rUY
aQwM/yPhBI8Tx2KMdm+3ay1HYn2iutGqYFQ9kqfzvgr+jpb9xfZ9Ovu5WBMGBC8XqdctDkl+fUFE
UdFmwWEYuew1s6QRuTA541cTnRLbFOMI92NZrB3UqA8Q6p1gZaIY86N6vkfhBJXLmo/waophnULf
hmzuG+8c6neh5g7ljUT8SBKCaEFBpClNESxGtUQzxsZs709F3u01Jtt+4B7/p+rzKZSRsfyibdg3
44+3qoE9565WqnqAYS8a/6bagfT0v5pwxdrNTq405L4NCGdzB5b0qddaNHeGAxdzwYHmtodr5FwR
ByEoYJC/FBCDSK63S3F7ee0TRnwlPCjgP9brzeSPWg5K7y5l0fj3QWEnRQ+4hNk/UkKlQRU743mR
o5UpKFcGT34xywBxgKl3GMvjdQqSgojHpxhDmbgFhWB1AY8MgPvgis9i2+3f2jsTqdchs3Os4SOU
mrVq+ZqCZvhWA/+oKjvbUpP6QiGp9GOzgPCTmz9SYISM36CtTmEMyUqMjTJFG94SUBIgi39TCRDK
puzS//Eg7zGz0db5YJIgvHgt7kOd0u14kjKjyzGL3bi6qW4Eo8QTNqU0Teuw8iTZw1F3ISSowKB0
Gdy4OTJblLz02py1oo258BUIPlR/uII2bl6CaK4kAI54320Qo2bIJEwR72uiy/RIAIgfE1RfAU+s
A+VLM1a3VKD+e+I8uNXGI3AAdkuvguvBUNSFLU3ugEbgKgZNy4MpYXkyKXvM1xDgU03d6Zy0bPn4
hm8AoHlH3Nz5BfX2bLY20fcMpGiVlrZWHSxpKscUTRekyyd5zIbgRk02sEA6m88YfA8pTV32NWIP
XY81AX+Zxk4wtrp24EPAHig1votQ7Ikkw6p3q+m/biGePC+a4+Obe4f4ScBZJTME9QOM7GVN1L+6
F3vPDebco02h2jWFZ6MhDMq176bodG6crPBOSlNLx2n+0GTk5hQjXwdck8C0Njx+/FPw1Mgoc6/T
CjPIIKD+h7qm20mgqF9JIOTXDmCYNFxbfc/5HvW5iYCO2krMthYJbdgeCeGScVIPG2UOw44z57pj
CfVhkXVYf8yaaGOiFn6DVxjcCVOlhygyRENEhbVPpU2p/4EAqCF2it68KrKaMbfNy5LLpa12MeGQ
aZTf1QfnKdbRV83R2od7J0KbmCYfPbRcBe/S5edWv6YOF0yQPrQp7pezOA1ByH66Ex0/oRjDHstA
1UsQV9+1k2jLasJ1uulDBDXiX7r0PaIDxqjLL3fTG6nPiHJg/DrqibOvl1s33bDEvnUVl1Qel5hv
bGGKaoXpSp10CQBqUGq5k7x+iZI5qB7DUHQ/csmFkIgsitbmLKz5sjoS1tQ3/ztOJRV9puEM2NiY
SDPt7pt14ZMQUoZH2Nv1cHYX5Bz9L8gfLlB4vULhf+yyXNAxSLk2VPEfvtFrFlgGEyTFyskAw2HP
iHElhn3MmgANJz9x2xFLUklwn6VAzePhjdUHZ3i/E9tEwGXeZo4kzbqdJd0oSbzJhM8u/guQZHqI
P00TCyho3exDWLN88SdmjZETAm1UD1U8V4lay7m7J40nEFaWLyv7MLAFaNH8IOnSl62dthOIEo69
PvqzZnVkdqei/JIbc2gIAdiTsT299K3bAOBfhlc07oWLGRkPjh+HqK8uk99kDtIy6Vl4rJBHVksE
5tFcGQ6SZOulYn7yfWUbtCpNKnDKLcQmhMDrTs3beBMIqNFKI3hPvjTui4e8NYN4YAL2o2++c3XI
zJZ+SllEYsQvKtC5j9+4OIMDOmgsQipgaGzwv4x3TpW5fCGVwPB17g2VSSYtvB/xysL5aIxZu7EH
mmnDl0It1Z9dHBM0eKa+2QCnZWh43DRpwxFP5sHfq1VJmozrRn2W7ixZFv4K140uBv0fpzkjf2ks
zVg86sWVP3zfCdEMBvdj1o8da4PxuFfhv7nO6Bq7RxdC7P0/1py1rD2VC0axPZszjDNp0m8k01w4
Iyc3INLNa1ltfOmeUCCLB3oKrpHiC6RDm4lVCKxKHj8D4/sVUAfViGHZK4Y1ZWkTlM2qmHy7QJEq
1JnV+iddDm7qiPlc46BUSJo03tCZesecmUiAj+FNXj85630ET2jPle+Oy2hW5AYchZS0/JFA6eNe
jBnthMDT996oann9kuQ6ZgMjdsdWzYX3QsrN9n2RL6hGd9rYeXsO2kOjilPDaBodqYdWaJH06XOj
Zmx/FmwSHr2CX9REVc2jvio8btPc4p+HjAuNq85GHJYdzY6hiv3kZ0gCzLsyb05rS2DdMd4goUOl
D4TK+60gv4Ypd0BcAasAVS5nxGCA67Xvy/6obv93Z7TBH2g1vgqL841zOB7GqGlQ0CkiIowR1zmv
cHIYaoeWs6tqXFSuiuZaKSSRwEwqyeGWLJc107AfPzgfQNEsewwF4p+Cj9xginfzZWRc+R+S4ulV
Dc9ms9D/Wq4PECjZAS5/j9X8BtaX3vcKXcHIEk4l8ll/XsNkAtEfwVCLzpfnqoOHPGfkn5ggkFFo
XYoJ3Ge5b0wv7mYORtmGKOGZGjdMcAdnY+44WJ1vTYBg6tecs8Uy6ZYcdzQm0LCPVYwUGQYzhbBs
FMvooeJd2Ayuyc8r90b+5cACyTebh7bGe4huccRad5R2OhaI2G+ZSbGhGFsa1zT21hZGMzD3OL7R
S4xdyPo5Af6uYnUhj+n8M7Z6he3rhauq6X8gzHvzu43qVtCWeX6M7dj/W4EzRVCRFC3t3X+di/yO
udeUgZPEJdoaapcfbnQbzpzA0NO6k86b6MHA1Ajhjt+tgZwAjQvjTFAOZoKdXUINBu/wJtFYbRez
bdD81rbgiivJqXDPPxuqUB0ZEK1L29qLKeMTP8Su0DUKudqVq5uUwFM1a2SQ3x4j5J9xHNx3NqR4
v5eWTU5aXHt3MJdD911MDTXGfnghdtHTGeV+eav+YIEJBRREv/KC7SniVW+MmwHI4xirmGOyvlVK
oATYurht6FTOVD0IQti5InLrNvFTv926Yq8pt4NOUFsOGdIQeOuUtfWQiTljGJKWBHTH1OEaTSm8
caOKgAo3zY8rO5so8D3DRNjvvDTwrfh+q+86k/yrHB6b4crSuxOvUHq91fjGk4raXq7ffGXv+zn8
b8PHy5Nnd2Md+a8GO1JMjItPtpxOnPz4MDUOYlwg2piTLl2vZHDS2SRLS09p7JiMW0J9ci1NOKtl
iN+9OB1GCYDuy+AcXUI40o73Q4Qc1MDkbbYeryy6UnxfRb8yfuWcmFHQpfuqUeKg+dzFz88ncdZU
DJSVEVEytFxAGrGQpb8H6ZR80VJuPBCjgYDk8n3qwyKbfu5Glmc9NuI5/Qx3HacHGBNFC1B8EodS
pHzwyHlLjdHJ07CIQAiyB4jnv1Yb+d7HZ0RXfoWy4kuXgt1rJGhbWkx1yC3VWqRQ/W9316/TWJdt
Txe+reM2B6lQuya4osndrgzru/HoGaWNez5Pgg/Q7a1t2SkbKxW94InYoaCRPbzQzMismxETTF2G
8M7wdx2Fnr6FvlyKHavDyy7pIeaFrM2muRfUIU3/UbJEDg+QtG00L01QoIhCZJEVlRzTWRkEogjK
5FjkwA0KU3AxRS7M+kDHn07V/lP5ZViwiMN/FIkD8emC8JG3tnY3HSOOxyqy1zfeTRJ6Gfd8NSZg
y37McQdwGaB+yCl4qzGHi8xRcniPlSNI7kfygxY/qp67SfdsVXC4Z5kacVsdg4sT2vtqzu2gKXqu
qIZSVzO0zHMrlGrc9trP1Q7qIUDT9nIl1E5cItWIOMPp7iN+HptGbojGASJ3jAkmF+ta9moih/hy
Qb+MeNsBZrJZFEPHQ8q4psRXENRlvpwxClyeJLxL1yBmebyEdt1HHpNWOoLt+UVjqorf6kBMjeGi
r8glR0Px62gdaD9XqHne3M3xmCaEmaNsw4Wz52LP0W4s0eePMXTukhErfGscmIV9261VYr91f8OR
9EcjLWXK0PkDj5oQMVzqQiepbc0IHHaWsIEn0muGvcZJxOUmHTlqOk2cXC5HYN62Cs3NQgvCHWlf
JEL7MzcwjeYIhGh5+yI/KalfmdPHSiqQcvEoDsbaIlGMB0lvQORIgrFpW/ADctqAkdjnscuQMw6/
QWFzfM+IilI1nLTmsDC6xuf1KvQ6uiXwB5LMA0Sw84qjtpBiEDVoHJymTAkk0TflRzzSUZRna5en
uWk059N/CuS4ZxvSWXuRIgsLZLnXDrZ+OLIkeuBok+/XOj3S/A2q2+BQIDP6CZi/NkSJF63qSuVC
S/fkzLrQglRQITaJPMiabIisQLF9JrfRJKj/SC1abKAVxI/n3jHTHCBdNB88nbxWOVftM26kKpSx
3YuImI9YZBk6uVzoYAyZU3WNoa0427Lo0MvzNgCQSRaBf5b/j0MCoPIb4kO7o9KeGxggB5Xrg7Hv
uuKdT/IqdFG7a9+M01Ibwlxfs9HW6UxjHtLKj1UPNvypsgmJ6TU8tJic3yCm6sSCYP4TnRA2dqhO
Igr5i+haUYXXfrvBdxp032jlZrmxU9SY8hGki0WONpJwAvg9xXi72yC0et2F8WgPVKKm2pR1rnI4
LUWz1xpvn1dXPWsDATGr9aMv3G2bkDKjEGa6IACCJbNPMirgIhOmIQQMWNB5R6r4u/GJwleDmBZe
P206DyWnfxATktY3PH9vpa++Umpsbo8kgbNqxHgYskymc7hPxaSISWz8VgeWPgkICIMAkiwjYZ07
y64cEjU+JkHKq8XcMC+qRez8X289E3W2PADUuG9TQTlzFlajmiKMyha72XV35Zj7xpg1AGxj60YI
Lncv/Ft+eTXzLE3zoeYWySiMofQLsPIhzbN5H0PAWAI/QgCdZRzx+vN8lb/GbW4u9PzCKH9CX57j
WR/V8seSSRBZRgnk9/dfMwJs4eW6BzK5oP+7MixnZsKHLB05+JFUvmTHYbHcwNTcXPNw4w+j17Ts
kJK5rdKEoPw5mKbDCivsIrGJiLpc4nLYOX/fXiS9RJvshBpolo1Wo/AhOvEHybauLG+W24nXxVq4
n/Epzcv3Cv92QkmrwtOr0GT9ImrjBraOvk5BVuq+FWbn82m3ccalk36GadTmER03ZOl9CPuIEOhd
fTaPaVmdW7UMLXtneakHN89edIqnlzB8wz0ZKgAbOq6ClIFJKNKaGI0I4luL5SDnhq/+MvAM5RWI
DNeTseY68Veq6H1KdqRD47MBawTdhLBt+SAsrvdftcRlbZtDw/QxuPrdn6edgi2Q1v84LdBgcG6j
Kkuwyzp1vVD+aF5Th+FaMrsIU9wPg7Oopg/TKDRidIWzRYH+jAhX2qzfFlflO/Z9CrF+vlQC9aMT
gxvYElZP505KLtTr7YpXSp1uYCxJCwr//NXDSkhorLIizZjaI8mb59NpTCUNLcGcc+Zw5dWhR8mI
NG2TqsBWtY98UAo6V2S9x/H7elwMl5o1JZ7DpeXZHof8t6QUdYfbpbrhOasnJg/wNrPXDJp5NRar
mnS+YSo/wEhtC49eXuLm6xnnj5VTE9L/6eYmbDeDQ3HVaU8x3xv+713WYRNavQLo9JJRUHBX3mlt
4NeHxP21aPXNPyT7Ra7yduEhojzS2htNet0CHL+RYkixIShkdQkGBJoeit7Rfg/X+X9/kkwM/YsH
WpYyM4JcWWqg7TZXbnsfXkyUKBe7hkG1HDHIEHtcNEEN6eCopJtEzs+97vhrxA64W0+zN67nR5Rp
5h4b50byIX1vjdeE7WTSVLybhGXjR+1ecaahtP4Vx/0Q5uRfydUfVrE4nTmfRIy5i6Mc1Oef8s2r
yvfSzZ/YiZbAsASdWjLqzn6ci7XQDgKmGHdBXJo3vXaeHKXS+IPnEFfiynK2j8ZXoQ9qn4XZ6eQb
RnWxmdQTm7r5ZFVw7bIhjDGC0mH7Je+HJPp5F75r2Jh4FwNLP/xrTVIPCcJF5A6e0IA9Eg3Zg6pw
i9gs0/4ZcQ+AC9WOAwjLUIn+K6QlQOvVBILnLWs6CoUkUmU7rPsStY0b6dgue+5/y7jb/xm9NXlJ
u6bcAKbNk9rxXAAWmy+oM5EB+1qM0Ku7BAbbSHrEzCKCJwX2AaehlJMiYfOlVeEewfk4l17PB3Oy
T2BL7X4lb8zxK2BJ54Hvik4ufwNYmNYudVY83gxcIS+gvJxklGHLVj9ZxbTTe+JhNz0oqBbwueID
kO+0qRaWFDlQuK9nvYvoTc6GJ1knxlFnEWsMPW7QPOr4nKHLeBTYzaLazws5CgeA0gag50yk+nnB
o71mgUtf7eAFsb1jznjNhdPBEnD6IBZRCvg52bD8jjsDkgzmckI2Ogfm7sRN7eSg7F1A5huugVyF
Zp+Y4x6DMcGy96lr76vj8FY51Lzlt1jLAA0Vy+G5AKxwKZKqc1Rnmj2Zl5Xr/fqkjq3XPEs+ivlE
RTq0Xazu0+950RlLbo7FMPxnvUaRL0zAnTu1TSptFOfG207wSk6cFgIXeP+xTtYdbwffYPnHFWVM
+qTpIe0CJFXSBd12w0sXIlMf4ACu8v0Nk+sdX+ooD9ClRuFvHsjJSMAMhTMAX3k9uRkh9FfuBRCF
aIPFABKO9NAERO8oPLmLpbSda0Se/l2azlrsHTAoXiVK2mXhVZXEvrrsQVee5PhWrXDTFOrl1H8C
h+831F9RQWTeFLksxNYZ4fTspsZ+vtyotcbFwqdzK07P8wWVduhltelVW3MP8veX4HGBeTxVZ5RF
AtgFf7uh1mfBC1k9+7WX/NppsC5AwpU0+oIXUo5B3M3htGR2GSH8ktyfrrgquxZOhPLpNqVS6rds
H7zhsINu0upiAuf/ADewKQ/Yh/uzfQnPvk3umEgtKpyLMMe5dAJPZ7lq6uk9wy6mnPb1+rYHrGl0
cL/+mJYOSdXXFI8cNiNp2b2dFL87atiL/r8UMSOI4niZY0qgbpJHBsg0hndiem2ToWUyPbvpX1rK
hwuWqJdUtO/wDnHy1GWph1Li6oRdIkstWBB3XyUxerNu2672K2VVBuhQNfIp43Xf0OgfikwWjxHK
Qdo8J/Q+KGtH82qT293wrdt6gIldiM8b7RDhWE6HjX1YrgJC4gBzt2vZtqHw+8H/ap8er72JMz8e
wcdtNiKifJS1SjJs5zMKRLRnyOgvJE33jdWB63InSAUgNvqd3tmiAo27p2Q54zZV5TAw1cGcOBXm
Oq/QXdIh9pPBnDNyEZLeKd/5+bX8kRORFgG7RUuTtOgvApxz9eZxNqTGisNRlY9jwO7G/Aoq+Ngg
If35od3MaBnqXa4S4WucWZl+RuM/P7bVUB77VtsSrj5kqKZHT4goBy77P8F7RVsKrgBpCAKav3yK
Zpbfv63CvQsRsZBckkjcxskeDO3cNtowyuZXAUy1u3ToYtOq/xtQ1Lk7CiISqHbpC+i3NPeE+NzV
obLqR9pmm6otk/acG8cfRqVR5lmqq+LRQ5DYQYugXrdn6Ha0TTU8OhXdbnydaBNzZJGPpBSPNUjv
MXg0jwy94QsQHAgIKfBEdRj7ydwi2ZDlaCicdZvs34EnwvdrhSpenbNqZXvFWBbHRNPGwUmdVQr6
Q6NC00gyRWQ+lwPRT9d4+2DJ3J9Rzib3p+4PvLoUC3Do+D49IEQuwRi+lL2MfedKQXRG0iwwbjLX
v3j5EaNjqUIZNGB9eqt0/R6/pYvwgcjVSnhfQxj+jb+n0fQycliFZ+wNI5vZw3n+z8vab3Qp58E3
FZrwxPMOAA6r8FfxUyt/wN04Tmp7R2pm/p9Tjy0ec+BMIF65gQQFmvi2xtF0+HHGlvs5/wPdbPkO
PGyX0H80EIfiihvueE9QCwzerR0L3fKMR9tUMDOnDl4dbHmbwbfb4EXbD6Lt6ZoKQ1z3GXfNPbQ2
OpdEyM/JxHqYHophkCcK93GbE8Gq8MmW4ip8qWMAGs5d92mGhZ2D/2bneVf4WeDq4jg7THOc1E/t
H3yk1Uv1wYtWH9vk4azqsH8KoOpi+LFhEGp93tU9Gle7ZQ8UGSoa0X02R/npOmeQPrvJnvuMA5Ls
fe0nVvwGMHEnh408umg4LAh+V+4LPk9As+WBPTp/ApG+1LcWCjdL+stSyUiwruEx6QTrxFCi8IRv
/XXwvPmEiPNFyWV+/WuvhTqNorqNct0C3+V3roez9x6dQs4rraxfZQTUNoBMzorLudUuG1XP94bR
ju3TDDSmjusHq+cbRsy+XaHo+KcrI5xtUTOzOfx8rhXPXkMUWAVBQwqpXamWNF4Q6K/xrKuUqOPg
R5r+6b9buQcIcsKmZ1L+eYIDnlTh4WcgZEYIAfMff6JpqF10JxWsI38xqgaSKu76UJhJNwTLNeJj
4mc+HJgarnR63EU7mZce+m1NM2gczyKa04GQBH/+G0km1Fk8jh5YbsEFaqjftjCWX9MGXj1PjQAS
hADjTLPtOvr8+LwpFXzshTL+tizM5qDufmuykSB3rOMLsC2Zs4BSeIr4xRNaKMQ0rvsENd6BlsfC
H46uwaNmj5GxHQ64X43fwHE9xCht/uFFnpM0T5CJUGKoKOoMBWXxbz2kH18YuLyzW/qK5gnmrl/l
iQ0+Nwt1BxO5sGUbmrMSK+Xe1FPPD4jRm/eD2xY+dA1fKmO6D2TxBa8QYzhUaWo5q4HfHyrPipPg
zK4hYtymAh2Huc/y3eFcf9x9/AHlaLWtGnuBc43gNB3PWm1ZpfhlvtNE/juDeaFDdMNTTT7QUawX
7rb4UvLzXpdiZ4KO1uOPL8cy4LxqlRPJ892yWmUbpEPo1J3kkA73PZ3kwyfwbSp/bv0J8Uf+0M2Z
eE4zv2PRWEy0fk+LBier7tFEYw4d/Q7FfoYz4Yw0qaLtHbMWbzHV1jbW1GW67Ch1ER3ajMlRC214
foeSGJ4aeg5rQUStyaUUL8RzUD09n74pcceTt3fVpN4RhuCcdlTQEjEIv46i+BRrZxvRshaAemG2
60TEqJq3S2r/+lLdB3iCjo3x4ZWHccGqUQr3J3Q4SwC/yZKBDS7FY1pnfJd/AMNNjINkNH1bW51z
FRM3jBQ+eL0coZ1xbtJ4YqEF4JFZoTJJMHNFT/FjQlKQvJGOmw9G/nrKRkWDayAdAirV/JkAXaGs
tMiT2ngXkFcR89NiKrXTOwtUtEY1eN2dI/BM8xchEXaUvKjlihNsDdGfsisVeAyM8S7iYa4m9tZi
pNqlnUCFwMom9fqkcbTIYS1HU07MtlXwtrSLg3o8oeOcIBBp15JcqZ9z10gJ52XxpTj+RV6N02WN
kBZPmaDQ/qGs8g2KYntsW979AGU5hzEj1M+9PLgIVCM+HjzQk1GNdl/I3CZXWJZXeHhgRdiPe0p3
4I5UENDBgHOYGGhDvPKplf8AEFVmBVjrTxvksfUCMw7RdWnLrLXQCdrELqMB87bdGHASZgnWsxRi
gK/d2BCz8i/xgI0nU5uJcgm+mwB/vURHgw00PBqquookp2s95cVLUu41aa0iKkuT6+m4CJlVrEHL
j9cbbKtaY4oLaq/mYmQyZUswA+xXhysDJxZEwnAS4Q0xvu+NYq+nzwOp/kiS5vD9KmBM7CrRMkBJ
HccsqKon12J9brd0n4G3RdE635cLds6/S3TeBEnvZeKFjrwO4L7Q3y1oeua8xf8qgs6oDEthB21C
IsDXaW1iP6w4wImRNq/gAnKzNlgedF4PnRDbMxutcuHlufGZrg8CMOMRgdv6qDWJUKxTl5Uexruw
TXekqWB6dWWywkyBO756zbda1zc1+gmm0k+rGWCOBqZe/Lgc2old9ChcT9k4XPYmNNeC1d2LGtL9
Z4Jk2Z4dPSqhWRD2/QIozdHdjPkqRUGzxrapZottY40o+1VruyvdC2yqQ7F+KMcx5GOB5OatZU6E
vKl9sckGuSLtj4OwXioE3jsKWoZBYuBVQiqd1ikLaX+5SY2+JVRcbNUODWJn5d88fggbjyBLqyQF
dp7oPwiagWd2wjwq431H0HjYN915wiuughZIKtLs11g79CLchtTmS3yU8/S+Of3kj1qvWaTCFHaw
qWo9unNmtHrTtTfSSohPcB9P8OZJnytg8NE1yBLViRkFK/iKXp+JzbG79JPj0AvfE9/9TH0XNIC3
Pyq6Jv5NVdu2xCEpTnoQK96wFkymOLaOau9p08UZmX/qNz1F298TZdSK1ObQzvQ2SIFihHY6ez5k
OEBaygeTiyuIbcerG3/Jtl4wHxwgY3KIKKcklVPa6OeRqRz11iNK6Jd9eBex+Y95EqwsZaBPH0l3
oaJoAOPjmnOZJWO1//6kG4BEZWT08Q2HJbwGscavIixrfb0UbmmsvpQMFn2liwYmM6wuKo4C7WU1
ruhfRut/CHQlZO5llgurVYdqp3LUpGSmYbucfNbYRDn9WWJiRMTBAwGkSTwikQlJL60xkui4ctR7
+boJ3fYxOBTE8d1u1Lkc8X0jLzbCr0PGPz4bsrYIq8bscw3iBME+SeXMZadNKw2bQ7EoOF++UnoN
WQ1X6Cqqx7dA0P7V1Fc80DaQMmZy/EhHE1US+rAh5A6uMCRnW1qHKaOnh8vU5U2A88LNpM7zHA8y
PaAxEBoETT9gtpwFXBPYxS2/QP0Bpva1usuzf1QLT/hMAXu9ZrXBrfMgp0wj9Dlb5Jw5EqYp99h5
uLIFE9YfQa03p22Y/wG5IVmNkGM7ZeH5vbH96tmpoCs+DMILNNbczNQoVoXQgInNWXYH5wAHq8E0
NYB6fTh5w1zbIFqwYjQuXXFxS1CubMecubIOR/uDTW6VDtIhfW2fKaRAE6JMtWUwYauE1juhbZqe
lyV+K4z6TiAvYKUY4PwYV7zzOsOtD2kzVJbx6nP8fV4xfZJNEzeFENqHbM/UcJGGo0MVvU1dnIQi
KA80T6Hz/peEhIxcFxDV0dpQUGLMNxrBDN1X7ljsKvQEvJpIYdpSigxK8k1OnWSNX4dC2eOKYOfy
Io5I1bJTNvtlUY1euRHY9onY6XVPs2Bnyey95gNg/BaOfTG6wevdIF2BoLn6Y5wpb2RjOtzTgu23
HkEZZ9kjsGRh9nlahHgpBqVZFdv6hKttbCc6KnbE0iy5V//wIZJUgs+KIZaqIp4wW9E+fNis7s5a
GtmIaJAc63oZEzhZ4TkfHohYd6JYQeD6EIccgmAEecwILCPS6PGuYVH6QfDyADLk7aGfPFTh2THT
boZ9K7jFFcyaxwsXfF4fkOeKQqV2TfuN0VOjFyC5wjhfA+rMRy09GgBT+EGwECVjBkSbW0ulkA/o
hhcpqa2TNam5qLvJyRHE4q3OxdBGPR2Ea/8jTaWgw/i8ElGWsp4raxI7SxpWJLCJt5HmC9HU3wKK
0SpQUOqOQ5M+jmfGH9RW5bCW2Tp+nIegS+QY5xPAukIOgc6YSAZ3+qJJhRpQfVo44uNaD+DqjEg5
mfBRzkJAk8mBh0cnIdTPPwcf41uL7S/nQu7HO81iNyLJMwq+0afElpTj/rMA97O27Qy1UwOYu1P5
uf/Q2n2q7vQvTJifiLWfpsMt7ym6yqZIWyiBwFdnDiH94rMwK8jfA94JbdAn8WkqX0woc5aqa7XC
tKIBp7WrXhaxgrf5uBr2FKO9auD8lxnj/mKm+pqC29cf3RoNE70LtsWCOeUcDalXG7HJ5Yv/ebD9
Ee/g5qGriaMn8hJk4FFeaejr8XqsBXJ8mCElggtva4Ahv6Hql5uXhkeFJhJjpJfKCQ2oPCzoMUt7
AWQdijJdJjBkbFFhqjPhMhqeY1bneDC34N/LKdwedGRUXxAhvYsHbgDWTIK7/XRC+zI41jXk3WHw
zRocwF8vl35sbw6W+sbz+UUXhv47NDamADoY+f3y9l+629lDYfptgPn981FwNKb/nKXYOXiX2KD0
SY9BIHhHUZXxV1+bFLEXBQbWBltNiUHFZlLGa9ddhkK2cxvlTuTy+JEGPxwncEENfq0XKwF64cz7
GHyvqfis++nyBzMdDj1QdZbdB1d4MjCV8sYZA7wj7NsiospiMWMQ4NurAPqhxpFjUseoJZ43kc75
OMFo8+sWZapIwlXY/NhkO1R2KuwiqBlFXzQXjbAc/TyTL4iSLtZ+Ip2DK2pHUEamCfllcU7BOmDm
+b10Fqjdg5rL9iKEG2kpxByFMOQj3d+LsBcU1y1ifR0Pacf/4xsgqZmHK9W/E4FQSs44gHHjZOpj
Yrm8u0vuWvWPBuHq4FD3xa+7fRo/ayv5Uy2y0UDajg22A2b9OGohpZmP17jWdGEebO3XIUkViyWR
TPwH7Q/PSak9Kifg/HWJ1bJwYNnKUeh9IjIe/lzXbdISlFv2IkwWoOLTPX6y5HT8zMMqPgYcu+v8
YFsPBMJd2IOScv3vmxbavgqFS8zqM7L8pnRPd7Swj7/LdzHgPGm1FjyMmGakHnXMIsUGQjnmM3Qe
1ifgYvgxQUC7y3K0wqYnLpv9rz8FCCBGWNIorK90i88WBP/pGKvrh5aiAqzwwlk2nAzXfTLgln0C
F/n7DW9xQD8zkq+SOUIkzlVBYAukaWcphBpQMSyqqq73O/OXG8UKTegakSj2CZ4uSu3Fd8TLnrrd
WEn7uO/SDLlGnpFxxaoAKQqIfVx+fApa5gbX332uEDjPsMpWy5xLewKuOAtXUgbGpIY8GHYGFcjl
1VGUN2RSnpnD+dit6ifXyB6a57/KcK1NT8QyGbTo95vycQh/biX36JF5PfH4Ei2OmC9LbDZy5b05
jx70K1wHOHXu05b55VgSYI5seG7AgrykG9B08awHJVbMxxWkjw/nbQMcoGd9/rIOUv58N0HFMjb+
4eH1GObgpX4LsUcCP74jyUyM24moy40rG/2TmYtQOaozPkdIEE7VOR8pljSerifVzFwp0mlfDC6T
h5r6ySORHKLBYNi6mZeQK9Nn9NUKHxuE+EHCvGVbRKEeWl1gTZLrqXjdnhWnhefmGtQctc1sjfo0
+yi9r8z03eMbaG6jGX6a124TjS8MJctiokjjldLOR7yvoUKH3Bi0KcyYCuWH1plx9msMbYvnAT7p
JfD1m9lXyc50fcdFgMkiNUAKT4tVQhJL+CdmtFiqtOB8KOXNBcGazP1Lyya+sAS/dzKYaIYXas3G
lnDLTcwI3WzyT1iYBF4Yh4NH6ubPPcsVfyBFZi8z8oMmAk41glQSRBOYfGyF3mulz68AVw/bUpyF
hXdigt++UJj3PgScTktZZm4mJKkCE6ZGgPJB/3aTaVmeTnO/WCIfrCPp7lU0L9KOu67+CCdYG5bT
UpSZUoiZxGsul0JC3lVVavH9sX8gfjLuuV06Y5lupgbdTnC/xESbLqAVtb0wXd0vlqL0skbhnAbf
cN4FRpUvuc3SU9NlkNW3YNrUjiNIB6NasI9mhnNqY9HZk7eI+NzmTxkod3g4uoxh8HivE1xfjuwH
bKgGaq//KptZsy40spQK4oBzL45almScrLwrXamIFa/pjguf0oGsSVDQMtNxZsrz2DiTXIww+s1Z
pzpSzw/V901QHah3AUW9X6zIgXy/OoBP9wYQMW4XeP6sTS+Dw54ljQP4/Blwq5Z/JrTF62yaClJ/
P1wPN8xfl/H5z89OFw7djeDuR3UWyocHECh4UdDlJaQYogIv5mai90YfPzJmB44+r7ndzAWkVBJq
IrFKAcCGE6urmH6fnhH638ojEIUFVtTlDHA5if5tW5ucVx1mirEWvEOb5pbyuMTtRgXjXLpvzsWO
A9iMC3/BU+DxK3DlpCkwflJpxZiH9JCfTD58IU03sQi3ER+35QGV4MeDrMbCgZLfWYdvA5Tcr6jG
JLO2n/I2O8Q8PKCfreXtgNuA5wGBzAGaFmBQymM5kH159Yxu1HD4kiLf1WairCHGWtaC543LL5Il
4Sl+C3urqJBTrH+l5BwV9RaSCgRKfku7QuiXfh8IMswc4a0aC536mxRAibIUQUNsvmZMx+aHc3kE
g8vkbLVzF+fr77pJ/Zt7MATsTmrL+ee1+ik7GbzZjrNhfkJbHw2u2L0MVBCaRimfoKCihYBmBNHF
FG/CLC30fTZJXUe3xJGo0uvgXSQQchTndDI6T2jiGVPwWj1OVYI5nYrludgJSzgZkhC21T/RuenP
0DqyVTwWpNwt2i0D0/b/hWY0m0QptieyoQbYIga0+EI9qdt2jrYwMwYls+bN2lgLDifhI2R83vhx
NCmxB/lEQ1yXqbFCkEs8y8Nr4B8auE7wS/L3EL1qmTCM2QhdPnIKceaNl/RsVhA7j21EwN/Fhjtj
ANmoVJxEtv8c25HMbddRKb+FPSidEjHCcu8KWxsmXR/RYIwasvs+2o7ytH+8/eCyIVUn99sCdZ15
I+TFVKzOHWP1NDWmZJNgc7qHBF1y7yMXYvbuQ7GAnNMoqGXu/DhhNb73etTxbqhvCcL6DAWsUpf9
si6inRhQQ5QsXsKF/HXoUfJJNUv+4G81357sJNSwhAILoMGoWs+HZMlG+Eb/gXWqeusz8HmeaveM
WWGjVsl30db3sOYotQpO9klTMqvK0NO3kosX58knMbYDsfQyZWjB7Ymo+SWl+uArLg1ILGbPjPqD
bG/tUMpAsw5byc3Craa5oAJUJfC1yhdZIyjEbhQ43brgqj9nipeT+g3NTHMILtlrO+UIWGPgeS3A
8fGIQbE21+uzDIb5vLkxp9dplsCLGq8WsT3QTc+gH4wRCbSsBxN4SGKEIHG4em2D4ALm6MEGuyd+
MuLZAvpzxnTpKHlO1Qmp6ETORCCoyxIsbMfMvJMUYDmdoW1P1g0J+QOBfnJb8FFEcj+M/tRE5A8X
+flpymIovY5noVH04coBXVFWqEAHhWg72janI348FM8ogcw+ekBSTTPhY4+usRR7qW5Ur47hrpjS
PmutS7MyaVRF3/ZbftXgoqvEtWpBQLHyq4RsXdZLFnerI4u0dQVnGQQ1f1oFV8mz2hV3Hwg2hoQJ
S3aOxysivZ0G4dZuZenj55A+bjgsBST4jJr0GHcX4ocwF2Pe+RTwNiSV3lGlYercSDDtxVcTCkXb
rvh0U/adluZ7SYtYI3dCRbLqF/Sqd2pw4oWrQ0msmToYohd6QXcMXtDCznY11LjHmlfS4xBeRSbv
fiyCbUQ50JK1kaTIBj/xq43WaOuNBu1A9hAEyB9FGl4PWWuIRRh11R41EJfKEzrDaOy+g9Skigei
HTNPTSCFlyjkqMO43MX+EGheNPqO6WtHpbPw257kePlvmDsZbocil2IjqfP5p+qctA4sNRH8h0Ig
JNZN+S4o7OKoJZJ1s9/E1i/Qcd8G2rnMhtqIZuB/PBf+MO3BMjxM/LPWWYmqN1LicPIVAfMUGL8I
t5wjk6A3UlYNG8r+4VB8ChHaXJgpDQx43REIPJMxqgL8bTpQ7GxtSK5W8YS8WdhRUvqoJUZ7SBFU
CGi47ny73pMZleXmnfknsxbRX9M6Zp5ky61FD96701+RRryjeFX9QXwfQBgvVcK67JoKEDLT6VpT
HShUiw2RTiQy+C4Bv7lCZZLORC4ARu5RDGlUdhKe2C2mQbVATmltYGv2MWGdKOmOgZTB4L/QP+Nw
rzB3PS/pxki/5A3KOCcvfPbmmme8kBu3zx49pnild2MZJfM+cS0AL9kyWTe3dxrDtk+Fp9cZEb7X
vtYjjZf2KI/gKiiKnCXaYzSE1L25TW7l4y3bajdd/n7HjmKr4svnZjXEIQsVFhXIkAIderhrVGbc
D8npgE125qJIL9dSylNj80jaFF9xGs/2Wvn80v84X2KAfdO92GpQDM/JlsU5u7RkCplGUr8Mk+yu
VsnpiemdlTSSZqx7+q8MUU23DbEnbuUAqAoxvwh/Z3Iz9Dy8XOqwrGUVhmJGiCazsEiCrDo5xDNp
z3dX9zke56shdkNU8l0KMKBY3yVq32FexdIFN6QB0K80tTW2sdvkf6wbQuT5MsU6yFKP9xaudfNy
s9jg5J+byFG3GJ/n6/7IffrOycbTFUUs7NRHdkNngdhOFB1BMgpCLtDrf2QqdZoJyqp4pl1QZGVQ
Qmv5x8QE1DMSZ+Py8Gt6PvgQakIvjAbzbFbHZWUEdzxPZPrJqKYnOagloilbc1O+pwI0SMJa1U5s
IvtqPywBimTuKxVCVZB5VPGzt5tnOaghBPgj5WYvUUUOt9/JxfEBuBdvR7/jOZ3C/AK/9a3+4LVz
n+LH9AuWrWXHmUxcfHgf9WaozE0tM7+wR07UMcKZ3exYcZB9i6Ip7A+2wOGNXzyJEmBT78XBu15/
BskqZXepFJUF7DUik8uIogDBYfquYMvkRIJcZmvwlY39FFGCNPEmt6ugsnpQzaiVLfcTIguaKLOF
+FVH3R8QPd889+tpk5gJdmOi4r0/lOJn7zP3mS73sN9NNQevr4+FFf0WLwSh+IcX2cFrVgvE5T2c
FsfMB1I7etVTbtKlY9VIdunNPG8msX6UkQEJptVEVCJl4XdGQmCpqtD++ZPTkjEn7qX08tUY/1Dk
/dDx77SjpgKO4nmM26bhag2y5IY45KuyvlS1kHzhMcICJTz+sArYYYzo84D5DKL0LIAOsd3suD3P
gyWje5bJqoxZcPSOApXPfXMK3vi6VI3+fQhmL9n6sju1Q49snY2k2hRDpzb7ErWJuKE703ySn3IT
LGzuKBYfznX0WsthrcmYtDUdPwoxd05WgFG+aeFQJFnCIme5xTkwbZfEPtyENhK3sho6Am9e04Nw
giSop7XLzGyd/gjqFVgYOof91y07HURWMY8MvEetiRNRg+IeRseoHB0b/jjHQ2FlumhKO9r6Jx0x
Fc96BWgNgipXIZ1c3gcL24+Jjx2RVe2gFpCHl2rVg9Z2EUixkHG2Wq3KhGqud4GhqxkxvkxQGiCU
gmb1xNOXqG4vfcoqg+gUExOF5Amtg24+fKDyV0+fbs6M3Npa+DdsA0q2KV+T1hDp0XC3/IKI8WoG
57RUmcsxlmQBURQMdbM63nNY1RGO5qEWJyqZ/JVH78FSzlBKjCLY11fbOQCq/T6YNY5Amy9X/yxx
i149Th3sKvxdhC1NNkuEBtjk5G+ZeNlDkG3piqVFsr/iIzAsxLA0nNvdW4YpjQs+wqR9O0MdRyuE
KMISLtQCwUaINGDm+LHyAB3N+LHNXIeXVaoV1EcQi/SljaWv3vBNTN15OG7eKuKhGz4OdDEPD/x/
Z2jtTGTOp9N6EzhKg/kqt3RIHmRjOsQ8jlTd+Ekhs2PBI80p2fSSqTbCcFYoVJdwZxYBLXJAQhd6
K+wdgifAJ51216bNmVhT7RPTVVIeF6SJVrE0846cWVemRMhuotremHS/y1kUB621G9B4zfIQ3scg
fUKAGY/oF2nTq22DelMtnTn2EJ0nVikkAHpQ65rdp7neLCqTGxq5rru5RdvRMQ+Ttsd15uQfBwa4
icUzqbk0qOluBTSxH+LhintqqvH7qQce+jvEdx7t4b4MNnp/zpv4PqEYi5Ewh5pl7TaeEADG67fq
B05cp95GIXzggRCUAmnRtQ+LJ5O88IC+7FUw6P0Xnv9sdb3gk22vt3At76zRHfESzjO7rGDcXNTL
g8j93UMqj8vP1UEWoCUUwgPaj9XpZx0Ixcv0mH/of9qw9U/tWrOS+V7IPWSHAc9hnZpdGeMlI3BM
g28NO1mr9Xg+hbS3YVrr62VcGSWEJfdC6/oHs5WGxBYBJ0iN1KF1oVQt/O8arVA2ER/1ZvcL5t5A
JFmGBykEoFKLcJCSTT4cXw282XAnAmo1au/1CI8KFs9sjjw2cSClaRdVTgVvmflxyE+hN34ruhQK
OOg60ZO6m1sWlqwMMbw6UQp5mdpR9ynpV3nenRMtsq8m5/izAxjFVkIPEOeJl+BNWJXUsLsK8z6N
dtsGt0IoA7nc4+IwPO0YgcN2sVPL9W3ex/S6m0+AYy+3oN78txD8KTEgfdAreomaJqHoIgLHyxOm
PA93V3wKeAwTpGs/VO1amKDJU/zBK2Ofc6EE6+9p8QkDsca08becwHMVwE6dubX2nFDAIG2SdiRh
+fgSGmYYHQx2qnyUK83mELACwX2W3JHjqfy76BYW5VQzvf2SsOSqrO2A493DJL3oM7npIi7SaWs7
uOM5EOvIc86shgXF50o2xPoeimUlmfXjP39mK4iHGm98cUfePWHugKZZrDw0jHtVq4N4h1lk/SQg
yVPd+IStko2gbfsAKB7wkA0K4IrQ9EURYCu9VrBJXBuKgSClMgwjZWtR5EeWrBPurAYcRlKrAopY
rQ9BSNcl2Kxyc23U88ck/qSTu0YTVkVqnpxWdWAV9H6s2kRpqvgBhodk5WaIvGiyUsZgPFDN6TEb
iWeJhSjqBG9WxG2eFAzfbbxmFa/k2BPmsqYYk4RfwD+aaQu2rGRizsFipymVGOvkxL4eYzLF16AH
PREs/4qGHn1inhj7hgRKa67/PSJTecFRGYWZaUZu3GFUP8vOVm0f3SgjGcDP6gJIKzffKVd9yyo3
Fy5Bs43VIVwD6Gck84En3gh5AguIpPVAh1xeBeyvHEnp+y8PUNtHjSTLsUx/h43nHeG2Qhk1ZTCU
Uncs/iTCs5n4zD2gaf4QRu72B/+fBuXLMDSxyfnCB6f2HktBZ9oIZgV//ejooSlLDkmbsrYHIXwI
TVkZiHQcC2o88rX4pX9pSB+EPvVmGKD0VOfqGZPwf3k7pyJ556UhyW+CYx7HmtbiJTGB+x7jsN4Q
BW6nsVVU3qdtVtY/HebgjBmHmiyOq1PSEL3rsJxd7/cPc0xDMfdbqQDfVRvLY64wWAr4S5C46/Ai
YbSBIylraDqp8+Opu/CdGg7xORu8U/XTt1/MKbNYhOb1MiOSjIJPCV3sFpvPXA+p+NMaDPvpN/8y
SUQgA7v3VcZ8MHqnShtRzrurvYM9PLjVV6lmgPcTYC/5rHHWbo8KfDuTJPPUIwpzu8mxRYflzUiJ
HyyLmQyP+LpG16Y3/rNTy/luXKS+746IiRPlklefqUKJ4rjbVmzvsuC7qy2mSaz9rVaG+SPWazty
XzmpVwr+y6ripOcSrHxpOvK+juptYlspkN37bxbkWz1yP+EeXPvS6xQr9cGJh39nifxejGrqzG2b
ju1t6w9ivLCV/um0kecJv593GDm3SUQ4Xo67McZ2ivbBmb/w4TRPBv8D+OtQGL/pZsPivFaSWUI/
NwOcXX0Fxf25PuEASZ7V8kT/yeADf6ROUisAupViSWSzsZrVQxMvr0gYIInNJ4yoTQCVHGVA3b4V
32iqeoU5uvEHsaDcpSIYKrrjNpGpCWi3aLcMoVuGH1mfq0l3r/c7JGbfwZxjj0gIGBkLB3zrRCpq
faQOVsGKYj+6U07Trt7zO5rqwgznciK+3N+H4cIeuvbE/+FkZLLhoLWuroMVNPwdpGCAw/OsCDUz
D54u5nd8fpzbBgRxy4WgsAq3KR3ZtO4XkfP7qJtYzSRCwA0xX1zq6kzia8fSXB06sRR7lg5L3HrA
LM08yiY4Ls34yX9/C514n05OJvI2HqT/j+sDYVzzH40Yu5yMud7UGQU2pxYL62COU1BWcjAeZdgg
uvYFdJfXknAUOSA1/1m5nYIGjtXfixvYTjytfK5S50WLKnTc8Wb5hn1VI9KMGgIuZpIKokjkBIb+
zh7Y616JHNnHSon0mXIvLo7vS6TC6pf6vfC/FKeWoQ4LQE2WZLIHWW4j8gACs5Pdgup8LGgHq/t5
kxwWRD54seUTnw3kYPAul9JOwBUzFYSi6bLWFwAxdO7fFoFzuEOie2E8g+2Pj0JPDLHg/pFAPrMs
4bZI9w33RC5HAEpITzk2p5J/w9tNg+qYhhMFkk9+HMBT3Zm6j+Zx22LvuIqzIBb+xd03fwwZ81oQ
566WUWgjbr0dq8bKpoFWxmQQirIZBvPoY70gHpecUA/8JNRQkaXAEeZhephP5aGVGVDlKch050SK
sas474CSt+1GmUJrH/uLWxDcLm8e/f3wb5J5RU667YWmWP7HSRzXmm3JL1rGYE8PkwKMtmgRsSWb
qjpn8saHkqvBbUkvF+r9xOf9FKP3mIxkzEt1PXiBl/0KHRL9KlxsDPWKA5Ss8wJT7sQGngFRXj5Q
FkNYnOFTmaCvRTaW8mp3CDTk6P5IqtEPPZZw9o++DSV/1n4UT/8CMP4W5/XptQYz9EqV/GdJL+qZ
PWki/h6BS1N+WYsFOcRy0sjjaQK70hR7AsYiHWRkTrCpQP+uvjBT/2ocZ0JfWs2T1nx4ZS8TNy53
e12brwlaVI3hoRalNVwx2xVwe23/KidyVndcdnzH02HNwx5Y7yXewruz4U8q8/y+x1N4D/mHnBhJ
mT5Us9k9pNq5JPO37rQCBWBwnptn7jsMl7/tjS+ywiO/e1MMX4ohf5FXgU0Nj0yVaiQIqyY+mOBo
ZS/NFMirFb2kZyCatBPwlGDibC8zKQOu7tqrnjx5Q8nz1tGMfEmLLsbcYUftXWzp8x3XmNWuNb+o
32MlKC8PNaL9Jhx29PWpS8N5U9SE+b4NdmhhXDqNUzgo7TBsu+uc0DmnkOc+CcJW2gv1ml7ItPaR
jdAsKDXNgMxB6qRI+Tq8wOkWDaksHelyRJnPiTKD4u37NZBqQ1ki/UD3UOQ37ChuGJ/w2NvlrM/3
eAx3H9gesvDT2/wlQVWX9T0zRiI8h+rYzozGHr5l2ouz3CxaP9DAn+igdf4ivrzdbAR4xHrVH/4s
0kR+QzJZg7Zgp0DxYMO57qX9HaLgJJYjtU8OaL8GRTtJAknDyma3WOt9Oh3GsLzRxM4ALdIc+sUr
zEkCebGXyjMFEQPfoyPPU8HXKlM3M4y5GsOuz7D8dBuO6rd/Y5rvtZ5pYY5uAsfHOThJ8C6barC9
1MyWGsugWsPOaAx4uJDqbMewj9T3wRP4PqWzusisDfY4XAWGmM+q3XlWeF7r/y4WVJGiCVzDBCfL
6KT3g8DRfMbFxnwHfYHX/6TRVfGff181Aj5OqaxeJRItO7W1VAvc0aFVCs1fDKoZgSBW5JwF7ZEf
KG5M9ZkHOfyBXhud7rSocPGSepMV/hPVlAaJENTVtWNm2L+o5nXJoRUWIfnjK4hc1a2H5lsWrsTD
vGl5yn13B1j9C5APEnBttdyR0qP9DxoY6yGtc1eAuzg4fQmw2f2sXbFAFqxUuroTWpgQeZqMM7PQ
Bh6lpzocZk8paiJXdkA+3/THwMq533QQwXV/SivKeYwUgetzxzDKpt9O89YTT4rE06e/Q9Sd60pR
HSzcGNPEe0CSw6GNh0ubczpK5sgKQmguGCdmFbzE+arGOZiCWMy7p4YUFHhHDmLEam8oa3D+faUB
+mVnvTSvWJMpHOloZlYDh889Y5ufQKk9DyXeT1ij6NonTSrr4jifud9DdndodZIXQW/oYSiyL/RT
ILaeXaf0X9vRkgM/jalWGZBXT7vUIgAzckh+FGqoy8qiySVJPwjTwZsIVQ1R85cjLWjgdYtzMeQZ
q/+95st9CrYwbAEx2deUlD10m2nhgu0uRIhSXGl2/nv+CEeYgqmjHe8A6pF9j27ZS/FbSsm9JK8P
iSi/oqqkLtJKlmbXJqfkJuKzxVX9esNDvU7PzE4wFHugRId21k4mV/SmCw9R1C0R8JFzGiH2NYMY
NW2KKrBEJwTQ80zqMSlnX9PkCPrLESG+n42JUiaMLZQjjPUxfrTpn8TnlNFiynxqY58Nfm2iv/D6
frAbCMXvMJwmKqDJMJv/cf7wZOutdoJ1G9V1DU40nKLqIQfbNxeGtuMDxBR60e0S93bu5UpC9OGy
LzA1MOQPfBCZtIxW8N3QJTepul1C5VnhwcwUijrBkTs24oXb9iuLTqnwwJyUFgfftlP90ggqKn32
5V38rkfg6dTv8zoci8v2NaP/mndH4r2Vn1gu19rPIFiqzjlyc4ZUTLtPj5ydqXtwdtuduzh1jsgN
JXWAE5i9KbpiUhxtXVJhgokCx8croDLYB/x12JzgBUDN73e1eInvfEvRfmXEP+YzDqi2rWIHDCWu
PxZ1oeLSGJnipS/0cXWt3KpKlDaCWGBM3KwwPVDJMlhC8nKZ9bFgXhrJ25vDLeRmjjIbzJTdWoT0
dDpdadG/CbT7R82InD2+gB6/D3dECXEQ24852dn4UV9BXmAj2nxzILh9UUYjj93ESy9uWFsKcuvn
/5y2MB+DRJlsg0XfVZ4SR30U73wXeeyGQB871EcjayiD+qu5zZf0VYVy2rKjoC4oNJIQabDLgJFy
ukXTUds7o9uHJA8vRfzSCNoykcfdCR/M/48gqwh6e37H9xfJnOKdgEqdPuSKPgyWVQU9pKc43kNB
Wf+EV2JS76WwP0f41GpD3N06VNIRWe+MkY5uCBOVeEZvepgB89hyuopx0ViRYjxgF0e4IIRxLnWK
t16yWIpVtaGlHkYtFBas6OUxX3vFNi8cWvmCbWIuK9UmmBaZK1L9zj6gFUHfE5/npNwOmtaLFB8B
InffRpqyu4DOPXhbTwtncaFOcYXpulemrq1a8jQ1kUSYASSrZtH5IrUQeZtXsVYXYuiyfA6JM6t4
b1M6wj8R/xCE+u47dPYuDnoR2JeHdsI9wiKuTJNfeHFdcGSLtTPRpacr4mKpdIdazqaIlxfUZtc7
mayvwBh+xAJX6hNslxgKqnZDBRCaM/0RgTn+9Uyz7zdiFzK/otQ5ZMLNYKoX0SlFHOVNz7ZYSxJ1
jJ+oHeDcZPvdIO3nRKJ14gPqs/0Mu2zQqkFa6/I7SPGhZUMhxRrsism0itJIFgNiVLyYSKV8r57H
EWV3Opdl6vQouO2i5QQIFCThsmzSeUMIWR3th81jFwceBSCVsCT84HL07D0Jevp1vWNUMM1yNmy1
odo3RizU2/BvWG1aK4KX1ET/YhhlxvfAu9OZ9kXONmu8tsIoKKSyQqbmp9i9ggp7JoQvkF0MYQRM
9d/VY+hvU/peDLPrF+swCzJBzMmYYP3X3AQ3rDwtzNlOPbkqhctX2N5BmmMhE718lYjeiwWHhF38
eCOG7gbonVshCSBrlQf4xkaDX7rB/wzWYmDLxR4EfLKizRmMd/YVnp5YI6quAftc7SAJxzR7avQ9
EhQw9GTL8CfVHzomUWDQ5psEvM37lE5gjSnIP+ZnBGeCDFr6oDJubALXUNj45armXCfBNRidffxA
pfFXaCARljjXiy4xfYLW4V/eVgwTXxMjnRrk/KRUH9Uvymsg6PlFmait0cX8tFIqiMDEnZG8Y2SC
KhsGoC66DXSI7z7OZU7UsZH8xCZYwQng5SjW4DV6kNYJijrmArQB/Kix5pTepxUI3z18YB7ngt9d
CyId6vXg3K+Q1uNF4n4Fsik/gm+/f/vdPhFamxu/kwBvov2vJ4X39+kEF5eREnkb/aOzTaRlxpv+
OHgNKMpKLRD8bGfy7AV1Npli2aBu7n2CgiN8cOml7TYIvGMTPGHTMbONoAonL4Aq35QNNxMZ6wAU
gLWRvUuQguO7lhY24ZS0RLUo1hUfkrKAzz006P0bKpBnB2qtzG69eZKUm+5ZvFGEexo10vHi1NmG
y/yoZtVs3je7rh7tylHmbjvxQRHyHy228R6oNLYn23LblNQ7qKmrLh2puqdcScnomvkDirvHvkBI
y2d5gSGGnVVHUVTsjEAnHJ8lbNrYsEieSrFscQCg4QGD9LL4c1IiitLwvDDEJwi4Cjj5/5s+ZsXi
0DuJQOLrGYx7ck9T1DOtrTVtaPLAJ/TcqHtet3QWd92We88u1OP8MMb7rtxVXY4jJHKI96UHySzR
PtGPAyGZOCqUz15dnt+obIzVKjI2nB5lbt+QZ1WXHmcTmKa2z2+zcMZvHGqTRt2h9sxnRVPo4nYQ
VQWOuJla+vm6P63728HOfi1ypVsUy8OxkSKpMMvDrGk3U58SRGUpPUx1/4/YaK1771zn0YK1fmPa
uPLkxbZUdqa6ykjnFu3guzzlPOevw0Bp/I2cvk51esnoXaADEbYmOg1IJgoSzQYB70/KsovZFues
NAFpcCjCS4Lu/4l2lq8mcKNGHUEyjXf6B3/xZCnLVZzI6z477I27wu+y9N5zIsa78cT1MUqc5s6e
KITON/8iHLKKQqInAJiP7c1xlys1Ol1UuuB0zpg123JgMqNLmiaZHn9APg6ShjUMvx2Va2CdrxHL
7tiCTdYSBZ674A96OxU3VQjUf9vBsTRyHD7qO7WGyIRFmrS0mCt8iFDjpA9/ijMfEHqzFfL3wf22
TSRgTurd6/UP2DFiE5J80/myiNbZaxukbCGIsrH5OgsvoXhzv+8VadM4Be4QGbtQseMuzRuTjJJ4
GOWGHMJsh0sgRKbyOgjsHPmsIZWUrMc9H9WqMoWCv8b7krQFK36uckiPsf8wARsjtLldDw1Txnwh
1qu3Vs7li+JxDpmLxF+uVByLQbwFnvKnqsigVKEvvWm7Ey7u799kpcqwyfPx/IBBjlIMWkFNyJgt
ZmAgNKiIFd9LTI4F5ciMziSE4iXC2DP/UpnhFHB6R78Mgjkx5SJ6KEgkv1exaUC3Js3Uof/xpK0Z
4o2c+36zgX3HBU0tnkaAQ7Jk+PWc0yBk1kyZY3WcLpk0vdv6wq+cywVd14jXvZ1G5feEpQKhhb4j
mjBOb7yUn9OxigJ9LBSzk8HaW1bWGJA4xIjwXdcXPM3YBCPGrKAyhBaWeda7O18ARdDYwUbEeNXh
OxieHvF6xfCoG8QxRGvqgpDzxqKAUdPZ38ITnDgqVBlU6m+jdGPHmnhrPgRkPeQJV1lYWO/I//cu
qhFGK8Tqfotoe5pRFaAMRDJp4QNpylGhgbiVwJ9EjDiBSsakaV5yC9G3fF+SY0iykKP6+8YuzudZ
WzH6achwag6unU96/QjJtkE5sLAYjjVytAXau2NvjhLg+1DK2jxYpZ974Y+WRSAqTfO5XZVzNJb9
ojAsFopeySIGdLwoduEqz5Po9AmC4kVNJhaYbn2zsfG4rZ09fKnGa2B+vbRqTpf0h1eP7vxh9fEA
d6KPw7FiRQ+8AYcEK5x25giqnERvp3aLjd2/IKyEXvoMqcmCSnVG92EiCHgW/q+wrSHv+x+cSbZA
rFCyEHM0XQhmY0ykjDsw6HlDY6cLRQsqXXHuQZInxPiS2V9zN1Nr3+hVPl9CejmEE+X3Zq5hV5BP
s+ATGk9rYLlbgPCL17/ni//2pBKFZdJnjpOm4IphmUG2H1/fbB4/ppLvsXRwQHMSNZ8yn+XBMS8U
K2k4pjfjPBwG3T1GKwqPnC1gM7nBge3w3a+K3XdGRUZdPixXjimeXCrIMRs3A6QJwe2U/Zj1DBtV
XluXWEo/7HJeqGIWHVv4DXGljPS1++NKJ6rUtIXiIqUxOx6ilcCiJ7zZEg9a8dgQDdyss1iH4gBv
rUdbETJ1RG8yZ0tSFgFXKFB3ZbonCdO0/LDMxiUv/jO3eCsSMoMfgYUqrN1qIerVGvYCAAIptjrv
7hlVxLCis5uB7LXaIxIX+edPFY7WlBNPgzsp1I1TI7pSRZCKEkNa2AX+CPXLAi3fus+pSZJMqVK/
Pi4HVODdFgYXXtmC73fP27YxNOu3x22kDZjsUwWEJp6I+8upiawtOOgqL7FX22ia7wOQN3nph55D
0xU02un6M0LyS1e5Jn4lMXEpgr+n1bW218W3AZW2zUzarqxQosmxEfk2JfI03H9EO0PlaoHryJPG
g1VQsivH70so+7v3vjgqV1WR0yDF8B6kFPk3MzsaQDTuNLOYHiLHBGLxWCOWqPxi53k72J2WKvPd
60OsOmtKwXYpkkXqC3rhZXixJxnL7Y0AP3OBfoXxnTL5JXpaVLKFdagA3dI4puYdb9u8phoXKzaY
zO4/SVOjHXsE8SZ1CxCKYiUBfPmdBHI03i7m05ijOsBZ27b24rn4cPaULpY4dz3pdsp1Lkk0XmkX
DVu12oIGfVZonhjr32R0FGsJL2M6RQiA/j/64urS7OPqoYrZq2lugy24RSGi3ffEhr8dEXjpuZL2
Z6fXhZM1Hl4JLcxX14HL00rTNnFyaHbn1pQ2GcRRwfO4lvz3Aj7y2v+QDXgo/a04pW8kOx9PCtJi
PnTyCLZ82jaZ8wlyYOqZhYlZHrwH+joXGSocx3b8aCLDHXPJBqDe6by8IfdwrWWsnTNRPT5rk8ec
GAyp9FDAaG1uT4kVuzIcVFSXAs7HqfFhpaWffh5gFqBu09wqIqezRfwmEFvCFv2w4zAXmbOMLKO6
oqwVxEJ2rwp3XvYZ3DmImTbIZ3TyEC0XshZxeTqT+FDVhMOGzhRkiOgZag2p4GI98wOluOlfsUYt
b8E4rItfWh3EJUKUb9WgWe1fUxRlOP6pJEhAmfSUyXMBbejpLH89lX3OZP96IA43yO31zxNamZCr
JvuTez+81NSwq+PvTeFfnuUNLW/5rK9LuCAsjk3t5Jglcb5N16CU+xLntK9kQzcTJZhKX5rL5kfb
o0F/K9HLjvxOXcz9Keuo3iEGe3YiDwO3cmrYIGQNd2VkyPD6sT9PyCDD3NfDjT+T6IxaRQDYC5tE
NgrySw14IUs/Ox2g+BQtZsLciMiMsZYyXbhpDzOB7aVWuOrhIQn9h3aDU3mev0es4ER0ayU1J1Qu
bM9HdBmJL3BjYolRqAOI1te/jfg9q+AmRMm+gFjy+9sObg5QLvUMy5j3Ff+IGzqa+1PWGqITCf5V
9KAIcWwJD9TVgblo/rPfpei5/e+KfrGXfR+RW8N+4KiLJYcN8jUnkSmAJ4995sbzgM7ZqCiI+v1j
5ufw5KmQyN0HmitGqBwLewZQNJX8MLDsi7zrNKOZY2z/r9SZ9hxfWwBseMxb2qvwR0WcskBBQfqB
d1SNJsK6qBp8kdjXcp4CjNNf3q5x7xokJhKcc5fn3RAa+/UHy1HOiX2AMHAzuVT6tGxt/k7LaQ1J
lXibAVKWc0LM3cOM9ghp1av4yvMW3a1nSuVXM4Jy0ZygBe2FnvwbZjqP59uOLJlfpOIOt5kIuCrq
k8MM4oHEZH/2CZlbxazPKjtuQBBMKgpEIiJn+rdXE90kNCzwtkzwQlEn3HG1r+EQ/NGvO92UaI1/
TlVB9yt6qo/8hXCWar9XDGmavZb4WGPNy82L73ao50wBu+8YEXrNwdXer/Pj99dUBGHarIb0ydR3
I8FUmg8ipTPTgPwE0Boq/3AodPDdTBOxOpL90Bb3xbJjyi19qq6qjOJE9cET1JtNdL3y/PJvTzEu
/sigxo24Y6fSTHD3Bi2+lNbfDpvm2DNlpmmpizjr0nsaT8adPdqoq8XjztrpaerE3LW+vj0C1Www
d+8H+NdfPrNLkHtf95F9UYjE0hNp2J21GHmgrsqGDc0bi75m0NwPYvVU7zJ8fKMSH7ixE6wnuuYf
bREMdCGyFq5YXEMcrqMTiy+tGlCeDX5L2ohxp/8QaiEe2iaue6+p0jXhB2kpVIXf7grpHUDnv+Ga
/Hl13CoJPXxxHRZX80nzZ/qSSN5WFEWrmtftL23A4wkbL7BYsVhSnayFMk7r/jfpmnqrIYaXCa8z
vqEYfSCllPAqIN7mN4NU6eAvrWTRQCD0zfa6cmxVw99AF87lxSnINBYSLbKStHXRIZPECUCE8ypQ
1kfOuLlM8VoYr13umLAwu2RxDQf2URHz6UW4hU0hFJXlgln+btUHWi6GL3Q9O3uZWyyJTzsrBcoA
pfjW4z5YIeiLmZbhCEUF4qKCW9szkvJi7P8pOAfjhxOfg9+EAOMEkDthMZTS/jS798fa73Iqdh9U
nKsNrI2HKGEtvB+Q8zeLCbp7RCUumfME67f6/nQ29Q53kIGgd02tSszJOT2511ZW5AgpekIVbVA/
Z5ZJ4B7THTl1h5NAVF4U+MZY5k4JmQcR42hxn2hi5zP9dC9GojjCniCpHW+vhZ4o0atQWdIAq0a1
9bt/X1PCbH899IVhNE77ewtOvfEaGQD5An0Qnc3GQs+vtgoBH9nQd1N60c6ueo6XDOxZaGdcpKXd
j1Kh94ecddEjI8/IcsbWT5fzB2IxxXD6ddVhAbgE+DyteT0RkA5X//A53QNcAewksdyEHd9MyosF
FkYH6MAkVYFkB/c8ZTRDKS1rg75eYdHZErcRXBnmYdjzpLD3Obje22JePgWBCF4lvLFIJUPzyx3d
9qmVQi4LgFwO1eiHfUDVwZIpfxT5lAy7GbTeHb6/qhafEX6UDmI73uYb0/Qfb0aTHecYpi3PpeQz
0VxIJGaOgOifrALac0Ek+djmtOnta8iTR+YaCUN9Oc3+A6DR/YtBwMSa6uWCqSUa5SnyZ9K7XARv
K4xbf2cr+U96a+if507HdoZyr8++3UfukDBk8CwiemyBEzo1sTlZOUjpSCOntB/7wMqSjg4tXZgd
gfN4fZ2UX/oRrWjqY29LuNqd/JAqzS6tR3UrNcb7zvFaNtq0A0xaDlxCjDKeaJHB8z+zEdPjp+Xa
FRaIVRBzvdTnsPT9JjC/GlxQNu0OlTql9cRPLMHUtpw37PmwLQ+Nk6IheaubsMNbnkMLOZBOuKaz
0Zi+C1Ii71omS10d26XGIphYUYwucMMDv3ZD8ur0GIWO7Y1cbZTZMjtzlyehuA089vAI4KNeTVxZ
EJotM2aLWcbUYxuG9ybaphlWuK12SMG3Hw/6iKqnHvGIKuW90RCw80NFnTbVDcVd5ca6iySGRLZh
A7krmONwnMztOBT0ukVMiCDq98GJC+yKXM7U6FSUI9q189MB47kKevoq5WVpbXM22vJf7u2XiB6C
JGxHWHzrl4D9A4GkGY2NhsrGebIfLG6SWOHNanSQH8NvXDlGfdbqqMHwvG7b/1984fUvDchzJrTe
X7nK67TD4cI6MAdusNives95O8b9ZEbjyqvp3sYI29ttGNtWhIsM/ye/EfMbhO8Lf0mNgxmJCJ32
Ts3qCsFBv9GyAySo5vJ9La414RSdfzXkvAGCrk/6n/msM3x5JRKRC+aEdmjzR6jMPi6YPgTE/5pr
Wo5sK3QGrTs4A3YdmtCur4K0xCQ/6gPmrHMOZDzG73nkLKjYjjF+NrrXU9IDhCj2mCbs6Za1a0bQ
a3eUDdIhOtDYfp5RxN86XOVumHb8OZ1MAARCrIpDjLoNh6Ai2xl2/sbV2q65+s0oLtG7GdR4CDzA
GjCjLD9lCdnkifPIyo/2mHlnPpJPoCT5j9XSMArF7yC35FCTwX9Wo3b/5Bjyb5iFoLcOFYnQxTAw
vJc2YxaJZZHG4foX6wAVyKer7JMP8gpnzN1ZxnyA4jlWuUCZAA6JhKLs0Jm//v3wgDvujZrX+WDM
bKP7T0rO1JD31uaEEYO7VVDiOC8IvnOoFG6FjbEOoT5k/CPJbLHfKKhIpM8DK2xwX8asWXw/hjX9
CQQ84nJ9aj9qVExS4L+HUsCgiVTnLIj9FZBF2rQPvP7WQcE0W6aM2jMZLIutymiGdpZ3ldQelMVC
rXcYWYcHXBdnplfStPxLHwdkE2x/rudxJYS+6wIkEpggZiFPvwAQn1JR/hnfuXEXvI7FIFl/KPXv
ILmoDSEYvFqpSQ53Xf6CLhail6tp2e9rc+luYXC42D346gb2Y9PwJ1/W2LQmF24CSb223uEK4jGq
ifXXNq11vrODCYgBideJbkW2vCTiISaXkMfF5/dreE+kHLh3SnrK7bK/TJ5Ii9EaBmxKKR+vBQLk
YAnytbeeHhT7+FHdieTTJIK7izns0PHuFmfX19xja50rShIwuz6UTjYOUEKvbAnD6+DJCSDITes9
suzJnDM51g8GY3zy+xFSJWKiTBKURIjoxdEX5qy98WGR1dImTb+tqVsTfIN0bu8tIaWnhv+F2Qxf
e0lp670FV2LaUUD46kkqmAvjgEhM0Bi6JQLblAEAn4CXBKadawA89GUSeKpuIcw5bTRWScrsvPnY
r0D8Jf8P9e8APPFa6OwSBVls2vtrCpL2XYCb+MKu4FxGqqZqnU/CGRJG1D7AvYy9zD0X3zRvBWFk
FFsswN4hsAbFRcvs3nkg8eBw3C0RlbNRRrwBrsPpHNAB6AtHFyd7hvPOLfcSu7a8wv6DAEsEZa+a
M1UDQYLBbE9lloS4M38Tc+ltKJbXlw3UHPfUCt3rLez/gnTGoAnSqtdV+GpOrQJ5rS3bagcABYzE
24gxn+7bhVvDke+Z4B9jyv4PkZd7cfaJV0bKBa/aJPzh+MzMlHsCNUnFHmHWZx/bOmeYiATxG8i/
1vBv8O+h+OOm4R7uNTr1QKfmp0c/7m9odNLbeAHoY5RJe64FgLbBh7eiUlQn4B+n5v0k54mvtNrd
PTqnjgPNVfUXmGfq3y9WykZW3No2vjvlJ3kg9ZeFvqag6Yy7TnSvvoaivaDgeamHZ+FHwh0uE2zc
iJYIX9PWkrZFHvA05KV8cD289EaFm2l24C6gnloXvJly6WdAvg62zT/E+TtjrWSdd50fWAs0fZ6V
K1e8JsEWe0v2p4Q62eQfDQ/GImFyJQN5LTTTkcjaxqjCVoIO24VpTjUz+tA5N+VKJ8JaZsB+5t1J
OjSe7CiLTX3GrFn81303Yy+AbePj6agzxg+X+dbRpq0i5LS5ppvwgfA+yueG6a36EBUZC8H5eu/C
1jNZ0OinPErhUoeeHfzVsHa7j8ooclAi/md66nt8Xp6FRr3TbyCrMbdodbfpJVmX6YlovwH0NOnV
xsyI10GYWKUfo/OMGZPh6F1F7TS/6d7jjqKKCU5I+f0gvisu4zmvn+JA4ZzjD5WkUrZAsex/M76k
TyClqnkgAEuSD8SadI6u6K21Z533TJWwLGu8M1uK7CFwYR+2w8QFgV26F675whf4eo5rguTOGOnV
mnAVEdmbq1ECBsqQ98G9a6v7+f/dR8HfDpl3nxAo/Atx3TLGOiOHVHx4OzSq9H2BvQi8YA5aCg3r
Vk6BxhhvZwJEGgPfmuPBdioLjKEn5O6hAYie7ZwUYvdFOpbppOnkQJVq/+M7G4iaTRQGweTJ6f6o
KgmJvNHkC3kQuCfz7BZHvCOZJd8OZz5w9RpvRzdAvjNkn+SZnNCKjBtmmfXkb35GztGxlyLaSr6E
mEI4gwBDmTHDdlDT26p0uXRJaTHfnd6EfzKrthSaedHTUVqUBi1JRCQ2B6P+Ql0ZRWwLk//SOYMc
O1jK1rlNcNKoOeJyxSkZ6wakSZ7Ak0ZXk6zQyvNIj0siszGJk+QbwWj0pDAfQJmUietqwSjyh4Rm
dPZ8qKa46xd0bjK3Mk1wbzApWZB8I5U1gI4R0qZYcQfmBuP8dHAyxRoxwNEqZ6uYxVfJZjTAFApn
C0w+iNsePFv0oPEUHD8wjPHQ5OPxQuzCHP3FuTYg/RaJkQI9V+FIuLkxHsN9x6GXWOzgUQFw/fah
zlr/2B+7me65snrxNpYsMWcC7o/iikttDUE4FBUJB6vdJUrMhESeaahdd6JlFIiFHB0ztHIxM/eX
H1u+aYqPGZRyE9nfITT6tRXDKl7nSAgI9YnfqoOiARm0CzCNuNONVFn1AWM5W2NEsHKmzGVn16dN
e6EpnItWmOzXCmfBx65OLhwGqi2RXak1jrXy2ueq7B9y95QPj40e5OzRREf6WhJu26Al8nZkkzQC
x1cM7KW/anCU2rCkew9xKbawL8o2ltYprwzDiUKhh2RWxWcEKCjHCsaSJg8mqaCvOdthR/dX6/L+
5YZn4/KdV1QQ6tIp7rwPPYRzOtPbTqm69nhXyh8CIaXqlSAi9ohKESiyHGfXtD8jF6XW/U5Ep/4s
Qyz+DYyHbbkt75np4Tn9xdOLDNyVf5YW30KCYpwh0f5ZJp1l3xJJ1v564KngY6nDMT8SU/agMbbD
EJ87nsMNJMLt2/0UYL7D15049UzlBNoENveJQmIyvX0inVA9MI9c2MQtgKxEFrw360SdObNlth6y
hk+7yp8yQFirBRdxdZB6sciZyn+FwsMx2t1AR/JxfgMNt0pHK6IDKS7KRh+ZRbdDvHdqrJ0aKBbR
iJkoZhgzyRGHobttt+sRNiPg9YBqy+39cZTPUkKSRjHhaEBCnz5DSEqYFyVNhoJIhHAxWRn4hgr8
zhic/yA4UlQoDQv/Ksp8IWJeil6P1k90pOCa1UPB2OsmN71it9+vaHJDRlreogHZzlzdXhrhQJFA
f5pDP7zr1p/zu9dBQetvIXTp6CPTU8D/uVa1BVEpEPNYSl7kYmjygkUBh4zTWx0sxlYD8xoWk0DC
TvsigSnKWJiCTMv9y3zFBIfzexcKkG6MlZFvPe68w2mOIEybOziIVISkOq0bPBL4M6D2brdVi9zW
LKgjNF9lQdmBHJHWf0NvVYIsLrc36C1Im1Vp+uhicWnG+zN7CLM0jZY2+rJXG41zNqt2bew3T7CB
aV+lnuESmzfG9DRkwe/eitgtG3UoQ/2fbzpBGwy4G1IReg9Td3tp5owh5v8vATOsl7eNfyp3vgRI
jkGwR5ok1yF1siixoR47vXsIddrB6EBQY7C2PeTFw8CMnUbaSLsk7hOQfj+uY8CExs7IXXvdgVRy
qiiwQQV+vYZwxhlM6yDlaHTEpBd4c7BvlnjlMVMGg/bz3pP21GYsEn8y7+iZl5cQPlqpuuSdDK+n
GHUu3QnhBAAbJr3TT/IO5s2/hUH1mc/VkrzVsgJ4kCxa9vtCi8ECulQe4cTlDkUSXBusum8MDHai
+Kh/FM0QYgdZdAfUzfMyaVuubXnTjSMmw+OW2/wODgjweHbcHURkvnptfsGE6GDrCwuksec3JijN
UmrgduDfLyZEApkz2H4zZi9BClLZ7y+OAYCU+8hCptmPxgAN74oK0QfSuJoImg1UPRi/8Pxz+h/j
rIHM/zPhdBYgcyPMlK1ZZ47JTi1aoRMbCZgG8X7aSLOWqkzi9QFfWJRvBlOKXUvf9GzcWy1X3R7U
QJePFYnLhvT8fkixIu8Xps1UXbjHNgeiKCBeyB+Z/k7ueCVwoYx1ljFkIaR8vln+Xn2yaOhQAPcx
CnCLmAfIcD+NuCvLLAGt4daEFFPbGEQHRgTaTqqwEDaLKckY9LVLGEAji3V0fsPvWqDywtwWyawE
cmaX43XDot79KxU8WVD1WtB8aFfxuh6xWe/9210+xeZzap3bBiM9aMLzhHMB3a3nFXeocfEZ7JSP
CpYTXEHGEtiE33TS07sExLWzb5i7uC3aBG3xXvJ7U1u0Y+RK/zxpkIea1Tfg7c5c2bejqdmlIckR
M613pIUT9pRNf78zXyYAHMnhSsAQ7cxHBQmLSd/X6xCAj+CDEx/EiZQnrRpXp5wiCxtrQR7ZAPJ4
RFhqnV/RZg0K4c+Scmbn47P/S1VnPhISsBuflkWcQ8Z7CAvMxQ0EKZDaW7aIqdbCZe0jwBfunwjO
6zixMWXAFAa2BSqGF+e2vTwDvK55CbUC+jutJC0EuekoV0QiBRyWyBgMdxRgR5sIZiop4xzAHIba
hvAsfzALZmUOCXQAld5UDJvZ4CkvtNMqZcX+R0jAEO8i+nlxtiIbT4x+o6NLqCrYLa5m7QQLfDzv
xwEfthOxHExhTF6Kp9QhfKwD/6NOlXBnQWSN8sKvP/42I8G46uL/nBOduRkyzTJRxjJkGhpQRO7+
s4emr5JP4fNu7NMtxoEhpQdFxJfBD4ga84gbZfFQokDBa9G2Ff39oZIQ3BqPBCYHa2Owha+wfQAq
sYJENjggRgZ7fKS4CBQzD6404rfvv7z2vvGMRYUpcPcwZn4n/CRLQBq7KTMZ8nW0N8xcrM7zeLM1
iTP0kSZguZTmV2dWuytH9r7n6oB6TH3asV/Z0kwVOfzYKGyRJdudAbG/qcMd3Dd6hCESM+9WGG7e
2PQTc9IBRIDcszFnwa9fGhUNK/J3fCIdw29kNu/f7HZQk2K7PelEzaFNB/igFCiGWUHCL93ixa4+
O0v/QSwyAK63F1uR75vxnzjmojtczMQ5o5MFyaBygklrgwKnGy7WTnFsIlMM18S3B+hdV8IBolN5
WCmCT8c06bxg8QJMii/gSoztVDxNi6rSIzym3N5jjT6kiHRZqmi6C6/qio2LT8kzhmZGjB3BiNlp
S/rXgOESBSp8SZgYAfO6YjFzTtD6Y2f5EiIy9YidL7QWKfXGpoPeklvGZqtpjqq3c2XCX4xoxc3G
VzTZQMr3KxrhuxLhUzQGTngJVGzGMgt3Te9UI5FF3tm79/MVWfxTshHvKuyYcMqH4uQVipq69/7u
fjWcGWRm+gU7PLIml3LcQA+iEysRHrK8jXucexN9nxyOn2mpyqIxNkDPaZWFUJHG4bPX5AY19iKD
SXSscQJB8JOpZb/QTPpgfzF6MhQNx2cK9s/sURkQKVjfwz3QQ7SWNVHvpAYzOh969GkOhs7UW9JE
ElrDXnHMaKs2uxvFnZfPyS0Y1gzEAesrGitrn7yXREDU2BklQi4r8+g2O4jMrsXa7P+yDk+9ZdPN
W2+qnjEcQaH0wAReTzZuos2PHdvjD1a7BzGMcLjShip0RcCJoYgkoE/+FrtkgDOYTvZcZWZMZk5m
9xohSyv1Xh2ZLZFgQ1YwJzOOpznOehY7jpqO6NOKLrv2j1Qm/xitrRfObyGkONeSGmzzpwo1goPp
9L49WyA71MGr6Baqcvn6gTKMEn/2HnLHAz23o3q4Kn67kj22rO3U0tM//qihF1VwR0M3mOCmPQh6
EZR38H131M+W0hy7Le3/I13vbODcaOFuzBS5ucnKudtb+94r6eapus89BcSX137OcWYAH7LaRuPl
oGKYIKp+lXRUaJhvVf6x1rTq66AkVBc1sAvm2id94U+L7Vcf75twDCNYgR6x6pK67MG8msS2ZEDG
1Vu1Cv/2ftLTQds9OzTfOU0q2z8s0Yk2MLgFp84/sLeU/Zs3wRvtpTUMCpEm7RXBU9X8BDDg8yqR
M7nGj7ef+Oha942jF+w2qehL1l77teMn5UPDmTroPfUrekTU6+Kg9OYEt0irwQ6C3KqPQbCYZ9MV
nBDvV6lVfZWCsdJLTspPMVqtLUvgmQk9xxyin4GsbfRcBNyeT6Ta5KGR9nQsLi6cWg+8N9GIesie
Dfkz0vwibTYajfUzZDL7hDuL7ygrDkZTiBBW+oyeIi1wfn3QxTUIZdYOzDsAA/5NcBsDkyoPL3Ku
ygHEvMS+zZq0dRjfkPJXamQaNldBm0CDonUMFSabkQrdibfKL7d9Kv2uepnwSC/ShoHcWFrxDuev
D80/n77q9BsTA6HLezWXhNU5Jr99lfi+J1dOeh931UQd+d6GWySxIHoJOtPYYvIFtPJhRQzqhc2S
h8PsxY6M5xvm4Pm9EFWiuvjHuT6oJdpIZGF+O7KiDCj0+1ZkzezGWPrrOIomKYKkdA2xQD+05bVX
kvYWuQfHkkoz5j1Mp/OGfqMnS70y8Gq6DHDhOaTySZJMi2TpoYUl2ItTAmbaJwSPTcJ0kfkcdxs5
01yd5VbAcQTOpTpvWLaeiqLhrCQjnXlj4HNXdZ4v43piawKkb5FokBAn1NEha3K5kZ7Gj69hNdkb
W6B8uPrBibsLED1QAHo1lQo4SOTUUZunkqaRRMo0d59Rn4aNX9mX3MG/75PVa20nELvYAQ2LqtN6
eNLvQl0UBRc7QB1MEkGKj5uOBDE+Ku7yasxO3vmJZuqqga/QhbBnjV/l0ZDqzq+Q1xKn14YYvXI1
L7e4v/nMyo5n7vHMWvz5NRY0yV0FDKwZslPIkdFpJo579FgrXAuYCZWhBCyRlZBeFxyNG/0p3L5C
u94JtkLinkqkFPrY5TC4cAANu5uQN607Dime9ywmTAecxeCs1wh89uDZTkpP9TuJNYZ0FReqvdoe
e1MK2PnrfAS7wuBa0q+9zQL1wvLzU/yNZg2cyNiiZnyuFFT7u8Tx8w9lkOoW9a5LxiU85rR81U2u
VZ1D+RaOPkyjBdCOx0W0bDAkzm4T4cjRuLLHt/irlGGKXpmRzYHSDC0Z1Zvv25eTha19/gMC7gpF
MLex6sTm0qzNDSX15cxAn5abFahCZOIdTSoNIQw/O50CeqA1i/DkPyRGT+BeM/n2GIoNd3ziJ3hl
6rVrrKTOwquZYVJBbRXAV1PdAAO5jvHeWw6wM3dOINJDgcqC+b84LiaZ+o0kCcOnv7QuQyYpSwkl
UsJ17kvN1Khneqb1OEUT2cCb54WIeoG/CErK6D739zxd2k3LONJYu/glkFynieCQUPH1GRrJ1W0z
pe39nL6RCes/2k4F4UD8h3nYgEkHhn2bLhBipVWTkWWqDiv+QunhVDLJ8sIqb2aJxfiZyRVsCqNj
c3u4fG8AsZevfckWKh6DsgJS3sNYvdZGr/SN166f92U3Y/XcMx4x7dEZzrR+uVrTZj6uhrsY68aw
rOo2h+OFqhw2+MQGUpaw1vwtPpzevYcukN7d4yQtzzWkrgWlsbPe1f0jm5QR+AyY8yO1Q1YUnBAB
A+L3nXviV25MMLQZmcVS/L05t6WEtNA7PQul2J5bfP+UyGzj/4q54ft32V0uGvGgu9wQ/MeYsjJJ
rOqP+JM7xCRN22CoZsml/wdvuXcjr4UczB/G1DYUKk+RW0441lT4ls7ldcxzmsGpL5fwjMhmC6Ua
QSvZ6fXCTWnJ1RbQqi/8Qig8Y6wl1P7Rt9uUkzuXL4fyKNKHezKq/yBHOxRwTX1Q++Uc6fa0z812
wHNXmW0gPtjeHT5wfs25Me/E0mUQkbYWUmlV32Pu5TF0h4QzeADHZUKydPRrhjubl/rZ/wHWKecr
PPIgGOaD88ZJW1QXuMW3/KhmxBh7PzroNnz0+11aL7Xm3kFdsieHTayQNTQDksLEHsMR/HrSeTwp
8BVDx+52gX729Zis/ALMnyeIMV58rcmqyvn08r6CrwU2BR8neBPpnmEYtfAcVwriCZx4u7q8CkV7
9Puvc0R/85VH1nTfxFfwxNxgF9TnDDY88oOzkUjMGtydMBUMwO9LyFou2u4jLW1wutttTYK1vpFQ
qaQ/wPGwpcyjmzBuJDfY34LedKr63rS3odOdAxq+WNwY3+0/l1MRlwmZ4a+ztJyApZBcmEggJ2gG
GuZYdcYl4tMA5jWAYbDZxDDM3wSbqP7lFHtrOPHRIu2jUiMZ5UNesURE9ZnvtoXtavER0v4Up31r
fXol2GF/364dS2ZngZPNpsox0T0Dpf95gvgpYqqnuwld/XH+ILVsj1HkwOFkkL24L8s3bk5k/lPb
xr0aJ4BfHmJ6pb+0rYK82hYSuNAZeq4i/A/uv5t0+XXIXzHNV3h46D9gUbgXhfQKcJEotgadKJFH
NstYna3pyqN8xaecZwQiP9t2YmpC3pMvuMawBw9Z/E7aWua35f2TOi+MFsVuNx5H+PaCle663cq9
ibCLDfx9qyqInHo4qPQ8KZ4MYsY6KKyQy78A/KZEFvmCqpE9+d6uDd4o56+vMQgg7QTAiYNN+Nqb
vLgFWUeTydx0PKBpYOZe8oxwjQ2F85is9VWI6YBLhAFNoy+shmwjZTk5PLQtph8oyUL9yqqFuSkc
eQAAGURVYc0VCp25Vy/qEfLCJ3rJEqUhCKNXmjRK23U+IxcgpNyAw2X0B8gAivKa15O1kzeLigON
ZBI2Wl0z1xYVgORyAznLeJRr2HR27rvp/gFZ+4EqDq4VfGnLYsEq7+igJjExTL1G6ouMYTS8A/H8
LUK9nUs38oBYKKx6/123I2HbMbakvzUC6lgeo7smJhpj7LHNErEDapAmR5U/WiKtKoon9bi/6EyX
eD/82e+FRiob2V99+9PF8HYWHkrXmAGARVeRvKvkuz/k6X63alg8VJtnO+ygZHtjJqo/45PJ+krz
7iawBPiQQn+GuFJn0rWWFTbpTY6lFbCcGMisb0oitLCT0wquyO74ic0oz8BEjrBYi07wCpiNjmiD
J4rkv9bIAxsYOzhcnciEm73b97N3QxwdgMYsUJPyM1zDAIJ3hVXsfbu/H6M3j1w5GKkNaZWCB8Qi
aSNpeUYfEvPxiSBE4GLUC+aHuFwfrUNvaLCSha41/0MNQkbdp8jkajyD3ScS5kBQ0kcRuo/yB83v
Rv4fX9QgMr6365FVk7rfztiUe+D4VvcDCxvtKFPwLzye6o+m+NgG1G2uO6LAxUhVPgc1XYOTniLW
JXfiK37ffDUeVfYhqL7MHX/Jc/6aGNkeA/MPOI6yy336fszE80hpUszWTODG7BiGvrwydCgYseL4
3touMb9EzHTI1CQsc9mEWWVUje8xM27snGs/+QxwzHyLVOF+ehWj7ztL+TjsRbPr81vfNEr6lqY0
C5orilljJlHxI2B9C1/Q6ShNSgBrSqMsnotHv6+2obkxkiD/Irn1wolpUgjfVJRzNPMtenNkTBys
gO2yINfyhpYzOx8Ck9S29ltrQrtHXVHQGeQaviDWjqhfPthgsjmV31UVpxhMGmaXhRefru8mF2c3
Xn0VGfIEljNmrbpovZdU/AyRHerAX2Rak9OVOGLxPsCVXFybyGks2xJR6SYbFB+Uu5VsWAEpy4Lr
Qc23CD/N9kgwz60c4nsPceJDq3y7v4guvrzfatQNMOkOq/KxLC8xQIjrqAjjH9K02xzqUjipmL/3
ofEIfiyS/7yGsonj7EHSvepABVZ93Z+3T5LFD8TOek1bteaFMkDzv/eMa26QI728vfGQwzbhH5yd
HS/OLmPFJgYk0+rPiR9J8WFDGWMjoJ2v1+a6gZcqYeYSHraN+ob8yLKqVC4eTRLE3P8M/FCOoGQT
fBAhDDfYKVGqlS1OmNsyranuV4DU4r09YgHFUcKPEyssp+go+pbtSgn3TstKRSGhr4UDH+iqMrpV
fHKyzFiBSLpJ6YxC6j1qJSPUizl0WNDiOS/uZhtOKMcyVbQa52vKOgzFzKWgn0NOrwmDbcGYa5NU
IwFgLEYOlrlY8+ZIwh3SxB+zxT9gM7TYKmiIjLt8rTbg7FSNy5BmYSDRM74qaeovJTlwRvNMARl7
1muRLNNKwUpGZ4UKK3YvbmoLoAWR9AAFhxX65wGdBluC6cNrrkN/jAShrGwQZRAzP+A6y1zyQRgZ
NW66bxs6x+bP5C9B+fLMHUlW1Dh8u3Iv6AHv5Q7Rkcbk0q8DbCZjwpuM2dPpoMBSE8ujbgGj7wkB
pDUX+CWd2osRlgp6eCmaVH6INbnIXG9QSFLY4AN8IPByd2Bqva2fmNXDXzbOrh0Kvxnz9gSdL5hS
ud5uVW7keg6O5LDJ3XYk65rvX7kl8PQDZ2o7NduVgkR6joJUAbh5deNfNn1LwHKR4Ol8R01BI/Cg
0QcXJaIzqjC/k8IDpQzU36IRkdY26ZlqYtfdV0+AkZvOkQ/hhRzDBsEmUfrFh5SzVlIKB9nO/ETP
FuMrkosRlLCgaFIdkI/GvOLN+qYqHVO0DxwlOjcqPzKvhHkrL1VTyP+t0mbeuWVuN9popA1Kkdvq
kdYukhG/1iR63DI8ziXRuGBYy9ZoYK+ergHedu/C1aifRqQzYsydrFGlQTOOoVDtUns/C/PiKq/M
46FogJWbnHD0A+5l3ge0XLgRj4RU9Da168ZIgAl7kyYRdJenCtqYUiuO43jT/pLPJFvPRQMZtQZS
7XE+QwJtlTFfH6sOx/wQB/PueZzQwRddoDNWYh5hO9S//vDYW0sA/5wiwOEVL7K5XGCMYZ785wiw
zbpg7bTCCV+JUQ+dT3t5phwWwLkbQ+nQCiacps30YNHH4KOmvaWcC6SJNifR1XAYTAfnoj/EEk7q
7HQTjW1Qr0X9+Kmqn+8KDyOSnWVr2IaWh+PBGoVol11BlgMDPCdWP56Ox7gss11/lf3ePklzhVV8
8qljmMNXSlUbluuRVApGFCXOQ8pQXcQBKFBiUahyBB412mw+Ryqju7W/DHxDVEDBJDCs/UOh8uEK
0cRAfAC2c2kD/At1QbN7ScUSmR624LDHidyNlGqOFrHPip/fgJv/97C0h2rl+qf16JPOvULcSzL0
jT5RLiU3AZ4prmGX9mqOKt95+c8b3EBOxW9Tso9+n+QaSI3h6jj3Q0lwJfq76pKztYT1J1h19Mva
TeOLjXnHbbgZJWA9sE/YgkMeRUP68LIXgW0RCVdwzVNPhc5N4DYa9LUAQ3QpQmUhdSi/XGw2Obi6
R+jSWKaU6eMtcGS64X8jXq/Pzkl/RCiv0A61mnxJ60Kf3vVlH3kK+0dP2PNT+jq6nHQ5KeTmQo+/
B43OZd3CVzJtozd2Jtu8Z0FdwVB8g+w+wRM5guraFNAdgwxUiRzdGDwhXdaYdRNBl8+X9xgJNVZ3
P0iG0FkfIco2YSeWUl0PGe+Tkmg0Srsc9of+Fz1+kOALPfak6bILNAT0lS6jFRSRURPA8HbGmdyO
oV9qiqQqLBREUaz0xu1So+xNRMXsUijgynrJXyFjvV8kUM02coV3/sxaMJb5giY2tDmK7Rs7Ksk4
sNN6/C60VkusgFUEuXe6rrf51eDUowKWBIeOoLzLa8Zq8Fsia7F/1WlZGXsMX5KHol9ItldzTIxs
bPqUrRza5DjiA+jSgbe/8n4SupiI/4KckLNXr3ufqIGTA3jv5E0MYetvS3UjBr8htZn1vWcB+cu0
RGas7Gzlv+/rdLaogQMnXMx1UBlZBkO0SRbjBFHgNXVRCOTwcI8cr8tzXeLDRthYXraT2jwYQhHX
HW6iNOnYRUsHtqt3s4vfl9F9rtO41HjXmKOztLhy95tzFUwIlXLgEcgdVu8auhe01OFz/Ibydzia
UF4X6SfrUZmcqvZTMLAi3F025VdvtDlsa6bwXDYY9w3wnEoGWzG01B0ftP+u276ibGH/zp+wSs8g
BeOxfqgsD/MOxvZqnsicscWtCxjTkOdzz0NAkaH2zYj1bD24Wip3ryKTzc6RiIopPba05OCvtmFa
I2ZduvmYhy7EpO6abTZ+UbCxxCvGB9u8f5lNXtC+98qN1EG1TBGb8njKAPeUhh8xrjJQJFu6rTgg
K3Ii9RX1NTLTt83mULfySqFCuU6tzrzQ35n5ARQ7oDjQwzgwLutZOIwjWRST8FeIcKhz00McMzpP
NYkyYp+pJNAezdmF/ypCM1IT9YWStkO0xUpFiwRxOvrdqYvFd/k9gGsgkoUm8PM9M431PzwBo3F9
qPu1+KViqC7itSmiqkYzYxFtFG20Artk/CHkjUzv0WtXqlrrBvU367C1AYL2wW26Qlq2kQUoWHfk
fxAARJd6P4D2jdr1OrLPlmjIJ/Cp6ESHXXjf4UPme+d1fdm22oS30h9sRwyNpz5rYdeaqUovtVQE
3he8/xxgx+/HmNdRDf68PIkeRddsgD4RTTqNCJrbRZJIYiR/aaLvQ352q3ATeMhacFPvJBSx3mOi
kYRJAe+CJxPemYGIktJGSuwsSosLKUH/HgpEV71h+T1eGsjDfd7bAuC4DYv/IEd28I3kgM963Q1W
XcVq1xw5VHhFm3OSGyKr2sBE4FbTAnD8sT/tHrFgVTLRA+zlbzHNRLmKclQodyoHWKzzzpyVjC+Y
VvCec1s/a63hE+w3AynDgsXYL2Z4rkImQWq+VIYNj9TGvaTsDdC0hojYg8ZJ8GsVRvWHhSzq39QQ
H4j6aCVYsU6PIZA3v7mR/fyQ3PNSyXYGeQIRVQnh8Hvcnv/o3efhOUmgoiEvwlFXFbmpV797ZIPC
SWHLDzqxavvARTQFmOYwfmm4KCT1z1AW5HcH2BV6OiEkp4gtwS1CX+5m9emQje7P0hHLpuTZDdT/
ftYm+Qjkh+rzRABmPRU1IUBMMQK++LYfyeznwkKu5I+D5zHSOW4SGD0+g72q56BZGwmECopfcn+4
eEfJYop6//kWuTwFs0Vs/fvrAlGKkiW0tctB3xMEzzb2Ug4jFPt4C5/v2VAYHX+n5orIKs5DMi2R
tLnrnUURDggFui2dsFzfJyXE264m0sEXSGYhyEA+e5iLBnCfH5Oj/K+DPK8AsnToVHICsFa7xTOL
JHfTwQlc5eMYltsfMP+9Zv0MSQFbpctcdySqAYgn3Nn3hpGu6Z6H8t2bTL1PzRfXqTg4+Y7T/YpJ
rXaHTGNXeR5IB7I8yY3K+invfCB2LTSrk/VCSaq+0pwe2Yw44hGiAwd7PI8+zry3XWzZthc4Vzn8
vFlzPs30fLulUmGPISGAT1N053zRs80FmTJGW1jPcVpHxi+sETJjvC1vluVAe2VIItgOTKz5wJ4g
evjIJNDICU5HMw/6eP03ED07chHKJhYK1FgttO/OH4s2FvpFVjDD3QOZedN4a3ILG8A6LRR9c2x2
j04qIFpjmUe+D4f9mFVbzlmHAujUkXAZtOfxuni9RZb9UQhf0OLsXnlbvzkoQxkYFIukHWUHVZ15
sKInevEgrH6M7NSlqv2Um6YD2S4ndG3qwhh0kyWfYa/4YGtDirGS49hvNqyXwSMDd2Z91ZLCeNau
hQtYWXomf43DjDbS4YM7/lfLAQIGB3Sph3jVCS4tmLAGD4M8/2/ZMQYPQVm7URuq2cvlSiSSicED
iUbSoJoaMatOj+l2pgJtj86alF5mDxNVjkoDxJR4lU2egkEEVl2GzmIsb73c96Ckk9oOeq9xUqGa
9yKDrFztbb2peKyiPkVfYxL2vta4inWX67SUYJL8rslkk3u9yibYMc9sDxBYTnH3LrHvzIcfR9vr
ZZJ7M1NJ4Ny0eiwyqEdgf8O8rtew2T+HNiWVufIZxUU2TzpnwkIaWtgNTuF/C6iuVfjPVJnrdavi
rGn6CrNJMY3q3fJjA4xbJyVOGIJvujnpOsBvY0E7Z+iVOlHxowpP+sWyJctRwJtRECk+18Ugh/9R
AxpuQ/JImtISEvAhvWUGITY3SkVIFZEekrdm7OKWsBUT/CenD2Vjvrz/RTE7mYISqnXRoCR1JyMW
P+QB78251lbk8ZlaIGJS9QEK3369tj21VfiKlssorHSCvnCIjZVDPhC53IzoZJtCnPN7joaOTP0Q
yT/+CgSXxAVH7paf/lr6wmmdQ6r8mcHT639y/ks2J656KhJ4adf6M/X6pQeD8i8vHjWmdXxonx5V
xEspDFaVAe9w0RdIpBpGlLdCmQReW+AbuTlOHyHyzTzhl/5w6XImHSZoVD81FuPfESjz3oiAbsZ8
cQ26meWzDrd5avK3gm+WCsTcIcsDmq5W05sx/zJ8kKaXzIF/o8zY5OVQyuNXG8qSGgolUK5lGLM+
v2bypsWRs3LuvteXyxGleGuy9P6jnCRcIl9GVNeJ8DWvphdiI/EpvVzK2U5RthD96M3Sr5GtjZbn
H1hWP6AtHdn1iJLEZT/9i3OeMpvAjdxHvr1/Bh9vZZviTuKXdYondlzI8GsJej/ZnrU1LAdhhCdw
t6nljECzDbWRDYYZ7WxxdzEni/vbEsx5GN5v1Pst/CTNT2/RiNj5yn9vIPW2zfshDdBmSJ/Jr626
e5Jb3qMlPdjSb8h/knrBtZurGBMii0tkE2i9ftrdMgloVyzk7DUTPFTEnKtgxJYFi8PlPDeLIuG4
iiU7+6oFzsz2m5k5T0ZUMkFdCbhusZvagqM7qVDcTL62VsJk9Ack7kBCU4i9g3CZ6Igi1+7X+ul6
qdct5iUoJAwDFWwrfigf+7P9V3xp56CqlYAEFk8LMqGLKITaFL/1UbGtrjZdZICkZt5ouaYfbTyX
JLrPxf8BirBPI/P7yl1/pJfsk/2bq7jihRDt3wGjyE7Z83EdQM+myaXZjvGxjLRf1IuPGTjtGOj0
YJ1jczWiU0Sx1bYcFwIBu1dsfn0aTGIt7AybOAsp5TCbgPg1Ns3yhUhbuBmp8CmuazLXAOvdoMkA
GYPcMI4VXEEEb4DsAHXF75ZZqVsnNtpciu4L37VHZQV6xq63strAVCiAUtj/4PQ93o4mKgxV8yFI
Z46/Iy67kyvPaP2PlyuBK/VC8CoLtgqCYS2txys5OlTzsNgEhCg39JX1K8+k42l7ikq7kAXCBAxt
ptGVkc8XEFLy+HZ5xQ2V0YN6L3e5V3zS5ZpFc841TQ07NQKFlJy03QcdsHMUVRCIKPXKyOYIofGM
peomc1nuq4b0ch1AbrwXPxeYLLKaGmZY720SNTG3F9YZdFmhbobPGjFQNzUeSHpuVa9Ithn2E+9x
nwvomEhb1byASMIAafKDS0n+QzEviZZBu7WaKWlACxq3nhpG65orjI+g+VMepMLCBxY5B9mododA
2YqDpWZkWfgwGNSOTNFd0ETis1r1FAGRr4jmOttqacuuh6B2VGMybyfKe5okn2NGaxCgkSAQytYL
ZBgTsyZb8r9OaLyoItP/wkhHxeUcbXmv+W9tZaOfe6VfdU1tLa0pSjYQIUPeseAqnf1pv7cm2zHu
oKVDIsidTzZzBXBtpjqMJY8OfX2os5W5pFehmLfiV3+zjmT8U+QJtGX6o2rJm7WqtwVxs8wsVdv1
MZLGWsLgm4eSeSXW/w/uINlTLJzrAwIfXtR17EOLqEN2TgMBSI/KgqnxHxE89eL+r5Edo+CLMQ0j
WgwmrgSR7W2VYMiftRw+XuO5BpnoaCUBDtxaSE2/dGv/vcJS0DmPSe3vuuchzbPQYCr42awlGoSP
pvV4dxAdT0mT5Kpr4Vr62etW5eqip8B7moqmF+QK8CJB5TR7pXBfZgvJ9L+x8Qa1eGk/U+3HkYhv
5KZdJux9jjAsgMQCZlzr4dYL6uaiBGuGQp6Klco6WyuFgQS0Ub6W6Rh+LVIs1evUcjB8H/jjKFoc
CsAfEEOB5n1pojatBun0aJ5IdY9WEGK3f5i6Fjier/lnMTTTMYOsHndCfVbqveJAqC8GOWw9e5eh
81wVEjNjYcVieVxbUQlK6vNBFCD8e3kz8PwdTqVMPqiQSsOIFVja/29KWFx62n9hGnJSHzJtRGaS
LvFANk7/DJHlKILTsSkQEqoAXTilmkI4QD8M/PduqsYtYJnvoXg5JDWRyoUREql8/vgjswmzXVWi
IoZuM+m/x2O1ATNGqpVq+8CGGCMmYFKmxfqVBGuNjDdzwbGq31rHX145ryD5LlFKMsZZktnVFPuP
Q0RxFDvtLop+NLyYbRR3TwgtNC/24kplgCSHFZe1pig39iULPGDMecBlRajQFHJBcxeS5PY+kIN7
HAG0xWvYanGKwF14T0AYEv60yUNqIYKk01JSu0t5hN6QlgeRjBQEaSrTNo2/AY5CxLad80hxUKTp
5EZzbKRKpLxTZPB2NbHDMl9+3gox92bMz/vkRliZpZ+7kUOR8i8RDRwrjmgITGUcnuvbJSaxuGQf
WUknIv5m6LLaGQsgYJVmo0MWz2f2+Q5JGr8KulkJgz8Omt5Sb4X7TLWz9ln7eKid25xQodwt4L3k
8Y6pW6vHX/dulUopBuw2GlPHEwkvvdeTreXA8RayVVR1I1cA2Uw5CHVis5Iu0OZ+TiBdLqB/Z0Dr
3ZBiNtRX+04tBGEkh2RWOzqxf/lZrpvEYGbAzx6mssnRVbFUvrqBAQP+VzsCeDn0fCUlFQIQuw5s
a47Lew5ZfpVbbNfujIy/JQy8TUahzGQMgYLDW7ILxhdjxGzmtNehBNkITaHFs0FtBFg/RJz89Tda
9nlaHmaymtNeGmI635Jy7KEIQ2viP6LZF0as/GNu5mzAc/rvXGrtUtvuQd8nMZD2YxYr7HNHqQTG
5iYy/Pb0whRHHqWKNwflsrYpG3j/GzoU7MBZ37Z1T+QwHyUKygkiOWtr2W7E+6xsaFW9RvFXsjGR
MYprYkuQmp+A/Qx6FszpNmkB0zV448tHnuB7lHdiegr0g0o3rMdct+Fei6un+vslORmVrdnTcOW/
DUokLy5yBbFPbFgx5sal43LgIpJj/YC1T51g7hfpsMeOJNPOFf4RUX2nP6qP+pGnyK8BMih0TWCO
vHDsoSYuQtNwbK5HfA5PAwSwvI1KfwKRt4ac5NH0Z5ygqaUAQGJuxAwKIQLato8a48oj0JjM1Uop
kbKEwtfpvIMLjbVjG81P2mWKSBePzLgROjktjdsblWnNMKwN3N4HGqRmTJ5TqHI8FOs8rQmB42kO
aHygUag8Ol/TWlSCmF5VUToV5AXUwCwDdVEtoaOMxzGInkMT2Wy/1Q+/8kOZzBhoIiwhF8OZWGvY
JLxP5fhtHWNbrN6JA8cTPXhnDB1JIPt54wiakVbICht5bxnIFU1Qqw5VhYLG5+fBMLTRIG/2mlJl
BmpwAKDW0RdE/EIR+hEy1mXifleOKVzPngUUEv4bTj7tnoLnKd2qAVFxavRRKm/k1v2PEesr0Ui6
VAn3+0CnMEYdaqx+5noYbKfWLM8jMTIdpTa0oFoXj9m/gCD2308Gtg0yw3Npi+F6mS1lSOAcMrGu
T/7JCakLWk9XRmSqrTUgfn2+u5iob/PGT9QznTioGnLXUGSfNMS3FjXE/hqwkzKrUxNf6i/nVecz
o6F+ZTcTOA7xk4mzSI/aqjKqBA1GtZLfW0BDPfomzbak+3NGhWODtalo7W1paxMzyLrcDdp39EJd
E+ZtF3kd3vm0UGGnTnNctVLYRW4OvLJoJCRGifDbOWZKy026uvzmxOOjR2uMDS0MY1l+Kt6QKMOx
iy6A53ivclC/kYrNVPnvhbYX/1iO8LquUbptICHcMGMgmj7hzMQJk6m9AxXHlzWMf/ST3U64HHk/
h2K1Aw/GUe93J4b4yAeokRr3gsPr1oPDdsX9kCWCmZ0IXvSkMF11+4ke4qljXupLjDoJKDVBG7Oo
wn81IJPc6iXTIrxQPQYADs6j2xugXOtfWV3gGWaXT4i08Npklps8tWUKExnlXMk8xKAE1sT7QWjf
vF/CHVBeDI3tHw9XxHG+go/H8hvrjOUMCRqKX2XqSaAwMdDZjznrCPLMTFmX1XM1UEhO8UwsBgKL
ByVnexN07J7B6DYF2CmYq2vZ2Icbjq1IzCTcppU8eeaoKaoDUFaKa1Uyl5JupTcO+s8h46GHqB7K
TDwCP6gS1TDvYGV5RPAwxC8Fn8R/YsXHxtN4JCzprIBhaVqGH7ekdFohmcBtT+iP2x2Lrc0aq+vk
Mkb76KxxOFw+s1yTa+/SjVKVKIActTj/uHTHlC4U5Fr6aMgieIpXtb2qVqv15TgutFLdBUJh36H3
PSI+GEGZ5W+6SdJcTrWvRBX0bSIRr9IP6ThkFuCh1tgndjGNNY6A69jPafPIbDosmpyyWSzOdWsZ
FH8kmT9AfI1EMTdYUZpRXNL/c9zOd/WVs7Pr9UII3ZDA8BRLgz7J4vwoEzkJg1qqHjyWqoCNMIOM
5zRBbOcHrXXptbACwWBEbtz48g0Ny1g1VDDc04LYbzKaUWxILa0NjWB8vmsTO2e/KZSMkyS/NghS
iK7RwbV+YT0bgoO/8PopNR3PlrS/5+qelpadZVDslzIn6Qfi5/i+Ui7rp4fB3ExNVSwbLRXEsXXZ
J+OAqH6f2S8j6bKF4/xX+6YodcqGlpwqdRvEF9FQG7CKAMDnJ9FW/RvnNjHtFFDxnMutrx8eY/u7
4N7Z0+K0yXTZmFN+rrIEX0miDWVzVZokKEmrnAfel83wgdhdreMc/2ooYHwAWOhASbPGKvjqI84+
/2LYY2Nnn0IFjkzxO397slpVCdUlzN25rZ73OZCyLVYgOpCa6LiE+7pYR07e9YZHaUjIKctHfnz8
oxpRjJ3B2QIaC5dz2mbnznYLoNiiRf6A1jAWrr1j1k6yg1kNA4veKmXKE5SahXCPOujSmwJZyIsJ
qlA7oYK9OU82h2Bj0hZ8UIW+2lVaAbrMC19pNyTmcD4A5OVXy57tmKzC9te+2i2oKJvOlZuMKXaD
dBQ8zysEthTUzFAH3/S6SOvuBGjtOIbcEbLSwkNDZc9zV/MBdDhHlTW4WtKYwEZPbVxGtw1DhWAU
KqdsR/Z12o9mGb2m3PfP+C/W0Bbh116UxVXJcgd9KFvk5+ow9TCLq/IwgG2DwqSrReGGWMmdnFRv
bwjUp3n2EaO3fgACV6YPD7FGduiFIRJ3q6DxXfVOCfwI9qLTwtwgyjkAKEb3fJ//VtYzRT0oNqWU
jDmU1TScEQ2mJS2qPpfizjC8yS9nTr08RBjhFodR/Oxt/Ea649ILoB9FY65K+Fx9sVff7b5Kzo6Q
Zh326U+FH/sK+eUGcSIz0FZopLp2e+YY07GdS2TLoHA8MRGH4qh/GDIbMVQ52r4fpnGvbSuDqEpE
94PcAbhbOM2ENk+0GZVjk6YBCzygHSLj+sdM1HXjQ/faU/Cz6xm4MqVB7hMSehvzY0PJ9m53EPcO
FVj6iWhxFrErW1ie9A6kCAz4adn2PDSB8+hABj3Wt5e3NB62PAo4jEor406hTT+lZlL6W7I4VAXj
c5cYcBvK1Y4HAONePwGRgvwvAi5ovoEXRv+WzuQVGrAD6QlvsTtQ7ojQKTL8lwOWUg6iAcC+yDeU
i2t+1A3rodRGJ6G85GZKuaS4Q6PqhQs/U/+wRojAwiF1PqLoUSbOGV2L+EU4EjbieoGgdY1mtE7Y
ES/5UNArQqGMa/DIlxA50WYMvo2YzMs69niDoTi0VaXN1sWNSNGgO1fSBJzSckwg/hn/mCDFopp3
MGzXP2At7tJlMrsBq0QtOZExRteFfVZL/pyTdV1pKRZDGKike7gk80d7CSNdouo98fJCChBrFcKy
qeQKoWCGNdKKLFCPP9Ou4N6TpBPL6a5FPTQNzpDt4PlztSUDWImdMqsULGZ61PjIL9maSFNLE98Z
sVj9wMXM0dfF81PpWSujQzxYUvQOPGrNmjyehFFuv2fUdoNli0gCEt4xYBufRW2LmMu18rmWkJfc
1p3G9yZniNoc136xYVcWZqfq+9aiK/xg89kbWjrb+ffQJkuxYMdkAB09Kpro3R4A5lBTHV8p+6m+
I4IsTY4yxsi3DFND0WHPxdu6rGaaK6VMfqesUlAbpiMB9jWrHGNqohOqdoAvyjigYUU3rjwA42ta
EgpLku0vN7dpMvrRhMdg1gQvzHBd1epXpHDtZrYOnDj/x01blTtIqw1vBPORHebvihrrXEbkAU7a
tRO0d1JTcRbLY+LTgwOTmX3vFxiRwn2eiR7pmHmTWjiJ+Bj20ksahnrTCWy3sJJ+T6hHZLHdmFe+
Qxa7tF+u4qQKvp2YEXhGfsgN5ypX5zIGs1bAKkbHA7NpSZwcU+lI+98TNPHX/oohIXxS5CO251cl
wdGELKJGNaUv+0Q2i83NKuGcUtDU+W5bWXhsc78QYqoGr7hCY1NUtdHEe7X6yBu2FI+qC14WN+Mi
9i6SvEsuONnwiwfxCrCV154csqZ36y5ano5GzBGWpwnn5NPjHH9pIL45vhR2KArag3LdQKcyqoAe
0nREy8B/pQO4dyYOvVJ8WJU/9tW5hzldHZdaaJycH/euhgKSFBF2r/rRcLJfHFMk+8/th/WbZwI1
+2QJiz9hVQsVRKpcElprsDHlBUL028WnouZ7KHMYi2fOtyjG73xdIv88+rGYW8Ew4dyBc0ad3Gri
mhd+TF/85ffsNph7LFbJWrXGqPgy9+kw49sw40rbKCZQXBktEbCFJKeX9aY+yH3fs7VEtSTrObcF
MtCCvPBCiWvs5boMgMLxEz2mugREjudK3tPCf9GNwXLjsibNEMOf0DlXQRunh1ZlHJYHiSw+VhH9
TdGcHLmLW24XDETjxpQdxkN1HxYQlcsBSz3MmOmSnSEOML4xSUb/cyazJs8R9Ycx8h3dqc0omKCE
OYAyCFUGDz9b0DYSNuYPT6KXMnGm978pHr0C9JXdX/hFkIJ/Xpt3QL/YalHXcX1ehr0UdJktVpmV
Ao0VCRg51Oer7ZDUmIZTA5uNQSQvKnsKuSFReO2/iGL8K6qtnP7p9lW8d3hiCxMMin3fx+mQxjIg
zlrok3vzBWvKNiL+iIYbvY5wHekjtiWENz+OiCamfRT/SWSEigt7bz+w6fNRd902KLcPKZo4Qnnw
OFintm78jDAH7U9GWIaz3SpZS3IfEcj7vN5GnXlwnBL/kK2ZdW/HCLxv1Ood6eFKqnGNZeyobRVs
Mtmen8AI5E4VoXlykk0pIwVveBUUvjD4vb+artTW/nsjgtUY9E5UtekAS4Jy1eITIX4tvQDdwSVQ
dRHmJZs8GGE0Y3xDkiyRkOa4gLkflLSgMe/C2JyuOP+1ABypLiy08H6brutngcOaVpuyG6BDxfP4
N1+5nn+m27gpRnifmtZcgAR8gmd1LGOltuL1+YU+WiomlE+JeYKhy3pCAggTX4KI8rOrVJvhnYme
qrMfvTPbPDgRT+MglcRvc0r07rNn1FvPMaLANLZ3WJkHOFKmpbtgr/SCCA8uLRXJeb/mXNQEavIP
ONqEbI08B/grj5lFfUzXFOCX3plimfAfRCKj0p9VnRjuGM5sWDNsbTmzt/3jwH1oq6Z1a4v9I8Or
FYRXHWyo6+B2XPM7ht+9gUAK2g93fLjGXTyAWXSMRWPmAldxJUIcnxWhxZdPiBcICSg+d2HllNUI
k+gQbHb/4uPr+SnXPIaAp1JHGMnjp9pmpTnKUdagiM2jaKejRAYjaqhdaD8mNSGC5hkNfEafgn5I
4hraDYoN5rL4EudJIDRFeXNS733LT9HzFg7l8imED2zz+DJrk4U46Ppx5G4nhhNk1SrKzwtTdvyK
5nO1egTk7es2IRxm/Yg4vuV3XpNqZ/NFxQ/fK/1xhGsJLN692qpUxfpOL2OpSDvqUosdfiTK6Qwk
9d6XUKydumemKaUwEJqk+Dg41gunrNXSdCkMsJbnkcra9/JXldFo8MQYtkkB77K8PJWr5qUTtqOn
cmWAnDNnG7VbUvxH+iQlYd+H+avQlRY1ig+q3Bim9NyEduXQPpwLQ5hOGc8tvwvM4w+27zakpcHz
r4NIJsH/4mAlZVNhYVG4yahXef9t8oJMhZfDsJq1pF57wuzF2Z2zlrxf9RnHpr+G0ZTrOG1KBCfX
OPxSx802s+3lRngL6hKv1UHFlII2//X0oDBmcRZTGKf22v6iD5ZabJ+rVL4pV1j0Moq5TvMrD/xt
7KL76AmJ5cTRPGftQ1HZQmg9mXyuGF/rZgdNsWy8rACeJnMNv42mpjI0wuVpzVW+0buBLuAqooj0
iU0oqeBQVBPgcC3WGGApDJgi+LyJw43HB00sUWIKo9+y2ovnPeI2btwdAzauVUXwg4uQx0N/i8aa
GPQEzcWco405MO0qAeg9SzqKYQiVwKA9KPhMvSdFKdpjkZ9vEr5M45mYxzQIvjA/sUx+Jpte+F1L
ZTcPLZZWn9tv4gsKScXizXXDjh0Z/n1HkpKHxJf9DGdzl5qkgGYxjL0jtNVUOq4WsM9vPF3ojAlD
efJiUI0ix+cxOi4nSn/EraQpKN30pLmm+PF7PBx253gxOVu9nfwBlEMR0DjQ4yTKqQA1lAqnppPL
obNLZ63urjCf6VA+x9sYNIskitYWeKiHCPo27RSuc4jtZgxPlMc03OitTstFzDWJaoJRHrRCuDCy
lWL7fdN7rJGBO4barRWY7Pb+HQE2Xv0xXFIxZ1Wv6W4jFLehc7G2prBtMWx//2bXF/jbRT3+DY+r
TKlSM/3O0OTT9q95EoJA8gY9Glz5WJfDu/r2MOPqBLz0rR3lIWa9OJrI2gvrAZSqRTeJVAYgyK6X
COL9p6KniCnEq35zM5JRzhWUbzQc4WdQLY8cwpuZw35IvYZYb+d9CQHs0TFrkg+Pn7lwX5bbGUha
2GBcuG0GWkQ3Ig4iTuVvYQDiPOTk9ktpicRyIA0Ez1XI1oSPRvpG1HlUkyredxg8xZJytq4GOaKV
8eGGCpbQZPT6Zdm8fKlzPtemSMgi5VlEWTK5bqJMHRYo1T7BXy3qwqOo+0dvke9bnKCDWXfAv5i6
2e/bS94V/4a22RN1ilWQ24SpFcpv51ewtJOMFiNDU1GodtDsVmK4rwfgm+c+ouwo0ZcfXcCgpzCD
EjZvLx2I2nifKnRRGJqmbGhSTK5Hce91KtuFY+v8mfbnIFpPcIDRyDYLATvEj9xJ2t/KXS8Jsuus
NB65/rBDe5AzlNqKM8FF95NnjURgm/x78Z0u7U4JfuwLHVE7N8OPR6jRwZDDOIB50mmBqpD+3Mg3
/aqJTJ4Dd090lGZoGQnoVVX3P1ulPgFnBOWgU8GC5Oc5ajvBRKWUS92PVuQBb53w9sLSrLK3yefT
4Gm/YOQouVhl129sDYWsFngl4sJRyutjeuH8lFDaRmX4IQ/V5zvrypwLFyBTlAagV17unXnxoKd6
58mED3e0v+T3N4iDz0+uofVGNkCGjkSQQK05xNKGgP/wdrffOQpjsggKLx+U9j7JXtlh6aWD8eW0
Brma9syauHGkULE8PtqELkJXos6+Sxnc4Ce7bdE54v+YFT8CMG5N/zmJogEbtXzbMq1BM0Y13OEK
bjDh+7FicIq6dKzdjl/wheierCuZgoDF4C4igd2H2HX68ZxdJ/PdSHbn1Qt3Y4WiW3gCxF2sW5PZ
PRUReL/DeMJiVkrqv6DeaoynaQ3s0fUatamQL4fZel0W+WgUgvcGpKqSkXH7D69Oj0HmcfbHTIsP
9hsswYIqOQDLeODmqTM0xzvBkJ6J9xISlR0zoJDk8/A9aWeTFCXuQEeKu1hjl3P5yZMVF99Ly3j3
GUCanwnWEh3zDqeHSV1howKgUr6KGox7B5jv1Bdvdcc3FDstwhA2+JsB4oIifQvXRDQLedq5em/F
e1MpKeApgM5bk6bsT4jd1WCtmmxUYv7yQvYaGO9cLa2BfWzuqcKtTfwlVwaKk3YF0MSh1WePexEA
2sRDwSdD6Uf9JDNinWGecW0kWtQqhBJgC6O4/c2ZOlEpJ0NHDrvT0cod/tP938QWANJBne7c1nWg
m4BFyP/Qv0hpOH9vINLI9sixnbcpYofioy2rF6O07x1WKCKcsh/gjySkL4A4+lvuqElVJfXzdxh2
mLIg1frPf9W/xo/l6miaAfSIx8vUu+5SxVJnXuWmKm9HkGexBKyVEk388xmY2tXVyu1/aDRL+LbX
kPso56U6A5sGt31tmo6EmQEEZYdoCHzJXy2+t2Oe5ZNaMnli5o+fTV5G0sFOPBCh9UUC8wCBk031
+lz0yYNT/+BnJPhJvpREMtfihPUBnQb8JXxoO3ms/RFDwDwSGPReFZaMKIHBnbGSEfd6uMd71eMD
PRG0ImdFCOVdtNQb54qXz8ZGpZki30DhRW0xAmRrWYMfVdT2rypNBHj4orkCcPhghrDP9A3rjPKV
dYx1nklkH2sMjR4P0X5B8uhaEwIxts69y1D7hZzJ+QEb8bbHUrQoeUDeIAHuN62M35XnZJonJdns
VDww/WYJLb2Ur6gmeZGQcJDOrlPgaRAdZbVRv8NJmGju6s80wTIMyp6BnUVqPGNW7BOcsASkDc0q
PBENUlqrEyO7G+UVWmlGn0xRP4cv42nS6gBglgygX6BWGGjppoYwyQvyCsgATduv7S31MxvrAmL1
hmG4CyjPE1c74FXOtFOLcv4/P4f++y/E2w6XhQQwbKRyicsMySsijZfWMsAmVirc1PcSpZDeSGAF
eZnduldtGwceb6KYSE1H8HHHoCC9NzU5sRwlsdn1SMYrvfSwP2I5LIwj8PyH9pKT58Wpy0lMZg0c
hv0zfg6H8muJFkwaUigYDttOUCcQWfYqq0lf/L2nPLBT+96PkIWGgTwfg88ZNOkfBItlpSWLolNK
pdDFs8U0e3IjgnyW7p0jmlaV+dzWz6aDbX2SHg6Ut+qVAc3OAbNzKP6HOo7Y15QpFDLpTQ5ig04A
Trk72x9M+8Y1qr/9OziFyoZmGiv7HdOThb4I3NxlJucrSPQSOcM7WQIE5kTX9tzHFJS29jNRD/Fa
DIMD7JgUhG1pau40K4j1QQvSu1eal8+yYBA9r+C8b2tuhhJyaZ5PpiEkSuEVFE2wFrGGhCDljq4L
I7b/2U5B7z4dMPzsEZKyGpDI1Rv2l/jV9BiI/f6eDn4iHDOcfXr7paKDSByVgZ1Lif6RyJsOc4qB
37m01oDHzssJxe/N5JHsDL72jQfm8Mwr1HzaRjOh3AXOU6HwpHJu8DalbW6pMORCq8wR+ebaYT+2
2fi65czzPfdZDNHeGc4RYvKrkUlILffB8YSVHmbRngqB9z5sKhduYHisWBNU2oZYf7udKvasDumH
YjllRuzquHHyEmGO+bc+JZ76GSBAmvlR0FJKAbMB5W3Yx4/qs3Ok4d0wuUctSf5d31NEN8/Zi0zJ
GIrgDLn30F98Cnrq0GfxNimsMy9hiRqKuYMf/M83lRaTdyyswg0WkooixmSXibV9bLnUdPOacZ2I
nRcF5yYVQAXx3rqweYXyVw5zeI6P5dBx0t/KT6Jy3Slx3afiHA9offjb2JFt/k6pvgPwpAd/Xjfp
WxvdIFlAO19r62fpGa5O4hdZQwgJAQSuuP6RtJYIWyux4ywbZeJPCOtkxj9z9VxoTMaWRPe+UeSZ
QwlsdlWpTCx7Sv8XioNc+WP6Esu/YfEEyCQTd7lSvKtW5AlG3zm9aHNy0qnlIFceL1HPQ5pGxMFU
9l6ZA92A7i6nXlqGncgWk4BZLVoMNaNfWEr4ftgPsAtZKONbwreG4oeX+QlRSgczlRxt6y/uJwLq
wokD9cy5RuGVm/iitm8KLuUeGmH6l5JEc4K43g3Pe6h6Znhe/7hMHngVsa0+LX8pDKQRhS+UZyUp
onj0hMulrkpSTrXdqgARP0ujyA3QBSRz4B3ufZtiy7rJvCpdThGRBOYAMconfN/xia7t+TTyE1px
XaHCOdxqx9Zs6iFnHmrYqSQhD9yH/zpNWXwSaYkizz89sOLDp2s2/E3ySxzb6rnpBGQQEkZV1hcO
wwPjWMUxa0bG3l4MQZflHZgC7Foz1sJQ6V2IzkLVWHle4QRWQMPXcmE0bbR+SVR5ttgTtrvFegJh
nJT9HEbpAjM/gT25zsl/DGa59U9C+awrm6wWqmTGNFnJ5P3mLLA0EEuj+i5UsZMvbsJyOMmsPMC6
dZApHviz/vELNoyVX2f7gldZUp2IjUx4sErOMdpwn4m31AYJnYlOKG8a95jktUMC9iK2uMboJ0ma
wFDHJsx23CdwNK6F4XiBTRHxQluFtnpUMbNS2qx6SlzjDn0uMuJPQt/6hv3orOhCSnlcD9Il5PE1
fCzugdZFYRulUwoMNuGpezUPwbgYDRq21Z4ObTZ4Q9aOjFnxaFpYS5v22yrXn8dW7E4ftIK0QmiA
tQ8WMg+FUH6cI2smXesYm52mduXwgJhT19V2uLgQyiBtyvIJYwWJwwUs4XYwdAfzRrBwuRc1Grgo
ORhScAQrhI6tFelwC04geBM5CFCFE/zwASOH3Am/pyTpNFp+248oc5k/86ppEs41tvCXdM6AaFXK
Y7ydMIDdwprb3e6+YDOAmf7LZ6+uDKGBZIY8rNmfn7vcBWbPk3+2k5N5xeEOxKP54rdW9XiOus0B
ry8jd+fIRM8Ru8Z7hxpc06dTw0Q2FgfKNLkVUbk0c5jbSDwvV74UxKfG8s19/pUvtoEmzOWWGmc7
ygshcbmsJ/qw/IUPDTA597NYRmzOYk7tRmB+6FVIyZoyjBvgjJPxQ1e+yWXY+qnqiZsNYYzQvipy
VOWs7NG6+Cte4O9cqfvI3RXZGVVVLivuYUEPjwvqN4QGfEptN85T7FXINY/WLhafEpLbXbw6ge/J
6sKGUQ9nLdsa5nSNy29qrdlIzmj0ehI+xyKnHmbSHsH6HDVS+k2aZboV8YAuOM4GdQEnQ4nV6Kpj
JJczAn9P2jdqqV4OO6HbeWYihPXgDvuNaMIwa6uctBCZGFI3LQyyeIv7s17MQF/R0Kqw76uMNphD
YP4tMVfm7LkAWFx1UcJhCyqq5RfVUbpx50RQfBUkhldaO7OT6mzzsbNgIbZ/HCWtAKvD270ely/0
b4afw03BjFoLqaw/e3fHlD8dXLSDhVuq9n9wdKEFgzxrxVm4Tw8XwnbGnlUljFnsgy/mqhhj8Y3T
EoS7r0IZswJDe4ntdlUKSSODxW9+EeTmRHOhtdPH30UW7w1FN3sXmCbHnBOwbsvmu1xvBGl+fJz+
ii5n8r5VInTAe1SUBLsF7pfmFgWtLtHnfPSSezlhRHNy0M8dEQ4oo/W1Fb3ejMH6gakw4EPdktrl
mPbfHlTS+lVKaxkbaRFw3w7n9LV5TnIdcwXZSvJAiuGSpazz1UzS3oqefCucFaalu+t2LqEbR2pG
usoWTaD6NahPvbu15bsowZt2xliJf+l+LkXzP8HfwyrwsZ55xU+0Z56OAxrSfdcCwA8FA4eYfcAB
SVanGC4KCPMdLCINvMH41JDaUVklftTKgtzXfwd5yK5hsJTkkF5cdsyPbMEfpoMwf9MtiZZfy0+U
tdw4L1qAEC+sNn07A8GrR2zV37Ru2NOP172QpNkrTiKi/+CD/mieycQzKtS6HjM0h37nGdE1vshJ
wkMJ4isIytXRxD33dVFjiM6uoh27xSD7O9Dn7Efa/GSrREPlILjZ1m2KNhgkSHG7tAmxsle4zpCx
3q5N+yys1stcYG34BQNudVJNab0BP4wMlTXYXmY6edF7O9tEuxypyUh6oH1BYlTiF1XzNun2CfPn
Ce/mqQU2Wp+6K6QHhJJWWuwWUNCQaYmPDplqwQyENuLIbLSqqGXgXLQz9Ol3jWHMHSQsi9vCg+4G
mqfW1PnjiYYmuF73Lpd8tN4/TEUwb6Nq4ZsSlPdGqyH2lK8QsVDixX1d/etDwiXHF/b9dwzYVv4C
9zmx6v5ujMluU/7B1deQ80R4H59fxo3QG4Y0dnJ9QBHcvGdiIH/RsUceX1b3J0+3iYgXtRJ+HhYF
BrIC29xTb5ZhegRXOSyvLjwoMd0rxipBai7Ho74AScdlkvWnSgt6ylpioqq+WnvqIIaGQ8BATHgR
qWRNCdiloawNOrjFk68EujFr9GWtHL7A83ntCD8Ad8sOLlJJ7ROPBvkj/kJ6I3N6Cm3B+sZ9hps9
qtITurJ/Q07NqoAS0xqKcBslcJoLIZH2SkTxFRn9GnQKWI4wB1OHyAUd11EpZ4M00PAxE3vmTHN4
NJQX6wbwdmi+TY6Bg1iHKkBrfbxafF1jBKJr6JBahy3pyAjpWoGFM7tdhXEWyz5SxrGbTtjZ0JbY
Ldj8X7uTJcqBfIxQ8wDzycqhvv5R0q5gYvQdHZgdbha/O6H/Yk2A994QQgigg0k/tsymAMnzp/yE
XVCI4g3kEKKTSzlA9ZkA1tAcfel/4c/G9Ta5PxAAtoP7KikRK+OzexQjnPaQJdZ/hqfLXCO++VHM
tTkNPN/r+rDv6RghrUQfOA+UlBEACmfviYPriwFD3usATr1APGKq4rvLJWIKqaP4bxFO92Wm2REN
vpvhsxhQuFjuCBGYx0oQqmSkWNLsrgjjCo/h9EBn8ISirQp7bl9yJbRvqf8EgprwdhODtNyZa5RG
rf4vlRtF2oovSFFKi66NQvFvCCF8oLf+EKK5S5rtHfoIhJIt3QjtH2iKCaHL5CRglbS6wXgYRXQ+
JFsE+p9UfP48adVyg5DFZdrg1SqdvdZ5KhHQTfzrV0BLLjx2oEr+EJTdyuDUfWcbMYkXgWEmqmbN
f2ODz3qiFG2PNmWcfjviGSjzc+DYlU+HXCQCjzd1YpLjHLVSZ/U8kt22Ow/PqV+p023kX21VxPNN
B4LNE/vlUJuc1PZjcckJa71bxjs5dkCA16SY3QN9O4oBqSOcFcwSMVYfQ0V4f1hh/lX8atZaqbD4
aYHnixRspWqnC6VULGwfN3l0PlDZrEfRdCf9OJkMGo6U1sJ+34ZqJgMwRN+vCJxXqqm2lF7eNrPU
djOJ2Qx3S06Yzb0wA9IM0XunFu2FbmX2PeI4EmKdUp/vgV5rUmAqA6pcorV/GbVULfg5JRgCAYrc
dfejEFThoHYMCTnGfvtlNy6eKVw09W10V/QeYOnMOIhG4o7OUmvfO0lnqFLxnkhYdVGuDZ5b1jKk
PLNCin6utnZqBHtBk4salxbUUjD6+XTyvdIvzWd4DSFjEkFHanFkDR6VwHJWAsk2cpD4WQfZ1p3e
EaVDXwMnyQvHocaLF16m0RlNPZJi4vJRmOPZkpCmrVwpa0y/8aWKW8bkuu+R44nJyz3C5c3xrF0L
AUpSUoB9+jURnqj+NHWdK/li7XbMaIV4DLB4CcLxeX2KFiTTqzG5piZQhV9IkPHJslt5+UzdSptM
VfksyjdTHaXEoKR75RZH4toxQxVVa8fd9u0pmBqzKV2VVp7FADgAc9SSB2qkC0/viNVfPnyo20/B
eHmcTofqyAKUMxRAwT+9Gi0bs6+V6Ow6XH6pFOWHSVhwxYdD1B6Bs6sj2vTOmToQ5Udzw8Orou4L
C8QR6ZWKYfZxnirlVtQ9VgFJEc6q9q69jqYKTUje/pHFrGzU/bY8ExHn1uhJ9bP76a4Y8ScUHjgu
y/PNlD4eINyf5W5/1/yNzUp2cTNYBs3J403KMeNfO+xXfXHFC81MqlJmqfc1KBg+9n2DwAE1XUNq
VNYonWBAcKn7+MY3xgcSpe5xnMHg0O3F7lzPuZPu7ELT8H7jLyJQb/G9m0P/zL8PyKRRNPCOUtiq
mpFpJ4QtrNwktQVR83ywq+Wx3uQwX/uk5b6LqtFUi+4oqR9brlbT+gqj/Kz0KWgHQVHCCM9wdrhj
7q6tgLU1d70lFO/KBhC8fmAeLp8BmgZ0EiM26ZGtarBmEimv/3ZQCbMr+K0Xf6nJVVCilqaTodIj
u97Sd4J3lYK4w+qndhSbRJAh2HXTrdp+ogQa01N7cqVG3r19IBcjhkuFZHoGRC3Nf46emljzp+fb
rOaAg4zfJ5WCdpXKEP8zYHqTfNTV/LoBBSYvfXVRT77OH/S6Q0X/+QewgNImdRDU9mpctZxd2TF2
tOA7O9uYyZhVDR38UiYXNlse91nRkrBsPCA9Fm2amyB3t9Smp1QNoDNoGWEGeAdfsRr3e8uuskUS
UuQpL16I8Dk0W+qliuwQ4dxbvkZnv6FgHXBlXOybn0hFqfDJEZ5x0bxfCYCI8LHtvjjQp1qfHcsi
ZxI62gX6pbaFedIxwO5tiiGedlkpEQjB4Ih1CtO77lPmPWX5MZlFSF3plRvFrFKyANRcoWaHq8Bc
KTqmZZsZvagWo/ln6+xnPzDlHnHdEPc1SxQvO62Xgs1mMwnZCWrNFBfP+HctzR0eMX9sLyZMuuur
vBM3J507ZT43Mmnbgmc/R3/qc93R/5T7dZGsBgVpt5et4sdOopPPTxiTVhCjNUOh2NHmICC6vo3q
BZuwt91CCsK36smBOy4TT+oDOG++ePCCbGfEhZc4jIaiRL3SwyIIq/zg1AubCpJmJxF+HJIqUh0j
Eost/JIoxu0Tk6avN8Sn3s50Z9jB1j1iluNM5S2krEix8tm4/ngpAEJDNgWyCL0qbUWaZG/o1nVt
AiSF+Tf1nPI1tlZZEDjJ7rHX/A2dHv+1FD+qdRFVBsL51ve0ObwhIoqr9brjaoK1/ERy1nktHxl+
T9krxZyV7S4VQlVPla/fbeAY9wUCeL1VemtkhVT5Jp5tgatlJ7KEuHhFRrDA6VuLyb5btO6pSjGI
EWpP0Rc5pyyARsoyFE356vQMTv/zb4piNfPXYDUgnTCG+SciBTD1xsr24wJZ0bgnpBBkDHckLEFL
eruVS833Z/bU0OrovhBdJQsw2eGDf1D9zWpGLrxF+mhKYsebHEGiqGfJU1gKXm/gNdYaFVrHqUUB
icy0PG2iq/ECKlsaHkm2JC7pE+xWRuCvLdeX9ys1s2fZeH8Y5pJU05+8Gt+qOFGv9RIxrTcFk/c1
BkMS6/Q44bXo8Jc/UnTjXrNho8Ts0hZ9GLNTqes/IginLj5hXLQk+4EytKl0tx0W3sCe2pmA5dsx
WwgyVrH+aI5TUYUuumG5GmJivN8cFwADHupiWCN7a/mMEWizzuCJhLnp4xhhKxX1G3qq/tmv4QZ/
ntEKAy9Mo92Mr31Ae0UIEpUiQQlo1ZrzgDzUc2egMHFWnbv0uiabVmgCt0R0Bd0lIrcZPRC06109
QpAp3VfuvYkoQUIjxyNc+MFGvkN/pHt8RWb6vRNTWcZy6B36btTCYKv3/3vY63jwL+ES+hekNOew
YLFsABv0drFftC8tbeHugKXxmWZWAVXm0Eh5LZuZURLq+BMOKYLuj5TXIYd/4klquJ6uSrliQmFU
QhodBRgUkWslVU+jz4qZAjQGBDg3uLpTIRG/AHtte5fUlcaRXdV+ksyrsrKkdMb19/Aea3xvqoZX
6g2mpPvKUTizKUTlgr5ShDu5IrdPf6WinUJzB61cmorFMMQWree3ixSjrrxv1U7ufWTNBzdXnrM1
VKFIh1ATqNGPCv0mSNB5PDcVxlTMqMw7xvIF353MPYUXBMcsHEMLfTd7dDCpUfoF2koocDYYAGrI
Q+PjNLixyI4EM00Y/W/v0yziQvLSuiOXAm3C9F5spM4JH6FxXxkxnOdtuWVh5XDs9JEl3so2PkuI
uRkQmPNZc9jnq42g3s/Ms5pyhzBolHx7tUsOQNsjVN+J9pbiru3WTWWTL2VznI5ASbgtbjNhRTz0
WliD7sGNmDCXZbmh/SlHRcX95VRDsYPBWYnhtKGdb3PfU06UeSnv046Dlj/2mwnHMb2t4k3PH+WX
vUdFXfagW9WFTaIUFXpguV3d0oKZAyI7lbjnj0PH1QwuriLcR0IU7OABv1MqGmIGfpaDNE0Uy0ri
xd10ka+rAJx0rxxDGyDsMnwMqbhcpF0R0Yk/9jUZfs1IEK7EGsYIpSVbvOPwh0r/jYhHnbuxu+k5
f4wNYwFTlgYZe/aQXXKw7rDbYpnqiFffNla2lRtp1HLgeSJSRY5kQliMLuYdSUTjAypOCty32c18
lWc+ia5niXChlvdNw2leMK9N9GAwCo3UqIqc51G+yO5CEGy15WGeLwcDVizB7GeToY0siOvSo98M
4Gzuo0mXhjsYT4Sy3jylKcWVaSVhDUu28dLgPOQGO4lr43HFVC7c8406KEEgoHD9+LvcPXHYpVCr
khK96qbMxCDPxRQ38Fa/+H92L1HISK/jOMiQ0qc+CV4CYwxMm1jt1RaCCI4P6cvk5az/jDaKzaZl
qmyyIGNSqjUNft62Xdi+PGrggZpnA4MJN8dAKdPwFodt9gnrHQ+l4vvdkqLEgLhbMMfX+Qnrv+XP
Yx4kfKmYpo2uugJkS8hePAT7HohrxKGza0YaR4Jd9VstUhLjYyESS0wUm7tIJMT2mGj6vSByqAvI
spW63OxV3HdZXCQZMuUzoHnT5UcC4HagZAnzfrZCyQOkrPDS+RrjyjUj9Dk0utmfYWX5gX6UtFAl
AuBVmxZ7cdJEio5ZHkASnF3iuchDEE0rbwA3Y0+buHYFztU6PSd9IzpZQ3FoPcpowX/xyl+cVkxi
NcYzxHZjyvsGH/5Dk/FfIqU6rrMzIeR0+6L2DaIjHTNMGvXWBq2JVZQRQRY3fvYUgg/hjPMRiVH5
4vC6SWF6HA53Bfb2YPbGuPTBpCkD8lD96D4JUoUmNp9IG2Ghcto4odHWPS7G+WL7UNrWjWkDGFcf
f8+LtlSEcvg6Rg0PCBCtIeY07ViljV5/4wqcONy8xXDazxld1ig0s7iIOmmsOICxab7BpbZ3vtnU
OrcCE8nYV9bGpiTISye9WwOSV1HAp6rcfIk+6MnDe5OLOIGEdkHu2xB0JEIC6E28yBSCEeTObaWS
yCWxN8avOtlzYtrArCThw4JzZRBjzZ4ah0scKBuOCO9FxXF2o27xq360a0eycQ0PxtjMZVmwIQ12
QGe51TnsY6LrG5pi9qtrA7WKOyb4/tMALnvyq/AJ0a8zKSN4XRaQEg/zWCXvizHJ6/ewaLvwk2Gd
zXzAAmYOVidWGRBkkxWeXiX+36jIwlyZeRFes8W9YFEMmPzmOhkbyEr6tYQaBFHHTBfgj0aIcNVO
SpISJ6VqEzPnJH8cOF+0IgINsoepp5XRgXdf9c5UuQ2ogK44Kv/3xi2mi6Cirb8dIj4vohD0boRM
9y6qkuKEaKfir/UdRQEHnq5+cJZ2lpmr4Gx5FNgEkVzKKwr/Pk/gx6MYn8x+J2i7ytnN/LG8iiw7
K8ynvtrXW5fiMew5E+nWa2b2f+FurBaYJujt0a2IOmbpvRdaHBEEkkigOk1yXnmGazIGaT2YymBh
xSBgBoPBrBKawZJyryADHvFgh6NZjs2cPWYkrqKI/drmuIZyjPzLunDn4VEHaoVV7vAhJMQieH8e
Qsj04/iIfoRpP1quoEww0xjghvKQrxuTTYwmSna6dcGbXtTj2jb1RvAo/4NeJBbKtaYODEjyEEUc
BMGMjOD2zO/12kaJOT0UCdNRdDwwearGDj5STZH86cURO0W88SYsbstrDxuEnktJJc5IeVkqiJFk
vrSEJy9rUI8Z0DUG33bwW/kTaLwoN3oW2mDtM5RV2sWMIMapTvPz3KhmandeAeAxiRHaBT78ixzI
sHi6hmhAB3Hq/rHIzgzMlVMuqtCcAyO+yj3tSqxBytwRAYrZgBRXW0F/2HLvD+jBvO5Ce0uSJZHZ
VISIiv+rIhEyMPsxDG4tVsMbMEaGLhbxMPfqgfdqB/I5LsA71zEtuaesQwdvk9kty1qlkNqe0Ola
HVQqJIVpQIGOs0UJjyvHJwAdYuNu8sHnDXOp+e+KK3epBjY7jlpd8ROJ/ejPJ4DixLLl0ZLjmJXu
l1Mcbp5n+54Nqdpxw9WklIQFpGHABFtxtScwJmC3ETr3InExbFc3RcHxYsp3QsHIzOAxcw5FCHlL
o8JQiu01FOEfIxUaEt9/CTDzjJG+Egng71mdpt5dP3c0JrKTHIQvG7HGKbgc8CGggQ34ksTLsyqY
Idy6GUm0v/EnmWX0X6TUwcwZSpr+nmJRAbwYRsOs3kr7DJjGP0/KOipDb1a6WGV9Nxqizxr0D33+
hK1MJDUiuYlU7poi08apuZejC3oV+65GvCewaD1r+6pEjI4ThfYwqE2j3qJuRsXpn6Mu/CDLIk6b
XgF48dfCvThLPpgzUdZ6IKN03UvKheBAmCWqiFpeXzSuv79CsUHosH9muCYtJz/aFg8breBd1nc9
4xyGtjpumyokjG1SGgkPM4AI/4TffQ1XYbitPQRCOEYy8jaCWUAbq6rbT8KHXbGakFH5bVuX96nH
WpeGnYUZsCW1kLSuV7jSOwnYQtjwCP83Zetrlj/5W8ypFuBQ6Mw9bJgPwFpoGVbMmQd6bsSnmMBV
Q5rEqEkBY1Z3jTiftjvMYs9dW9XTIFdLJmfArl7bHuNpslN+/VHSMG6DsA87zHPIv34ivCQcsJSE
jHq2CeOv/8MKaPNLvKOj/Da15XNXOKmF7p/mkK3PEF0yytcqKy+qPOBw3hRTb2iZ2rtxFWzEBMTW
Ok10z2B2NB3XvngmCk8zXlHepp9bKZbBoWsq1ANCH4r4CNEnNtuo+uDJaXUd+k5ZzTSBA+1ucMvT
RUegaAteLFDXY4XC9PwH4rnE9Hdng1hHahQtjgXBew+6o5UnkOUoQCJUf65UZpJWqWC+TbJBeScU
lliIBaWVej8DRIjYYarItvFUyV45tnQrEXMYVBe9IOuprLv+NspKUK3SspJOfSkgXRZHZvMrmgco
9lcfeZw8mW7LT8tRZ8ZDDosjECztf1qfXtG1w4qywvpNA4m7f5JcIM6mbMO1nLuhlYIZaWefNMr5
NIWb9XkEUxQQ4N8we46zaXf4HqiVqhSyMNKYR8PItCXo7OrzUwdCxRLoslQ9Uak+jOgiIUhQAc8w
lZyLD/Sl0SOaPaz7X+okrVqIaQsXfXgfzNRsinqvzrjEzL6x6/VfpfyFLF75qhEt3Nzt3lUh/O4n
Sbhq5WRTCdbjod3pb/B9Y8CoLzcIXnQDwoFMIyXHUVS0kyEYv5+XRuEnDi3QJi55pGLtoorJW80H
mXH1PHoouZKRLSgA0zpYRE1ayI5FdYC66VGstE13OGiKGqBRGnhJSlNOfRzVO8aC2DFM7GN/LGay
1sbEO++Y0ZRyA08ldyN9XCzcoeq6nsVgoUnmDYN2yK6sHrRaV3uYSpZ5cdoKm2FuWvC36mrqKV4h
jtzF0rshEKcAUNz4n6ePbOoMK0G9TPfSxl432QXpQEgkQ9bvWXg8WccRSF5iPoI8Un22VSw+Ct+I
Je2HACgTRW5JIzMf2wMF/+Ww8y9x/NEEtxy7a2mXet7R4OYgq0dKx/MYdfORfWX+Radgms9/Fi1l
5+aJpbDa3DCU0a0a3qPQpWnnQWIObi368pO2Oomvtx2c5d+8l+Icik0F70zQAVXWBsQPbnRglePQ
Xd1vVp+PhzyCa78sQ22I+jVAzgKLMjK/fkOxi2XBXJIa7Dj3lu6Ju3OB1lF+ltRH5SLY6iv7YYYN
0hIhliEATLgwDVEiVgEMIvrGgmnoMFDULJA+1Pt3hPwGrXAx0dcd2hYAolQxG/eAU/McC1oXaMBG
4jN2pnsyKCnIURziP8UfrnnXevKVrO/ewDyNPFBzQB7dhvC6TVw7PB39wcFvYvnRWBC6X1UZfYEK
WEWkl/tuG+8apAGnLb8oTImkJPnQ1O2P4aH/bxcOuYe5A0JQ6wfAQjFpHkcdzle5TTqjeHYB+XzQ
R8ymUp6UPxY1bCpBWjP5rK2SdjwOKY8Z2Sz20cm9DeG+gQ5e+GPsdWZ0qRC/Z+6SkyexXtBdzO25
qpxNnpy0z5o2eZWqv9HNDpODDk6W7g1rJ51ZU8Rl72Yt9MOUqZsEw/fqxSgidmJ/iuPt58DQW8tE
ohawxLqLbfL22wjYyeyXwjBGetoDzyry4AdY39IY6VHEgtMlfn8pGS43MczWZ9BP1mFKVcHlo7At
BlTSfqbLf6LkwrrEqugs/YlzpeaqL0k1nWtF86q5EcNrzEA/Rk3NBTme2AVqRPGogZa9XMkTUyTq
iJ3v6r/DKwsfxAOvUsQs2ww+BJFFgmOjcvEr80po/a9IbJkVIQVUFwJkDsFEIWCTi66XoUhaWPCL
OtjyMwO1LKFIaeqcEVDzLCf9zQICTKNysZdFoimLFxMd+7nsA12xaAN2jvuCM2UKApSgvaPtdmr5
IGsPmBAd4nPNdvq6dvx+IAlZlr8suCJxjiUEhmIMrlWHNmMcXlQwGzl5M3Vee92Wy64asdjhWB1n
H9AotXk5x4ChO6OFh5DdIRiQ3XPVFxaGwIdaqdpChLZormDiS5x4UI6ayLUg4ShIQI01m21Hu9qm
tK/6TrG9zQo9IwvniihFgMApCh4jmbsUxYC98AmscF2Bet9QcFy6uG4v5JWkfPq4wdrXahc9x9Ja
/VKjhrjYqH5/g+OdH/yi6/vMK4z1legPzfh8/IX237qcy6vw2lRuJaDp0Tj88BZZ5Av7YKbjhZYg
BQICXaf+ojchaYslFfkzsR7x3fTIXzFL8eeedYnzXmbzOL/hgGMKGgA+b0c3Y7pg39qcHT99UWeL
dy2hdqPhcnB41nuAPwObxPwHpIrt/+lAbOz6bIM91gp+9HqIlereGq3wY7LC8i+nzPGg5iH5RA0E
wa+IIf0iYiNY4kkhxJE7JaJKm4hV8AZ4s8Jg4R1F4IZXr1ryKuxRXST+N/z9q73sBIgWkTzJCqSU
Ge8Cc3HyvB5sI40Ef68M9A6/9YtNmJ6LaqWZcOP2L+HOym9dcfxT44Qc8BWodDYzTFSrnxLZpCjp
1LSVWXiQ1M6DT55V9V/3BgS0vtxuYJTNJdEWAcjtKAqGJM2k6v2aFmh/fTL6UjiinxUDsTljEpce
5muUOGgc4RZxImiAPNrQApgiwitxsFP8/jlSeWXiZnNM1VSyoJppY3PG4vt+bmXx49PlKjbOz+Qn
Mkg509ilDbwYV4zLLFgTBZbv7cXh70ktyj2nKCFLskGC8oW2Z8+/8ybaMf+dR8hJNERz5u58ipQM
hhQ98RPFSnWMawsSfN8+tZO4Phd8/fntGnQpuROZ6vmKi4wJrfhR9cqcKR+tbrhCOdfdGMw1zChW
QKthguBpuk1gnv3KDFU3gLyEnknSeUEPOfiAiLOT/60sDKRpn1z9e3irKcnHRChrkCxsYkNFYmah
Z4+dllAWNqufwvTgq95b1+v6pY3rouPVHXtF06umUHz6AQ8P9/0vKUE1HamhROndLLp9ja45MFh5
3i7WtOhKf79OMvWtN2L2mMn/kbqaK8jlZbBHKtiYZkcSeFulf4GTeX9Hl62k31JxFcD7Hnmzh7Hb
caYVw9lSWMIhvpeWuto2765aBuSChY5JHgMq/GC3zXzmRQ/PxYBPYHjzVqkmlcF8wVMT15AhDkGo
k4crT79umLQUbnmJm4C0eZXOZaWC1zXt8sPhudKo0X64Gc/tNLKVy3GPRfDEv326hOmhBgkGbvuN
VrYBRX4c1e/xv9QELhmcvlJMFr4dGZeXiap2Yhi5iOBzCYenPERTcqqjzLA/1N1mr8kRTTzfwzX1
3GiNqRwGQQGzhjoNvUA0RgBUEYDQBQ27KQwMnAr6i5+zwr5xasnCcM2gzGRIUXdk94neqDpTiTrC
qagFyVZ/FPqj/xh08zzjDaC/j6tkPNoiPpRo7gJNKJbVkz6Sq9NOCXIOBYpmoe3nimc0zHtOpGGE
Ngh4qE0IJPKe8UuXSI3Iyw25zWM4B1Dtt9zN6eko9yP9khtSA0y5a7zNQog4EEV/Tb4hSim28ta1
8LWosMoNuWv5AC1sbycW74yBSVdaRtDGEEEVrC2Mtq1qQhV8dXKwajqlgLTGvN1KbSdm9BSVfeKg
WZQWBDrl3mSRvmus834HdCxFLkelTUcTb37ESv852MTZo26zi45/sribTFFQYXTX5Wfm9hwDqvKw
z+U9Dlh6z3xzv/6UurCurE0BYa+q160ilakWlT2q2su9LRwX1N+2Yu9CzB49fdBQ5jseDzxeKKWX
5mi7xDb22j7xtZ8C3NWp68+vEinPMXt/7gLiXZTsmYCPyFT0ij/DHniJr0vgAuVuUKw7dfaOu+SF
9CfHJDnaJ+SbDijU+nRNOFgsWzHkUthP8XyZoL9OPHvmC0Xg1zqvR9/KrNqMW57LVh3vWaquLFhj
L4cmYRWdvhyOEDfBduMXIw5vL9qocMPFaUXH1br5GyRx2qv5ASTBhWPvUaIscpP/e/YXvDtnbf92
QASTMu3BK0e/LyTiNxbHmMZ1mV4D9BkYS4QncKJ6vwCXoDLZBNwglp3VJUGq7EKSl2KrX3HWLH+B
7VAOrtLyILJfYlsoFps6qZDrMb+dPh11qCyPlefNHTZ5jTtKMw6QQE4koxD2eca6pXFWvyQesY8u
IdAr8ZDcx1gTfqbLm0zRCeI3sNR41WMHS+jFSL5GNDtGVSHcKF9jXVd6lF1JepZ0kjEpq58/kGrW
pzxCXffvHxCrXT+hgyS63MhTyr8Z8rZqWWYVLlCHU5TnT4BIttdCPEGpDHyxWz6gNjOOX+HgZrHd
LjyyfQgA7YQ8LhyKWUBRUSPbJ/t9HBNMubDDu3yGyFVfJHn/j8JqXAluhxaZLPO6UP6sItB7B3cP
V+aDND17zPrsN5e0c/cTutNerdgwLQ5O8C9WjlcwPs56F2JPPifm7pwrNJavqIYtnPWUOsb0YYDt
J1+7r4WlpB2XMCQlqE6OVlZLdFDNHwlADvHyJ1Z1gf+aTom9KeUTPf8qo4+YgSoXrM3vfHis7krd
cyxr41QxR2ptas1tb00XCK2YdCAQ/1X/geQxfqZfDopaptHT9YksiFSffXb+/iXFiSv3v4Wj5RHP
NONOXFsk+XkfqXcEG9Zod1aVofvi4fK08bTIYdCqX8/rtBY2dBX79ypMiA0mv1IrnZzwhFUVx8ZL
U+qpblW1k9v+Lf/RI12HHcRXWAzzEl1Pv1gq+xcOtkrmY00VsOGSijZ3/31pwBvkusU++NziGW7Y
BAKvn3W705RG358jlR5MzBPVlY1qycuMnLvf3yUY6CCIaLWM2Fs2ZSAsL/8zqUueuBy5LVsq3c9o
yj8UWMIwp9oFXWsi4e6p9L7AariYtzjNCGqLlF2seHj5GSh00Uw7MrYARH92x4QZFSrSFTsHLdbf
5eqmA2Kolwi3JMaVTFzTZ45dtXJrZby20ZSvyaLvZF+ti5f9KHcn3AjMY5yGLK/VTgNgL6Ufwsqm
RsqBHsctFvTwu3Gq0aaywJN0jq/W6ltNSuASDdCXnHRqmKsH0OqF5d/6h0MbW1jX5Dn4r6insvAd
oE6XC8+bb/NDG3ONaq09oiYYnENQw3vaGi1aWsfpm+gGzvs1Ap3i/oglPnUQycjjhtM9/xGdPoqT
/XKkfjloO/dDYDXMMrXTXldOpDueYdxOlopQ9kmQmt9Xb6YlCIAskyPirAm8Xbmj6lvtPt1tY3Oa
sD8Ul6Oe4vsot6qK19lUCKhZGY6xwyTu2wBtU1CiwSsfGs+FypMFzDMmA7iCFOgm+yWFR6WzoHyc
hDXhdOZMg4N/IyFONUGfgU2oGsZxaU/iAP2YZ6NrFezhWlewqdwGQxSvPKe8eXf1QF9ggEWMiLhC
mnTByHtmfcw+lMGnLalhwZmMCpCfTVXzPep2BKvUdWpCrmiBhLyo1gCEwAluAWtanoz1xH2K7Ox4
v8sEKOnbeZVe91Lgwj3DucabxuihZJWurzVlRqZiXUTx5m3uHQ/StO0A5Y29o7pXvTYABWN1GIBO
iaqFkh/7wUZZo4MvToWcp6cdC8s+xYsUfocKj5oiV3SwiQ8/MXKkFHdzfkF05JT7hNSy332PX2Nk
ieW+T7UTHiayFlc9wasqAdxYYV1byApMImRF257K781f1dCi4ATmyOSq5kpeP1J+ldfIgqSYPNy4
Nh8y/dd9z60srh8BWRzc+Kyu0/Ga6UoQKJi3zrpsPG16wEK/U5mrvTTMZzIyvHpPSkoQjLLFqiMe
5l8aGR1CsxHyBdcR9qVzEbmtyudMQvd8aWe21aHlTqkJB+U3/T/TqZ2grb31nlMHJKuHah4pF7oX
BIBsroWay6WdUv8F3IxdVC/+/JYfsuwL8djOrCbOOvZSv4tt8yCmAMzjWf0zPo43hC0DhiKqV2LQ
j3Hghnw3CeudTD+eUOCtbJsqw18JduJgQuGsiYQzl1Q59pNmNC8OpgEngD2Icei8vIS5L4iXaueM
l3ZiSJ9ZMxVJPoe0bHK377TtKa+lsOFe7YuVdBNY+E2+Y9gJs6nYeirMlPqU6+pmwA6H/ZO0I2Op
5hkkbiqDFqXIpGgUfuQJ/sHQaV0UsYkA+uYqFUsyPafEwVl3T4aruux8cTypXq30vqjhvAKio7BL
ybAChhpFHPmJGVU90+roeatamMrYKrhQb/VQfMb3+VRcnf4ZxUNHnWHjUhWDib0Jzy2WCfZ5TcvM
cS/wNyWaxKz7ZZ3+KYWRzWWemp4kaaX5wlJI4sS/6ZW9rOzhUcROBBxaI6SvHSjTc7lH8CAs0F6F
dR6pgj7yIU6opOM8CSboOyzb+OXXhJzKBpMj0IAHlvucHKuU7/xWkKwSQWIAc0duPVdfevucpQn5
XcUQF/GEzpfbJwnZkB1j4TP41/5GctalDwaI9JfEAju27nqjiBXG31MG3FVjBgcdsKi9vwfbFWGo
/BglUG+sL25mIYceLKiILvgqVKcuyt+KgsGjeVUD+jI7J6+iSealx5qQfpbjKYaykoRcB8zJ6kg/
BqoqXWuwQai9SIkG7lEV7p/59I0L0mgmJwsd5BW/LTGSdP/aQ5dZZpEYaMT+d72dyqpbRgy7lUS8
osXB2cZqX9gM62GFnrUaJHOV31g6oCoejdMeVd5E9cAW/XAeu3NkQhOVzBnJiochJMSdjVStwECx
B5bOBkVl8yorcXeVjsofHXNIu00yzd2HkpXviQ6F09zLHOJN2N8i31VlD52ODp/b1Bg6oi9yLYB+
aqYsacyI4GJiue9d1B4EKHXw7JPa5eyohywyH/UWpltRqf0ABhab2Xp3NX5WTEq78wvJNOruHQX/
xsxc8mpJgnD43qlez0CvrHYGK9LNOBo9uUG4O0JXoCkSQpnVUM/NpD+6ogkh1fWAyBrToNOj2h+8
9AEoxf32k4PYzy6vLsX9YP4yslgppUfoZIvo5y+hvHLz1iZE9rFNTmQafLVWTzdHIMaHfaHmgPxe
UKa5vsUfer6UuryYkpycrsuOKWhBVv0T8QrT9qmUcxUM4Z5RPXs5sFB5rky73aklVtCaeqxkbAvh
+amE2F5W0jNMAH3OOvaNQQm+1RPYU+J2ar2/R2/MOMocpfmcTDg4O9Wq4UfVQmXXNblsnIOOmH9k
zzf/9WF+nffTyxshIXmPnnj58EmBQ40TTg98pBY/JwSI1kMUdiap1sY2GPTJQeVFxOLsNrEgM39w
wCepotrPQgoDjkWjmkiuTOQo1PK2fkNMZRKUasLtE+ve4TfJ/I3FPXplkt8HJIXltW67N9LTNYJd
xklV5rk4rWojp35WfPhyQ9ac8E3cdORl9g3l4+prCfs05xhuTv0pSWuR9pNz5czAwMPG/oc+Jzo/
xim3BcbGWzW+xgLZIBaA0Rb0um5x4Dmq+zasps+YSsvELTyrR6xqq8bjQBL6mcVsPAOZKH/Lh2z7
vBtPj0VRg7kuewm+ETjAMQX8+Z7Xl/VE53XAwBT4zkq6LFNxglCricDurB9vteET6n5epckq60n5
Kb0qSpH9UauC0yCw3XTCkOuZnJqIsOibXqdFXZ1noy44psdrk3uvyWIrn4dAKKd4O02m0+0eMhQr
rlukyzLAtpekQw6jQuNGoh8db9tXtTjBKuVrzUmh7Feso8EGji0Q5nVRnS9/TTwZG0Ac139z+xV5
eA7JzwMQjxGKQ5dJfdMBGV92/b4k4dFleh09aKKczffj1dmOz4tmTtscG95DEjQ7qprfzylwWG1w
A1TMA0Z93rwsz4BxLdqdLXCqrkLOnAZ09dM8RxIvs9An+o2vOQVUpF3vwEfATnhHSJ52GAEgMYRJ
IwayPznAuxuZJInY6GEozMllqwQ/U16O3M9jA+kadsQWm5G0CTj8ut6uJwEufiF+Lm+pscbwnnnb
YJJhfkzE8vMpQX6PRxPsaEsHtU7HCyj/JyFjwzwYVOlAZ7lb1lmPquNpfzt9jva/taeCODs/DPwZ
1qIR54dUfMRMRWCvBaIpE/qSMKX+2BTS/2D4HAMpo6FJ7lC1BFlFgPyh4gIXyPzrOweHYBHDiOjS
iqberqKEOlUc2isHqyvj/1QbPdKmbtQQ/GLjHLNSuMPwKgUS/IDmuOmxN3y0jz58oeP/KkzJ33F2
iytRL6A+AMRzgLjY157BQA0katCFAOJrvYVOoinor8L3TkZofvjuGAKd2Is9WPGPMhE5F6FcqVNm
nQRc3fFMoejj/lP1N1rAFqbWK44wpf8s6rGMnl1hPEv3xesSQqUDMyMnd67innwHK1p0GfyPimLY
zq3+5aArYf3U/5w5vgQG1kw4bzqVkYCjm8PX7OeH+lqOKMcdxCTXFf47e5tGjv0wAMuPNMhy/xQe
eneo0QPc3Dl65+korgQqHtCS+U/ls5nz/mqyM6j6NjND12FMCmijU2drL/BoMKEDj/85MdjDCCq+
zf1eciLAgG7NggvVP9YSVcm3gf8w/UYr1mmdxOT3GPN9cKaNT907qZv6lnHe8CXes+XGzif9EBRF
uqIGtqugiPwUAwSWDt/c9TmBLvdJ+WawNwg/TxXYJP0/zN0aql4BJNowlNwKUNIUVxwcchEgspZG
pLAgB9cSxtVtn1rzmxZ5qlDmjBz1k1lJ3DlkgmbCQKH9piRJDFVLAObbPAQnt34HV8vFtlTEIJ9/
JH09hJ7JvIzL+sAmldedizNQveLIrkdelMvIwoFw7oQ+cD4FILKS37eV5PTiWPvzw/BC7GsD+rR3
wr1W1H9jEQW2vRW6zVebxoH8QS9G0JsFK3nuYKn3xZCe/XToV/GlMhIxkWBOH9DnNxqo1ANA+yf1
6kQqd/IrWUO9/2WK91RZrRq2SBv+X5i5xVHaR4BBhASioHV30TzRXFodyhEvU4AdbZI32I+/myBf
9VE0yZXCW/SLTwFefQyUECVmmrXyWNKT98Sn3Sz7KMb8wRLNuiUl5XltH4ZzyGni1DpIU120n8F8
owfWUoFmaB6SC2a0NVYuIO/sJzSVC58p2xN6XmNUGep0NXXFn1emwHzycv5YB0R+92NcTkac539z
xBTJ062+LhGB+WtRDmKmdjdLnEHwNABmd1ql2g1XjL9Qu7A0u0zzsVv44BKpglRHmKW5F8Ejylbh
ocYultF7ld7f5NWU+NTeSlLTvNyb9Ot3qjPqnE6TNYFMPusvSMnPdYqR8egheMe+1mfS4XfC0bRU
JEImh3Hk2YS2OlaMSKLPf6rB5FW6yzfV4OgcQpEd5Qi9Kzv/VfmeXM/dpu9kDiiYYnEyeaQBApCR
MSNkK0uNZZT+Cy9jSow6E/WAVmSeVrxUWf7DhIWvdzdrLT+yCDZc/hKVc+IhFXT1Be0EI8Y1mCl4
FKCuBKuz6/9htjH3RyKixZrdaCH8TEC7TlribXp59utsqNPwB2sgz1GFntoKxHB70e4nAJ1Vn5d1
cnFW0hU96JS9rQQB3anLSxNcWcccI6Q6d8vAorbSN5pxePZib3zDQM4qWzbFzARV1HsA2B5nvCuV
qzajuF28GcPrVSlKad3QQDBaDbs3FLsEzXJXz3keYmqbOIYsUlvVipRSR2HtA7MDSNieejUpuBfp
X/StOAkTKFV3I9ohkI7hTLFa1EYaULYavynYBkTI1utoWv20z0q4RWRhSWfgoL3AlBqOHy46Wlny
PkE5G05iUYlK/zMhTVPWlyhwlpuFKmDiTbstIeVTVrYEHO8o9zdl4XanzXxIxr7oi9F9t3nh3Jly
zrsc6WUoLQUPg3gRchHDQI+fMLzud7OmGJg8K/1v3dMhHFH7/EqApsRZUyTIYiuJzxEUsbh9HC4N
38HyTS7pAm9zbfbtiUEZejEDx/tJeEfl4OHmlBcl1XNPoBfaIW9MPB0EQghvFnFyU/U1Qm+wZSWu
DdEfDx/uNcienIbgt2MPSyHdTIF6eKtYirwDu1sU+Ghp/gXCoB1RhgQmrOZ+H2vHm07o17044A9v
kMenwMktg1J2UbfNEKYZlAaNSoNneEQOdR62G65ldkh/pShLxYFYRprmVyhGaRmf7Hq8qDrt2P3Q
HIrvFbyS7ao0VEPVHDxOueV/bJS2h12FLZXhToCMXVkC/4VaJnKTjJ5VPH4P7RF6XpCe98EvEV9Y
Xtgzq5Yh0tCpOlZwvx/8l7Gi9cYPa8U2Mdw5QksKgYxTD9+I/SvFjaY3FhfBxfytsaIkQIcYM1k8
vLqZwVuPRKjuvLZPTJpJ+c1YUrAYqiZCU2znu+Qna8mZSu/FvjRdbzY/BF7WLK23BiOqEyxrXUbm
9MybCHSwpetSXONtqhBRXy3itpHGgPAs/bWbvD6tO9UoQn96uTHTk0CW29pM/CO4ZB0MIp7MgpnI
9r94kCrEbu7iu9NxQgmmOvtYSVU0f/Rq7C0mcOpVeRimhmW3Uil8FynlXWu2pOu5ch8q09+SbBaW
1JvxJn5ivkFl42jRtLGCX1AaQvIsPbLFO/yhxBp7FQLlPDVHPZK3AnYahf7WLe2JL3wQJQmJdOnt
AGe74zInRfSIPSEtuyJuY4jfiwC/OXFPF1sE/CyTBFTdDtglJQ4si0sKEQUX1crEjTHDAf1ZHGqW
Z0TUtELq0fUXJl9uUwSmr42n6Ih/tQCbZlQL0cZS52hIREob6t04oTAm+V0zpZR9alufzKRjqFMx
j0A5xprObfdaYrrkaWeaykVkCEmZ702DmqzMyXaG/iRCiOoLFWC4iCBGiHlp/NnMbvZu51bjEQSB
PCL1qxjhzoJALIkuQYIFos+kJaAfRjqogms0KSB0KvMan3CQMh7z+AVyilEVgSsYonEokQO6otcn
ep3yoqRBE+MDQ6WQ+6JeASd8fhjQDDokzdsStcbDVOM68h5bJ6ulOhH3I6BwNCEzbKvo7Kw+qP/L
fZ8/t4fKFccDbdUok5EW9TyWtDdylIEOwCpczB7fIO+0V2tfpbGlkVNutkkqmDH9/WlhqfPP3j2b
bK5Fm8WDv3wBHoL0+FC2iHg1AcD3vxYI+AZo3I+12VJWyC6dm0H59pPPbe1C2eOTKhxl66jMzxQ4
aHKP7Q7dkb+rZOdANzRoGnuB/3TgpR8rXSC9ArNwlASQD1/7K62PI1BGxrVhBj80hVFfcy3N58v8
JIlAhzO0qIVxzAzO9IJrkgmhpMfXabnEw1Yd3yEmZIOAxNEFi/5yje4n5ST9c26/NBfHT7KwIyOp
JFe9o5FMrcsEU6ohwxlHfDfpaXO6bBndp4sGmMYghocEUOBmMt67/GmjWIQf6ZfU0xJAfsctOk1p
kgzdOV3ouiMdzQp/VW8UtJq8hzbt/A3E23RPLsWOa0TN+zFipQy+V7UfLxJgc0I+p1awEejjk5v4
UHyPYij8OAY0fdT9sqUulQ/0MIgx1BBUGy1e2D0jyC+nUyXO+NK5ZZDD6wiXUQVyVx+abfDgMn4F
DgykN589rR/dQqIRWZu+I1F0j/vUgJBJ+WMLNivdQ0/c4PPBLMPM3SLOIZ5YYqEoPq+rWnGF7Ow2
zA0Pet/f+Nf74a2ICnDQ24P0UyWKvIgOaiTAyUuxDF08lfvJ1vOzZChfEdzjNZhrKlS+d1YqSkqu
OMQJYRZ7hjTYsiq8mKuN+WMscTdwsJxb1uAVRawpJJ9fXfnBgQ06zs0V6PKrU4zQ9qa9MPxxVbiR
UqmTSbeG19aNG7vaU8K6GgtVujKUqjU0sZlVPcV1kJ/u9XK7QlcPf9UVP/s2owjBQycy5J7PsmPY
z42iqhiMg/TjkSphMO9i0+Nq3Pt+Wma1K6i3XNVYfAiTCIecRif4KQqirqLUU4n/AOu4Kpp9DXH2
9GuJqFOyLVd2tTO/Pg8qsbOIX/XTtRaclBXE4zHLgdRr2Xxl5aXo2TIYywRse+WuJfk39/BV3grq
Gy4AjF2vJ2+vZfMvh6W/wUiPVHCYQpF/k1Kj38+/jSvSH0KcDEVX0QO02FnTYfZO7wYs9YJMVQtn
lBXMulpJVi3BwAf+v+FN8BlbsDhej15fQoBmhHMVCZY7SP+KSv9mWjwJxBez2gmiJMVJWdsJt/h1
wVVGwdn/M+HNJLeH/TwdP3v556R4UHQgy7JqOfcmY/XIx8PQrSVvYwzOl5N0YNfHZ1qOtvkDjSJX
FUDsnNmszMTJvT8+LuQqbsWZ/mPLv6IM1t1yzH/ljebzHwsfDFlN4JJ+IJYhCKOO9L+0kyT31+Qn
kpyBHTPlo1AErWKWqXq0xfFvQWJCYzanqySJ8m356MVe25vHZegBeefeISIxLx2U9+Cr+g/NF+Yt
URHy5KGFcVe38loZgtaZJ3qp9z6dyVm3HASO/eGX/qzR/PWb+o/lWXR2QjLboaV196rrZtnT0ENK
vOaWShleWmpTQxXQR3vP583Ll2q/WoJOQpgI8uGSQMgYle6h6p/Ph1MWQ4cgpem/yoFCWia41Ny8
1ziSaslEN7PIarUTa3c/ut59XWC4z/an1Sa/KMemc4WeikqOCIb3K7ntrlQEjbqrxkcUNNe9ausZ
fu4cmTrV42kJeqkB1Lx9bg/WaRM+LN/xQbiTsvWGN+p+ChvXiJApm5WB/W308/2PpE1yMjf2yytt
XvECBT+8wJ+OWTuT9xcboGJa7ykWekz3Xhqshpt1SWzJ4swqu9Tq0emS1wTwO8+jg23NEs02NuVG
7D7o9wt5NmyczPi9v6zoCt9cWaafHVmo7ApEQVKLXg5HWRG2lr5oA5g1PyICJ7s6N0AQkBrUxdj5
1zsQ9Jc9xSP1WVuknHhPiyaPMde6MinUWoko81O8qP6PMqCesQ6NdcwFwXJ1c9t5o9T3xxi7iqlw
/nXa1sQnu6KUEqJGgjEGo7iC5uWWtEqn1L5BRmoW2bW0DnuWiZAVIZxnbEX6ETAurQebFHU0+vE3
XRxYTR2znszkCJRzFBqyAAMIdGIeQodIShrADoXHRs2T8yTck5aUe6Cq/oDoaIi1X5wqwijCaRlf
mm/xvn8Hd7CyVbSr/5sD90Ibjaqw7J7+RMQYpB8PVbcMIXMyJclz0DIJOurOd8HGoptWTWjeTapG
ZvavhKWsUeSju8iq7RDqfsrufrtLTycqw604h3pzrmLZnBkjlF6gwV+wmpKkajZhLxMZSeSQ/U6I
pO+DFOvYZap2sNpOUBEG2GzpuWCClicbIC6onRMo5KiIOawPd52NpDfJ6yS9/9jzNEHeehHaCBx5
qEeil/XhGKgVyRjQcEAKdrzez7F6Pm7Wtr7J3pSKbO36fTtZ04oHNrFxWz8z1UIFon54yY2OzSvy
fSN1OO8WqDT9X3+zAGSs7XZPpSJRzyh9ikTIiTaMTxjgyBgZFzshcOEUzLZ29+YPidbP4jeU5wwL
RxwajgBfgtYRRo2m6awJv73RDgRBXGv2RTp953iTUy61bnESxpENiv5YnT4zJqFHSGIoOWYpfCLX
fnkE4HJSnLJUpEo16iNZRJSFEY2euMHfLMxtHfWL0k8zrcRC0P11kd19vbChVBad7fb04E1kWQpL
ORoXrcnwc+YAEqWNtuT0h82eH2Iw29YOn7OHmXdkd/KqKZQD1TR70dBklhzE3q5E1j1c6tYmzPZz
SwqBYpcL3kqKgs5GMyom77izeNlyaEXmyJsBydkFzKXwFu1p1CiEg8WHKmZHdzep/LORBd3fVOax
CojDOw765da5joH03KQ7TNI1IoBUjcODPFdX+CdFOiRE+qbsiotJiabXjYujN+1dB2q4JAk5odxU
0Wk2Ybpyr66SKbnIlSMw2xX3MzVCErOu/5u0izTOv+1IJYZaCea7zP8iKVLW13/Ze5EAFM7yzVFC
/FzDjaYLKATcFfjSX6hlrMj2CR2LdtVk4vJDM8q4R31tWlNFnvJDk5IAdoe295qJ22JpEkjJW+k+
ha9yJWtYI4QtW0zvtiUAb2j3+4abHLIcc8HNJAlUqcrTE9ekbCwdTyIQPenPnXjiq0zkiNtbTiy8
2p7ybAFjLvFCG08Ttyrz7/Dvedtlrcu0TyuOkQmsBAV71/GPdavHH962IwcvPCD9/q/YaLNcCvVq
w7kqXJqf2rSYLOPIClwOCy/DS79Y38BhwhoqSpx+zSvqbn1MCYadtxEGbLX/8uOEgOBWOUG/lKB4
+u2IWMNfFfyTr53hYYLxf+HfNBlX8e4qzUF9KyaZB+uwpiZ8N6QACb18ESaqEXEVImIIHFhgI5zT
gbDpBOH/n5Nwai7x6vR2OlFRjhX7sh3Hd81uZSqd2fd+Hun9nJQQTNRUnduDqUpy90/tDdYnTwDn
eiWwATJ6APmNkP9DGZBOm/NloGyqt0wneT4x8iJuSWV6f2GfZqn9bMzHZPqcxiuVcXFg18zuVAsw
DPQVkMc7a8o5fCqUX0syFbzjQap3t+OX1ptBE6IjJj2xX5r5anyWSo3e4V2YXOtJ9uZKcMscR26P
x3CU1scAK2cqTc7GV6UWax+VscayIl1vDZt7PRNtZnq5Zo+Z+yOcBOlUBEaKT8O1h2a3xrPux78J
9Rtuhjx/648ZP0Z2iUgzlp91/OX1TvZCR2uV10B9zN+hdENcp9WUQ3/34Z/xtgLyUmj7wmgUlP6A
3lkkl+NnWRIlFwSVukbarEmavz+pUohnYg0Kp60WAZHscCjCUwJW3zRSH7+gDpvSsw52h3D/SSYV
bfKqCuAFSdG/vaTC5oghyIgeRVAmZyncdP6b62sQvIfR60mbUNllobFzRGkNCU/HdNYzG3OSSByw
lJWZHgoxgEweoPRqlvkg0R4HZ+fri8niXa0gtslR//5QzjEuBYgDm/FXJFJYVFZg2ttHuG3kOicJ
9p3nxNOT5r5Htk5C9TVRVaX2j/x84YJcow41aIalQ/ggSoSpu8vXaktB/QrrC+1gKpJCjw2p4ZER
BuZxnEsGKTvolQlPZTSxcyDwpz9r+1RBcrEDO3I4UqPAZwWgBaZzRf0/2pYKkljKRu4IhlkW5avM
c63q2vXm/JHeNQldzo5mlYaj3Z2RVPWiGFKOevW9PEb/OKJ7U/j74VEDNVFXlfzOgl72fVgZZRuw
gfDoF2SxjS4P0h+94kI9oBayrD4bGtbRPSNb1eBVP9dogP2ZcngZTyHHrtrDjAQBRzVqxfV16lfQ
K4KEZOyaJ3mJq4lFG4dvWrcOyVnggQLWLg/ulIljsOs95ZbzUixYUHlZQ2JjU1hOPBLgMj7CMsxR
0MVYD4kgLk9p+/3rkElaSPz5a/pwShIXwGvujkXxgAwYuAZnqOH9kYxdiWQKSTqwe+d3N7CmQPsK
QpM3qCSIeZVdveDhqxWGmlj5IxSkv4awWXAYV4nBtDICP8RX+BZ0G0BzGo01lNcxetoiBq8p8Zvc
xepTL3L19PQP+FC5Sa78lGf7sF1OEb3VTvCymiv9WH3w1PeyymAPVvLRT9W7In+QyqNyNbBZxUzD
vLWohcEoBPCiCuRqvgsLqUdQSfkZg9KCR/997oFC9jMvbhfR1IwM66xWHOPYiLkbyKh/hFa59+Au
1jk3GzvyF9W+7KoQSzohjNoZ/vMi1ekp4VXT54SoMnwZrmZkY4w7ulHtd43tQ4+ipeynv8ta7ciR
q7+5l9dYhb0iSkKInM0KEBHSqsyHqbbN2yAyQqxtngB4nIHDm5HNUTUrzu6fwM0bBZY7ubNKg07P
PVJbVvYGMOtmD4JI2t0xbrUFI8FFiuGNX92cmjNOa5QO96l5C6PI3MMYcPCVr6UKCCSjuTIdRPMg
LNBsmedWw9TwYkU8jNC7nJr6ATZZk/GFZYBgAzkTPF3g8RMAS46wD0lL/Vo0aU6pX30aGIYAL6Ke
/Jmb8lYgRSxubRTSoesFzgQuLgsEHSx1Cxr7tXtYwzrz0FGp6umMb6ih4vS+uHQCo2Wq9K7oi3gg
dT/Vx2icMymzINXBzQPqIViU6yY9H5SJEwA8a4rarTiZ12JblaJ5R/j2ViIw2kfZUURLsVCXXOpI
lGMrnJi/6XpfzzFcJ0g+jkTWoJamv/bonsmlOIEkmtqoEsdVcM5OM00RcbdWgVQkTKWlSypqirN+
OYj17BkZA5hWNKMA59KhBF1W4ID+TMT+kVfuSouxwTv7sPA0zu2e+iuVD4ajRNqS+R/KOhf4xRm2
f6mxQRanNmKpn2uLaG3NpRwF19NTBHhIQMWO2TBo5pt8Wmkq0imPkQOhYDqr+6Emp4cp+EsplKU6
a2frsf2RxAPrvWDBF+GPFxAtBjrkaYq4+K0Hl0IbyXHK0jeq7TmxamFfEnsIFZxfCCsXq+5WMwNM
MMS15wQipDgOJ2Ah6hCv7g04YC5Wh80QaeG4QUgQzIAieDjhhKv1OHI6fLNwdhq4q2RxUP1JAzNV
QKMLcO1mryTbvEIHPTPGFqDZwu/arwI7nlc0N+2uKPcndLj+6XmXjBMQ/9jUNpmgqbscZrLPTWsy
TZklncKHyQ863dWvRouoAsOx9rZCUpPzxWOQ/Y6Dg6fafIbYu1nyDQ6Q/reaPAiXtHUl5Oon5Ysm
ixBff+HknnnrgCbll7IZIGm7exbhlXnbvUSqhhUWO/eXXWp3mqUaEcKDYBJPbGNQ2xjXpA0IEvKa
7bwXVGJbMnWCHUcUMkUb0cOQ2vuCDukUO+Iha6AfNZpdsy3w7CyAx3FaYdJPloNhr/T0NwzDt1RQ
Y7E8uaxOQhMV+16bqPZOvBG3kq/4n87RpsVkCgM4K8PaXznEBqOmClSUG9sGfKK2SATmOnYH9Okn
6NQGxqlmn5e5bB/0V7kFotRG7+8SdgZzz021AeP1nvhRdzO9g3HAismQqyOflKTKf++3hzopWR2A
EAhq7GUoovraHANQcxqPuh8oyOeqW2K/uC2dj6VVhcOSl8hEJsUA0ehwSIGpqwKGtbCan1lH2JJl
uKgKeD+GTGcy8F65rcSaYvXBCPec7khmwt453AFMwgeVHFIwy9nYZVXjXXRZNgEruJKKDwo9qqH1
ouZh5gymRNvGscZcDHTAM1DyXYuO3V/x3GNAEbKRP5CASYFjIc2DxF9Q8ZQ/3XIZf4G5tLDCxKd9
DeTFF7wSGjUhyZxBDrDJ0G2dUiU8YAoVetyX3rR80RlFkuEeWK/yvc0p3Ser90T0HVRTsiAduCkX
d3NqjIygzhkL8ZE8c18LYDfZieOHZjPKRXTJiAHd1D4mx4sZLZmNxhkZg+byQ0wF3umBQLzF0ker
673SHvruC7076qX65ZhAhxJc0CN7x8boDxADEQF3uWK8qooUXqvsnkaIlOTMDhtokjDrspFn08f/
UujJLZLziStQd4COXlFZROp0jAGEY+PpJZKBwDQuXgYB+D5i6bLjDr/t+0ihyeESXjFKji6hQqAX
mzpjyldLS+GKIOcC+dQuVaUlb0/bi2/JuEu0K3ypaGMy8WMgZicXJPSuPVH/wjfWitmTQ9BEVSEb
lw/dxdOyruOb6vZ4lCy0yJ35VT6IasLJY2wmW2Pxd2W7fwE3ZeIUSNbexgBC3lCtnXZL35KN4Te0
sR7F7V1rU6zPZFJkxt3xibuEMI+OQAN8uVGzY46KBxSdH6XLtCWh9bqGyUAtyKeiwiLD19Nt/rXj
LmJfM1n7rlu/y+YQT79Jl19cN+r1YLdOAKEkIArN9FlyJMbvxcWV+fHpfbaQ+GVO/7VpX+vZ0xzW
zuNiAXvMD7oZZBCLU/A4aLzDFrfeAGZBXAoNeNU8FC/HsleVOATv4vf/zq9zHUMJ+i52iYeI5Pii
A/OAb36BzrjDacPfzDZiEYYGPhZxRDQfEncEGgHPFudFACdSTM6NEfMHTWA/mYiY8krHnpVxQd76
pSIBwcHeFwZXp974XQNH1EE4B6UA8EUCt1tqrLiaygPcd/aC/W8SgM860VBi+RNhP6SB1kVOQrhI
vSVsQSlpnO6ueR3nakiSGKU9YlGRv1yhYn+Pf4l56REtI71cMSzDX6JJdxbEZOCrd0KMo4kd+xle
jqePRFvDHhFLyZi6PXj7c4jCxsXqmT1Oc8I7QAHzRgIE2i6QFxQxqJjbjbPxEsKdaDmUgA5XRQym
Bb/M/XWUXPAKGCk8pkXSbnYCwRKuajHDl3wNmv4IirgVv1WbSvgNsR05o8S3WC/TJ1VXjN1Lp++E
GU5mGV2KJFn3HIE+qK47z05EWy9nVGkWW+1GC4/0mDxXsk0M5gMz+tf8W2nDbfi6D8FevKEd/pwG
SCSE86xUKMmz0TlIn3H+dke8rgQSOm5ZhzYYJiyoDzQh/0hrX7PYLNFv7PFZx9Gc830PaUagFG3V
sZxevOR+xoAu0Tu0YWOZhsCsUvr5W8DzwXWxYLw8yMyDSB3ixSgBJTgBBmy5Hl1V8Y6+EYI7+HnX
xRPfhGWPn/1KqZu9o9xpk5o5x6z3dYLNmejVWMkBnf3VfaZfS/OLa6536baoEOR22ox8oOxVoJKb
xswqOLQ8BzdL/Roqae5bxhSPcO8ebNdBJDWkIq3kGcNkOQT2hQMxFhu2xCjHIJYsnX8c4k1WWyL/
Nq+Mm18LSGfIhyY5/bNbtxk5nGnkGmvlOhSu0nWukkgZ9MKG2AOL0N9BQD6vA0KZ1hZHlHkbJUK2
8CqmdYGFDPd+vLmwWm+k5YlO8lS5XjDFyJKt4tF92suuNdZ1VLvB7qsfyjWhbk0zi9/4f6CSJf/6
tUx/08Lqgw8Hamr2NUbEhkhlkgup6hhjjmmkU2bVV+CcjdSrs2UTIRexJ2iw0lom9OaCqjLiRIgo
iJYaHn24RlNTnHZ8NKvpyQHkEkgmaRR5knx72hMCgtFG2+0aq6+5iMLaBpdMS4BHA6a3xbxBIpAf
OmftZ0sVIh5CaBCg8xFvcwrVHxi0ukemCjBaBj4pmmZCr3leBWpLvXTQUCsvl2mWLTZqXTj7BF+a
3q8FqW0yPBnRzjAn0lau2nc0jiEaucq9FhqNNYHlceMUzxjEzf/hXceDJwUUeeJLwTf55LA4OWvo
FEWmfSyuLSp0rR3mn4wX7hnWX+yWYqCgqmr0JNyb6pudAzsP0+kzEN8YDE9+IZrk6QgpWtPWraYV
42qiuBXrAlQ5WdCJu3iOugbrCdqA6NXWY1SgybL77q+vuZSHkg5ZBgwFij3fUcIkgPSVFcp7urGr
HjGGVZ1h0U3eFWQauzeWh5hApDo7e2Zy4D6Qc2ynXjLAJQWHLh7wLbBfkOfClGihdUuS2kVaNmly
ACB4S/lq9fY75xquL/8k9L8AhAzu5BY50UsikiNp5+qTjdII6WjlEZJYEnlG06Xif/MEezcCuZSR
bqWDHky61CsJEYWKhFjBASXE3pcUvusDoV9fYGIKaTVD74+yeiyu3khSb78E0Na0beDOvq20WdUo
i0bQtZ4ZdTewMWWW10xbyQZLoxdCRht4JgNamzcs1Q/5hCqQ+QJQlsNyxBQOODGA63tGp9IB9geU
tmgqyag1+iRE1jKq5aC8VdeTyeqQQA71ci/Mb5PTYi1OMHjQOhuuJZ3ocwG6YRaNbucnx0ewvK+f
UK/AnbygeeUM+HKDCBLLIPCvPQO+tYiY9YS6E4AZxsm3SEC+5Dqg1v5PdcioPX9Lk6n8NngaOLxV
wdyfx4GriF2iAETiYiUdr/4bykmXn7XfHgmC+CAlkjBDb9uKX97ZpfrQfn6RkUjes0behpPKofEH
leyYiSNhUJDcK+YH0BfPyWzWaIAOzBncuvb8VAR6GyCR1qWPxhG70GwPlaCqLLC6hOZX7DFo/+yQ
8KgdfAWCJB7mmz07w3V/YcM/DLodgTVJhlPcccd0mXQZfNP6Lf4rKexqg7RVYkY8icpy0NZASMFf
yoPHdWdwH/tZv0HX/jxJFcTIIflGdLTeDfa+hlId7y62MVeLM3BalHvyH4MI7zYo2kHKfi4OWUzu
wg8ImoHuzPoluXvBTnVefRwPreeMQlqDkcVsfjXn6EJ/jFeIt+RyE7IEwZRlGEo1bbWDt9TuwIHA
jmQzquimy3QigVdN6GDIZ5o5DkrhUv7Vc6u4YoFNOALM9oDGK/7fxybQFMyy1VB0hVjU9Q9i/sSG
MTALDcF1ZDRdqardl8HzK8EBI9aUfQTXdbmF+c6DJekEKRh+55oPUbqKR2bm02G+cyKGquNilyRw
igbD8VdLw5Fqlqou0nM17emiHFrKwtIV3NOtZiZi1SRcRXA2bPr6KHTeLB9s5cBPPi3pA+ayrsA6
2FNBa5XR62E733cHHkasq2VEEZ2YaaqSb84KMbYzKpqWdjI6V3EsS5VRndHtz4w/xYSpmW9l1RhO
ESMIT7l4X2DkQA4DyW6MFyFCF0xMv7Un0lgbhO4n6LiGAarzUiIKB5g/e9IsSCrN97Bydc8Tc+V8
V/OB9B8cZwFHPxp1CPDublUzn1oIc6FmgWpZhjD7X7Wyt9C1gpSPbkfvy/ZzjD//uItFH6bm5M6X
p1Aq1g0jl+jFpJlY9zxY/nPQQ4oUDs2vEmpJLRtZOMInsldtbE3g+uyiEZvL1ZcFFyyGDDu5cHcW
juPZ857dx4Pz7ikR8flUOyXZf3GGUOjlOCbumwbSKaAu2ZTDuWTUc1hWldwNkLfSu206sJBETIX5
zsp9hUcBUzeb1WIAagYlw/z23oC5I9qSKTT9C2A4vGwdoS8KmFxPcAXS2oOBM6nK62twmmgprMiM
skuKW0tkqiXlc7nuE7yCsXpDHVY55Hk80UAK14WG+uoBqGh7YE/vCsW8/7XPZC7NMrrBBeOSt9TS
ihD3g0jCLEiPBKP/NXp1YU+9zNe1aYHxg+hdv/VmVsFKB7dlRUQjXU4RKHe522omBm0VF2HwfTdW
t7jfYhiWiNKbRmi9kXz4pUQiKL4o8/1c5BZmYA1WkFP5/W7EgkP/7zuPz7uhcr+UOkMIW8iDLeZi
UV8+PUnHWprF93+LyiFtBvQAgzDydtooJ8PuJjqOP7m5lVjfZLuBe0AaRdHW2ZDehdnBwRjh+/L+
55LMpFu3i6o7WK5bGeRfWcxBYSOUVoHVNwFA7TS6FiThCMYrrPNcQU9WS+cj7ek/VA/6BgmiHr5s
xm9oHUIJquVBkMHhoAWunqfFl7Vq4Cob7SxE4YakqrKaKBx0/wl87mAQO0amioyvfm3ejWh51MQy
Mur5YtxP7vP5fm0+t3Fg2oX2B2XwZMXMIeS7tAjn9HxOQ1ClNB9i5vNC2y+VAquOR/M+4XExwxNP
G0F5HZjCIuWXZk5+nuMWxtbmwhzMCdwvLN7uIGlB5hgCyw5SI9Ha9+eBab4D7VTVwTJG684isO1m
dBGwmARwNnLmDczGPTAb/pCKPdAA9JU+6O7pLZ/id2jL8b3GpAde1E857NPEhnLBxl774S2G9oH2
FAtLTCYWjyFdNahGYyscLs8S2nxAdEZYiIxchTvLLmMuC0WOnzUcdtGo6x+6UNYiAZNEeGqxOs9M
PuSobYJpXOg5WTDqF7xUGR4bQnNzjO97SCQkoLBgVLZPxG7c63Fm97b7eXJUllKJXCu8zvA9zg69
mNqom/MarLK32IZtFXnUmTJvh+MdN1ein8LTpt5DuEDhUs2MiDd/Y+2O/XnQ4z05O8LreOWbRqtB
kIxg6TryJYA5py1Ef94G8u8EuWAFhx37iqYX5kNLnbp2SnFVG/ObU5CDO+FN2sI1QCXS5xvadVDo
ad1NLShFXnmGt0NKZEGFNBk6lfPs+RkdDQDUt8bd/KyCZsHLl0J7GXnr5u703auulWV+jUV3WiWw
2+4dkiratDhcGBXAbMZMuSXahpvlhKn0HLFhQXnGrgQhCHvHieQlBYHTA9uI0tAiaak7HWNTomkU
WhwerldWZqlGE7kYSiwAw6guu5AdN9DHMRBraaORvbWpxhjxkVrwYBPe4scTWcl8NoMCudspLvtb
mKu2MZPAqu6qyz9atQlTK2t2BvsLG8GRv/geTBO4e7tI4xIWnNlJ5sdp798SDAkAnOvCNrFwD32O
bsJ9lH3EZmE20dh/1MfbbTi4Z4jrxEEFFwP6Tyb78GDmalN+iLf/6cV8eK0nuD2WCvWNBvZAPCGI
uo93JkqSIRNlNQITuV7McW9+9eLeovX0YyPZ6JoJhlo7sLGUpWGMBYCbBbZMn5kR0hlHvGcPWO3i
fb8zg77xnAGI77ouGanNKZmC+z3DrlGoFTQxjbBdmDXbWQKBR/+NARC2EdKRQEyg0Dudryp1GWfW
jwavucq0CsdykhxkfD4YxZAhooi55krIe60vNzZd+P39MNOP83aT0iUpjxy4/pJtdQ6V2vHjwwyX
l5lt84Zjm5TnsbkumZHgLPIv/F82SQtQXNcvLMcRIaj7XKVGhvXnETU7b5Fm64hPbA71C+QKQ5o3
VedD7Yq+5xkXlm+HHAAg0G75/81L73fX/Bf1ROMvkf9bpcjeULEjXipIcV7teS2kySCOxCT7vugF
uL7O9yhSJQCT5nr3e7A9TvLb7GQ4FM0LuMXLb7suEPPRQfIWsj0/5/enRU+PbY/BN2GIcb78Ckm0
KlfCFTBFzA0JurE2qBbGGrFsIL5/rIqkM1kPpt1tmyNthsH5h1gAILdKJMykEyr4qYO/NGcZ9rBS
vm2WnNm34/ze5qi/YYYJRh9K58rsUp20IYCweYSJbGfVL/acHOfPcoHGlsr6KjaX2g0vSe851uyt
yBTPhxE7nyDy6Vel2xsYC33Od6Q/9V7G4Z1ACKVrsA/feDzy5zTrZtXftdfuFNtxCZwgfN8gWpcF
KSEu3dkqL+oIxRwqKB41ZOUDw3jstnENF1k3/PPSIjD+DPKW6+FqJ9sWaomzAPxiZvz4jt6OJHIw
16Ew6rixUhjhdOLFFXM8DKVa1JOmHtmsx0MX/w7yhXew4OSdkOvDT7M9O0VJgL8X/t/znF9FTwMz
7+2+WL6PR/u5lDsv92sr0cfl5i2q7Lw+NXPUr7YARsCZ3wy3baIvHO/WL/W82jhc7T3X/pLBnQp7
3bW08HPkqLBj5aIk5FGfKYKDYMRo9nXDvT4G8Ot3ZjlzKhHnx0nZJN57iZ24xKu681VvxNTVqGqS
7bVerD+2SfLoA+2H9EM3IwWNK3uDHvwlFQ1Vm6cbisv1jlVZ610uUhsvHFCZjbVW64N0xe/Qu87A
u6QFshFiW18iaKS5rNXJqQrRIoDjUhBhdOwFepfrk15769WZUzwGw047QVatAXQ+sg0FzDNLr9EH
z2chNE3Yu0diI9GC+I2s73axyIQv4F3Vio4Lx6CzNMP5MNAl2jUdkPNRYOpYQNsAL3BerOiv6Pdm
Kum35FRec2lO86xqkyo5dZsYpEBlD7NjcoISncDd/TkBhhXSw4nanTescNNTKBb9iyF5lrbVi1zU
GMKp3NjjwVtTtmCU6ir7Z1JhDcWzXjN4PX+blHl8LfpsVRmVdbsfKoof62+a9IbjKrPy8njpNZEu
SfQm+bQX+/ZHto+QSvz+Cw/jciphx6zIrFp0beZ+qGUdbXhOVTzK3bbNKy88Oon0PC4YUgHoF902
+8QgFQckahYRroY3nvH82dMyKkdkGrk/VIHhN+OL5MIJEJ3vDO4RcCwz41Elnb2aSlRyFrFAuDY9
EeknBF0INF0TZGmGX2SWeX94RScEA8XykXYSU9gtrirsRM8nkcxA8im5Dk7EiKw9KEkknwl2bxlo
8WluyJQqRhZ9LU1BjwZnUejFZC8lKlbh5yBLJabdeTqeEHUYzgXVusdTb1IOQ560e3eon0BPUAXT
bXf1slwT8uYsbZGo6pK8UbtvwxMipGLwN8eNLiJ619knEyAcypHz3ng0txPgUpqerIe0BPKe25Nl
m4xFmYdoOxjXqkvHET8+EncmWnwSSAoFAJtmKSc7fRw/ptwoJ8RDybdmIieXGE7NLX1eUFPI2lE3
L9La/RNVRhUtdw1B5XUkgdyFZTX8WtwfC6tFFn6dWuyC7iSsUpqaOdmWGRTPEYwTFZAZOeVM/631
aDgHYm0ZLf7zfpXDalaLmOBJ3VCfnFY5bvBh3Dw/zappbUXvEey+DWPMj0caHCkRgpGjXft8rDz4
wNklmBg86TOG2LsUH0tWpbCF3rhv0ducs+OMfsm8alALEzUeSqmejExrXVgAKjPQQaHfFbKob82R
AgGy0ZxgKbBxvefIMQxqFkaVUdxg5ve1W0OjiWdGD1vi5d6P1HzYbV0ke3VBXZ2oezUadUG9QRw4
fF+mgYigQH7WD5I0KrJ/jtwNJi8IBBU7WNB7qXosHekPe9QLlmA90th3wCnA7QMRmlq8O1UjUe1O
gtjF60uOam1QW0tZ9hoX7nuBq925b8Lz+qJH0y4duYMPEMhnxJPMoBfwd0QwVDRw2Ci7O07MQb1Y
+tbQpEpV1/tW1XxoIJu3Kvob0lieRM5q+6YrJzcI3Hi3/c/TMoEphXGAMjIK9RsLmqTilp+uczS1
dPcRGLgQBCpU3GQvPQpbzJjYZC3TCdvp9b+zLHusyRcZc4xp4rKGhqC+xpfpe2MULB1jVnglq3Pq
kSplPX9F/l3zQlkpS2MWpdlD0fkyfzY5EJD7q+BoW8Bg3lCWvxlrcHoW9/K9cJVIF4mlUoWNV2v7
BEpNA3YV8+3tL/XfPooX4NIvrXM0uDPlip/dpDEqxHkznEFbRb3JzQ8C1PczT6Vy4R5Pqb2lAjVl
9irfLOkCEOvJVHSa0k9JmoFUhs60JkXEz74HozR9CRzIzej24t87EYJ0YTmeb1UMEmGRosM0yPVE
sX5XTc7iH9/5kPpbjZIuJcJTX0BeIGrqzySQHs1meDfJDGahMQ+zrRL0+vt3RNLlFxWHxNtU1STe
k9YH3mczLXFd39j20J/Ta74VBidmIyJ7fd9475Lm844d7ktUYIQiAPxBEOR4IV3xw85Mc8R32eSD
6vgM39NaYREsTf0pFniaV7XKex5WIJYQ6pLhmAPRfEosStJTpnttm6DIxbXVLzI02dREI/ExgBBS
dGzp8dJQFtCM/K29U7ZEe/y6o6O3ciGlIcJGi1hXWhpC3Lyi3pEu1c8M2QWgBsTu4O1phxJtdPgH
ZTqMIrgKESNkmgDccg5VmHueqYnAqeVPKH9if67ODYaKtVJbMMJO4zN7Cn/4SzUD/VPadOD4wmdj
73P+9Eq6aOV7iPGlt0sg5Dr3FhYSvmnbz8vzsQqoVmv4tOsOLzzAiAVESLrO5AjXxo/uDHsylRtB
Ftwlwb2/I6hha/3SoVUv9N8iQrsPCxfUDF/YcaYyHe76pbpv9YsSLYsIsjNLoCzDl6nFBPxAu9dY
2gt7IokOaCosq9F1Npr1xjSoKa8st5U3CI6rLHcTO9MRbW5KThzFnsZ9zkzsq6msdO6xUx54s13W
O4Hvzl4UdILziLGRDFXo99IVRGmNr3FroRbe7iYVCV5HJQIR/U7ia009/4qO6Muhxb5OWQBjOsVh
wudiG5dbGUkJgrDgBCt+oFdaGTIdrTv82KuiedqOZ1ACX0uoXLbPgMV+nhh7RnLuxfTbRWtc5l6X
lfqJJAIQGYrUiBT6ICw+YTS236ByIkfmN9tyiigMDlGJwaDAZBf5nQ2brE5bhc5D6mV6KRB/L1rv
oVNvEtivV8ivK+ori7qrKQYvI51yJkPr0gvDwyQB9roeXp/kNhm70eQfNFwAyKd4sNGBK/j558Qn
/yEI+l/DWpsJypKEWEETUeQnRayyYv2QbIfiJ03jnKsu5VqynPjsSYU2P6zAJk1h4RjME+w2V7l0
f1D68+Ov8IBKVywRZ72D86Hi6yt3AWLxTs0LIZys0YGXjbK0eRGeZwht3bBh9VMvzrNUK4wkbrXZ
0hlnECwUvJ/JB0tyrveRz9ab4Y0G+LY3tpr7fC3aLVEeFL/E9kIZK/YLlzlRPYxJ2oEHroc/qHQb
UMyEcbp7QmYSQs+cMefOD11TrX7U9+MF4Iydmf04onvj8/6oLyCThlubB2KcYKt/T8noEzTdxeSK
jVeqwkEfzMrSrnDm0prYVTPCWJIGxHdDHu0GyU5OAMFU1taNqRp/s4AFUrXff/JdM1NDUHgmNEbZ
G5mZswXXDCGdM08zpof2738MGPGHb4oZUswO4MI+XHFPxxfEQljLQPY7QKTRxl+dVo397q6PVN3j
jcLyg0q7hsE9ePZm6N0YTY+4vYyMRJCpjJUc4Jf6bvuD16dHIk0B3K1ELZVJlIfQyTUODpjPKNon
KCOeAEJyVOJXaLZaowpgepw83YwAqOwCVUPkvEKYpBtmEXOw0Km6L7kIOj1DoliYz9mYxteAgxAW
0xar/+ZBk/P5yvQLBqtGqKgtpezWo0QJS7JY+mwTJP3NzXeue/jKuXyrcrk/ANVytnTFVDpKND91
46xkH/TP+gm2SYOQDm8Lq9iqgIm5/Aj/aj5+TjcatHU9nFKdVOxbSAm7SikJGlnO4gtJkrQ6nvTk
ZlJzTlYVdoKknJamwCREhaySMCGfNLOlgkqfmTl8qVHPwF51kpEo34HNZDkx8UR7qDAcRs/l+nW5
cMWYc5we1z/sqK44ubE7E9P3tR0QgPzhq9/9w/Dc5ta5LG517G26r/GifPLnHJsuJYcUI/LxEv59
DuesT68V1zYsNV79eZI2DQWVKSLVGwaQ0e+CH1pA+q3EEJiGWu1OkkQOpR1ElG2GJqtNa2qTuanO
HqFSLaOffgzy46pVgpkCaseqa8/ksqW3MS0QKLU4M0bTQs5y1tQplwWXuKYKSqNzhcT4Sr4S+1HS
7XrT+3drYCv0NeR0YGvNxS83V423T7Is/aVr6OkzB27tEpLZVYClXk+vN5UnpDpSZ1ytp/6boetF
y9+DEuAgfj+evl5blf6X1RXRCjdALwVHtlTPbCr6b8sJ8afbamxtmYij9AD/FwOm3UQ3LIutqIkw
NL4Vfib/5405QOKvMabiFBRbQgMvUaQVyu10JzMdigeJK8CUy6dZBNsKfA7VAsg6U+6ocJj83NF8
h3700fyZILh1ttd3DpRjabnkUmYtir2dr1Ug+0Y13Tb6xLHVf0aumTy2lpGM1XBhrckZvQ9MSNhm
yv9SkcWe6G6xP98LlsYTiALLQyEWygXOiAmQRzOEfgbKAjyhpeHcomr807Mbipd6VNqZktq/HvPu
q237yT7X8+JRRZ3V5z59ApjChhlVhn6FnylU/ID5fSObWw68v+++tyPsRPAdDhdBCBIvrK9x+BBg
TSlovs3Ir2x8RCsZ3gmMhhs+xS6hrHRjlRMgz6wZYvAvQVGrIKg4ADtbff9s+Gfu70sGCVjtEr14
QNgTrTblCfHm7OeGLvS/L+0DTxqcSzgUZYS/7QmOwpXOCAKeEdXlbjbiNx+tH/RBRDpaDcGwVdjR
/SzPio2v2GPIGyRswqgL/eRq6QbqLng3SNTQccwoKi9T4PhfooqG15JHTR4hdDmjm+gYRzylxCr6
XLJ925IeXiFBzphD9TE0PZGFLCFCnIlAHoGaqABW7+pgoaY27Q9QenXtitHA5zV70aA4kp0+72WQ
pm7w8W3p2uRl7zEQrxX9LMvnM4P9eSjN9TJygopQEmzWV1R5NeS3sF3tp0Chl2R1ccaio7XzZSHE
AA5KwqN0Ot306h5biiEJRhmy/Bq8Y9gRVTpK2nVsqmwuHa0D0g152meshTqtWhpCb+e5JKIYoWkA
sgPggSQ3hvjy3MRjJRqNpj8Csw+AEDrHeQMd+RqlBDHV0p1LvxAnNzm7dfUX1OFgnG8Li6BFrYu1
9raknyWMcj2pUgkqf9RtWhHwFmvB2HTp0tmtG+CaVjZo+UvcEdEhkE5PFRTk5m689qEaVXvkhqsH
XVsj84669OiNkCgX+MvpZH0HcSQlKYSYg943rOMLbYyArji9+WrCBdfj6CJNQKC4AvQqHSwI23br
Ss8ktH0A6qY8cLZ28rpiUrhL3FSCo1EzPTmA/0MM+P54F2x9DLrWP9qiYD7Pq/MDzqkk8if0biGt
2V71SpSj4Drdnpl/GcptVuU8gsVlGXNPAjX4zbywC6HSPwFZeoZD3r+rJiLDTN74qUrYArQGv8WP
6/rLSjvfDP8u1WKIezy4xJSjtuGw7PpC7N0+Rm2FhBEHp5K/fePt3eVufWfnNFOfDlIE7igBtkhs
lBgry5BglPSPhlfvkpofpTwpLASw8vF1Ngb8w7FqdIYzfHXiqF3OzWELeJBslL5fzkcR1rUBzl8G
gQ5i4bQ82dOfKMvIzvek8ucsD6qyiaNhGPkCW4nI6mYp0bJvTsjs7aTb4yYqZyURSu2YNp3ZXhor
iggpnVSh/yzBFlxhGjqa0f/R4eheLONm0IMFpVOGmKP1kXJoQ4rFnnwJ/ztWkk1funtkRavVA7ci
z25e09n2koTJy48egR0qupv8lqai0jfV0lXy8XbF2942m4KXNy7k41RIWQxSenaBWqZ66KL56dRE
dUEB4dHHOq8sAFmvWSNyNOWDLAITTUL8z4HkuRgjCp5n2JkhuB48QQ+w+ZVjV6dSVe/xty4SqOBt
B4HoVgUduELYrjujZtE5jRLqf5uNVU0IuPQm9/f9r3sDv7/f8nsplzTxUzsDRJ+m9G1RGwa4W+nh
AN4dwyLVvK9ehBJvFxoNxwBksZ/K0XaS+dxg9AIpcNzdWhDxzldD5bjBL9MX5NsEwbF4D3i1u23c
Dn0uqlgkPlRpze4OhMWCgqUdziNK+YFFG/bWM89uD+ytq+DD8AG1NKWtF60Ara79F14ihN2ZooJu
8V74cJJfqZXJ0D0PSlE4i8kkU9qHK3U40RrL6qBhvdFr0cmlMEcbQK22Ll6FHxHJ2YjPZpqUkH4I
/IOudN7ouPlcJq4XwoROUmp7Hl3vxNTiCR5lBoTL5lOhXKIOl8H1Y7McmgrFxuyVALVqtELgpvso
j+4V8oSROyk0rbNvmFZ9NXJV72+9PLz2N/itILa7u1u50+8pKtMZbXyx+MxoY9hEn6D6LN3bqvvH
yEHu6TxHMGjrvCsemreY4XrA0zN5vjD5J922YKoHUB0HbEFjt/HPVBKLyohVu3yQSdqY1EyZLlrc
1Ri9x/QWqRwgSAXlx7TllnBTj3tvN6hOrqaYRI2lSatIkxWB5ms8PQw1N7rnfUj5UI24ygnYXX7Y
G5KhbrULqFhBfXdIDjCi7B6lQ0Avs01sbAjrLb+K91DqUOfo2Q624Rq1nxHqKaFFlZVSu+YYU28+
01IfYDT/g+dBGozsUIZ/cr4rB6fuP7igw5ifBe2KPS8SdOUTGnxz1zOfRlgB66Ot1DJj7R06ocLw
zYxZoP5+Se8csSu3tjUOLoo/VsyuEDifj7dHXncas38gOR6wA4BanbAOgr0a/IEeJi4MV07gsalz
drIEeLOhXM0IAjHpEHLca531kr/3EfTf+6e92IeHVML+6U/ihjIqlKjvOuKxcU0uAVKpmHyYUh37
xgq2BzY433GmOwqa56+2PVKEIwWoDaqnzQAfgABhjrXVZvwLWSIl0KOtgK0c7eE6c1j8oiFUF8W7
BFa3BHbR/0P4F9cYyYc9Pjl0xckLwMHOQ6c7nAD833jgRiOneYpJOZhBDrLe1hFy0SQN0YdROP9N
5C5eVuYbO/8aJQxpy7zJpnr1UEQC1BTaXXziQ6vEsFQQuuITbJh7Ch3CtQQJQWxdDnO1338/e/QG
7IDzIfyIANaMy742xUaAnA5MWk/0o5SHykhel9LP33G0atkT0sAk1hXOZk131Q+U6fDtKAjtuiG8
w0GvQbwnwstiMTBqU3ommp8PJNLwmqZhNnwP60a8yzCP53YwVZgdAdVV5XZi8Z8cxj7dvJMuvMWe
UGH5Pkj1Pevg1abFjQ04im2RkcidQcfujvSs3x0cnhFU5hPzOWW8yHoYd7A40+WxyfUSetEiOHR4
r8GhUuP2Ts0RLyQTg19WGEPu9EvBkk4aL6Nohw6Te5dpuzngXkN7sV/NYdWsZr2DzGjDhtUSPw34
+qyurwdVZdvQ0qMyvf7NLl1nYRoAhAA1OnO2m/GR6lzNwEsg7CjdxbUEWJT2iyDOT7chcDxNLTj0
BMkOFOXPqv+3Iv0pFdrHsH3fLGeINZ1D6DMF+W6rEXRAqFFdOq4BFE2FGX6A51wWAAMtJDG0V2Rd
xdjUg/xuFdWEGmJTMLDMdNq2EbZ9Y+wVh9WbKDuaPBwSU5iF3RbHFPcT1EZbACTNWuP+ADgzg50y
U/TPHQGM1hqAcBLTfzYv73YOObw/Nv5EliZpRt+JRR5Em/5YbUn7fxK6dhGC+U+TdHiWukzHAuxP
bXTAaioG0vqe6UETg+9x+B7/EMH7JfUCvfEc9twD45XqSXmb0g5i8/ovmfwgmY0USE2SzPO9m8zk
DVZxC/qEhY+h8T9NoRhCdsFp5B+9tw9ovraVjXMAUkQSbgm8yqV6E1GSrsmWpU/3lna+KBbyhytP
601PWhHqXwqVL7I1Lq4Ihyt6Wlpoz1BYaPFaV1jF6e4sLjUkqCeWdHQcO1kvOZSlyqrUwtldFWXX
NRff0m4JuD5MNZL2nI0bOh18eFmLPThoLyhQur4mOSuk3VCGXYF7rP1kUVe+8lfmom2sD1D72FG0
nOLkTLpca5mPzyiXcCNo4euw6IWxxN+eacOTacQ/e98K0Iiwozpf0dYtmGIQtnK09mKFGamYQGjc
3ML3n7RfgXrgF5y2bsIwbVCfcgC0BfFTz+CXFym9ML8oSiNVYClKw4xBizF39ixvuBTB9HC3qlCc
Qzs5LcL0KSZUnXQQY9Sj+g3fWhbGfk1VAevFX7lgIbmBFVldx+VlNGqrpnPKkH5c/OOVLYtB2Niq
jUSOgd9Q1Put2FXbio55vHOGWthuYE+6Tu74q0bxDtDKj6ZPEAUmxC5kGCrvmrr+jy8dYZsODua0
K1ENahHmKY56YtxbzyMr/FTEMv8u/v/obiXlIM+LlM3xFB0snWgfA2j/DoCCt4xwwrV4uGql6vI/
/4vxQctHShIAQ//YuhR61O9mvGKB7uLJ6API0l97tO/r80CO6mNHZxZNK1AC2qWBMeqYzOZryZFU
2nXgFjrKK+sQlcwXdsqI+AeZQEmJPo6GoFX+vcvb1G7ws42IbomT3Dh0YskZ42n36u/S9qesiNS0
tFMvjjtc5wMbdVwgmYk1lCMLp7E/3diq+BqvklAWk4SsrmIGvKrzft76YfzjvAzN0hla3qX/SliF
mH2K3WMwqdaMg1s76cQISk/HHuGuFa/oxr53SMDYMsbSzXw5Ecdo4kjhSPAj8Xe+ZkwJy/fhHfRs
0twH4DOh64vkP6b7+SPY7AIfGz0ROmZczgavaVpLjyEgVNLpcS2aJi25LmRKbnJM5Rf8QrDQEEpu
tIH7jk874blDh/9rDSQCkCuCycZBjPzoZhIVZmZwDANTkBVWmfdQ5uM05eMxZKDfE4skOYHOdBye
s3lvh4+uVIgY5OffRYPkA5tyKbB8FBracRiN6zT3TIVRZRtrR1TAiDXrk3ZGEWcnf08mZY5fvyMU
X8K2b7pV4yPv5TLzS91yIl4fSaHdkT5BNqdTNtzaGfpzUIfk9YYGgED/tCpQzEvU8K8OHWOg9M8x
wXiHtSLE/WTDgIxqEWZ7tzEReOSRDhYR9mQcvErZ+AznvAtFPQm1W3WD81yMmmhCf9E4jMZ9ltNn
19t9NTPZ1/LxCB32ltquKOCE7v5Co4W7dZ/EwQaqDF6liBx0pQpuGdzagCv4QPIm0afwLWzIGses
wRjo1L29wRCFiQs68flkOv9CVEsJsoWq5utZ5gzWZteSnP277XtjMjzolpjL4AQUKxQ93BO0RSPM
iuIV0BRNMnyNqd2Tulr0xLqDxvurvsf3vOd2Odfk82mbCi5fOdGZK+T4zRb3vLmlw0T51GAWGlzb
pph8lHRDj7Po6hJ3DfMtyTR3oITDf3OvZOVPl28BoqU4sZ+VryUXgx7bYw5UgvzUT2OsCa1wmLmz
JE2cEpzSR987+5xpbrqilUkZTS5ELUTZfgiAn2PmzBGMjg1BtuBc464xttb4yQvxyZUFzy2/WDDJ
I6CdMhmZb5gTXfdUDCKja43DjPVtj4nP7NL1u7WDSXDmNVyRg3vN7LOx9e8hDpKDQfvcCmA2ALo/
ZHBMihYJKo32KtILaDEbOyWcv+dwt5QuMsC/5pAq7qvpoHhYUFKtivhF1tNkUJw7tZtk9hyICETe
I9+eu5S+GLxd+0Z2zKTjUqsrD2oKQxV6HwOI1bjXDnqiY4rfzFFQLsPChSg/i+g6UOeqdOo8XLEz
ENwlpWv8fzgbJrnaBl19d9RZHKIEmlYnGbYswy+j8V7a8VT4TgbXbyaT6tFwrAH2Pmwvflcgys+O
WbStzBAaVh2sMhHyPnAKS1cye8boL5Hw2n1MyypLwyv9v8Nqzs4bsjOErf/aNKT2Y/h3jyA0Wpkx
KvAcdPCpvvOIUQJQnbOToJw6fl0Hn2p+yVZRBRy3UTaYQy3YGOy/EEa5mUZGJkMvObCWwrX4NAnO
Xq0sBcQnreuEeS4ysmqF6xuJEL2JzXatdglDn8ljb+K/a9ISC7iKKwOiTmxA3gtzjC25veSprL2d
TXMzocYkSqvHrUr3J7smVjHOKtkj0TwDMxYqnhtHpALo+lCymr13DdQ6+reKg4pmqDxJIiVR4Jw2
nksmP3qCz7W+gr1hjFzuCDCTmTe0sWxEUL3zWfAnHWbUrg9Ge2oxeqauutOZWI1Q9mgwIvzFv/k0
LVW/YPH+csBmPzuA7/qGxkgROtyBVQ5qpqNPKXERKv1ftTHlOaNbtI25RaU46YnY0d9oX6E2TfEe
iBOK2x23UBRD5HR/mhzy+wGEUfG3AO0Jvc7ufFQtyk/UdhIFzzHx4WB/S7qZJPmcDKVgm5TqBPWc
qbNFSaJqUvjPG+hjReDxEMaSWEvOrs3bwmhnCl8AtkYW2i6apkPLCIkpBYC9QSxNCGNE5WHrsOLU
Zei+S1uCPWBxj2maScMXrGS3w+rxCXuNAzo+AlJWDWldcFJ+2IdIGTPxtgLzvoBqZAAKzKnOYjDP
0+j463fNoR56hjWnLSM/TukIKkaDmYwpnQutXeC1u5es0N9NDlePFGY73AMV+w5A3s8dC1uLehuA
0WGkm6crjGb6tPr2hWCi9JJi6AawwLGronwk4gnZNJ/PtwJ+U/ObBP6yoD6cx8ompsTRL76TQh9A
YG4mwa7dnF++jWY4o/N3HHIgAUBK5fcsEpIGMVDLK+wBhQ5AnBzE70ic/zimfQoWhre/L9BqHwiA
ZCeOUOd6aD/EF5Wm2XtyQbBVVzsyKn7TycZRVxlKHrxIT+bXxMhXKCQcmBeJkQHkmlWwbm/FpwdC
zBbzLvNRdWpEJAtnvTk3REWrkri99wbJC+8AkywqUAJHLD9fhd4Wv2WW7EeM4OnD4DaXGXoy3yev
XdoaNXpOSN8hZ4UB6DLXjJ+IRaB6UV+DXXV9AAyCJAe0eh/iqHjEm58GUVg4dX5ZyAiAgoyEaRiN
wP0rsLFeuwmkdEFvXQi1Z6Djyl7TmE4PyVWrS5JqIJIMUzqgNPW5jDd8A1ByEGGhBMwfyGJqWQn4
aNgJe6fPpOXav8uvPST7NCzu4HfRgXmGu495CJPKR/+9WhIth6/Wvz37sZ8ai8tkyKnjZnQOQdAY
bTSk/qCDnSo7BhtL01ZY4j/SMT5uqVUnU+pUsUlkoTM/EdTSO1+BmnJ2dxMBaq8JzJ8TYw1pWgPC
iuaU6RenOVXXLloQI0Y69daI8NHRLWb+BDTlxkWrZNhfpjV0UKFsu3+FqcVXY15OfP03ST1qPRm/
juqbGVZ0VEJUfhKW8/G25qeKikCT8ahRPKQ6RR7ZCDVGbFKwzuj/r0leJqsoW4waue9i154PioIU
QpKQvPCAkK2lsr7XChVRCGKzqoFVvJgPfnjfyh3JIAERumI5M2TAo90YStWHGCbaT9BKxhLZlbc0
uQDGJxqah9rtqytMmL0DO7JLg+Vp1/841+w/6aoGO0Lb4U8/vBosEtLF5IlSzdmbMjbBieVCFvqt
o/H1L6YAY+6V/HJnWByCiUfxWKPtO/htnOCUVjHjLdgrMxZ9PTZ8pqdEO3b5fZHEb1VxB10xTL27
aLOCevRDZSXjwXy6hzzrdr0XFiBF/yaxfO4jiwT8FtOoxPNjIitlpUFGINDVE7zUsNTKE+vox41r
Hu2iDbSe5AXpOC6dg6d4XsKS3RUXdnv3PInCjT+Baq+c8Cw3sUMyhJhKGzqPL74BJ8LP8VWk8R9i
RXOfRQ3U2uY+To7hmD2ffGp4gzGUleKtrX4Kju4zwhGmtyXqDwrU7NcAzIomX4mZaJVaK9lBqhgr
FnKGhQVnWKYyrSzA2UZgLx2+t7XFIYagmu2dz4GmccSKF9Sizg3hQ3UxOJ+HbcIKimRhvqAJhtrR
v2rhg2W3KDDplo8yn2g2Nn+fhJqJE/k778a1yaHMQs5qKER3zlbjXUPzdEJjvGTlyxSCHQSa+G9o
MyGMZuC/xjGqWmioybxf4n7VzrU0meo61qUKNFHyHp683Mf+PlZ3e30/7OxInA35lSyeoifDOdjM
3viYOVmv5A/p0pDi999TBpE9Sarih3h+Tt4PRhM5YvS4lSj6f/EVsnvjBSuirnp1uk0AWo8H3cCZ
ehFGG5oA0uGAcnXzzYsQ2QGw1UfX4MC2aSZPSaq3Aja9bGBcCGtncXFvbgBZ2oCa6UHsGJlgVaO0
PdX4oDC8u0ln9hCRr4dMFNUqYspbjYQEILYvWL9Bfol6uXvXA9m3pr5DCtYIBwVDmjoplFXVYvN6
0i7yPiUuvW9L8/zbCg+RY6PElv9gVgrKPZ/+QZg8BkcmGnBs1JadpizYTPqUU767NBQ84UweMQ4y
vwq3+oITLlNbnZ+b3Lbil6Mq8SdBo/0czYgMDIO22fujJyyKJB/kMT2eRmnMOphhS4B5PKxWM8du
11Gii9+1hGhVmTrgztRXxYl3l/CVTCLrqND9NVeWsRJ8ubguQRKdY7T881qQpIcTXx1kghnGyaW/
NjSoAL7MGT5YB+hrLt1dBe2LXSFh527yjSEgenaNFDAT5r8isyJAZWKlhHKqUUyHcAxq5GBBeuHi
AVBWIsSFKoRuqXAcdg4KJ///hNF/RXu3AtgK2jP632tWiCygMET7NPxeR/xnN1haqjis78j5tP5C
VESNx2SdScQtsy9i0rozDiRvRlWjbEplF6iDGkiqf5IbIsfcHYuVukrHAIPKYoDNnW2rjx1vHcv0
YhhAfkw/+YDpocZKlT2/m1/gAV1MohTfUAl7k5GGD+qLe23EFpBArGTJbZVn/oHVaqRfuq1syvcx
MqqbeuIe0VQjQg5ppd14sPip/m0fD3ufe4L8Yjcxy/WN/eqBYxFcdI7ue2idFMNrdxyX7cZLzrZj
YB1fSuM6eTQ7f5K7N9rmmPrkQMweo/huu30XTdqNLQmuTrQ1nTw38BcL3uOtjg2YpoH8yKvEK6Uc
2XoZAYAtd/cqarQTB36Ku8xeymHYPJg7wFC1e+XeSJScURO5f52OEDaJJ4AzCj9/AXH3eXb85iaO
HuwETXcxc1s/RiiaafuHjms5K/j2Cw5Fw8WuTDScHXgZw/LsKpAhvKX7B+pgVyWC8nuMCN3IAIMs
lT4zsnbhgtLexaU8uQ+Y4sw0vHWci6QgY1WaImQQnyMsDi3eHD/HZGCvtwQGBLoB+GhF8zER3rAr
fCESQLMck4bKKeU9D5SBacvPT8RIzV4/uZfxeX5K77Prr/jJ+fkdH3pqbuX09QEKSpZWitGByCaB
G+1tsGnIKltCH1wmi4RJEzEH38vGPaI7dLM+wGuXqnDqUVBOrp6zENJH11l8WHxC91rLgPeK0KjG
oolXMo4Bj3mk/zeuJxHC79GHafNNEl8cWsXfxgTu2GZheQH+jE648iSSSofo13LwDbY4tI+X1ZIo
m5ZFtzmyObNd0nPc1rhCSkGdofLg01eqO5yGMBCceall9TkHuZCofMCJ6lOo7tS4ck2zEReFMp2S
BzefCJnh+gssJP3whbN2vBrnkrk4932fmkWrlEb3S9ouNeFT3WDwwmP1ok2CBD532pb1NjSpmQCo
660DfroVT921gt9gHsRxMIazBIIv/mSjtCPDKW8L4ai5J7SS4LDnDfjxU7Ys2uS09qm4ECH+o62c
h8gGQkUnxZXmpMT1/51rKddGTBkFfboFhRXljRyWnyQSjNZ8ARn3GcP6rLVGkFf0dY22Un09n1a5
BmB4CGHSI5ldF8+xJeogc+pmVpxA0CqX4oMZhstdlyPfwwUFTzx91EReyDa1txsdKdsHs+sV6Bsv
2QUZcawvMUiEvmb5x1KY6O2TRJCJfTWgOTl3wvrXqrK2OiCvYLsD8VkOYk5P7Q/jtCW2w9dYxmEg
NquiIYcva8RWB4pS1Qz3P1JkYQEVqi7ZuhoNLiEAed8xn39UxlOgySxKKYNVztPOalbK8OAjVqxn
8Y8APC/FNKc1vxWFdlenhWy2d8qfAUQaGoL8RPw9Jt33ZGps2TZiGjI6jMm4MJDdNGAkGSkPL22t
kVALFGkrGcrYMXAU0CvoP4uG7Y4K1EWItnXq4XMNMGOLKH30IvjoOiB6ccrXaVuQfEUcD7aGHXDF
OlCiCU7CpiVnnguVafviv1iKzg4imiNT8WZrzE4ck0YX3ULX8ZjBPxzT7wsz3sNHmvMwdCCfiD/B
TindqHlBoHc4U8RT3G8PZSQXz1WR4r9GJa9rWddVA+yp72ajiTnP6EuWQx7gTSg8aiqKcd023h42
wUgQe77edAl6+KqomXlY20vijhih3/JIsi3vwCUJRXURM61B8LurqNOMfx1g9VkNX3dj3TsXaOtY
EEBKYZQsD3Ko7VIJqUhLnmT3+55LlO5rm2ihoCs1kUjV69hziMLy3Mk4eskyZXXm9T5wuhrK/WmP
f9GDpIili5YppK6gOJqlTyAJtw+cm5zmsSUWn5ZFnVlds+yj96qvJDPunkL6V48E2GETstY1SlTt
hh3OM9UHSr/v+I8Lj/J+Qr0DsqoOMn90jM+Z68TBCMsRl8F/qDnIeRsG30dIz3WNoS5zNm0ynvyd
o3jsz/Osdk6wAKxXkbtsV6KRFwkHtqR0U0TkjpyPMeY/pVx6qGg0rge74d9/UrpR52V9dyQSMhtO
oS/jYc0AUonvhYQJMjnzuB7Z61MWbx6b6537+BSKj+exh3yn9pdb3vH6j6RuXxZAfn4eIomUr/1u
T4ykSOzf3/7A/Fhlm0UTd/wHAgw2+Iyh+Jl3TMx3gIhG0YED8rLuQoRS5QG17Ywiyu1DGfhXKpiT
Ms/KbvC/JkyntGkaDYnF4hSsSGIGFXK003D+qTAOA7iccG8IWQMBv16rFC8/GPXKIspZUtrmhvgM
OkE9Gv5N2ZCvR4N4R5YEW0Dlk9rVedvPSxyyE9pOWtPmSDGQca8tsiPSQYCTYzv1QYpDbBdrx0p0
OqLpZtLBhERGj8Nr8dTOVjQfnb5Kt+N89IiezMG1au0zbCzuSf82MuBbed0R/V5lSCyZMiZaTq5T
sofqZX59krD1RHmCjDUW623OOh7ddfZVhp8/t2jC9R35WPzixItgab6yxMygU/1SJW9hOeTjoToy
yV8IK/3PRTqh4Bn2BqcLIMTZC9iI8c2CQ3fqWn6W6sCbijedzVRtRqLdVyv3XOP5DZn7KA8ebhNS
KU3rzjojzz7/zk4PB56+GcTKsrZBzMwTDeT8PB1tBrtvHjMrSokvC7fHJiSXSOwcDo+6mOxMfxTT
PIYRJd6tPeE6etBnRkyDOJE0J7uKM2rOdnSE/I5ItFGFKrYeZRfUPomlhAIN+T5I8P5pBnCw3eEc
FVxj1kt7+V0tCqmxurnSE1PBvkd9GbE5TfyBPHqski8N1EkzLihSDFvdYo0D2KqE6s12bB7BG5GA
ZQd/eCdPoxf/oMzibM7bMX57KHMHfJZobLIYCjMrztQbfPqhhzgvocumBEf4rSm03u5SNKzrg5Nn
TGrDnJ4vr2YzfBdyb9Aby8WrhysjAHU0ljNLg5jo+rZsHH7qH6d1Zzf/ivaAaKAJJvnuAApygEPp
0N3QlC4oddZqpay/FBLLTBEPLP2HpGEHgqZhOH5KgBTGDsSyQDiSlUmxKFD/yRHxZsNEOukEtFL5
10LFXr3EqTb1PlNqULgrQncKbRZxUBxSHmc1a6+nTNfmMGE8aa98XyAWyap+p9xE9SJTHLXsVqzP
7DGZl7V66qWi7jxnikqu7onpgqYcxpW2Ep2CHKWXo0TCTXWexqp4h+Iugq98qHAU1aBr/DIEP5iK
itdB9e/5X4shQHYmKFTXVYMELg3Iu9lETI6ykg1qD6HaNZPeH62qjC7/Mm9UfI8tm0u4w2BF++P9
Ph0O+8Dti0f4VQxOsfp7mluInHQYylYjj7hAJOEbYo+fVkttC8PZRuL1881KUJrFwVw4NvXmhUD5
fmWOBCMzQSwAd/bNBM0aY9eOyQ+bPi2lOn/pQX08WCkR32hc7uYnRqeXfR93PxSSYzJ34Vu1ioUc
dcTGpcFA+9sNjr1V7T2/p4pU2eiVo+Ih6zs1Oq3keUIiGAfTch2clrNhQ4dXrCwC6iC2DI6mJizW
BdnupXnRrH4IRES500vqigijpKqn1I0R2PPjfaCh796MF4qC9cBJh0Wv7N47OoaYPk1hEXMii0G9
lgH5AHvzrqf6zTW0ppREZ03+Jzy1vx09n+qNiJevcLSMfLqw1yeB+AfoH3QEJA57R8BG5c1HoDYy
uXjdDUjr5rKj1HwZsjo2pO77gy11VSBmrevu4pETa3fnvbwSMP8S3ZigeaiZNSW3VN8gkrZAycRf
T8M6iauFUco7NVgLCwC2YZtlfX7F+/dE+bdFYi5ABkFM+B8SRqg/PtutTjocPsbcP+onqhwT7WA/
2iv6YWrI7ZilxeuwPi3kycqhQt349T/vEgedjrhJ46Q3g6FDaPPUuxQiAh2/JT3mbP9EeCztP1A5
/qgLBitnVijcxxKswmML6L6t0cIdVHI+O7cxr35s7x78KKBt0q8AIOwDacRSTvGG3N820VVvG34e
tE5W+EkKH8SrAXtm78hLE/cEfuLssPhcx6dd0DKxLgvuHq+XH7mEhiCVXnr3bH62Q0lzU886niZ4
dSNtD/ySJJMFpjSk77dBgrAKObPZPfwwlcavtvdJCxZB5EGB4DRauO6BS0iJZGtxNXHbkZrR5+Nv
Qzu8PpJQR5HCZ9QFaQiUKRvqyd3K7X4UwgAjCq2WlS57LQ3U4bIskg65nOqgy+1PW/fmjO10BeSu
0rFuCa/hyfEmQRZ8A2uqdtmhnTm7blTj6i6SIR/xg/0aC5ZAoG2yuf0Q9VsLI3ia8HT9YEp1SJDV
9+9qWsBnyNbE0r5PrV/NJRX4vZ3ybN8enl9a4hNmMj4ORXLGfURyjGQ+080SyTH0gVMHUCtpHUjs
xFGZc3QLIuxEtbZASvIBU4Mg8/NfpBWVh6NUeCOj0MAOAj1Gf2LBTPqkOKC3vmEKPobrZ/KB1EzE
JL7j4hAfFvSip7p87eSxoG4IlX311azGxTvhwcHjtnvVEH+4aKV3fBaNu58smtwEFQxlMGDq0JWL
lx3yhuVgtAzkjGF0nloftHKBmHy/MauwkCwc9obsxjXVertNtdtiLv1IXJmyyZAKxOuPaRfxoAKm
rC9EKy3bX2U3i8KLURuhhDA9vPJyKnbcGUVJGVdhr25YpWJIpa4Rkk/o5N1SFHSBKp85ZEh5d+BA
aVCgtMMFl9iQHFwVCa/I6ikwPf/kZvIw//pw9ZPRxg5eHvy+SdAkHoIwYtMTOeA/9u4w2Sfg/G3c
aYeMFiij0HFl/oMcjuqYmyQyKYZuhBxlRCveXXDN0W9kJH4Qck74PJiQYny4E5UM3y3fwpbuAMco
AhOFki2UEFPj0qdG3cVKNGscUDeR3DsSjyfuDAzq7gRivyzh75Eu3qY0LjLMH8V7B+0eyWbyoMJ6
nobkHnKxma3mFhlzF9CXdgGB+eV+P2NjkD/jj9psYfBEfY7yjMY9/sFPCvlP9IoqmNvA5ilx/LOl
5RKBFqKHMjtlWxB6xpS0ab8XFYq/BfaS85OGPQ6ySp+lXutQT83xZcgvyRyQwRCMZtnYIAsVWZE4
GiXXOCX4+XRB48tmf84GIxXGyPO3QMWMz68Bwm0/U11jQtR5609D7gUTwELcd0d2jEjTXzQ/CNaz
pCJnrzQYkpb1sMUFRjz35rkmV9/Dp5mRFNuuKjB9wpBhUvJu9BlCUwQHWpNIZjmBZDCdPcY+tcvJ
u2qh43WPg//OFxIWI6ggwZTJ2TCHQszKuyG3uaJ004OG2p5CXD0D9lSVIGFJuWKaL0m7gKIMX6iH
DjZMuTXTAAF20BCwQRySVk44gxZfSRv5sd0FpASAReugg+9QIOlcUN6bqo90VZAjKDSzI8bBQwPJ
CqA2aK5afyJtFhmC2M5Avjt1ojSf8xyFmxxk2pvZAn/dmSBm7Hn2M6vGu1NYmEIjf15fhoMdvuIQ
i6eqSRzOU+uPFixDVsxFjUAACgHmFmKt/8TojgVievLuy2mwS1xnOBMiWrkaAFb13M3kBDrPJN7r
qRh0NHhaM0nXIqHPRy/rF1uCmf4o6QOBnkbWxiwncTTGJTWi9DggxbTOoOwLvwYpN7ZQVjbY5szb
+ltp1zEJI3TY8DaeXbIIQ6y1OF2briI9/QPXMchaDki51dMizP/+40j869cPpiBonBw0W4g2uLNc
C6YqzPOYPa4khYpQQ9XE2MXxbIsZyOQA6I2B2+R3HfiGaguRv0gB67FdmEu2yqEG4AbCxUOFQPnx
cVS215W5WYBdjX6s4Xvf63YIcryUAGYneEklN9egnkpvWW4bTnIF6kiibZBQbM4K8arSbqP/48Pe
uAmPZQT38wEUlL2CjwV/L6VxjUlyyl+hPWpwzGNUXQ6b9kMZ0lHBkfj3D2SPE6zorW8Hxi3a/lUg
YEnw06jPwu2AsInDwk0z5GSnF47+0hrhhNAPdsF2D38gs9/W1cm/Ah6D7LwEowym2PLVci6uWL30
mG4gU1Fvu+1E/FxADR+9BHe62DB4kVcKZ77DTYVW/I5WK9m/n9ij+YIt/9zDW6qsXsEhCsFK24Pt
t6KmNUZ9HtGm4cWnTN+DnHzM8xAUqLoxyA+SPLZa46hMPsDrA9JJG0Tv3PUstClxxmQF36Pmhp/H
YA8uHxcSFDRBUjHLFL2o4yabrt9w77PyJS47yQ6aYLs0Y3towhG9LIBUuAWgjRzmLK1yNr5EFL8Y
RljMpBmbjewM8jVsqPir3NZU4pwl9mlpTvjuB9S/s7Hwu7x4qxoqGyIkgRsk2mEscGwkfbpp9BCP
zNLMiygpKn53bjkUpUH5lUOeTzT1GGoXPxcCvnlwJcbGTpJAh9qELcbKJlgPKZUBNHMOsafK1moJ
SkNVdlXWeoqA4OpoutdxdG27NsNfeQlP5lX4ERSuZZdySGlOD8n968hEsjz4a/9mIwMUEcaxnxGf
pz/5UbemVPGcBNnxYfYEA5t96DSMJm3VLnvg6LotGwuoKWWDAqXJMReTGkUREk7ByMzMz9pj2LNI
3aBjDlHK37EJSR+r0S/9BmKPjTJMX8/LqskWyb4aqRBTKFVRtsFLpIgvMoTvq61fhVVlNEh0Jci2
gRayz4k+CyQgCq/xlBFSgoxdwVK4NELWCjaJNPJCrKKaoHrBMT103oi/S1nLy2E6VNSG5Ya9BDr0
ZcSGxRL8ri/VI/rgtABW1KkVqyu4RZ/Jh9MRiFhZG2s2Q4ca9jeR9QD4B3NGUuWUsnfTRKai8XUY
EnNFBdvblyQ16k9CNhXRLNh2/jP33/3OWRRgx9CZwnngazdFlps/HweVsVmY2YR743JNY+Wi5/UZ
6YRzF3Cjy3i2HkQebNslFA/+vcHe44qmx8Dp/oSbkgJwCPP1xpbO5jW/QggznYvf9gd2PEgrxuGp
hHOpyvWP4+Z5+ju+l86kGcsOmqsLOEtaAHRMj5MWX3ZDbsvsubxur/SX4w9W1n43z1XjTtaz/FvL
fJRgRXz4f+wMvJsRZzk7RxF3evyhGAaPsCL1fG/AKa9vx6swwI2xdZNLQni8CRtFgEgN5e3hw9A7
I+8b3P0qoOegYgR50t870JY28tzCo/+tkHP/86ItJirQTeipdxbmViI4grtjuIBDzmgZWFu6ZuSc
amedC5QMNWhxExB16DIeY+tQA7FMSuKQMfKrxh5ghqWfAy3yuoR6D5KUVbDeNvuwgD269LCVnHWv
+8krDLfZo0azDSnm4U57wn/kbe/vmK3GAeP8YC5a9de5Xhzb3a48vkzzWT4VePmjk0zK31yVy4HC
Cgm/oa2ZwPqnj7Rn/KHCsy03x/YvaUm42yOC8mJIdQqszqFAN9DfOO6tN1u6n+PqnvcpmOzKTz+/
mBiG9yHf1Ke3t19wcJ7NLfNKjcWhqs58gN62joK4VEFgATXYn1CGhP/gmXk/bn8zF5sOF41utCW+
Qz8qL7lIO1Qa4vVFeB6EXou4Uv3peh6UerfZ7hvoslYpV1Mh3RF2Kxta2td+Fx2oM0ZeQMY9bpw9
t5nS6Kg5TmHcCJxtFSkwtfGMjjnJMG7iJiuJGpjRVVgTZZkXeLvF3uN2sD4d59DtzXcxnOa0By12
H0GTDmA9iOeoLjwBZc4CKuhZ7h13ODBjdZejUtya7aP8UNuDdFL1d4vAqTOuQEEHmGT0qG0J0Jxk
fnrAKub1X0TfOW824XpNxSztZnZSZ8ZTFyYeqmu95InfGzHGwULt6Q9aUWhe7L/Q3c/I4c2vE4g/
phinDjDxx4/w9wvnB6+HNMLPuYM0b/9ZbhtMzawISMp5jJSUP0QR8kqynO7lsp89eup9z7vPioUj
P2xSl8vbXeSYskB4jlFxA4VJdTe/BhuPVkobFq8uFPgYxh+bZv53srNH32HL9SQbYVBj/GpVeiWG
ugcOz4iy0oQySQwZH/IT8qynjutWBXvoq191STtk3s8R5C619V3aUe0T/1zS0ZPFcd8O0Tf5sbtK
li5FCKtJy+nuXAxgA5spB6Cse35S1mj9ae7T0qPtGOHU0Ihg8yZDaK/SjmxoIYbRHpMyHVhe6qNy
0+MFudMWMwwaEoxqxJy7yGn0O361/ipCxEIyDTsHTsC28n1gcSAGgIj387Ac8OTpbdcQDVaLxuTr
QHmIudq9ZenUtO0kLr+QyPy7BkLrE+7hJUj+W+0PF1oV7eJr36FNItWvXFVU38OoztVJO+fW0OkH
RBhSNQSsSdPFA0BUVzSklhDKnYpjPKKQC2yvWvkz19tKYteWAVtnz9I6UWhDJ/8EA1X7XJoXoBiu
Qw2Lycm7OyjPS6bnEWOK/iVDQ3vOv9fwfir+Hh9iJ+i0GI8/Kp2KCTw5BCpuzTtY2r4KursEw3rO
F6PipJ0SVHvNRpWNPd42gHnM6hY4kfzZkT0ljyM8AnfJaangJDf4wsq8rMKAuJ17JmeaXjN1eQmW
8hDzGXuM0wA3yA7KfHFaKOKeLa5w+9HoMt8rYnZJXfltrk8Z9HUASBg2RRX54mqVW6/8WPqwLzj/
LEfiqMJw3y1Ks5eqlWxIogUZMSYOB50ysK54EbweHY7AnHAPIn106EHz4i1vq3FIxVal73fRLy+A
f1yl59JzNMzIFQdfVwBTOYQKAKBo4omPbVVDwpH3yxHQXO+/pwy6FlmRzQ+REjab1szYsUGLX7ih
3SEq8dDINwpKChwfQvrrpvZqIPL0oNEYeHiepdb/PQPj8rChUCqcDxXZT435KFtqfdWJT3DOO51i
hUm3iAhm6phL5VQR2cmw+AnLTb0j12YBvW4KQ4TXxI0egJmqllykJul10djmWKGaTb8t1t0qB9it
uzH4VP4ho6tU5+5A4i8EZKXKQxtjec+DxaIJ/BBhHHeWxOG33NA4Gu53IGEvD+Un67FBceajocDc
WleeMyfEybg4WA2RF6diRoO1hccOgL13+jJbH7pYTm1BAwiaW2oKbFW0sEkWASYvskWd8bA/ii5m
GI3qOJcCL04TP8xrGgzbkTVasGgM7gcy6/++fQ5GXYisVJ11V/2czFPIjpdA7/PBA/2kHVS89haZ
Ab06AQtPafLVM0f5xtE5OJZuBmKa2ze8Rl+bLG/fyDF6eAxTQLixcSBRvAubuvzpw5Wb6lpxnSy6
fAOrjTJOQumfiEWAGhokUOQ0E6+f6dPFNuMXhlPk0d+pFWUJyeRF9gfXCXeIsc56QmzPpna4raFX
B5ztNoTz5D2k+J6Yp6pfBVOFhbU9R4C/V4cm8bAMUPsS2EiwpQtBdxaVhCEK+I7TJIEgoPT1cJB2
rP+O9zldGZnXA0f9dpIPkEWR9dKnX5DvMIdbO4fXYdstRlNEyCJoErW/VHcaMzoeeRT54A1xny39
w3GQVLWpcM+fuE0wmEh4NcgT0eqhjF3ve9r5KD4VFevFOkZZB3KTSlo5dDkOJSFF/7AgUMAz2OGM
4a2iEHLMliSvb7ITmz0dOuSW18PIFLWZgCp1CO8DYCTm4F2rq7xVs4oc5xY2Jb8GpX/QrCRos7ON
cbOJV3nTy4/S3xsu66pVEK2rMdH538WARfL+AqDm5+J9ZBoj9xXP1wwzG9vGo/J8Oo7tWOAfvuam
SstmrJvv4uTcW79vdDFT7T6zBpN5dSmQIpXtA9Q6IK11t22JuQsYZDgzAqkU5tounzJrMMb4LaeA
n/Re7DPMa7Or/w0JM3naoL5U9sk5Yj8Uijcwf3jtx8WNLgz2//TQ0+YKZ1RK2P1XVQJwZFIjJ71p
vwGDuUnsHKxPOqBpkeEyF/7dju7z/W+5OIlkAeK4XaBPVQYVl+LsgYt+cwFb/UcpMZoNgclYuZJk
WgTpGdPJuJnjbGOnygAffwQcc0gdieUgZSsCaA5b26R+euftotet8dWQzoK4wYNl9gbHHDOEDfL3
YoJqFSwDVVz+oF6D9KZ4p4h8/Bd9/eonPyccmRUdemohKmbDBjT8xRtOjcoEjFGgyJ5A8EwOACrh
5OCjUilheWawCAzRNVRBZoZrfoJyn9uvLP4R7Tk1O49+ZTlum5WsSWi1J9uC/CT06Slg5kWW9rMz
xBUyM/BK9ds3dVjbdU2u1GjW1TF5svG/t11tTY2dPO08+BVIPsMLH53WvxYIqT21OcRInXPyRuuD
xIabndKAckbJJWW9xixgcjwC3sK9rQexJ0w4MmkkjZGvQYlv2HlgKi5/cRWwtIbh4hVS03VfhS7h
vD4+nHEsmI0/ERhmEdd+VZhuaSKPqnrnCDMeQRcwe3ukxD/RzddCKSx8QcApvysNwXLwatNxWnFu
+14pFa04JLcYWfWfo9d7CEUFd7aredJAlmiKWN4s/otU/Chj0x20+IaU8L4zfkvW4X9E/ZfBNhe/
ExiMqH+197sI7ZYuqCCzJFrpjL4O4iTWr92ozwQnP7JY6gwqzM+rwxYDryiTwdbBJoa2EY2KKrTn
KIXC5vO7xe9Bg2QRk2ESaO1rGNZyNk8k5fW0eD21FkxfAab3JaztrP2LVLeRxifAjHhQaqut+OVK
fkl6U56hXAqKH8aI+yVZkGXrH7a3hJJMKlMFXZkkWHlWmqOpcdP5OagWJG+enseTfvBs2y7sUeop
5jlztrCIa/N+YuBh4yXUR0znK64axcTF0IYTiMioUd2LKfF0XDH99IpH22+30OUOSKsxguxzsZWf
QmdPdP6d/trGsbf8y3KDPIsvZhAy6H7qAVOeCfMdfVwHJfY64792JFKkcvzpPpBAMpHPNhfmPN9Y
uOufUgoWU05qHkDLJdWiPRqDmNwNLfihkPdo5POWiJiXW1SwVM6Zkq6BIjqyX72rZKG7rYWzXtFK
AMPJlnSux0mKGhHJmRuU7vanQVGtn6DjJ4wBJGyiM3Z0hwnV/MP3xoNSvUjhx3uF03N7FWJSBwgd
Yl+wskex8uHmwYbx1HOA2KYViiHjuui1x8WUjOlmYZs+vf89r355pqgP3Kp0M7xntLR7Okp8XSP/
puqnr9VWfL1yINZLRjMOKjYqpDyfY0yW3uODJXWqdJcUYlqAaRnUPzd6Rx09o/cV2AvZjxX3qphy
tkFulxltDKxxERuBc9xpTuJ2+2bzUHDHeHe0XEgIyKGrU2WOipsx56UzJRAqtwBSJaaHUOx+lR4i
JEGCe51ksh36l+FO2NUya2d31fT3ajAwm7x1Ty7yDp07qCWGoXWMSOKNj0E8PIHFv6bw//yc3blY
A9eAtTa7Af4NFobNorNuy+3GuDuh2b2swLjI3xxZayedYHpTADfF4jXYhbXosRMohiolhlu361L6
wigb5sAIh3djTxnOiq664xMYaDSdXTo71K46vxYdNukGy2fJf636WPPTLsCXxHm9wglLsdZh/y9X
0FBl9nuwz7i4Jqomz3k3uyuHgEYncCa9tFTNheJVwWSv/LhH2mTh+12RMRhcuq7aRmuZD5s2TCjY
UQo7ZdXZQVrlLteZZpAXEEs5ChV7NhjPrTq8wS+w5GNGGDDBh0/Y6TZEVcgk5RnbCmT81bjU1e79
5JUj0dGcBtcJLbJVAxivWu74tuycAmqTgXGmvmmCjxkW+y/CAtbifTC7M4TzNqxhoXzfbzc58Gmr
PEIErCnByM73TV+fHfDgpr9rkpBdEK6tjAdNH8h80KXBsaNG+8mJbgXaNPanYe05sE8bEBbB4DSS
8ti/QArB08GD8aDX4pTBFOhu6A988DANqVyMKc8mLvtj6ZigLrg1d+pvkQGygOMEhjP7LP4rB3C8
P/znvx/QIKywqpOBXjYN7PUvWCbwJ6fDcdHGO4z8I00DtpInl01nUIh/Lq+6O2qGvw+WO6tbNFX4
+gv+rKzE6TwAyf4lmub4stlyEX5tB9NSaZCBYyMytAkjs5SU4BkgwZ3EZYqAepH6XiihTaj0wZHs
R7Jrk7SdyJvBYH0MWzVCf3iYQbjBfj+eTkeVRsysF+1Wy/zQVhAxTc4O36Bh7cDNkFVIww68khtM
JL5v1B2XlehPWl2Xo5WnW6o522y4+lcsTqKV2BJszM7akl082/EslYko/Z01koE2eSOfnOiWSCny
pElZBm3zwL8Yikl+Lr+bCsQUNNdyRnWBPmfiqIjv5S3jkTltlcjfyJu5MuUYSQFTQbm4JN5AP7yb
nFbr99tp6wseOlv2mbZwIEXeBGBXiPml+QdblWlbmc9GirujAYbiaATE62EfiLutLqoCfBvzmz1p
k9jLTOBkcJxoCR+GS3Os+rxaCt5OHepDCDjGcCSwkBeQyDG6GdMPCZmKl5yRdyYCRmXGlJSM4Z+0
fL/WA9LitP+Aw+j2NvwcZFuSi4qK0dhnWe5ar2m4ERijccddJV+yYSbzQUfAdiTLqobic51z/JCV
9pnPx307XxEiFMFc/L48OKYe75jMFsGeKX3FAx4ogRA9vrFDiCBz0NqkIgau7a2FweP/fOlsKkRA
uvryR2X9rSJijVdPpz99QVkj6ss8QZFgRIjECoVXH0hNvIYUm9lPPNKgy2acxlNEJi8/n3LDv9FB
xHa0fiYzftSoRLJPWblLY2k7Kh2DjuEdWlCe5maE1byhQXzcheYiyv0VOid48mk7kHgXYHBGUkIV
6Y+dh3frtnIJ/I7r7s5I8YW5ICjodYALEb9OLVLKAAlBX5ntnslxoUJsTYvT36RQYPr0vstP6DZi
y7gwjK3U/4YRVRKzuW+LWfWmPrAfVTuZvdTJxe9yOs9IJ6YxYv0HGf4OAtZ+cTeRDMi9lfu0bAUG
Z4X1DrfxQrt7uKAv/ZLCuev4g8xKwEnaBRHYi8Uqov9W+pdhJy5BSteVNs/IFksjNEAFK5u+7emp
EPmhIrCmpTWK+gsdsvVT29oCRGS+gFu9Ir4IlFPs9vTqGqcCpvFGKoIiJx2NDVZ4phUWQpBv3Rvh
sn86hmGTnGXgPodFuGkryv5LBLlD1autT26+7XJmtMGGN8TB9dSRHNeQ4VaZ73JlBNTAEWC89Msw
xNEpRDfh69o5nd2cDMkguVPsWz06vC2GzfvfKSO0M/MUyApUs8GyUoADb36mHTZvsfuSE0NohvgC
vPIjCAfXTd2iwpaBxucyhSbxnQuqVnjn3HEek50GlixOmGDSyxLL+7rZ9x7mBrLVsjh/WdjEfH0l
UeRFDSIhfKNXG8kIRqBLrI9on2vzW5zS3kcV+1GuH7d4IHyNRZGuQJ3IJ2Gw50Gs5TGUISygMs5m
bDjZTZGaAjgySfF7v+mVw5THqZ1rq+lsbBkOC/kLVIWeNjltCNSC5gpVuxkmMJ0Ei5mSS6CbD0Rr
8/ZrYnIcc0Dwy2ve4ZBquvAaR4VmkHEcpKRPlI+8LL7r1oHOskjEDwc2FQcM5Wadkfhy+KbJtLRE
Vs7Ly+x38vJnRznwaaYL+ZpROHKEL0fHMeGaNxBvtichHPHJsvay1OaM5E6ytt2CLZ7EACQ+CD+b
rTbJmxBRKFrL4OPEvGnAYOCD8oAi1rb9o56pm4igPh5e6sFtlsoUAzwPnzMsPLuqyTLDd8AZj9kK
C2MxAo1moCsopKpf/JIbxv9JBPChUcuk92EBwJhENwxkMQ/sMrW1743IketF6awfMYko+iCV+RpE
+yJdrxgKm/3g+6iYR3d3bHe+50BKhj4ywnpzdD9FDi3iZQiY9+oFn/u+a/+y6j+5EzUQcFbes45b
o6s2HIAsaKZL9GtT6nqK9qGe40yipEBVvCoEpJxkdcH7tVAuYiSDdUYfoNScrRab8jz+h4RJX6yY
Nw9JLhGoBgfBT9fRwzwGeI9ty5pBr5XHvSowSU2QrQDyqTKMEG1dmzhWcY2XHepTHm5Pn3tWwx4h
W/MxjOVbJGy2tazYxRGsreW58EiQvUrBeqFLl1Xf7nIMf5bdi1ZBlJdkLrovkbHGpa1tSwzLVdoK
Pzw3YuXY13YZLSTJpRA34UHNj75IKqjUOm7jLTI+jbMle3pNIZcZKH5xq7PziRt7HRTos5Zm+1EA
Nbb+QryjoCk9iG18SeyG6X7RN+sgZaFiQ9RtUABB+iaS2ldDt6eaVHC2xx9I7puUlt9rus9kMYWI
eRAvC4NzI/fDX1LLVPhTwhtOd0AWYGR4LS1+4x1z2zesy32Nn/hQxjPVEGRuxEqiv2LO9xaqDRE2
0hFQEOCoeSoDkeo6VFw1TAN+Xs2MMFrQqmp6eYLsy5YMKq4zH3xS3/DcYI2EZmxoY/wryfclwqI5
rZKmuGz8vIuSrdeE4zC8JjEioWgEPBDR075uek5qjyyLMWw+Tqap++SqDjE7Tq9gwzr6jrUal76d
3Bh7aLEXR0Js5igH2kFuoBpx3khT566tMVj9g/ydylpG8SeV2QWYDE/LJQeO5Qj+D7iNEZAUhXbh
t7jp/8qULVRAFt9kLRksk9N1UUXBJRs+wlrfIuA8nvOmtpYmEEtPJ1Ib8hEHmXDPNJPAJP7d7+Cl
s/VlXqCrA1qSpq4EwzTj4wTec1UMcrBQ4qM+SF5/wk8OmtoG2VFUtAaWsFb9uuly07cZ+9Ba5xv6
aPNd0qbxZG1VibWKYmCyA2MEn6NTKwy/re/I4ohChGJC2j6tm3Tm3z6eEHs0+62EgW3YsbMH6l29
jwyyi3EhKYT+2ZEh/P55earn48OQT66HgfHIBtej93X6mvY9fUJxhTWNtNj1U5AYdf9DbUWzxsXt
fYEUVjugeN8nkHVEgCjxtuemkORdhcdvrFxjYfuDQ+BMGa8hGAaWMTZU7EOY9r/osDNCVF/cuLJ9
miwof7zVaer/wUOTNz9hFZjVNy5UGoA+JppqrYTfQy/Bb/+rUDNKVHw3XPc+n5Y2KmFMtMgIsPAx
04EvbgPNSWyyb/lIFuj3nomLxyr0t31R2yoXDsLaj28IXYFRXxOrryBkJ3RepRT94MZeg8BvIIg9
LfDbiNM8kfaICHcQ6gO0sRrimewm+wjRGlv0OjDFtNsDpJ1DNEhS74H0IrP8NBC/XrJ38XcEya8z
VtA7Xi8YZbap49AeIDmh+p5S3iotPzQQoueVbfLrsjv07GimWmhonJNKLaGMS9QDmvyXtrF0n0/9
lyX3n4lor5JiXUrEedTiQEn9NtxIU2m68s+9r1iZVR2jc28OKG6I9bMjEGRV/l3UkHd7tSIrS3tI
aQQbRIqUmnsRk1oNU9gBT2rCH/LsZAJjULMGSB0hZ8v1WpWVBkE/beu3KvS8N419R5GFfTx17bWR
pyHKanhLP/OAHG96XsDp48iG98tykaxR4TCW/Pi08cdXjyproOxQu+KRsOW10SZRffYdvbcYI/Sx
3lrOU44z4z1ETn588Ggna7hVHkkYBl/0yAlcZj55M2dO367Ce3qNQdja5/6SAlUaoMbL/pWnmQgS
DHP7cMRzWOSGSuERFH5UMsRnijzgsDw0peBEJNJEpcJqrCRtuJ214A6oYRqOxCRFy3s689nsaDQ0
XKR0ux/hXNOHMZ1OPcbjarHoQSADk9ZqX3ah3rzG30xLIlVPI/E1I1DJLyr/2YGqWf8eItgrRiH9
9LRnff+5xIGKBSyYeTKRUyrfYWxHjAyQrOWNvQ3mmfWII6Z/P+PdcU2jMuF32C9wabI7WAmAqiE6
aJv3fzdwpHdJ0jc6wMHoT/+JqXDyRgre1XgZUR29JvBxMS6BzNcTiTP8futgqlZzuSwMTOjJ6oAj
U5d+osfF81+oP0u8wZtyf0Q2LhcNcUBvv/TDkfxinsdLRsf+Zi4rvqeMQGEvKetEMchmrfMs02EV
h9nnAyRodNLfrtFTC+ab8Yal7+fn8tcL0eYlFW/h/UPMCLPr9/uGxLGYmi2MRwf0eL4QNjLE7XI9
NwyYIp7SehFzPAyoD+YMoausMQSGkbCg8FEPFdiV2UIEdgawV8r4HYU7U0FfnDRp0fc+H/GSPcZE
W698Moj0M6Sp/hmHgBddU+jXUCXoFdd786Et0jQRhAKV1/l8+St1B0c/kKnHAzUr6NFOnYAB4tgo
vcg5qvz3NL/BS099YiRxHNz3WZ3/MlB9HC1UkBlmN18cKs9iWMMc40i0czRUey2LdcwY9BTubK+V
BGQtdMMY3KyaDKedt4OoHkQi/hRgDWLc8vQpSDgtS0i5XHIsvkVkg7CnBK26Ye9ctgDza+UhOf4N
ssW+zG230jwCixfsufHPnWln+wqQIOzh0/2BCpeka4p/xCrg1EZ5PMduNr5J9xN9RFOE0CCjn5JF
98OnSaJu7tIHyb5YGAYKP3FJv1Ce59OxyB6hexnODQSy2KykPfGRJNlU/u1GSBRefur2VAhzZkpP
o9LiCoVgy3vav+rv8HPBd8ZWwgZjPImAfdH6dc85WOBJJd1Ao4+5VpzbFc1YinRuTpYRlIG+DWmK
d9i2NMYIwDJJzBRe8ol1kB7jqxino36cOdgaM8l0uHjrMl0lYRI5olMxl4yo/xzgxz8uLh27FTJ4
EzNC2f9RlGsHLhcpR67MGeWyyB8UbKhE2vwpoMgczfQ+eCqtziPe2+zkXa9wqJwKpTqE8DUb824z
xXB0N7Xhq2wDhcNP7kyZoDY7rdVHrE6m50YFyUVmfThjgotrmvDs8aWxJRth2wBIuucHcJgYCQDO
nKXJflhc2m9NV4AaZOMPEesyufYXKCGxJc+hL9xBuNUzwBhALRqdkG6NQMQxjH+yap+51xFHt+ZT
lv9b7CjECBYRx6ED8+Zq74snK9iI+GeocFLVU4B94c9a1hb/YB0QSWfVPuJhxmk7rKXDNasR8yc/
CnNgMS0XOt1rAGUWerM5P6qm3gs7aodKRQ+cU62OH731mfiirzU0NXqE8M03UK/jjF9IHwZiBW0W
ginpTUWhaV10zipOnBxBvPyfgnIqQhUIu//qZnpOOMf1M8rdkowOJcp4ODG6Qb1EpkeXiNTDqNpZ
Yw+pQMq5IV/EdRpDhxCdhuc47R1Vh80JV+SoEwcsf6B3cjhKwwPOcuyXFJ0zKBpMsX2cPDnsEpvn
8BO3U0YAJ11Ot0LQCI2yff4xa4YM1Lr1IdxGBaYf997NbwnQrTYUY9x5+2G6yRiVwZ5lx7ZRb5/E
bMJrANthT4SlVj0l9XFQnrpZFGB8MD0x/3Z7az7w0uJAj1/GpKm7UIrdy03EL0mbYPpdU1FyHMNl
vBnwLe53mFMn5hv+9O3wX7U9KsHbcox+akxGTzZ6RSeIK1chlzwfVO3HA+Oty4OCH5g4LGL3K7KY
H5Ci2SszW748Z5XU4D6xls/WGVKRFj5Sl6cwJTgCwuJ+jcYY2jgA8Nsh6gTaISBqwD4YY8RDy49S
vU6fIu0z8CIXiHwyQ+gQos9urB06UPpDrzoY8c8vOWo7Fd8lLG+qi8OPNqK3IzQgL1P8BFZFxYeT
ynR5ufTsYcXeHIwerRq0rt4J544ka9zo2aj+fVpDWOSEe88NbRHW/ZazDg8ToZBvoWZelJSPkOMs
Y8rvIMONVQ7gOUv27jacxvUZxdT66qrIgi4KTE23ByP5evXHa3ihpnawZxT1RQq7w+t2xszKWMZ9
IkPa4KN1Y5BiV3nSe0jrMIIs06lTLFvphHf0MHNUF/ZXQKllwPVjbZsrYTqCSXKUK60mhXeGmUdy
X0KXVYNAuqg19rmjKgUKgzJggD4Thlji6vvF8yUILM9b+/FD6hZ7NSNjLiGiBHOZ8RV1oKoeRw1A
9iPXwkQfYk25qV1Y29P350jRso2d60Hb5qtKSFkRyEKMlvCY+mxUIua2XtZW4ulQFxgLqSIaC/An
FlT2b1ayv5Byc99ufPvfZ5WQyysbrpZcfxWC1XKg/W0+2UFpR6DXKir+/CBBGVu/PLDUoNRbUPXS
oaefJyaiN66zkafP2tbWQK4v4CyHEIetmKtQbpY5wmmWOcQInAXl0oU2pI9MTS4XGhVnBM/Jouk2
jaf2slbcpemz7GBEClnkilACSV4kJkOOxXEHQ+7aYb2U3gC56ze0mfVJF3np7ZdtZfpen2Lb1f4a
wZRe9qtF1a16B0A6iV2E7pOXx06SFb00+WxqAWuerrLr3t0XY7f2kSPWpXuoYsIKLItUv46zuB5b
o0im+g5LcxOvOQ5cNhsHOaNqHOf3dcFWrw+AV05EhpxRj61ZHpJ/ef5HCKPe8O/xA11Kv131SGZ4
5nq9OGXfquQYIKWGZgPBmD9Fv2up0VlLRV1BHWNTw5IjJT+/APpI/+jpntFnGeegW3EksPxhJntE
u24bsRFxjMHNay5umkuCfmxJN2yzznLBqwaxi5r8zzvY4oFA567zozPiMkCBR82tLYF9POCFj/4M
tEY+JdntFOpRj9XbNEhr8BUI54pN5359+I1pVxwvTt/eTb03GXLKTH0mCsZqRuWdWPqXd90AMXC3
Xr1ABh7MZ09SdssNgnvgyDUbnKtXW7xd0biCultblhKbwcy4ayZX5V8dNl3iGbZSZQO55CkxWmml
iyn9eN66rFtIoXsw2+5zT78FhGgEHirkZTG6EGV6FsDMVOJEIxhr/+7z6ARLYg+7hURbvLxI/D3Y
iJ+4FXfgkytlo+sC2ugTT9eFPZa7ftJr6W49Xov3XTPPX4x9iNpBZC8Mp5hxKFHB5F7Amm5uciOQ
S1FxvAB5s97Bi58X+DQ+fQ4pMrThj+YKhkvFa49HJwhW6UyHEHu4z98YjbVrY5T9eMREJOyKzQ8V
n1UqC53VkyVePZpv3VZQilhBZTser7s6yio62W2vHF1PQ/gul+VrZ6LhwefO4Ry1Kso2uGHq8LZV
uSsevSYWRPbEI8fd/hibIREFsSv9RzHwyavg8OVcxFiSfSZnnduPUVedrAEM8KzTxKb01tf8m+8r
yMREj7N9jOm+tCDRrFJX4udsqEMvaT1JWwoq3MAN/KeNn4/OHQnPbfjwvZ4TmqQ0ITHC35XSt4Iz
PGg1pewM06U5vI614K4D4xW0hQm9olh51L3uXsHPZ9eR2xd0Q8ikOA9Av7olZeqrs/0ZEUEzs+yx
79Mh13/O5GfPeOhIroVDrFYPv8qZWRCUWefi1HZf1jWli4ohr7GjwrCCiN2ch5/hDNbflfUbNmNq
WqAcZnFCXvRUy73XJSC47ONjYcfzuZwTSGvIo4u6bQuKuEj1Ed2Qc+qHZ0Cxtv6YuZ5c/yeMtzYc
3NIcv2LNOGIrs7MIpo4PUxiPmhlb3dCLkz4zN6RVhiiswZjwATVTJyrdTfYSlaqJaESB25/x7TcE
0L0Vx94qtfj0vi66NHCFY4YvHDJw4zaKFdpKCbB5T92Ze19HVT3rKrwQwgYqeYAmnmUIfMhd06VG
8eTY8jXjG0i63YoEj7pRbgbteUNyH922D9jSQ732tYfpBtkE2ewNpamK1BFYYmwOC3UYJE2MNk2+
emZAurBKdGPTeYHivfzI3my86ga7mAJmiEqaYOoSHQnpGdVWYQeu5vO8IaF7PuJO3g6KSgxRIZKB
Jjo0bCvy6eAtNVdnOGVuthu5pyuoXJCo7ruYFzWQpxTeF7kJlrGkXTeWtUqbmEk0I9HXEoOE39OX
uR4A1ek8BkYX1YDtlxIu4bLLgjUe4j7d2envVyijUA596qjddG0KRC3VIa7tI6TVhQ/WOU4g/2XP
zO0IRCScrPCli/U8re5TJiliaV7vkQqC9kHQA2iJf2cEtKZqMHuvaMeM7wJAcssiz70s/33sXryN
7b7t/NBS1na6j2H3NWLooZq3TrISnL/MtT5k0VxgtUzQ9RcB0WKqkWQdJUVTEfEHsEoAeHkx/yTl
X3n/EeSyJ070v7Xi6pccC+suOKGlOLQjRQykj6Faxq4gvI/aObUCMCmN6L/cb4rLfpdycSfoKZ7W
nT+aGtBz9GXg+TCylNTGyO3PsPfr9okFL7o8T6lmCjBmkrlWr6fT9ArnK928ECvk4xRvX9TDsslp
ToF9twW/cnAHulssnZ2byNf3xHlxm78xASxhDbTWRE7hIDQiCXXlXdQWmi0vxDQCMaFDEaZvvZIt
OQuHSfhEmqUDqua5duzd6EWUCktCiqJgwahLko4hV8yTvSL2UhSR205zL8MCe7jx1sU6pE4OTBF2
glb46DaNpAnVKooKCTIP7++yEPCq8fuJjabiFEAL/+bhllmSNUgKwFn/DSjLvQb4WVZNhWDlP1kI
0wF9b5XpaktRSIO5kWLzLB886bIy/Fz3jDeNZ5XPIguY0vk+Vgw09sKTTHvAOwR4r0GXfSxTtuEm
yJtRmK8TKRYy3wajfLGvM27qJe9iuXfy8KYdIoyzpj+8kAT3Jz/X/cTty15IVpTS2ZqXXlZiq7jQ
rDrzrHPhuZEmSGqRBrr/Hq+nSqCkzrHKi+SUFGztkd7UraUavG9mkj761YLJT3FnZI5qWcHfzPx/
0ECXDjoQvb1gC785mkndJ53Sn7J27DVXECuglqno4zsTzV3N4rLSzaYPKHXHWdsk9THJBy7qyd51
K9ubgGH7gaZgLStfd8+SSecAZiKAdlgZ1bhcvVpyw7nh6AQjSYck2w5Dh+S/RzAYcukKXTo/dcb4
cwJ/tCRTfsEii2YX/yZvdwKmqn2Io9w/TOMexp+mLhmCUOgjxpjtRW6WEyd5awgShBwM2JCvlg56
nrsTV1bpjIc+S3fna8yszknlYrNtAxxzwLCtsLTmovKEH9DTunk40VZercOxYb8qlzGSZBwXar+r
l9p5lM3KZxrnf4ASjgkYiC8ZtJSMP/SGrXfrfsko7ZWt+UlxihssGwnLweQmwXH9OBBTY8AreECV
fdGNye+GasBY/7fv46afY6rSD1KzpN8EhnvurmbOrkVA3GqqaTZWm97qIXaloavL6um/UHC8y8zU
cRnwaegohP8Su8Ft/wXRih0Kx+mENR1Cj08IyL/A0SLCgU7Q2IEcFzbzvd0U0LTLK2DK9IWrKTw8
QcVrA7n6/KUYR+FSxfi3up3oTIU4iewwjCGxkP2ULVsqm44DBHMGy4/kfStJXoYwrYVqh3vdDY82
DIWKl5H+7ryQBW4XO2TiuFaNlSHAJbotCGwadcuuoHatWscE44kCUmOjeA2pF/1lP/2/PeD4Unn3
s0sHpaEv3MLU2+g6jIy5uUC+/b5f5vvWkpAX0VE29lH82Ql2Aon2orpJfP2UFLDVIGFmLq1fzx8F
OwMSZBfR9eNevawbV4bdfLqw7BSZLPEDZPQBc+mr2FSY8WZdrWm+rkFEvIhZTKZMCBc0eEwjRxHu
SSxMtnMn88QlQp48rHblFORpbs0/icuA84irb172kJ076Fc5EjMEkZoeut3zKwrGip+P1tTDm5ra
OcZYAaMxc2ySFLpelPFikgEnzsMN0qsL/RQ7LyRUB7XcZL+xUlIVjgB7U/1DEUf2b4xas8PHILBr
sIfbjqI/lTkdVbBn5zQnad+nJ2fYWKJN/LeSba46sdRxRJK+hQpnUiuXSYr6wf9cyn+IsHODUDRk
/FxlzbfYH+5PJEe3M/ZDUlcNc4eKUtib9V4tLzINzBMtc+80uwEWpuHRANRmjYkhFRFp8h5KJaOW
Hh4hVfFsLY/8BJaawhAw8JHH/efFenENqzfJYqhEnZjfdqwcpu7L8iMC5ibu+DlCLYuIMj/Sy2Ko
LhxckLVa9TEn3palYcAc/O2ceY3rU8EFmle7RF5lWTBkQlJfWxQi9LaHFUX1r6RBHf2INKnrJb15
U9D+rNognSzxifalm9YA1swUm1E0qySCTW7sn+u/sTmAzPoNHf0qFaMBp0XFHZ7eyoqniSleQho/
sWa6in3JBhdmKd4v4XTP40sEvmvIT1cRkEjxfSnCWAM7kh4c9TSW96rFTAm/9JHThI4/PlcuczFA
AwMWzZkyqdAupbSyR/JtDUQJwZTHyo6yZpU8cfwtv21xQY+6EnatEdWhzUZHe2k9fSUJQ3W3ICso
vGGPmt0gN1bav8dtzELw3oHL0Dstq9ct9Hzskj6dO7KS3CPU1xdvv5aR7T4sC21+ZNDYWjCGYBXO
KxAcFeaQK3FGlNAUnCTIYhjiN+nlti7Y+oFtdZZX28MudCt2Unlytn+VfuBPF6iUYLIP/Y3J7Ncx
szUQs2V4BGlBHQs1SlU5QupBcFmmQ+ZP6LD7oQg/KqSF/mAxoqitXJnmiF7uLc3+49ztnmpSu6bn
9ZsX46IUQzcs0RAHDESv4fMl0/HlLRU9P8MZPm4AIx6vmUD+XTKsxGVYUWDNvORFqq8xvrwucHSP
eTnClHT2UQCHd7IvY/nkM1OCXhuGZENTf/EsXcxOnCda+5PBBqyqK1sgeK1PYfVnLJF8mIdG6Uad
uKxH+OxCd0rbnB7Kgif0LJeXDXZzWFDG5Gf+MgMb5KLbJCcSb/7SBE7wBzvp1WDsuxhX4DL470u2
Hgqofr8SGPUekBLSzqqsNWf5Lbc7UQx9kz7fXtJ5tXo5T3K5u28JaLbpA2nxR99//qzE/UZg+hKZ
5HXBvRYw50C6zcc0bmD2SH88GpHgXsIgSxiaiFPdS6lJIMWMFCCs4OAFcArMbfI7SvCN/Z1PNxi7
3H4q3jtJk8yVJvpcfmB9dSnPu8oX/15C028kqvqhS32jKMgDxPDQpiseiAwb4wsUFu1iXlfRiJJR
kNCRWI0RtwbJ/B8DCCfr5NcpHrUk9cSQPp/0Mp2paayga7LgxtrwqF3b7+XyRWuqXfGZgqupAmn+
nKy0nBMLGh74kNNQFJTQMYVXj9YjMSZrRqIKnHeRovW3N9EkAHsQIVGlTLeixJBJQBkaB90df2MX
JiGZhIleUK9Y7BNQ5uT71norryXI8j+uC7tl+hVf359NyqkNlkXzcaXlBJ4YadXTfWWmc2wIf6Le
nR9Isl98mawpai8M41S7musS/AqPNbIua4kpN/lndIjOsXbrzQFwKbd1XIaGonRaa2HcW7uEQS2v
XeRkUN37EYjSvJ7TyIYtMhsjZdaGzf5Ss3zQ7fitQwbhHPtEI7DJSwIO5kX7JybbcOzgO83gmsu7
3zNQqcSOdxeaCR01mq86FPRrqOflzIND+8Bh2P8fJlR3N4KzKtjjpZechWJdqr7MOJ3RoMu1vO/6
nKBEIsX8wAYVUDlPSWNICGO2entqrGPR0BOVwgB7NVTrnqlKIYeUvPF0pBIJ1R4b8bLJWVsbIDNJ
qmZRhkrbac0Mp+haxczX77ORozFCVhSN2aeN+Ql6NAkwuEG/+M/UsmYO7vUeOpBw0pqpOjWVDFg8
emcrWM1NhxTu2F6YrwXrfc4VZbsYhYtk6lr+INCMGQ0D2vhhnGmfcaYqfQTRUs5ynWdim4YbnQKX
vtMfGZEjVN8WNGhXtww26C9R6fuggLaeuqzM1fpIBMvRz/GrDFd2jjA0HsElZTHnKKHHtGbLMHHZ
1RxfzQVt+2kYSpLz2Imdlo5wSzwoY16XTsSQfKNyChuzHkTLUVo8c8/1Cdwkmy7D8dwe77MPf4tN
Kxc9USQ8Co2YBP8qF5FiMsjG+sY541b+R1eB1WFSvsGul/23GyrnJet4dANWcRWb2MJTsHPsMJN6
QLIn2UNqohqZp6w3LiGfuBvxHUHhxVDv7uSrB5y4POgWM4NJNEZUVU5kmiPPcQYHqmhku5TEUdbf
p5LsApE88b4e136jNgGPto3poO5fz3uE/wuBuoPqoqcqOjkSAh7dHYGG01oYd68cmdK38S33MXXx
+hPi0gGrwRxTsvKmOiIOQnFp8jqjgfp2fusS3saYCzAqF1LvkpFJt/4jVJgXQR8zkr8Tj+HTpGes
uONmpk3pRKiC14QxeltadgfREUM0EIDsacue1y7EZVvYD/7e6cCHbUtGvLv4rlqHpnMY3hb+S/bF
5Bynm5DERx9x0OZyqcPtDPpRmB33gvrTd/3f++xB7JZpgm2F+aMhIGkrS9q5pPx3LoR1lQ0O4nc7
wMq2gCUJmuGdtq4juF98oGgcC0TA6ytIpXohQBwZT473+/azJwZlMkk203DRTsRB4xDwO7MTKVqR
IqOw12H6uadgQkdAmvpHLSPjg4KBgvZ/O+HscL5PZbXpqZ0VlNH00TQJyaM9lPEtT5JqLlIlRjvr
j7u/Yk8zzU0eS3vwNwHreJFusY177deLm2GwR/8FbDvK80PwsWWKmZnKpC2qPiU3JVkLiN3KSSg7
/vK1zofGO359BugQiz5W4VI/25wdvFMOUus51NcSMLNe4Dk1yUt3YgRWiVj83FN4kA5N2lJkmt5J
lFdn9/otyLWzBnGHq3xeddI9loAapQ+k+7qUWE62GaEdKX9ulaYQJROOoOe9em1KDppjUXpmEOcM
Hi9nNc82OtVsdrfyCTHu+XgMriFvxs3fRUEo+H+TfUZC+kkWNrZeG+A7uBMsJ5KtbdR+zSSTIor1
PwAlJ+si61bJV+zyAF+XVVAU2oYKgzxgHeUwsTdUnaKILNsFJypwZc5XUhKa8G6/PM7d0KNekBYV
myB7IE35XaolO39tIHloTZS9PUWFQikLlR1d4MB1QZ/cYYRxFmjO3gr48z5XnD9/pj/RoFXiDd2E
HtO1K9Rf/B/oXoMOeILwxld7tXauK5GcWOOUh/wMgNIOY7P3rklustHMRWnubbUHUdB1vZ4BI1ly
1sKeQ1FRJ6fTk0CdKugpldBaZpsOeQEhqRkwnxu9zkuw4c2wHIh0/rRI2Gb91GRm5UI0BzUxnE+0
clwcPzdO/vq3OGvjqdbFriv31TlZ6mhRAPfTBDmFR11/zaZVCh6+7WunEjb+rHcpTiVfsRF+/uOo
fV4vgbzvhy9m/ekSg57ux7AfSZPb/Vmy+4UUTfsrwMovRj0altz1plaP6sZDsRnimRu/GFXNIRZ7
9tRNoBdGY0w/LGij0g3Mhon2H+p5lCOSuSoqSVEJe2Hp523DWp+WLfhAtSWuNaE9IDI38NFstsgC
334FoV3ZfRoGpSEpWs0UEXEry17+yKr6O4lEGns79tfYgiqipcKvBF4nyg4A04QBjh1ka3Be9bLH
d87wGEzAUhSu5+dz2K/Fk23YmBCTtpFBbCqJ6GYQHA7wTg1noenJsZqVl/By7ftTqCVq3RozWnxq
C3TgYDiK5lnJ3WSbb27PDeuNyML9c0/OW1+yLGR0tveB4b3EHjeUZgoeie+OZvpSW+M/cSdRzIip
5twwwPvEz0Hb5911TNESxd1Ye+YwiaCUyDNjDzcwItoGseTsbEHF+xYEu5hz4wpobc5t+YHgzfER
nLEl7Y77uQmT299YwUGxf1+iFKAbut8aAXGn0RDGDCpSYESreemfYlzydAv5h7PMvgQBR2KYYbEm
M97eR19iGL+rhyzTR/qFo+qYKp41FtKU5AYZC1vkFNImwR9UcBDPNj6Rh9u9Us3CS2WWRC5URFId
YAvUgAFi1tuCl50MNZWKnkDqR+63qryuKpDsaoDG44bH6KujXuIlZyMum9bwLtg3AZ+BdLJ9+qq0
2qzUUvHf//w8EjK4jAWvPa+rEfGWTSSVj+aKTDsCSsVwQzjvDwox0XHbyxGhlMAQIrVIc6dlp79c
NAopn+ITl7Wop+R1tHlufx/2d1taNGps056Sg97xJk72wlQnfHCT7BBQLx8aZH4PIKuypOVqEuWw
Gwd62dO6oVI19hKC4HyiXZEYaeEK8mgnZSqrD9b7YkXdluAgUg3xuAa+vdP18FBBPkuJDJ55l1K4
iLwUhqncP4h3U5Lnik/vZ8elkS1JILS2EFIeN4bk+RHFX/ApuFKOa86DtySekjoJ+yKROmjbkPGW
jdPjoN7paof1TJPQ/vheNZT8Si4iXuvuanFpQqocdK1O20fnpUh/PfF7MT+v+Hum0SgG4vA8coQe
464eVDLof18Cg6kYZaOHU/2+DtxkCclcm8NmbOVFDVdUVxrKhK3mnQppj225rRHivfIW8bdu1Ow5
9tyPL0e5fh96WO8Ms7LXGVcaCSBKPm/tTCTIx/9i/7/8ZhQOxZmRz17F+KtwVFaHr1RvwsXHf6jF
2yOJAs/9vs/cGN9sJQwM7qWjhFEFo3XDCW7EsTkjWMf8t0q8aWMX5nJZP8kBmylTpvBzBPm5lSVC
i5Jg1WLnBwjdU8ociqaoygWalQbwS6y5HzD+D5uEHgPbrXNEp9LYjsDDSxy0nibIj+9y5BoesK6t
xUVZjiztmCA0asZG5HUClvV57MAmZvuuVGoTCRK6pcE3eie2MpRnrLDFCywMgcJPQyNmkVAIY8Ku
NFEPrmwA4kZBkB6W0qwAT/dGoaAcaSZXZ4ArMVQGc2tmDnzBOozfblclluhc267CSU+R1AepeeuU
lWYvirmbn+HMamAoxhQZ971RTNgp9Q3op0qdRco+QHMA7ML23k16f4O+Z3EMok2oXzqDNM1nZyNq
bvgsfsXowdEukOl031YxrwQQ3xnmbqFSbvxmQft2D8sLrQmGzAVlcmRtPweB6bfc+PLyjSkeBK7c
op/5Vr134Xuz2kXmwbE+HW6BfSR6EiwbHrlJe/u9MI4xVGbaaHC6J6/cT0ad95PocxZEmwHeVUu4
ODPveqgqraXJj0Xi55kkyndnkGpGdrK4ikQ+O8Qq6HJfzW9J/o8zC7rVn6CNn9NPvdPj9/zALKR/
k5YdUFCNLUHGn8TzXLrsR+tHo5LjsXtBIA3AYRktdCWksx3ncLe3+K+vsysgTziFqqat9YVZWQ7a
WIcj8swi8syy0gRBIxd5NleGTGr3G1OOeRqkfu/8r7vP/iiKiweC67jKD+oY+IwV2UPTXfkHVF1N
+nEEvp0MzaL2ovTZNkdHS2GFPPyCx39Xrs1fxmqX5fSbTtAbaPCkEuLgoC0/GMu+ALSrhrgbVOvg
Dwsc52150EZwZesWH7h0vmSDf05lqD4WmIbzSsa0kyN1B4TU4HEV8AovNE/phcSF4MCFdeRfqniB
pHppATQOtSxBDd1NWsmD0RBrMlqd+5xGK0XJdynE2O3LPpDXK6x+kQreaK1VPB+fwiwt6BsLGWG7
KNvR97WYyGWmk0e8MUbiV6dbxk93R/GsVuMdMEGVxDMoQl/tQtaXExwteqkr9wih6ZekCJXcI7fY
9ymuEredTcv3a1zm/czPdAExFjnHLzqaM8AwRVfXdFEyZFHRlyfvImFKx5HdeGc3HTVqfZYTx76n
pgIMEcLz4YpeqhKpkSrVMlp9TzY0Qhi8/gbzs8FZQtFkpJ+fLTYx7JlR+0u/SeQMnxDsg1z5xuux
2pZ/5YIACTCcMyIQLodk49oL67R1mvKgoLz4VoUA9lesIk3VyRj+BcFeIlBuKwKfw40P+XqBNQwq
UvDGUbCmF3DJpFzl4682aw7CTCrpUPPahUlCNHXOfXPsMN21Q24J+HZkgspaXd/BYjNOad/PxRkT
GeqVVF2jRcIIUgaC+954y6sP1tH2cOdhGAq/9l5/r14tOxq3YKMhAWj8gtnbhgV2Hl72A5LYRyuI
Mc8IwvqpnyEmXeMguPC5LpsfSf+eDuXHlz+7Rtcb6KQ47vg0meiSBf12WrLTEWBEDVf2SpLoLVzo
vlcD5yOL0mKLQ2u3MuDvXCbDHIX0pV6cU5W2q3Dgt7TAFrv8HCLeOA2+cjfLnOlpnE/1QCVFO27S
tIBs15OkLKEa7e7NqihaXY2o0+eATgXCsNWbA7KEVC41gbH4rRWG5YGWfO8fbI0kK/esWoishw7k
irJZ6pN+A17glXaILMJSl8AThg7oIYrdqKRNu93naShoegwJ9CPV+ag8ypGp9K8ncpu8w2ajY2z6
ADL6MUkArwwyhUFD9FFjRSGpn9gSrydJRJPzf33l749ow/rp4Qgp+WjstN1Kq1JEhgFdVq5oJrDz
8P8hiIphGa6K7F4+azETmmiHIob7QRjKwKW+gj1P7rsYKiZYKTjMPEQ7tmpw6Wck2BN6LD7sipdI
VYZnTwN66d6KDwegB8HWkgA+L9+0zZAi1moF4QzVn9Yhyx+MtkX/eUstADgfYIsoQQIg1Rdazz5r
fynd41NWKjWTyQZ/UfpDYdjRq+NgjyxAQc4JoHHNC6aJkKNArWWc/ECQVL1M/LVl9ZzUB63F4+1N
JRiBzWU08VKPy/XK5Z4N7+Bg83CdA58m5GHRwxpIbil8HqjIgB2FbnzdmriXtkrvatvEUH6MPHn5
WED9e2AQl3j/BFPi/afVAFLpYDqu6ghyCJEFn0ah+MiJjmkJN0Y2D2jXRNk9gY/Ni9TGUdfrl57y
jLatqtZ79l7jKTPk+D29RaD/ZdG4iNRMkFxBB+QKCLVNEZw5ruT9dS5zjk5UhBE9JmjLbOXWARAX
GvMeYd7drNpLpObC5yZBXtzrtm/c+n8ijvlSyGY1tw+0Xh+D2Rxrkx0/+twaymqvd+xWhE0xSRJP
nNs5SMGnfWr453KzS4flSCdGhA/TdEUkqqMdgIU7z4PZ0GgnqL4SBP1UcZYG1XM3rhcK545/TxKF
cwp8pfbQkvt/Okpy1rOmXTTcCo/8gWkXS0kiZNIX4LVEIZ/eULbmMzb6pw05Cv3N0yfD2F7ZFLi+
8rCEoZFJTp8Sv+p+o8/CopwA/Fi6rZotnSLYaB0uBK79yivz4EfXdojXbpAuTPzqmZa69EpIPazL
CMMmhRN+JWt3rjE74lQ3rCbD254aSuZh31psh18WRguaLJ3Z8Kxc8JCYkgoRFuA9hOR4X+y8UmM+
kLaIg7fXeKhdcO2xzT4Xpu+Yi0NUsrfjBXJyVx6Z3oGw9EXeSOmv0LaQSlrZdn+ihgSPfWUWtdAW
eQTnsMEw83f44DbNnZWe1deiFHYnfGkzciMg5CYgzjrjE+jMKt+5YLlMwYOwRbsRsOzvbC0keFl8
58ZnmrFhg9zJRQxZAJK+8tmVrioZLFGtsCe7S5NPPw+TF+SWHW+rSkvAp9AJjT6fOE4Q8w8HGrTK
E8a44r8xIJBo8VRN0N2oJnlKhB7eJIaGjes0d0mjy1gpQZbCkEUrsfKfazPus1LfMDDPzrUhfBhy
T2ThaGRjSboIs2dLM92+HIAe6sg3oJwXYoJtD/JPQsOuwPwi4M7vDTdTG0v2atw6Mg5MwFhVJk2j
zQ48oAQM1xB1r6PjHS9B6t5rc7VZBztBe8FWfc6Oftva2OjuwsESvEtde6IM7B1rIui8Cc5yNHOU
PPWeW8sUpopk95WHu+E9axNdvECGanPCH6qYG1/mezb5gKscgSfgd9Iwy7P/S3mkH0NpCjU8lhu7
TBNb+ucGbHBT67IpAu6kmAEASRiiE9fW3XlT6Ym0pUksywyxsLCesEygoT5IRtd9592GLKpCq7Pt
uUm0SFEIl0YZgZ6WHsJyotlijQtZDsk0UhOyqdEfYQAkALpXBjoxBfvBK6MK68ORzynoUuykXrAr
jzNUQJFfuz5Y9ICFvvGAQ1XyavFIz/xjYfTiiBBJT+e++K+iI99/yDyOmFPKevGDPJIRGXscXTwj
WnaLccSJ/YNFVJXx2Q79bsJmVhsvWpWjosBYZAcu+m/1RGmgU4jBKqQTVz6vo5Ia7ydMzfIDvqi7
XglPMmEAM3H01KEKuEQ9jeJDmon0VMPYuMAr2ziAbQrc/No9WjjHo3ewo9umMgAb1F/mQA6jtl3Y
0x9ipkmBUnoMl5KI+ccLVext9lnQjzWGRsFGxOc2xFgpwbqSSzZ/xU0XhECJJNzbaaACNB80a2TC
cNtih1KeMl3YeqFr7/TEj+TojrjUz6DoN0VwppDpWtlHtFdBnWTnAJB0Nw6csZLDXnIdZhbk6Ard
lvPYxTxq0F9hib9fcSdX16nCbJthZpkDO9dSU6St1OgugRMhSZ+1fyEIpuTZgyvKCEcIBwOOkx5k
aJdwdvfivlMzMs+y6l+ToEpHhOExSnLkXPG05IqEJKYQ7qSdNbfcUtskv4DqteOKgQO2Z7AoS3mD
S05DysuVcPgTZmTX/Hd7loCH/0FO1ed5wpoU7kQO1Z0XIw4PLNo1rlIe1d1o6bUse1TjYTdGyE9I
WO9WxrmCNAb5TSWDR5XX3hfIgAPJrTARRUkH8lss4oc9YHEiTihgBj5PZFdTu7Fe4kAo3/XmO4zK
glyfzt93MZQ28EuA2QPKquHqxtAxJ3t4LNmHOV1VBeN3fQ/G/MnSYaml6feOPcspMsQdVvyJYlME
g6T6+VNdoiRW78Her/z1uws5KATts/bTsLGf3JBcbhW2YMnR8GInqbXGrSo1mSDdtawcHSa9kBOq
bZmDJPEUxcU6i3BYyNCr6L1cgkr6fbwVw28IrMGjIW5d1pp+H66nKk64jVtmFJGHv2hbW51o49R8
NuD0po3xyPZt0NuOjStl2XJzzLxf7MeoFXkhoiFbP3Qnp02zx4f64gL6lby3UyiCe+h923cIB9sh
5r8+V+791dkYmWabiYxhO5H7IAkDbBP61t6Q2xXO5U2rLBfFFtqnhrA8m0ELFQnmH8BC1Hyz8O7y
mWxavIwlZSUS224dMuUH4r62jUyVGV0gyXB5yEZs+TD0HZwViNnulUuVUdAeTYottV0uYi/7lQcn
OWAU47qJxu3h2Qq/L+xyiHHWOTPubLzYJzcfBwAYDQj5kHYAoajr9OJh7GNrlLnTrNA5tyG1BtmW
X7YSRNvB09CX14kb3OxaE44UbATTR/j3dpiU6xOuHjFim5Ob87pjLoktHJFimlIE7Zm/6ANQ8/Ze
8ZiKuXwhyi7b8GXCWBwL6HwoEFVXvBxTTdv1wFL1LTdNDJL7Bn687BB2EyUeJVzYtHp0kgJ1VbmJ
zdiityNTDzlSHlglKo7NaH9MU07MbiV3Xl+Y9K0j32abUEm1fjApf3nVuR12tDQalsVmefwLNnDj
TmwKYQlywONQbuewFUFGdUvGX9pht9RDEEAZzCtWf6sbk8YHppc63REuQ+OAlcrT2d50a4j54ZMW
gSye7Faf37mQqpMOX0uHyQ1Qkmpti8nvREKqUZWjkoZwfdRNZI7Bk9u7E1STZ9qGmO57uph4OdMn
hcvDIWtKLo/TVOCTmwGG+WfAXIDiZoJKcsJP2dX58/Gz1DWP6T+iNoh2GzsoR2I5zJL4MxyATESe
MR1th2q8W57Mopg4QPFcq9w3aDOnU7P9bFW9wmVBrIirCAa836OfavwfE38RicnnQrea0V8l6Pcs
qzyNXQ0CeoeHeybLIRChd7nJ93AOgBmOQdsMlr9CEcgMp18uJjN4NnIpZgiZHSscsvJcWgFk+dVP
xfxtR5stI3syFllxy3EhSbv9xo/QroINSLGhHZJOeMCazZbv2m7doXOSyjhQYS+0jzvYXKb5yuUt
hV8vIqi/upYnd5DYv3EZg29LQsq3tHlWsZ+cEttlc+iZVgoCW3d/rXx+S64Tc6LDXc4wC0bS8qWV
RL36QrtyTpSwDGppOrzxMJLTDCWJg59XxWnH3PxymJYav0YTtRJwvI0Hmhbhh5n+BllWVwOCfLXD
51thhV6It57Gh17vPlI35PX2zzqdIvWCxteJJ3WWNxEe6sXi6CO1/SRDWeqWDs2iOhxJb9hq/o6+
EwGc+RvnfV+YSsFo1xWysipBoHNWuU6e7uXpInnnfj4yyYlpoJOiM2fkgKAdNePaiakmCEheierJ
w/eVJK4oefznK2AKd7im0lHLvSXdfj+lwW1xkHkIRPF2kjyYD6IJiZNcU9WxKp1dQEmlJmRJozPD
aqeKRZP4JEQHN5BxRAXof+q8FOPlAjXFNInMWZP1z3kY70BXWcdVEusgJgNp3ZRpuyIkoE/cMWu0
kDArmMjNihHAF65ux/oVhlf2KRG6bDkvc40W0mvKYQ+vTayrt9mxn3jrYpvoghbcdCGQTIPijDEF
8jDuR1WXBNMWOV26xiXhtLZ7gnXiDuJGMIpN3njy4cpg20mZGxhJN9vHqyfvgwE9Ci83IZoRHcgD
nnR6WUreWw8ije1CO2Z/imBPkf2N5qvegE4jyVR71c6lhYoqyDGwblNLztDg6Xew6TqVcViawHfM
FVFhG0fjHcVBMjHf8mCamAZYjn6hH3IvtykUGRnlOYscdfgl3McV+73xpkrxXULAuBmxgx4vdFiY
WSwHR3Zq5zg6UCFTyzVSdYsI+/VqQ2LOZYzZ/PQ7ce3s6XgS/6C26rB34sZ+Cq0T19pUQE+0rBK7
W91X/pAp/6HHKsxrjP7aMacfdueDtLqKmO8vmFY3uIayC/Iq6lzLtyoTw4N+Y16SFSOwyuznNYyD
Ouc9NEMEI8/YZlk+mZhIznArIWx6UhJXWqvVY4DSmoCG8mbAfYGULXHGF+zTeJJ0wW4MCdEmPjX7
FTShES0xVG/4/qcirmb6jwbPkZ3NXPM6RqCF/Dk9lyyLbJ/m4+uLLn3imw2rrcxCxeCyUSZ+y+33
v0H58/7We5uTu3tSEsrTgBaZv+FCtJQ69kRjsDl9QZEnR9NFyD8HgLb7e9d6enjDIQIKqW0bua2Q
WN9ZIqQG7LEYXKqS8coS1gqvb+t0UEYWyBYksObK09Ki845l5zu0RkK1al3XUuOT7MZwcAaE+q33
mrmmhquidRl+n/lGM0AxbEdiJODzZO41WQu3uOSxM8W2ijtOGOvYHMs+uAUhHdRO5ed2w7PZ1F5Y
EguPafnIJwcT39gFC9/ZUObc0bPezS+HmFG1xnDbtrq1EB1jrumq+imlYGXk5idGcT3kARibPrqE
7xGUmJOlGh4yd68O1zgBQhOZlgvc9QQjqN9/HUJNzVWy7w7xSrncJTnhtJdaPJi37nyBq2kb0AG7
akxrkQJ9zu+s2ALDgGDXRM89xLSVTJiDL5VVNfpQJXGWEDFZ5e8lWi2BCTcZWMXsXIIR9lS2H/qr
99ms2FnVDLEgArMcDtZlthmTQG1+sguLfBfbpt2HMKyMYwP716QV2GeLHqrvrzprt7fCz5fJbv7A
KC8mVW7BuOnDQNNpq/yA7eI3cTg9aHjeNcqvw6xxkh3tT4JCU+O94/p08fIntnzRIUpdD3bl1df4
NFWLzmLi5MDcp3KfSZHL9MRUodW2FAqbTUmVsFg+Z7hMgr3CP3HCPD0BpPy+XCKvP27QplLRYsfJ
Q2diR9OCJSy7MF6aSpXWa8ifw5RAHx9uW8sK13M99Vlr/QUzlFB+vsLDxy5bTHvU/4EsDyfFqimX
MhVxo1hjsSgYspTSMDcf0PsXxgUMF8Y2L058ITh2ahLnBAsp1OSQnlr7IflfB2rnARjOKd+TyOTT
alnCtcbnq1eDFigpQyIVb1qooV5S+gwHK0J2kE3q+LwW9fogifP9puJ+DeUQPS2czK4D5QmmGG07
OPdJWbSxN0aoDjcS8cxPEAWJrU3W9J1Uv4Jzs3HfsL7y/MFLaoyk7N6FnE2lApLtHZbCYOVYDzn+
UfKATYLO/tmCuz64B5Ixrh5muCbbyGzVRh2JojNKXdPXjrCRkJfE/WDLWO/G99hmLHKkR2PPmNbs
y0TfYmA3EOua1QDEdVx64cb/oLa94PqwaS8Lt8h/NzDMbWko+yWvVTwvfQtP7fN6yhotJlwrPqBy
ngBtT6qtj0Cl6GiACZLjcdgeFZBaL5K8TXIT+yyytSbiRXmp/I0QT4PhuO09YshJmmJTo1D+ZJTo
vKdiKRACkPb9xL25eq+MYu9wB3ctgLVjQKOMicKkpriLi98K3P+pZjrzhP9/bt7kvFy5omZwqx6+
ngEYTNMElMsopmj+3FXH0gAeAZrEPBe553q/suOpTuBUn4jhqS7x/tB+Au2LZlm/mgL0DEJrUWJq
UTAQGy8C2c61wL0dgqKOD22WMLnKUoUx41ztc0qLK4NIbV+NS/ceo/BDBokA+vCXyDvW4EElFJMy
ZzBzNOVQ6RONEi3HH/Qi5zTTYw5Y1JvGpxFuhfpoYTN0Eb8jmWek7arEaSIpDNb5upNQccxv+d3O
6N5ppjF9B3e34Kqx4URmdzqI5zKJ58UzprwIE1pcVQvtKYZbpRIxMi2ARYYfNdWOfX9Ytlx1yUc3
aWrBwC04xANJ+F44/MWu42B86V5YaFqxxUdrlgezHp6c+B38dzG4G5tgtifzi43uKl49j4LNPCZ7
q9alSW6lZXX5HtDhNz+H5rG0zLtOmHIoDoPbGtOi6EETWtVC8VAtmC46/Z7qxdyUw0pyg516UhZR
KmExzoHC86hSzJK9FQwu8pqfNFzzEZj2iv6ASwgj+aDjaMDAFbti9M8UAUDSD+NYVNVf96azYUGO
NHHGm7mVRiy2rQ82IQCb0uLHPmx/LW3yDfqjyYaLL6xrnGIUqQoOKoX9RKV1oGhKNQRKlUZIQlQY
zMHQ/JQHNyksrF3S1eZ/V5LkkVDBZzSwhrqfnHGRpj2frgTWnsoOVPiuIRoKfEBjEcXgqWVkMMwF
gQwLg/zurvWmneuIkXafbbk8PJiqTPe5KmKASWK0fcedo1O7T6GsI/tSBNLZTKh1JwZ/5e6nQNNv
ub9XPggZgTdlgwZWk0chOhSzaCXe6CiktmsG8eJxLMOdSURAgbS314+v/A9rHOlI9i3IjT4L/v6V
WPF0vXiGQ+Dp6hAQa9pBJxe0BLPYR7LA88l5lOt4p1K8dkaWlJ3BH5al+IY7Q8In25nSwvSnG5jj
ffRdyOrAkRxgLb6YnLFE6fvyKFaJxycKEWa0SGfQk8ZRQz+swZ0bp+IAj2QQvOHWNSJ0VSoRhQi3
OGWko7DnXcSp2E4nM3zWway6HTVzMcYCOC91+mVnvlk9MEcazc1vcu4P8mQYl854BjvRfZSgNZj/
CfsDBpxahsee25inPsBrsoREg+B/V6Xsv16+coq8+6kXNYNR3F2WrvOvM4uCP5HpuznyjD3l8bf9
NQuaC72Aox5ppe3YffXSeqjH+fEFsAHTBswvs5kBCy5mZ8y+KBKgAr8ISvA1g86ovnAoPCIOb/6Z
KtLTHI/SKOoHg/YVXx4KNGb8PLO721N5AtuZe9svsC4hIsBYruQpjtePNMnZ3lJtURyIyToLtHCn
VQfa2EXfu9cjwuQRL04gtKJc/O8OtlBWowWsS1XGjSvTV3Frvy0UUMuukib9L7TP09y+09ToFLj4
yO2ADaMvbp470NQGf7PAoXj7wsxw3qMVFd8lTkpjlpAn3NazW30lVjJO/iUfuLuOlpguO3vJXuA7
AnRFS1GCcls1736SrIp7FENi0b59rQCD1kJrAtHgHY8XggHvWyVL1CFVJPvZI+3jR2wOi3BlXD7g
mYWh9DXnp0ofS3iB2MRXSRqlcyEPJmKR0J4X4YRKwGLK4jTmuvBwyGsVuzPVO8G3GBCnoS6Ho6vf
EdksgB7aJbNtopDrXQWR5BsiigBKNU8Ot+go7AxX/bnfdNNc3qefkUpIaDe6pUsMILCroib9S8yX
sbUsFV4PYD9UdnDlAUgjHn2CcQ4R/2rusGXCzLKLlDpB+dpYV2wHZeUMHGHBeJ/N5pIx9JF3vFlL
zCtXV/NAivTqFS7SkU1m7mVy/ttf6ZVBSdcm5hL7z9/9cQeATUz83nm16ljJ8IUFftbG9TpQe0N7
LYEFNVjwNHC+Qjf2nFxoGQZSyGwBQ7RrK1Kn8+4il4KvmGrUs0dnbmnaZhdqm1r+A9l6X/izhWFI
AOF+Hs6IHfj1+OVJH8aa3N0PwkDRMrCgoZoE8jyO5uG+HS0kLaw31NZ5QCtq9vSZ5l0aJNh1PXZd
UYhA4SsO7DEiebEvM93GQH6L+/XZiCFTXfdHX48SkOf+PM2wvo4SNftp0YVroYTQpdz5HC77YBjp
yeFLg+AFJ3zPFtlcr0YI3KLVXVhLdtE0mYa/TB+hcO84+0Ye5eDc3BcXfLIa0Qh2ZWM5POUWayEn
ym0kDeWp4eYaO066Enw1kAJQp0fGfdlE2Tn9Eziixc/PMV7EIxKz6dvy4MY0OaNTCJuXNgOfbV5J
5DM7WKPNiOwRSmOoFtK1yc6JDpF5FIcc+rJV68pCQakGCAOwiWdynmn1jFsfMVK+PHuO4bE0atUB
dHwjM7rFH6f0KVy57IK7B54N20z6MHqX3Pz4eHViKyd/sChJ8yMhQ+H+gBy/Ua8jh3ySCUtVsHvC
VCb/Jwva5DfXloc6Gwn7RfwGa1GvPRjVi+A3MeC7hDVpKOWE9K55+1XrXaU30Yf6HgvCMRjtpEyb
JUGvGw66RfBD1YF8G+Bbi1N7/UCilcQCMKhMphNIUSA1gITuu1Ma2JvqhmTQPVukkkXRTVrepMiO
QRmfNZMg8wmKXanVU5F+/VoMwoIhbgLzP0+tX0N2eofPbILLGtinFcUm9BmTIckwIRScik++wvi0
m91uJhwAbQWeW8L3/Qdu3OrrWEMtKnnkFTbBep/4gM0na88kPA/eq7izgQbj1jAOlEY0vDyHuZnL
Bmkw/IDsHSKTcF7VK1rd8o8BDAg3sqtj0eCcCYP/xAY64EzvicpJNqkrrnNk2jGoZ3wS8Z1gm7LA
wa+5r722JiIIrmJYwHmWPB9yvEu5hUsWhn7mbK1IZW/8YbWm6lcVlVN1fe/RZpoRzRjmYcDSSaGy
1sYpY4Hxuly/U989HsqF9JQBHkEfgEIK2lT+yMX0xdqI176gx12r2i0mUYz6hLaGatiH4Atwdo6q
3booz4iuZHg1oFciYp/phZbSHyFPD9HwBz1TaAtfyNSRLwepi6+Z3uZrkyRQpqQLDuXbvM97Bd6a
/NuZn1pg0MYL5lLmlFWfrCikjHsAMbLAYC+EPbnFdgn7zMQHLOLLqXLUws25686IeI4mu/LCEPuJ
Dt5HCmcPQWZ9PpJoShf0bJNrLr/mB2MMIzsWFXZszXOCdx2alCecES0OJQ4CPuOi9kZ6siXpO4Gx
Kk6jDwbJvNbts+br7LeoDI+usMDYIclaznchSnruxbCFO8ks+vGu6BpK72390rzI61bHYV+bjEvy
NiYJ6MeGBu7OvIldgqUcl0u2o9yk/AhasytX2T/RutCYfQD0qLOt8uYe82adloFJRDdvtWv1r9t/
G34UBADxxfZWCA9W0KuVRhuJXYOMvYCCOvfawZB/szwdOi795lRqoJ5dwZZBIdqpOB+SLfyhUL3d
Ydz/CKXBqnJ7urBnj9d58qfQXNneogAoFQ/UHB1d1+F4BuI0gtWQgawbrjDheE3LcVqgxIrSydyd
3VyzrNXC3cOUSSz6ZzlM6PJe2ABcDxtTrBE5+AUD9TpqF912j799cuKyx/XPPvhiKHWA8d0pXxTl
Hi3bMe38nYLLzi28bcMfX/7eoVqRIqO6/fMazXHq/xbQ7DVkq/Ym5a+G8vBk/krIu2mBXzxKVVKL
Um52lx/O4ARfkhGt+zyum71pFqsasi0haFCnrJxDHRaZ0BEIwb6Oc7CLkXs6dVARbm3DHG5NYRt3
iHgU8H3RaU5pWeG/pb1OcMVx0hKSoItG/SN1Rq38DT5Al1y/RXL5pGq6Rhg2KN2px+BqeX9zlZVZ
ewOUHRqlUo7PJNFTYctl8TMNYwUeHpukBBy2E2tKh6//1hk7X+IJ/XoPpZWSWWvid8DqOWMv0Foe
+28HUJjbWiZayiP8zBMH4ExUArihZeqL1Wvn/2ylnkNua7kImbfS5/IPP5wrhICsVzDpySTxMUNl
/aT35Lg99ipG9s6RupT0yXpotrVLqH61Wjz5P2xjtW/TORA1MJivfHvnFR4Jd+cIw9yBIwXdDOez
Pc368XU9jhSGGnT+K1qpnOFVOnaxAyMBqE9Mc89SF5EfnI54WD+Tvw+zrbRBukCZ1Lox53ZHYsWd
M4HIniw2hrgAi/OZeHE5uI2nkdZwyifOe6EtlvtMATOUnfvgOfl7bGW2daGFlt8ueZa5BEFNInzA
9xPJ5qyOsyjRmDySz3x0qPz9Jg9pzluIkC23pW1iVgHWLIKDJSmaSJSTTmL272ZBqqdKrT8n0ZFx
f3Wo7ueJQKnjbaZXK9K6znnpMs0dHKbZlKzBkz2YaghihSh4sFnAo3Yi4/paEugRXnfQubeeQkdf
txxe/7W3DkxGiiEeubA8ZiNfTFxas5Iy1GtFdKgUd8BwiPYYqcSN4mf6EcvEG3L20lzOsj2K+pBO
oIRWsTDC//HgEnPYS1+LSBu9rfmyKlT3ReyNEp0Rg0TKjVfDgEY9+t7Vm8x2JBIAW7DyQWoFdlri
aWow0/jiyaQkA23PPabGlQhoj/9OERhnJv1VEcd9IMY9kQtLomRgRf4Pgrglepo/51c3DHD/QjkO
Tii589x6hpDPFIr59X+I0LexxU+xLWnJ8PX4yMHCQalK0e/scajbsOSFgdj4TydtHR/hkiRMStxt
1MII8DTDbOtlnWgvRKddPjMe9zLwk5pSI1XzPz6qz/K7cMdaq+tQVtNt0IZniyXp+bKdDpazJsgw
m0tctV5yEoXGuF7+oZzf664Yxxbp1Nd+/ILTyMEfWDT8U375ysA9znkmrBTovFHgm00kn+lZGj+x
jg1vKSHUQ/vKNiR8ex7GZGIXbjpONVDsNfGIrVJ0EeT3PfXM3gJLBJpTXI1e00hqE6Z1gg/dXYSU
Ien+0ApoaMuFG40Ib7SYpuy2dI8lQwvYN0fV3cPWXnAV5CNARDhy9jEMqXvxX9kCEFzRAwItEp1e
S3zqV5zIiRyHn21ncMrj2cSpPaXetNlWvpIQ+tmDognsd9/dQ+w5DRdYyPFEcGEvcolw9mSeKwNS
h2JkIsmZPq+sjQ9r3ohigUAoP3a21w1K3yzg+ogApBQjszoEXUIV/RLgmTZs3VEySfGkNE5y/O55
7yBChCVELtPekGPWE4jO9n3U8/g4gxrzWBgIjGygNfjwZR9F+d4oY4d6XjemWRUWHg96bbk+23yj
BRjjvdMRPbfmdlvlpb7BaVuhWbvgTUfz2ov36u/JJNR0hkkapX+gPc4ObA4QQLUzVBfveH9ZFex2
kwKGQo3C0RRelY2DrjICVhYAwBecopP+YynUETPYmseSzp+ek8LW2/H5AyX+LbsIciJ+ukuUkOdl
8fnNONPVyaRH1RnDZHt/syzfWEV6oA7dW9JlQyp/5zqnnKX9IRXPjXrjZZNPDBFg4kEwR2YBeTYf
Tcn9aa1raeW6yoiE1dbHS1aVjDWv/BmrFgx+v7FBCifDkRtE1yHDn5Q9gy+856OMxft7yzqZGEg9
lLhwV3OtMd7qQ1RJYxa48qUJ6UodntimeroaX6HFXF9nvfHZgydJwTRss4oapGXCj4oXuUjH/VsH
DIgAkNX2mJO5uhhI5Sdg16jKutVno5Pja70fUf2ViaYzm0uhGjWLrBM5GNeeoCjV0xuq9kpVVXZ4
KGikSZhpyDbplgjQj3fgsLKt5MKq6G+Af2l2InIURg/0x7Fu0SxrG746YACv7Xy4ODwMMTzTRlwG
VAuDHaLBURkp+fJ03eWfYrUZhl6KaeUmnZdWa2D010y9+vbH7iPag4w/zc+6CzBuk4ye8CzE2y61
C2f4wtXudMf/+pTW6zZFGTZ4+RFFgegvbWPEIqUABccXEnfnqqXWvtOL07kkZNW+QkexjGGFf2HK
0RJO1N7K8ACy+i/uqH7ooMISKepgQ5JNT8B5yAracg+XMltBj2XtPYR/F0lCaplhe0GglnqRjUXi
GHoCulADghLEi3AZY4Olm1W1RCnFF19fDL/iMepB2UqqKdNrRbSRJqJWp9f8XODUIaUDIG6cm9iQ
bgLoVarq+q/vHLZcDlRNw1VytB1yTX8ZJwgZlVjIzpVznBkGnIz2KhRIqsLEB4Y8pJoxu8gq59m3
OkWC+DN38Jf7+Rpsoejs6FU8YaW0hVD7aNVOt0MbR/IEeMOKoUZI8Dhqwnmr/UwwXrXSB6NZQ3Nr
uuQlNz+gfhSks4Y67nL9pylfbjZmaa85vZrraafBtXaH5JTyPCCyHPoDGi0YCYI4JnxsucC1y853
jEDYr0ERkBHaVB6wUuG9rekq80cfce9lZk2TReVb5eM97YB/zS6OQUooet+HfsmjlPYwxJAjAAt8
rnqs+NtYbuPEDVjkb/OxmbQbdn+aS2xMtitZo242GAGtC2vcjgp3hPH/nYS8LNmpd5F36jen6LJW
EPOTV0NRrDcyH6NfwRzaBQlBOXg6/+ppU0gLvS7ksPjf6bnb2UqsWZHGYRY5q8WMblbRpbNxe88I
MS60a6T3eGANx8O20nP7sn7achYR/8wAgX6lnEriL83m5QRzWqsBDA95U1ogyfRFjcxff/tT/f9I
hWcD4xXzkAP3kBKXOms9tM5zeDO75vJRsjZotLKvIR+FHntHe4zqnJHFnGJ86iQ6GqJCUQSqMXVI
kQXUNrmxl5yMzM+FVnLEDEEcE7Y9xi2xFsImcsdtGicy6JB7vK0mhw/EkiBKjYfyzxYTLbx46sss
Lkr8zbgsp+g45CEDbBOoM/Bl2AeK4UcdjJmLzNTxqylx
`protect end_protected


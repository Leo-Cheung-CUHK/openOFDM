

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mPx7gcQWvUiXAIlptcS0ga/HwxoglSwZPSAvh1Lja87QFX6EO1tvAtW3BEg2Vp3HivYkp2SQvnX/
wf5IwSVugg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
u4kYBbKWjVmoqUxGQIVLXWFveYVGjS8KXANLcMWW+aY7ihS2tZxXnk3ijjHseANEw/GD5bURIhkJ
wHNHgMafDMxk4PoyqdLtqxy3iP9j1MeEpH9OoyR56v6qcdr3P1DRazxtJ2ZaXaFvkJSsMWBDAVQb
EAvsPUwG/uWyf8K9wIc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rcZYcqDcW2nDRCEfMQVN/Fk1OfFW875uC6ei3MlaCqhRnkhzT3xNk2eZbf+e+AP9hFcz4gOesi0n
ZoKrSwPNM4QWWQUwJVjaO8mmjT0knl5bHqmrP5PtUa8Ymb8JvpM2TW4eZK2Uprb6QEt4vqyh7TOP
vhbgM0gvOVsfurZr85pM+sdQTj4K2NKqCt95to1VCJH/hGDMuK47cP1uzcMQplSPzUkPukYqc5u1
65JQDYRjOTqX4AbM+yyfDWw+pb5SzcyHehsXCJH0dv97fYVSVVRFHixh5JYVGcKStfxKGzXXKQhy
T709LnMhsbkT9A3rMvt5la92JFzNANaCQ4q3CQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g2wR7vfvAF0uDhoyjP4PFNh7OLccqK1GsJSoBjOisux//jU2ZxVmLxA1YJAl8lw4jONkagbbp+bD
DeKzRS2ZhyX8p2HqWKvZmJlJpU91NNfgEUeagxdfB5g/ozhVOyy8QGxIiIMb6WrYXhYmtrxZNloB
n9TcaPYLMM7L3bin109TK04mlunQYKeEo5HzUOQf5KJ/sqzhE+gaF5v9vGZc+iE5PyzEZmTRiFkB
DIKvHD3bWL6nrSBv4kJGEMbH66PqN/cEKc8g6Vp6Q1KwRoVPABYLyvfgScY5ycPGYtzU/pyN140X
1iUlGE8ESrGXM/xbywed16jF2DlyQ3LUN34B7Q==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QhX3pm1tgaFGdr2rg1UW3M/brT66TBguCgts2VP6sg+tkLIps/ZujQpBhLiiUBuZpY7LYUF6Ttcq
FSLxzJjaRAKHhwz8QfNP1LvV8beGlrmElSBg4WQ1vh7an1NBCIV9vJQ12Jb8lKj8kV4h1jtFHmSH
K9jxpumxvGxg8OkyiZFRMV7wxy5Vgb+iLbXznLPN1sO5bxy9oPYkEE6q3W2XOv/+6RQT7jrgsgij
Ryn6WmRS1JEb//SBh2n6mIErQ3VXcu4P5ctFXtDE8hGFBRyM1uhm92HrFtwOxkQS4cyQYHYO9iFQ
G1fTJnB7JigyDvGKfvwHOOMtLjFExIGVquRFGA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qAV9ax+P5GkwGl6RgX4q3QljQNwnp3qvuISp2RvaZBQjaPrHqbafHxa35DhyBrgca2jSUOtBUvJv
KqsgFgfZn9V1QbQ0RhuZfQ0A9iTYX/dan3GdDTQqO9dUx+ctLSRf+zGO6pzzUXyKS+BdkWX0VK7T
nlxUO8Eglcs41Aow9Bc=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ersNAxW2yyOqkd9D0cu/x1eK3Xnna2vZ+/lR7+n72DdUl9LOW14owvbVJOgkJzjQh9R7373dUheU
TJqG2Bj8ZCYCqOfOaa5QxsPGyvnovZkK5DNfXSZyOo52a3W+1/UREYKNJQXMoI7o0buPSR9vjzfT
VP6gcUF2vI61llqn4hGlzHjw/Hxc7DZ2qNeQE9EkKFRPZZAg3UFlr5FCYYM50n1xKXOPz1GiYZ1m
fQ6rbSyWQGBnCD37asaeCyMWyupLe9e2+ig34/lXawgR9PYogJ8Af3Xu1/jMBPPEu+9fRFMGdl/y
WGXnDPxDcFs1W3SQMXNmK4XHz49a94IR6/sTyg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 133280)
`protect data_block
rKehyzcOdEOTzVmMDDLJUF55wzvcVFMjmV6uh7xRiipjb5oEuTK/QXYUZYkL3yVWgnHxXrPSobza
YzJOk4epGQ9Ha9pkdf7TPb2qocZpqlpX51Z+6NHC9X+onZDa12f8OEkircdgiBodWi24vbX5BICb
RjeikasVLanivHKgeDbYJpC5JMY+euNkoRKCWMuF8zcN3ri9vUIAa/fBPl3dEhAuSxrGWRGO9Ckq
8Fp7xLKwj2VNnOJDpLRVwngT42FL+eikuD/WUDIhL3ENA+mY6d4lWcmv3LPCOoq11qbo/jJ16Zje
4Qnyx0O/DAHiI/uJH5f3xCtzt4j78fBb+PqA5gD5fkjU+HEldB1wHnXvbw5bFIdLtCvItOZD0QBU
uBZQirN3cGDl9TB/84DgQJG653kWtdJNrmEYxLvh7DstCjij2uHdVAGQYw5I9wp4rcV4md76idZG
O0cXcdDEVq+Z3WffdU4MViXvJTv1YNizoGKraRVHaYlDgI/KNj0gIPZ+FuqN1eZJsiDVqhN8d4Gi
k/uwauUT6Lo5Psmcvdt3ZR9R/M91j8YOqSSJnwKeAizXxQT+qMDocYDGerQca4boQ9i6Y9szWUh1
ACP1W4XMWkfigdyYhoYX8xTKnrz3n09ikctUB7nLeuoo2cxiLq2Qxq0U4QSb0Es0s6ZLcBM7kMMg
E7R/NI49UYntIDAiGor1vgAnHzC8+HGQotOyAF4jD8juxG9uqxb6dKLS3NH3Yv+IMYR+XuAtRcvR
Hidq4mXtxto8zkEOKVH70+W/NZwL2AKlywVUFwrvvhQY3IDyWfdk62nE6p0BtRozQwpo0z58Qa+I
0Zw/biAtxPefgj6sw41rdM+KTGVdhV+GqyuxqW5gKDXHKIdIgZUIjkM87pf19D7gRgNXvNGKxgZt
OGPhqjrdTeiOBcBDNd+NRei25dD/A21J4+7nNsA9aHX8OSw+3iYJroCIa9LnZsR5RHwNiu8445mo
uqV8FME/u9IF5FHfxCGsDcn6oBb418Bp+KyeOyJspFFImAE5lS4OibisULdnv3JleOTNTa/0HxNR
edAyDV28y7tpnh0bE5YGMguiuX2txI9IfiBPuwO7fagvGg0NBeJOTCQYF7ngBmFjpL/XSPHITK9m
oR4x7TZAeO9bel3TzIUwxl/9yu0MLlvUBGp39FR+RfQcjoQX8rmYKRhO6Ybxiw99AiEelkMH2mHS
GxoIt0FERv1eMETr4KBp2mi2T7bwF7m/J6me4o7Rb7Yir6n8fXkxac/xNkj9Yi3siIqwJKEpbRgP
DqfLvxTxjELO9SiZ5D2O+6YsaOdW5pQI7tQrF2QyADerVVQfJU7hFHiWR+wyNZ8P0DAX3q98m5K4
t+Xc9QAexJVve/RiVf2NCOxSMX+c6LbWTc7R0H0P7flyoC1KHHsZn5jmquawa6z/hNHt9wYyNmx0
poph3Tbo795MzVlryOoaIdiOM14YGOm3Ihzdcn0/1/ce/FsYYWDsAYOyLqqRHu4Egt+wgppI21sT
Vkv3t9n4S1mn+ETWDhqetaWHwrjpsdvrrtQKz3VyGAWTMMZ7xbm+TODi1qsjqXMSYYUnGdxwuicn
ZL/CPIznKPkSY6o0QddQgfQ0C5EZSnoEoRHCgYpnJUweYohVM54k5KHO+9m1rNNGW0iB2pmkw2M9
Yc+uzxXwNc5wQRijab2BJEJpMfDnztB+ojvPylxi0jIDcce8Bw263Dz4JV6+5mK0SaA6WOpnYR0w
pX7XE33fLYowSFZ3aClTQ9gU0YLE9zZYsQE8kb9MXbIR7YOAv518U5+Vj4oY8QVQLES4BSdbJqtM
5cTTDlBNZV7MM/3OT8QQYaS058qy7wE0017mPt6Lhph2B1ab8T109WOBWUSDXpl54lizXKmTnfTc
uX7To7E4oHKLTj4WSW1Qc/CkzRF+1AP+RE8l5X87cPXUMPC/u8OxnvwrM+RDvMLcVAJPNQ9nQdyq
HHR0WEHq4m6eSwr6FDTR6HHOuIu9AXf7DlUftR/FSAjSee4bCjlN6Gowld8g3B+goVE1YuSWUm0e
XogjbaoioAcaih+X6VKotmhg9F3TfgHLNpJjRxxrvOAGl/ucFNNv6a0OKm5dlqG7K7jRcVKPJwld
bN1d5BLGUWQltdZh9F9XGLH5BLymz0vZrnO/DrU5uzaB4axLnqnrMuWqCW702dkg/3xHIaH46uIB
nt5gwR3pCW8MT8Cc48WlW8iUJXZfXU5LuYLH39fgZDaf4x93HQ4ghrOq/FftQGtbfY4IGRVkIBxT
lAqnxbe3cL6l5IZ3EQVdn4cn16/zufVWEac78KnzSd8Tl24Xhp1dIIz+YUhN1gOthfCdEsHXUe4D
0yoZ5jwcP4RUlVYAZ4vRrlHJuJF3SNz1ZNZWuOUflo0gHeassDGS1Z/pRIaXQ6ERONfcWCXGVtld
u3uUAC8VLeQFEksBNwRHv4t+kRZMEfUhfJobZiZTnmxI/lW7eB2K2PPMU1BhMAFpXrHQrITA5SjA
l9PQkfYkyqIgdDqh6hAtomTVO/xmHv7n/ECZ7DRmCG6zLhKWJGBVqWsS2ZtlE88wEEDhfWDjElM1
euvwYdrja3hM3eHunPBORp9QVvQNAf9HNGhqzhrcGt3jdbAshJFadwyw5gGCZUoAu8fMGXkct3Mo
oEXZUq24yqEKM6s7m/iObvjX10jMy1Jkovq0d1mhNldPJDxFko+ce7tmbti3pyBJTsHprpHlbkvS
K8g3LzsjNGj3igCNNnPO2NxO2rCEPB5PQ7/35CxKlh+xB3XL8olpxJQUNWmncGcTraAoQADxY7Pn
AC1ZtYhCZN+jVoTN3PttmsuLGZaYK3BdPA4TNdaAbQoYGmUjGykTz+n89TQsuV84tXauSeVpzzuz
lYcFjNnuOwvWNJU3hdMlq6+Ak2gnIMrQp8LdyP5j8AVcqLZw/CreLE5QqFDzcNOaZdi24hqMs2OZ
cBsdblIoUF2sSAFl9H1xTgEWTiu5tBBZxUoxee3yeykqjXNRQkq4F4dH3ICuItYH5geHpCh+97tV
mugpB3GdeBQrgHRspeF4WJv6gwwh5zyAOcsGR0M1rlWwCLWAfrzT/mNgW1yZChR1ZWmn8/NSsIGv
euDeoLYSVKYlN0UlLQDT3P1BSmYH0qWcP6/EXOIQvqlbMo+axzKRsCxwf+HERb2t2oa/3amb6Hpz
zeecJIBERUCH00DtIDGDuRQq9aY6cje+7t2WJT6pu6TUieokGyz51o03gDs8qk22/qTtJemjyD/g
jN2fbmp9u0p/Q38oKgWk+8pHXqYDVLULZSqsv+uoviVLn8WvmpagBK/NEoZdryoxvlojAhe2vEuB
IuJLaGhWcYejwERlPbYNRAYVXgZsRA8T7cBI+W7fFJzhl54oYZnDMM45Ik1VucXVwBX2Ef3jHbng
U53cFJO+esErv6ybkzInxQ72WB7QkTE6SDqoI01q0UslwTJUnC2zXd5civTmQ1kNk9CfwkWeP1jc
TuRzk3O3G7IRY5OOdP3rZfCEIeFzNIPK9Pwhm8srib769U5HswX0e4ppdHpX1AdkSR+azawNMxeG
T97g9sxssuF+4ixQQvxmyT3xPruZHrTfpgUr+X2ZmvyG1EH53Uzyko93b7prMqTPP7+AyVmFreov
shLs+uG4MFitvWdgRK7252EYXLJZPL8kRPEh74eZRIijLInyW4w5EhTWv1ARAXP8Nc78ytMimiYE
0bFVFwlWsCMDvHDjNdjoRYpjSy2aMx9DI4g9WItOYXTxurM+V0s1UvjmGEF/Rqsp0VWrGCaP9oKx
ZN5Gj6qvRZJSdPjy+Iu4yWhXVjHPd/zbWpoSITJO1Q0RCNzJhVQDnpmhlDT3gaKwIAeRS5iO50Ij
vEL3kBno1qAr5akU28xY0lA/J8NrtmJNeCCVQP/8zLuGSu1oXx88HSf4hSDHAEAPw8ulUwf5RYFl
OFIU3SAcPZhxRJJsGYtozAYw6ow9UlTA+RPajqUlNv4KYzDm3kacCQnUwXMTph8g2n4cUzjnPRlg
aGJX9I4wyYnNxYHDj6P+pbd/hXVnW1D2chml2Y9FAO0r6PTaUWAXXcQ7fpzXPIlG8MT6q1cXR3uo
1piql/O7OCONMWwhvZrvDGXDZGFPsHQPO6UBNqxICGX2+F2SMOXGVFNzMSsM53LSTuo71Xfd690h
9WmXrSPit3C2pssPvzIq65FBKkEYtzWx53UzUXmkaNIbPG4FLunXIKuTkzrbXLpvxD30fYhSxWE5
JJ6HFtLTadjhQDq6PCCS1/pt79YROZNzA9wpGNFZQjCEfN3KWFHaI8uMEiRh1KjlGd8rt3cQJY/F
9FiSiKhqSw24eqwrCUXs2lk/hk2w+0OfSFn+xT1KaSBpyqmfkHdrJWaFwpZO+yP6ar01ER8HHeP5
ebaQGzL9LDSaof1mPuHj0Cq2lfwW/+if8XVRRlGpaViGlQ3zflU0FsuCHQ/i6fH3VSUleFpbF6p9
gNEtZmTbbk2Glj3hWXkIaMtG9i5JQgqdFw9wk3aCS+s0CUKpXwDNrd3PGxhbVR01IeXNB7vf+1WP
SQMt81V1T2odyM8hu/e88UU5wftL/BAJRw++tw56bPCR8ZsWcBTk7kf8goSB8Sb+x/y6gtHDzJ6w
tz11HOJaBqDqjygbYapPLKAwKhba/N3glC+nJV4RwARuTLlnEz4bOzXWo74rqXkpuscg/8vuzsnQ
z3shbtpgFTomRz+Cf9dn/Ga6SNo0xZQu3UfMgiT36QC7CX2ZnTjlj2bSNlD6Ug04go5su2Mk2I2E
pnH+n6WaNI7XeEI/mDTP3rhrrPQryeHVqfGHDjwz8Vywo68apKB0+jqeJEkY2IOh902JxDqe2LWh
eVBb71zZbm51MwOjPv1o3jAwEJ406Psk5g2sijMrzjY9WFYw+znQj7bhSumoayupGQ8etaqqDX6V
Hw6vt0wL1RphssUZLUMQEoHUrirOjnPDz/tnrpWGx7iVNXZIoVb73tbIp1so/DGqYAel3yzbcGEz
mHCTpI8RpcKr0w1T70qB1GjVLLa6c4GvKyX+bGsF9OY62buxIkRHxBMjN0zniO9Ld1nLZUwkcazi
Gfm51K9rTNwgTOA8CblgnZ2hKuG0I3vIuQ7a04Wm+kvKvLsOmC6lG8hDncPPienmi9IEbmjDBvRQ
OjAvGN7EWqM7U73j1tor8zj87FH8DZDk3AfF9RbGc76p7MLIStCSy68lT4Ynpmmun0GZG0D5rk2F
HtY9thCFynDLg1tJgFkVleiQ+ShlXWwrONsjFuxspA7/5xyCHUiL1rYvslrFOr9eJUFYQjjMv0Fq
50StYdJA4nzA4x9+fnZOGQJmZ3nCkgLrRcPoChqTnXVlbMMBA4Gc7u4Zx39Q6bZAkDRLysX4MnxE
af9m/FcwOZnOiNmWb76ho1H08KjLK7cTZDuE6s8QArlV0b6CviBJAnoq+HAuU9VOHBBG3pnJLM5K
EObwc9G2WMdfA8cS9gOP0a6mXd/9JZTXCUgkYs58CrYVlc7d5usjgnEHRRER8LuryJl+NbIJFiYG
hq8oTNhZGeVC3a69A9mJBw3H2WR34KPpJduWLHibzSgBa3FoyuhRT2yQcV6kZbIWhYbCU1yd2AdK
OYmYmuQ/bIPhOA0Tf7V0iovNG+UDfSPxuDxRQHu8gFpXT/zO85bfkazH7paI3fN/tsEKB8iw1Dsb
ZJOWcFq2hF7MQf2v51a47E8XbB7OxxoHJr2LV+Wz9LWKhHwyaZbTMamWBr6pOKNRSZqx8sE5m0kP
lrQ+X2Z9IzkyDpekiV+Noqokr1QspCywg2AUscWGm//8LIifXnkH0ibevBKdATmO7hRa+7YavpmR
rVoETyZxjwkM1cfoq54FX+S1DfJul37HtRsa+SuNMI+Bj4sq8Rbzl9melA20Vv9ul6FVs/AirG8u
ECjZljSMpIO36Qx1d3QLQWqluKd26fm97gWwtWR/fLlRfxCUhLkd3JHk2rivVzqopOj54Maq8POR
DRDYyWGqav3sZdxrPvorda0mjdEG1KwfC0KFuMwocbDHeWrdTjKnhv9Jjmmqpx7OBNWHKA8mnaep
MSWnrONrHO5WygOkhdR02ldQmecakqBzo6AgzcrrbZY6ramGQsabvRl8yibCGpd94unDlU+cOI3s
Qm4xZInUlRhqDxeYlDSHRA/jd/IAn4x4eVfMCf4S1MQDeKILCujNAZyu2SGYi2DnV2LmNBFHKUYa
nD3edbfW7eVOfZIligVdpKYEuGwg6+II4T8H94ogix/hmcijXhTYBRggi4DP5N/GIWmRalFSiur9
4X9oHmbglshlbgTccQZqrYMU9kq40WiYzUoTcc8afaY9k9DjyrSQN4Kej9irKy0aZoGNmvo5kpKp
EUu3vkPz0S5wtbVZJZDu24GiIJRxgmthY+DvnpfZqJYZ4py/GmKH/ryx5V23jG4cTuu4CC1/Gnw4
53GYg5Wyh+swxCOhDVXmyT/JCDgA1LZ2k6S4f8xBQghUEFeG9iUctILhRoa+NKWbGRiwXof0J0r/
kJr3DEDg5c+J6JNOxfQv5IWFo9RvZHW3MFXxLT5tkVnjHcuBEc1XPEa247KMCZqwlW4VfrMSRhkZ
hriXbxKlFe5vZ3asnfLudgaisacQnIKd2Gu4fFSGsWNbrH8lYD/X2DBkBMDnxe2PLNoceMaP39FP
fzP7u/rlUb6slofgW/uvBqH/6N7As9Z9HCTdS9tLjIzWaY2icCjgjLZrvyH3qvhEUAVsiZgI766I
UySWEPzwdIApXG9xSVigEMvwGsb3dlueGBi0LsIXIcSu8AF5jkd8zq1P6vX0ZGwGYbkGpXUQ/CtP
yqVlx9pUZOLKIAum1aeWitB8sF8MRkaaoFuGVAPf34+CtWkQMXHRCORByE4+liP+9tcm96eGvxv4
tf7k/arAk3Kcf4Xpj1NOWIoM6XalcgFiZ+e09JOjucWUjd6QFpWi7D9OuFY7ArN4KHppw8DJuxzB
0ABp4sD480RxJlO4+7aP0HeBjatQWkhp13Y9NXisN5S/L3YgIiuvuijNOXcXCWFAG8hjSdQ1L9pu
kyWreVh4Y0FOKDV/imR/o+Eq0DsrjsX9ELP09kF3Hwgkx5ya3LDSjR89HXftqS0NAHPkj8VXqwyH
TAA0hZEvHC5+coiRabY0IjUr6hR7H8x3NMg++HvLRea7v1c+DWc1T7Xe3+r/U6eHD8u7KRShQ3W/
lNeOrOgd6uswWwy991MADaC0fa3O4ChRIrCj2D04U4AyGM5QMdtvr7K9cI6/CIVK8nJpWmCIVWk+
nn8HPTp/BSgYquK3/MtcEmhtddPojIeRnk165Fi3VapZPejR8YwqxcOmj1PWwHp3lUuQMYa3191C
WQCh28dhX2BCyak1ebfKjSStF328080ZNDAfLpwn/gtaKi/rEZYGy016XbABV5xWHP5CSdplBcAP
2gB2B1NmrnrEyITQoge+Mv1m7CQoSfuPjEtcjZOBAaO/sPkAMo0qzI8M3oYVgIzZYua+Qg9Vw/bz
sP3ABbqjIo4PGdeNUpbKZUpQ+kf2Ku4+GTGJ62BbGVwUS3XyBXVA+P2kmBTj2gsFshluccAbheJr
2J5S4KjNTx7rLuenXBR7vt6ZrNKO1u71QlTAvDTaganJ1hsNbmHuD2WkZqHDKmc0GACpODsfDaDs
cjwpozKhJbQbYnN+IORkuztGMNcnekAIR/8aoRuX+G0a2e0o+jFpeJoJQzIIjRlFn42w/ySP4Yyl
UIQFGVRkwmJ9kyIntGZAlJFYlrKxFWMCUgW1TEU4mg5pA8iAVSu+kq+j2tr355E0CyYsZxKT2wwE
4NYUsNXC1WfMFyFeqjZOr8KNo6ne94pMRm3btfAKkfQ9tB0kXi3+PHn2wZeUuQS/l8kQ9I9kpA0S
Nue1dy+0hreeLiMeaBslAkcm1JGP67mrvvD3dgqsM5+6zvW9nVEVD7F0QhEg+5DhNuJslKNS1mH+
q/IYb7Dp++id1Dep09U6E4y9Csjllp5R+Vd7ZZTui75xF6ATetwFOKyou1fOIVzOWuniIv/qHAuQ
kny87wD56KfLZw9WG9IRjZOI8nnDydcu8l5DfekiBP4O8A1JCo/25WzO3t1i4bjhr7x5JdgUTyU3
th32HBlvB0IJZTnYPAQ1MyCvXuMz815RsvUUubnHh/OHZAaL3ye+plSYeRCfTVHKrAQ8G9pyXUbo
vw2EbE28mTGN/7pv8emWrA0aECi+C7gFQCmUcxNlrmFMue4bEksvtZ6l0XSGLQ3hKa597NS9ZLjg
3BXhcDXtrBzF3X2o7ghRn34BBGu/dCQUXR1EclcG25S0R3VvryCVrJ2u1kpKrksPlt0SZxGeQ0BN
nHLpP3tH4jzlP6UGrZFOK0a6+AOVB/YljkCoJGmpbCYBrchesZi0VpQy+zr2LnCsy6zlrkdoxXZ3
jntPRFOo9df332kbdErZxMyYI2fqgsC4XHX1dDCAgpAwknmgRxVErIUK6jXM7zyJZ4xuNsW6q4ol
gubZYmuATo0HkhgjgX3nVh0E04GitaD68Y59PxPKlCwAz5UPd3XslXakdg4k4POVhZq6nMAyvIuv
rIB0R+K8Fzx5kHwYKck4c42ePC4U4ja63gblyH5TzpUtpFbjBppiC+7lKj8KzcVtQbceDYSvqneE
Y1qLmiOzX1LO8Cm4WB4fU1IL0b2HCqOwzBPnHz/3qP3wJ+DDEJDTzt0fgGzM/S1FzqCcesStJ7B/
gQvgSEFpiCpFiRbp+Hmjlt+Mjk/bkF6RX5HwWXYIPpiDLEj1rt88aTxRqYsE+9wUp33MiDdJnSe+
fFGcGh6Pojfu294PEVVF8/rEDajnXuR+V4gax0CI1iwbPfr30Ph6XcnAkmRiLAMoXpDAXjIWvZYN
b/zkTNOOQtnd5RPfkSFQfpWyqwzHQiTeJ4Sc2UlxSAOoFJ025xwuSJOkdV0fbkAkdyXWjLy08Z9b
9FmMAwPs/qaXJlZB67KM+FXbJWcvJKccace4L89KApVKbqRVcLJlvRDWV/J09rx5w7js+yC5SZjd
7LFKDw6sjcmCa1vnEUIl7WjJmijZha0SxwQlChERsdcBbBjbyzKOAgIxY4AFD3ySgcx7E5XdvUjq
tSjqrt98PLez8jSW6Rv7bABh2qvCDAqkJDo8ZEdqGF7+M1h5s6+XjySJHk26xKHMcAtglAbyJIEO
jkrMfixVFDKngLcMFwfvznMaFT9RzyWeh6mir3IkquRqQMv2NWHlHu/v549V3uwhFNraB/lUhGda
mrixUZwQ5duKSGAenZi1GbVlZ2c0rOqaNhNijKOutSK8j+Rjna8PaCtmXnJG519RcVJSxxSyX4C5
A+431N1VsJyFJnKkCkm/5sDQRNs8d8NDZvOPw5W1xw/nB6AfyYljo21tUC6kZJnE6o9grQ2Lifrx
FB7IxtUFJCnKm+Uyn65/dqFMtERr3ychhDIK+XzLsPDNIgEz86YH2Lk8umLaennwREiKuwKSVgI0
5aUnOt8/JzagYMTQDXlqtDauYtJuSQi5ue5mKFt+J8DMeYZwL8Uh0nWLYM2cwV2jqHlnfyqGz1Yx
cVofYj9X7yjUodXPix9gml2o2H+JaiwA7vcKHlaHZxx9i/GO/RXowcQ5SJCWOaQXRpRTFpsAmKDm
bWk342isj9giEBHoFRrp9tXKa8Y99skXgLsodSEiBdxK19WeQ2J0pShWUjrzPc/mWpnpNB0+gK6D
OFm5fEnVThtFEorcV6rORySm1OcWtf67PUDSbO3FnxSHoL8oj1Vl8jl4Cyozl5vrvQHVToYjOlZd
3Q0o5WRHT6EdkLBaNeCLl62SaiRygeN16Zpw0bf/wFGJENUCuxo6tS9LgkuRybzQlEXUA/Ob4Y3L
OSVHm+EBQ8hfo5946rTHnT5iSDltN363x398uqjH/x4vTFFlQDIltVxgqs5LKoBRaSaI3KW6M5LG
k4iK11IoY0K3bG6Ir14fxC8wFzOCQcdh/90rUHO+dXuJ5CpFZHjMwi+PIZIykv1CeAMFQ1iA9iLP
b205yIfTFNVcYVXOAgZxklj0F/Hh5iBCgAJnk+LMnM2cvLrvtEdWU2b+Vgmv/x73kJtOLb2nmIYG
7w6+etwydF5c/bxiGBDWulEVqtKRgv2ewInd2uxqTxbaWOJHNC00VLeiNEkHAXl/Rao46I0qUv1l
p6629ie2apCpwGycRjvMsiJnUrrMX7//cGwAmnHMYeCN1B0RBq5RrKNNjJOt1ZLitvPAspSDh7/M
QSX0nLldQpXJRnVhI1KkrCuie77Y6UUMXiABz7MUtDelVFcY2CyWACbpeduOYZOv/KIAdA1f57Jp
Xh7EiJL6y4qLsb+OHFFeVZ2E8v6b7A7kFBm8vP4O/QUGINIyinNWVK3pgTVQvxhnqIglQ3iMMcKZ
orZNRHqY3Vc+wo/YiGuUyWAwILtHLiukboqMceav57qJtwJ8SGyht6O4Or8Xnl0YF6wnQNirQrDJ
jqVZ8TKgbICKg3ZY6WkknIiwesKbyD+MB9RyVTQ2gYJf4CmKzNFP+2fTuCqx5xyS+my1WgbGyKOU
OcmBzdmXv/0nvlj+QtQ7cFHU8o4rI2nVYTCQ1X6YDRn4BmthBhgHmezfUVpiTmjeboDFhL97Gv3G
2fi6hEBFRj5T1bdCFZF0T4MeVqepkR+CXlclCYD2E1giZnIXtw2uaOisxHEMAr6haO7y2hFy3xv2
14cLttlgv2Bn+rFcVq7GKMuzl28RxNub9/sreLL8t6x0K5IX5IHu07f+VO3ra3tPO3eKJDfn0JWg
fvOKs3dWZqI38duNaCmj4eLrrmYx1I8cT6317yJaQGed9rP2f1ndyiavo41IrCaJ2IiiQL6AJHhT
mLBS4pHlw/N9ytXtsnsmlzJodzUi9ewv8L58vNaMo5j38idDTDBlyP5eDTMwHKMg08eOfzAeQeuJ
puYJkwpaij7C5dCEt6V+IYFJh6pVVuw0X2ErgqxBd8AHAzg/6ugnd1ct4We810DWn7YGqvnfvDT3
x30vMoNyrGJvQ3zk5fn7xTI2UIXxINT3mWOxKrwiLt87lzfd/PxgzqjqiCVusGrRDOOE3gyNMx9u
wc9klFPHt8GvCxmUVuMwHT3FMxF5IZ9vdXoV5lazMgU+VzrwmNlUJx6Yjjd9yEAz0VTBygkRWW8V
4gv1HFeUn3s5SHgBx/CK3JYejfN7C5joYxc3NCgFUszbHlo9grd2wsYm8J/mhTCDVzrhjY3zeZWv
D43ypzXcww8k1D9YMXp/TOCHtxcgwPV3+VDjwsobr/D4N3Of1O6vRVMKyxzIlT167Fz1MahfuR9a
m48KZHKYkqqyT6DhrAqvclb6YH81jRI/YXVLKdBo88D+XF0BdHbpuaHYmlrSkTaJWylbNbNnXSjz
Vo07yzeeljN/f9jnkS61dLNrMOoKXxSc0SmcOdbac86Y2aweUST1fwHy4w4Z8bP7aywke0pelVrZ
ty3jxcs3wb8DUIcfQNkLJhLmP+bXagcJMi8+tyzQBbNol96Fk0yXOv7wxY7CgCvHRcx1fwXCl1Df
ASNh7G/+N85y5+513tsjGUvDcjrJ3ifqg/sJcHO3pDtLoYnhxc8974E0Ns8LzZUkSWGZNwzth8Yf
cORkgUm4wWruJCLlrycoRwynJHXrwsjr5mYNR4RC3SMSXOQBbVM20mYNwEaHNiITMEk5NyU9iYY0
Fg5ubMH9CFeP6YTEeC3g/QSoZfFRrPMjVWUQIRQzkbn8V/Mm6aNEivUGMbsAV2LQJZkvgKR4fsin
MkujzHKpQ/NBSxfeqLeMnSjlkejZJiaJYsnNqGzYPuhN7pqVFy1ffK29x5y1MMz8OnjMAc8lxBn/
5EE96r7lqLqT48zRiQ7sx608HQoHpwZeZh127qxTAl0bLW4kyaSmqHz5ugdHr4JX6GiUZHXHX6UH
IjcLSHquMgs2ITtYQ8tNwqjBrQ3dMI0hxt9vuLHm5x8YdDoFD2581F25Eo7M/SXvBAhkvjexk8y0
DSFVbrsG2ogd8fvJwdT21BK9Ci8fs9GrHPd67jzqqbhsq8bGSv/dm8zk9FxGU0EPdl7gJsMo0t3Y
PDpHq0u8SMiScIJ2+MlKABGlV++TvYMC3v38djCP920N6O0JAUJxsIuUsqadhI0eOZrZRzi5NmDv
or2MW9gEiZPaeArSeanBxIAmKJy6OM7rq9GYffmQo1S4eExvw5JLa0hxCp/KAgmQodUc45x6HHAN
YYK86R+Pow3qfTfe0MbGN0SyDQ+cp4mfOp61esOtyKcMjrnGxMdbOdb06wpHIKVeK14nvmqJAaaM
oB2jDWlpOyyWSsAzOyB7poyCcXpVJb88bsySmAbNYAj9oEZnuuaI/iPmdaI4tmiv1gx/1RB5Roqu
7GM0tyhjhRxM10x4Tu6yGPU6bsXhrMS2aktBQLJuWCa8s4/8ds98gPwd78+LcX/vlxhyG1pFUVbE
l3GScJ0Cw+T79TWqgK3AsZS9Y3i9fkow5xlBXeLXhEsAKZL/eW+5qkwYp2dVHeoEifJaI8963wn3
+18fDCxEq78tcNZnWVfJLYhAIhG3T8DouHeIGRs65myWK6N0i9xXXvxfYlh3STBD7GABCqeMY2qM
/X94vWRjZk1DwCHU8Ks1XPrQPrs3i25K3hMVnX3zuaMgfLN/KeitSydgeREhZTwXQ0xleVP0VAMM
LJKBpdjW9FPkE9UzkipD+18Bd/29h6nd8UcAaRpF3m1bwyAFebif4lmhg2F3qdnTqwhLS1F67wEy
od++TmuKdMqaNyNUQ+H0U6yCeKgX2XdFgLlqqfAwzHoU0M1V+75M/InPEt+xNvljFkYMyhpmyhQd
RyaebqZ4uRcMP+XrQFwn6uaYeMeBPoFlBX0n09Mm2od/vCGbptgHWxR+geZ/IjPRBaQca3FT0Pch
n1y4yEIvEloUzDXNDyzyZBeoPBaEtvQUFWT2xDPcKdG0SW8Iakstsgxp0WU1Jh//YNNZxVAe7m+w
w+1voHG+gHX0400rDCd99d9mN8UAbqJxD7S4ZcI3p1SDrif7REWwhidVY+J8kSdsp7rzdGw1hFQI
m+NDLKtYIn6eJtpAjRdSF+VNEWg4Az1jm2Z2L7/QK6nQAAcFBQABXdr0xB5Y/AqnhsW5dcJ35cfY
i/mzK8tccrA+77eSHJp4lC9oCuut4e9GutW1dP88m8fHZJV7w4MVRO+rKQzwcKEZdxGCdPNa4v7F
pI2vrXRgL5dCryqbfKh2HNGWudf5Y48QXj52RzTdSxn+PyCeXjTyvqfSxKDvmiY/MfuhI1bhjght
S6ZDd+15G9QiAgA/jyAlkdC5qelhEcVsIPYZLMjTW1KIatiqjsKJlaRFFxMUvUflX11S5zCHIt8m
dE3shbpwuzjuRjFYL9Xi2CXtjvpmGl7xYxIP6FJoHabuEZaNaoAhVDf1FK9ay4pRvDHzsP4ropsf
ytmTEF2b35SKO8Wlmae+24MWylpGiUTiPoANyIW5cANFz1crATylzs7b5zQ9+6rsxdnUZfc7ao26
xTnN6T6uBI6jsGObQ/KkStqXJ5ceQ5Jgx5wWPlKWgHpClttxKFewRQYpgWlgawh9Bup6anrSPzKi
7NALk9ELFrjJxfZDiL3KJTahO5LvlHIPiIMPbXnN1HfZBM7teWXucs43UmlkzWMCGK4Tc//Ng38L
WU/qsjMnS4Zk5uc73qJhGYmjKpbxhhJMZSK+/eDjwxj8utwdmGP3TEbkAM4dCjFZSlWvvwNfgJyN
JAnk/1JsfAa9JyTm4K8qxs5iDRDBDUihS7gblUpH8ljV7Ybdwn3RE876Dyya8t4ua9WRJ8uVwqtX
n3egkGtCamZXdPA0c8OtL8/yOSilf5fAABallgKXfQLu6XEEx6vCC/QP9VO29Yr8ji59V7QZ4QUH
SQ5pPKqdvRE4GfzgjlfeGWFRbFtomj/39+AJyZS52ME21qbrEEsEKyJURHhuGiyebUYwTNiX3W+/
ucRoiLdwVEbVsDeLKca3RbBUqAhJGfyJhlKsKj/m035ZqO+Z7qwlzP+lxZUKR5cxHkIBl14b3wHY
7jPRQc9FMRr/pkRsewSWl9hsA80n1P20eAjGvxJv1RA8xQxyuYSjElt+tunERfJt2Ki2xh2S47e/
PvdLL6q5tuwVYmIXI/+0SQlhBK1LBGqG9WeShSb5uiDstwOk3sZtd0vOrSZEeU1AXkhKWz98l7E8
PKkfWolBML5BGUVN38LGzTtYFIbv8WRGFhsvCC3p/nH2wDMC/BJVJtT7FApuyh5vjPWbSjJWRL8G
Ucq6aNE7Yns19sjtzpwz5j4eH5mXkSgNK+RCJXusyog9LKJErQLvFw0cTr9DTZ39TsVf7vxYsZQ5
B5vDWpAThR9mKAEn5AVBm5tWnAl2SDhA2HHiE80C9hAOd88dbC3s562KJBBLdPymQqfmwdLb9U19
ml8B0Nr7/zgDLUbqWNkpYdT9O8spufdA4LVfOE0n/crOd3RXLT7XVY/Q0KQFudt9j2o6Mhjj/Yfz
eQodPsaR35Z2m/+vscHrL39njy9l/a+pv2A+tAWqYIc+EgKt7vRHV9RR/LS4F2EVrd1c7K9HIUpI
UYefwVSbFfwAM+M45slHO9iTWGLXCkpMLm/avK5nq1QKGbmWDnf0TouQPdkM6ixa1u5pi0A4Zdy+
k+DJ4HGUl0AbfkxISkkuzAXzqP57GgpE99fq8ooPS9fWM5fmfMtrbeDY24hP7mGAplGjHcbia4Zm
QQ3Chf72VB5EDJdP+mJemz0+eI9SDVVQp94j5z+m7jvL5WsCwmOqKo//CpdVb2XfbBHz4w4M/dh7
LOaMpu6v0FjCAxvzsODek+Bqe40Og20gcjMKlb4fs5TJKXAiLdNufFVxVoNxM8G6plbcxxI1tCP1
INyD6exO60xY7SNJ6uNJHot91LWZmKbVXIJWtftpYKK7zQ0wzjAfxxPNLMU+elAruV2RDv/LNbeY
LnKU2nXv8jxk9CJvylXNRhFtyRsg34HtlD8JKeeWMHZuArcw/Jlxo3i8uZx5jWQ/pJk3xxFnENM4
4Ejg2lvYnyMJNaOtwQK6V0VId51SADTtbRLr6C4jVdbM0K9oAXYxEXKztzpBZhpZxROgKqXO5V+v
EuD8Vk9zqXxXdR8+Fnc9CvZhdPTeEemRlxM3iN2Lu1EbTcCRTiTkJ4o/Kd/0FNHqlQ31GoP0vb+R
49SFzf9lEStgty8lcIdhBXxW+3hQ3l6ZXiukWq95KDaVWF5MdzeZKe7awPUONZcJu3wRLWTvRE/x
nrkf4Tq1BdwAkHeIaioiECnRPN4enoZFiroFAATyGXuUgz7NZK1uYmNbQunxlLWr9BoNAG1IYTWG
9dH3X5qSUTiHQyaUoMo6MlKbcbbz9IUcgQineF1dpaA1sAZz9z1BL6PztPYBVQB0d6nTKM7mj3h6
vFx/AldNocTsXiIHKYndGuv/pD3/p225EaBbU3q/wFdEbfpXjJ1izSTMcIAU2JjJwL7AjymgD2Ne
SvLKqhQaTTPfSS0UhWOSnvO/urKBCoiyiOGxQ3DenxOgUsfJmodwARXMTDwgdAXY9khupt/PCJTr
XnbcRECvZH3UnBIud5wRADh57ooss6gONC3JQQm2G7hTHMAhmvM320JBpnzyEfAb+o3tpPE74C5U
i3+oeBop1+A9z7CdvrmuG5Nu1R0RfuOOv6bhArAqYhA8EOPEOzX606uH3DbkP4RqUi8D9D1rrHQz
roxcl7nCsp8Pk8gCOiBjghvDLTLSgDtKdP9Lj8vtpIHjgodlvjc2Cd0XNt+ImL6N9a4bMeZrMJ3n
CY26jHVlvpOqXg1udR9DaghoT0Z4z3ho7V4qhYICscFh+rUj3MYWFLPJfwTdsmZrCZyIMrMTg7Z+
YbRigpFjaJfJbvfCzS2QkmHhXL29446iJIiAqdr3xUKVPsu00KNYaptdrK/uZ0p4bz2sZ0Qd7db3
Kqz8GqRqNvhP1TjsWEFLhonckh31ng97K4W6zCWszeNYciFTqj9CFHeAOmrFUyVRfnL6YVBY2q0/
xIgb/yGEatgrr9rThJD4SK1TObeo2o5DLtwSgsxIkFh8LXks4iSIkLmNgYGkJRkbT22NYntPwGUp
GDpP+j13hFCs/hheJS7uCENYCe9SuaWgY765V1H7sM2lnRPuUKKcUagDsm2jLH98Qv6Pvq1VxBVR
4aOqp2hZiZBQN6pA4HsDbytoI1DAt3qJm7SzuxivnONsdNNGZ5DnZEXwINpwZQNtH0/3MYZz5gAr
wxo6gvsJ5CV6x4ajiY3RjyBpGnYgSv4RuRDmn19c62GhpRanHJ8i3mDQwQjXBuLPui89N0KPt61d
A1XI5+gNOd8Mx1WHrVpXnOQojtJHKIP8wewPjlLUy8TzbMyfu1Yg0eRiSIy2GjnDpXOxf4n6CIK1
/GqfcNU4Uksx/1FtjacGsJOgSnrkSFXd5xJNsg1W3GE35r/A4q4Tj65z7BuhI4cGe145QL4OFs85
EL7VgVDh8bgSbW/PsCBO7DLrN408Q479buS2PMmKpmxlNuui00z2peoNs5LaaIB6ZP3eG5EKP1PC
P5GGr8W2eAVx00dkAPTt0Qm7FWgacWvl+jhkVmL1YjEPyGSRiXU3u10Fn4IjC203YKol/ez0XeRp
hUdhkKLRmjKzgKN8tvPlwIM5HV3cGRh98W2zXj7a7HTO2bwnr4GD4vmzR9gFIqLHZDb7LXYsYR5g
/JTfbtu+th2hFowY8BufynPnWG3cbaJtJvLBm4S58MEy/Z5WsyqVFiCtdCOMWLBo5aKZLy137/H0
FHFr6rB/PMOVXf8CTlFdkZyt/Yw20p8KCGgHfCeyyVWh9eYkgWrplOxytiWjWe09MkB3digo6O3M
pv1HA2Fq48/ocBIkzLRAKpDAoVb32Ot3i2ijCqSuxa4e8yoTVPlX9oH7t9ohKKz6D/uG45FGYv7m
uvmP4FahHl4hVd47MaGRws+oUyXPK/HLH3ok8sbRmyOtIFRdvqgPQbPNjVnDJNjS1BCzYG8gcscH
XEQQc8JGH3GF9wpsQ42aXIN+lAcKS9LGExAsnpLWDxZzgKWyNBywJjbWbbcsGFz70gDzhQM5vpcO
++2rwGQ3f7rGXkv6IisW480jXcxirjNTGz1T3CIFnVXSIxZhtYK9jhFjkxRyYaoFfk3O3VU/DYs9
WPXFoQJzpoFBKvsPwwJanM3JIzxZQ+vOND9ly1WrcGvtFGj+ghOA7BYZTW/E+vhLsn5O/rfGyxmK
Kzbgwykk5iwU1KD1VYik6ESNFQGhX2IML0CgEMfGcrnrGP5CH80bU7g1OHVA1UXnGz3dvLhulrM7
PTKa1ILLf2hKLVRpSGooc/KFSsdwXJjiOIjMWVk6baH30GRF7jQPbI4WhVQlkWOryg3+Bl/CgbbD
RwI1fh6rSxXJwWbpqFkrKl73nK4K07JKQB8eKZnHF9YzOU7H3AhbQnED93B55BhlqmXHRo5k7uON
xENzX8g7F9VUyt2P5lMmYnOmnqKXwfdQ+Xr75whKS5Ntz9lyOki45urnOVpBuXWx8NA2XYCyVvr1
yze/iU4oqNYbAnGUVAR/a1ibJ5MGUNPPE/I0Bu+b6unEhWxRpdz7JXsSK1uQcHL40szYlv/DB7uI
I3fdyRUJIPdWlU8wLFBqXocVUBVh7EzYObE8XWtc12Z8Hy6mHMFDNF1kJaThJGFm2Tf5vvZMntDU
30ZFLVKcEuXRZpN18O0B2ErxDHtmKkKby4wSpyuwkSNibn9VUGBeRh886xB5HAq9yLoGnv62ISXX
eRl1cYkgG+6Rnvd5doWn/pR2GwSPZVkCCoLB5V6ctgzk+K2QzRMnjcXEeOtrOO5ZJAK9tXRNGgCE
4XhZjZRQIz+5Q7q1S3/sdh76eBaEeUM/pqHZWRZjlxJ75PIMbbd4wQ4i2W7sEnTvTvWYGY6OSXIw
KRf93WQR8mLuRibsZLtdQLibGGrShpd9+z6KvQhgUV/FYE5eweSzpO2EdYB9w4cHgvv6Wea6EVod
3uyAVARbBI90y00Cl5DtfA3OUmW3lAcsTLmlMyV+zgBWsSbBrb9eaGS77WNw9hmshR1CORTAkXyc
uDrxnS7YFe5xdSHaYftQzD0IP+D5tpeKQuK36ApauFCN4V4gd03tOReXKtqDB5NjliNBTLVKdr+U
VjmWa69TPfYG7FOakWOqUeEAvf+vo+XykDNtYNrQknAOTkZo1w7iXppFc+nxzAyUECepW+/1Iuh1
2Mq+gxcbj/Q897Vzo1mrMGa+skzv7kZYsrOLZVnA7g4AFsZAlsLqT4EzXANEjx+CihEWrM0Jl8ZA
arbNrsimrmIoKtqFTDe7B9D3k1kiWsgW30w/Mo699Ql2xuGPjHkkS4Kw9HPSzmQImDHptdkDZNwJ
OVVclYSCaTHH5JH6/q2fYUBZ69j4xuhSD+6D9JAoQeAFxJ6+Fe+L8VII4L79rQhmrvpgBAVs+IpA
6eBEArfBcFnwwWmEoxjb7DsqYDQVuEKdDynsRkuc+kdrpzBEdQ4IiQRKDjCUm1mhpROQ72hRWKsQ
ckldK/KZRK1gaTGKayjwk8MlBMFlzVdtbNJ15AoQmoAzCMa0uyVZqiInPcb5NaO2wnX21wsMY8IM
9SfT3rZH5FJCp5fGd3pQ0knf04xwwlbFxdtev3aIQySvcJDemnLG0kRybLXS77miPDTwkRciely7
mKxCNxj7Dku3xn1pYDVrnBvAl5kesLqNgSeGNXAccZfQJa1C9qXZv3dzR7luoAmzoCUzl7Dm2sMU
UcsFVgqMyZtttRxQUlHu4ki6R/BPrc/XJPeSnzy4PQs+6qoEQ0OSFlBtpMbRou5QzB/y4e2f82uV
amzh/vRUk92Sm5HErrsxCjT+v5uKa+IRNNrvDWtQT/vAH3hilJDWbyOxZAAP7TOaSBrm2G+AZUYd
sN2u/GfBfEWubACuy7fC2RDiwa8FgtP3xWK0KabotRRppteF+gcUi57y12HLqjWn6Wzf8m+nNIBa
BDwg6E7UNNbB8/b3FQ/xykvMecyflrjfv6yf96FwpkWtVP3q/wifICfn6KC46l10u/3pwzPczZko
bKdDp1h+8sgBc5IU/jb1e/plSkhrh1yXEddGz9G3qeZamtLk5YnG7iYV40U98X32hfnvRzcOR+Lr
AIjooUkELWVrnILkjoNMPcRovGUtcjdWn6g2BEPsxC1Ev2JRkQoJ8WpMXeHI53PjXRCQCtLH8zxS
qfCknGSr/9J/Zygn/0u9IgY9ZQFH0IRv4V9scxR/JxWvgxSmco/LWLoYC9sbMlrinogC/92UKu26
WLUkr6S5pPWQP9hh34eeV/mJSdMofXjo2E6QnC7yEhv7W7QXV8RHjZdY2ISfzcFuflwbvYjllWjF
O1f+ZkTQqGW1XLbWtzT0YY/z08efy/ITNFX3seSO4V1JhW27/jr71pwbIU38ce04PwBkxeomCSrh
uCYLlJO4oXpYmRjaIykLqcqC3o5fWh+lRJ74Y8ZRJv/0On/pGYKeTi1vN9b4bxlaKBu7zAZF8HiQ
aEua0qFZqRhnkdkpgUV4BuUY+cV8DnN42NuwVj7Ak9FjMNJJ9FAUB4pTCLoBleUbenlhrbf+u5Qt
PFmn1XwqiTA06Z+ZFbVUO8ijqG9UnWIiWvM0Tc7PHDqYxgHBzYxEe7JKNX0vpPt3dDTSwr6apq64
gVtZZcQXm6To2YdX7oLbFn5iHipVSbxA/6IxjqB8lJeMsPQpBxOxANGUojqSHn4eOu2QkFUfahl5
1NvmNSnVMAhyfYMhz54u982BZJ5Jqt85znzkic2eeU55WGVgkby/D39qKlKpc58uB40bWnL9kkYu
DgO2DzrWWXsdhzhidsbaIq6XPBD+b3y2fKaBD5AkIbnmq2BgP2lXXS3pzwkg2DdE2H6vYQMPBOAn
pKW60X5Rr5+ZPXQNL/Ql6IXqbMT/9zo11tbAYgbANoywuneTyOQVVCCxCsRe/FxDhRsAJOZ4wXJs
fuj0q00ANSQyb7UHVE/gSB78nhYtZiFlyX5KDmGp0lLRbie5Qgq8jiHANaynScSU0i2up+7xW7kp
RuFVDd6Us+V3P06Wt5Lj5e82MdBYJq85R6nPaxNjV9Nj0qkcNnp9R1xDwOGKkE91/mY4s9HuA1A3
TEfjF+tdPd+BI9jFxLLwE7k2epbcI3fS+cgv9/mYVm2WiEYBUQ9HObr9lKbTTHkbiOl6O5ka9jeM
9bUf261aBwajhGVxpZXptiTpFENnoX0aOwaql1Bz9WkZf9C9lhnBYrA2eISTAvJP/Xspc3u1b4AM
811WtiP63kdLSl7+U1bdQchp5iFgEqs1T9kga52viktBiSKd/aYW0Dbrz0Kge76c5MCSB4dl1o8p
7TepZKyplRtmlyIxTKnrh/jK0RqVROkiBm3FKz7bmWV1RN3bMFPmBA4Ws0SIXxc/JaER3W6ciRGs
VIMN563dD1uA59y8OYHkAOoRW+t/kIEg2ZrmiQlgoZTDry24W5+qkK65Rfv8Q5fDPGfjP2cSRuTE
/tsmqe+UmIkqthYRekOLD64/1qFNjK/3bCZPjLPbIrZ8NLRFNdiqDRv8k6HCVShxgwTvdEmk7CKZ
x6DPeKGHgI1lcjo3zlrZa+sNqwktcDpa+cadWORVkl3E28//Fhi3wSspitnm3NJLWkaCYqgKdGCf
KD6g3XnSACDZMIkoa8EnCMoOSOcdcLwGfkOXd5ArWUjOGJcEjjnAXyYbQ0kXLy2SpAsB2ckOvd0+
9l1jHrRcbrDhnZlfk1cpB64K9Xsu+pkH3Q4WBSkJU9Bpa7yugctNGKf//l5+Qt6Pu3HuEO6EEYf1
VKZ80rY9JqwFIghvsuHo2RZet+rfi5ZEj0QxDLyeLbm+huhy/zg46Z4Yo+LMjFnXytNxdZPZ/ReW
IPi5gpslspJFu/qbdjzbTQ4+z7QwDYXneEZxaEhxuNkUcUVfDTEFgK84BWxGiVqwkzendJDw+dqZ
xskQNZMb/pcGZE9Uvt/TfEgoaC+ztibC8WPoNv+yXBIbqys0TZ1wG8CM1psUTlRM3cMnbAoscPmV
cafolQSxkTIptG8Uy4VxTq4Nb35zVhdP51JvAgYb4RZM18KBa2F1bpAHplXyYQXUN7/BDmb6jkTM
r+XLLLSnlcALe6yGBOdI+3p39Hp+ebDquMOXqzPSARC+7H7PaFjY+J/dZUsf1f4kWhPC6DxoPOI1
9+qVTXvpG3PogMEjNN658BSWPdB69hu+bBqwFomjdyB0ElcVvp99+WLayXqYQloXGFs5pi/F/oDp
PZHJSVZuYj+qw5YrCrsQ7oofReVD5Tt2CDljtC/VCSB6JpiUXs/X7vJIjyB9R9m1azz9rOlzJ71k
1pAX7BjwdmLPFOVnK8868z45hL/caq3PRq1h8tQI7LV2hwOBOaweb89IDa2DDjkn6LSRSeYiOHoz
ZM4wuADCUt5PMmK/zZ15RFpz53t8DOD0sbSTbbhDyk9L//aOnVxocN1EwEzR6dTf5etm51P+1dW8
/XtlYSEms91w/0eMSJ3PyIpiGDNd7oTS7ymzV9pEAfHfRYYB0dqMZZxSnJVCe/hGRbhB3RKId50o
c+pMyqFk9zyIe7R13ZjvWazeoDjXkO7Vhvgg2ycBeeJ/9lPV6X36ssV6nu0No+AdLEP1fjI8hBpN
MwF3ccXHtAZ/F/Nj0TrvzV9qDOtGAeRxIxDryaTaRwOEYCkwb9/XLOm0rGWNsD9NQBsuKpjVi3i2
9uKQMzym6SIgY074/KyWjui3i3NBQjqzlTtegKRVPfZc5gmBuoHYUO9wMP/ZDluaNRBmK1embuoW
2xC9p2LoWkisrCRGjji5/x9VLHaj1aalKPjeBxkWYMOVqYz5spZl11WoiFKsiff8H8IwWOdGOi3o
IrXZO1Pocof5Ya2TOZIi6phwqz3xpl4POF3QrIS4CgUYxMoKOCaHOzXf5tJxHkkkBSg9nLHLxRA3
IrBXZBsgk5HUP9yO0vn8Epgi1vLssJ/5zsZtnC6yBhv2kaEq+QYflu5CsljNrxJ12zjkhePn+rmN
sTkUHdPEo1beLSbq/Tc/gzOxMWU402jaLhZ1HT2JPgbMIiu1BtXaYdB1MM/h2/2dLs5uveW4+38i
jWLI/BUVlcwCMHxBCEP0aaZk2HVHOIWmkwlBrbiMAyTcwMNkWMfFqx62Y8NwH6iL33mOJazRKm8d
gvutiZ1xZDxvRorFIfhE9eaMyq36HARt9Db2yOiQTA5OUlIKC61KM5vBfS3gN1lfVr5IY4VsYERu
LbjYkuZr0vMvyfW8u3M7qQ39zSvJTWxEa9/Dh5YN89Z+jA9jSC94WuHvV3NEBYxoVClTwFtKy4N/
Q/QU+PtWI6vk7gguN0NEt38nEN2I1cupEaOGm2mWY7xhA1KonxTWd1Z7+OEd3jdDdRLS65jFv3xh
1t2HxTU7iJM7R86wOCTiCNSxAjhRp0A4/odT2HcHjKY/jKPMAcrBUa2kfzUR2nKfySjGpKA8OoS7
HsODQ8ZhSMrTwuOh0Ep4MYKC8pTwCcQMjEY0Y5z1IuIOGXmM/GkQ/bTd8ExYMYbqP6ZzPbJvE5ik
QPpLvWAv9dFqmukpoj0IAZtoExAYEPuMpyAnEyrR4n8g9Ti3IN/hR8Yy8uOgSXjYesjtDavIBihW
y5chlpY34BtLxqbC8VJWFPbuQTmdAY6J5UbaJZsZGakcwwtRa35rcv4THaH/OWDMoRJomihbSOZm
W4pYZvxtupAPORZ1HuP/IMWN8nwmPJNiqzz1+lJjKXYtJPcZzqOfaDNJKAJMdihdXSr+whk/9JF8
uymdIJC8wYEwJa8+g4S9vEFumNDSTpJAA81eLSpHAPl3+k5JXX6DoZ0s1PCQ3IKoWT0LJxpLxuAM
AphAYT1a2yxqiqrwbzKhrt6yUKV02e9RUneaThkzGf0KGqjx5fTD88UAuzp8oWynhzkvs6ctoHg4
yIfzH9amHj/V1zS7arSaSacl5Ld8z3G0uIcouMHB0yPCEMhFJwLyi/RE0P2E/oDERxTT3OUi5LTF
nuPyRupLBtWtAQoYx8hKdQnLo8SgdwG+VnZAUYqy/f49JDgXSri2tbaujzar4ocCj36ux7TNRW1P
m2NYWf3z+pGCjxjyvIU2BabDpA0P3glwcoSVJq+pTlYBYiwQOXbBX4MNxi+E7W8X0NV2WpmPfXoJ
hnRIeyrFsBF2a6kn0ovnNrYO/lynraX8SjuBYQPkAr90hPeEkFmcCKfR5WO4M+Vm/itFgEu87afV
HBOa89N4FEXTZ8YvW5InWheBj5Wx5sIP7yLbknDiNm8a8BSQKntENGb3UoybeIC5UJVUbD4ZHfqs
/jpPbipNggbvOp4FL2fV/kKe3yJh46CiQAEWp7Mr6EoTqQBZFcnrnN2G02ssF0JAQooSelejD01E
ZimpmxwNKVgfXzYZi4qFn67/Rn7qp955o1wDgoeqiFU5GQKlhYatlBD1NBIl2uqVYS12O+VyaJm5
iwbUGQ1QUPHIV5cfYYeMlYcPuCkWUEGwdj4hPq/n3eIt7DJhmybc5yv8hkkknAwPQiMx4z4iE/RL
Avyz44o8ZFCOVyu2UPLvFN2pU+u913U3otAKJnt+WL/BU0EKykjtBDXydknIoql+b6+0vJF6obRp
L9JCak0kc0xexlS2bkNey/qL9P8dNSG8+dX7NBSJAJWCx5Dy7bOV6edQ3LGTR6CtGlJv1K6YHZNP
DV+gcnQ5tMhLdqdBY3ltZrTbbyzI5c/wQ4Yq+mWbfjgSqhkt7MkDUBQaA8i762JapO/j4RH+PRxf
VL1iI3Nuiaf5kZDw7KoWDUyTGNFsOJDol5eFUoefiziHfLm0YV5oyXqxkTbClzp/5+LZ9Jy1t/ju
ETrHwaXxuKE4IVPybEQeC/dF+AfOwoCKC2sdjse8+udbYHj+VoaaCS8/psdhsNI3F212hT4oB8OP
6x2/fT4Ut8Hjcee46TJqzZDZmgOPLXq0+uholS3usgR4kDlZ/MNpWSgsAq33816cJdNGJ2HseYsQ
rildgSM3khmxrV4DVucDuHo0xASHjPlnAINbM2cr6EQvGiUnWZJkXY/4dcth4nQSLAYbas1gj3xB
9bKc44FMtnrG2dVbG+d6zl7E5dmAmWayFnDmvUIRlVVITJJp7JF2F7EiDxt5OjtjDb9lYuYggfDV
hm/p0eksnfUke+vSn7RKNzp3lNBByAMw3bCjvxiDTCLDiPVpmZJmmoKl+SsK6joVPyCDANxR1Knz
McN/PH+OICGPmRKYxpYA0Do8ILe5wHyLMiaIZSE/DZtWsS6bFVDjne+HhuvCffNQxUlqNK8JIBAR
tfoIR/G2iproV3U8vO5knDDIjbCDlETQgGf5BH3v+rR1sUY9Kpav7bVPROkUa9e3+X7WTZUGx9Bp
pgDpKWRKDLvvX0+nEYSa28K743C/TnorbNAnFmd2iXpv0scUeBw3DzFdiDI4E9+Upjj9E3FilitW
pD4uCBev/7/WGijgg+KztRbJpK98vQlZdBsItODK4i4P81uybrU9IYKkyPAxILxA8gnv5BjmVGEC
48cgrQGzPrUkRwyDTOxvQkbhH1L3jNokAvRYQxcLwNGEUk4OPUtEMzazGT3wtl6JItxUI9TvhJtI
z2eEpceplinR10jQaH5Rhnqv7edQomww1tgq/c4lt6ZbfShop9qQCz92bAkBOKeG9Nqj+t4YrjI3
Xh2WoK/aXQ35cLGBlMW2r6nbLSrKr6s4gNYSo2YglSLi9E/KtHZxr4CcZ/AD9Cngllj9BXmtQqxU
/fd0wpz+vBHNkR89jSWNvSxVT+7cvLJo+PuJVn21ctf27R9iNgkGgRIrNjIHsMsYBvbguSOSO4C6
pRrFhcskons/DZB+ofCnKsTjn7iOI7XKOPTZ671/C+gVB6w+sB3Z+w++hX2gesNRMPV7SL676wHW
2RyAWh3Vsm2T9gscfVKILjC87+mEUb5jG0TtfqVsq3IeocbnOxKo7q/352tD9I4i2us1ehJRQjv3
n0DBt+ExDWtFP7TFJj+3vahycCsXjolkbAOJV9SuoYHShoUsNlr7EcpCJpDnCpEC4TldDcZIL0Lb
QJAnu4cZ8HZIgqz9C6DVMOwj1pziaYldmaiGPewWDTmzaYoAu/Zvgh35xKZM0EsSqW90PO2ZZCG/
QwpWAKNkZK5t7wZfOB/mfuH2Yqf/1ubonVBRZDYonAjyksZG+QyYuXjrUD9PhQoktxi0E/aN4m+E
+k5SQhbD2uf8guB8WeKf2BDgqz6+xtDKW+9NfjYgaPthe3A4JpyLU4eO5blUd30LdtmGCi8p2XJ5
s9IZBu5W3pHD56iHQ2hVJD2mYhDx06oOf08mS8a3gM9pdgTMtt1BL5gZhzXq0lhMN/PWmgGyKlPD
pAgql/22qfnaKiTdLjyrH8dLlns/dVCfoQ5A+bk5muI2iXnewnKc/oE0qFemSnKsTeCpD5BGE3De
CJrVUj5OtXMLcR0EfdzkoR/XXqIWEFArAHtMSybGvqUbdV3S5W/TwqBRpa3wjnGJu39pZ9SJi7kW
OlZpv3xsVodciFKUew/0iCGvxH4pAmP4bOEKCthDOfaaqj+OxUVJv7CkvygsPSvfY73lqzyHbNGB
rpEdgz7ALSqEAoD/D4u4d2pLBT5yePoKFBY62lnBxIqhozO72h7XJdcO9rxRC2sXomvQh7lz4p2b
JVeJyas+cXvp2ixRSDuwq8BOo12QqZSkTTpjdNmwLuEqI1lRuUH2Eefk2/N6UbA/CfWiAHdI6BtF
d8g/eZRdvJtz/L0scHQarDjJZyNEIKvP+j6aaF0jaGm/u6uj39pXGNGx87HFNOW0Ec5/QOq7/nin
OMUFSybZ1ly8SFwGWSKVxpmb8KGFvDiJAHSX2Buv2SX2+7Qu8LCLW0iFMCZKuabdOI6KNXP3t+Ox
fmHgHndWIu1Xmj1m+YzjhH1ft0czjjNjUdNJNOUIA/gxFhP2Dn1ZJhJU+9iuEiW8XBnuPgjmAOpV
jysf+V7Y5TtdBQI3/vDeXnoo1K3qiv4BMIbbpUo2+z1SZLhSgay3uhxELaLRfJn9g9GPUSx3QqFX
XASCFX90ApyT8QZzGLZ2Qq1nmcsxjyagfbru42wY3l6czRsR3t0DjIAAOQZSG87e9x4m17DbjRfm
Q8rRCspZVwaMOT4cyVAVGOBy64DsORn2vb/5XlPw/K2A6F4JgouI/wSHdljNnk0Gb7CjvvZN55+w
XOSSzg7rA7ZQcHQBghhLdEStymCxe1/KSVXWUSS7r43nV4/3g7w7c5+NhYyBu94j6DaSXyDR0rvT
H3WYshpjVsiQUFBEqxC1ldFcINnlzeNaJdw/JnMzgmc6aguIEt2vkM20WmnmkDdgT2soTAZ1Wi7R
gByTUp5jT5lY0FTLYM90fgvvkKrI2Laj+vvTw9bpBNfzfFmAXRAuEVCaNmoR2TQ1DChD8yIVA/ZW
wz8hIYxm0N/Zocr+7G+7bxeHui5XPRoJRwH2zORQqApkBLbdeTSBpwpFwrXp358dJ2pevJk/RVFK
8BakoLKW7mq5r8Wzhwp3dabDIpolodgMlZOHW90shvhupQ9bauaPPv/aeRoQGg86w4Zb/LJTdcOo
Y9a91rYjRIqeS2VHPbJThI7qRr06OxrEs12KAng859kcYNsai9w+126DMLicKuWz65m3qPDHvNwb
Tbtxv9mgXJ/S5ROU9bsa8/wcSVtMkvM0/bHwM2IFJvl4RvXJr3u++l4BZrhZSTix5ICL2z22Zrxi
QH3SdzOHzH8VZkXRdlYwu1JlQZ2ZF3Y6dLlh/Ck2dftfUpZ31gNpx/WB330K+Rq3EBGHUdfgslR9
AoDZW/NltIMvY4u8wNBpNpM2xI2QIqNSk5+YCMDPW6IWqflcXidH0S7K8OD+pQjXvrGBJdryBdKW
anJP8eMg6n9SIBwWy1QmCP63zt4qgBWP36nYjOD9NdKEK0dL55wtZnq+98tkSGopaJQVHnwp6hOE
muiPkPr4A83oNdBi+sl8mDfOW7ltTRzl3/QiA41ZthuOZP5bwZfVnawtLvmD+q/Fd++WjWGQ0QkM
Uf/FkQxmHxsUt6C8IU9/eQezMVzpGwJU9b6N680TeI2bqvmzgO35jzk+IOm2KxLv19Si+Juy7vxA
K7uxW9dUudha+2WM7b+wVdOUR/UJlzN0v0ahIZGic3GwxgPEZxPHCGtDMtBKfvDGg202BgVzu5Se
z+f0jKfyF3wIMwZoy/uItsn1iWSOJUhHgtW7iJBuTFFZXEi9o+3YcUNt77Nq/FRLNkqAx138o+FW
P2X1F5nfM12JZDwzJADES1XxicUhHzDZsLwltWm8IQKJzQ4aSwEUGClHFV6vyDiexgzL6q7WE/hn
1TtHGMYxex63d4+aKJi1EUKhPfAnE8h5vwWZf7xzHDubKWnKn1DLDFXVbe9ROu0Qdtjy1vkv8+lR
p2IPTOpLIjh2kwTALUB+ipasChoYgkW7+KHpInufDTRmJPdKiVSF6pW7ARunS+lekm0dKPbz9SyV
3ENxThH3OCyV90EyF39bzb1pu94RPrVhrsf5ieGYe7xO8bLHhqKva8F6N7t+9fA6DRt5sbTm4+VN
By/VL0VoECz+VR8wZ+GSr+2rbF0mYb4Ks8bjiug8mWn+UDC057v4otq5XdTOToNpkx/LefUmcz0J
5q2DIpRlCUHEIZYUHUXgmc9yvDgCsYypgQ+xLiV5LMTneXDI/obaqImHdqphL1+VhfKrMU7t4+ud
RvXK6hpoqhzxYcMZzpjra7SaIqjHM4NZqlFl1HlW2pRfFwxujFxmQN51PtbIiMTu9wf8xmhykEWz
P9nN3gPHrE1bj+li7Xta/tIr6yxofMovqd2WKn0GSkgztuPXvMrcWNvrqcPHRDZP3HbwOa3/PzqV
xGv+hrw5F9IKYipc7zcVK+m8NX9yo0cRAj8NeuHei5WYxZmJmUO7Pnb73iRPNdskVTxP18ntDSOK
SZ1wWYx6zSC+BmZE+ox442cLdGACa1t4EXmGswO3Ln4Zn60S8mYA4hutVNkGEWplDZzuKPpdhG/S
orFdeKfn6bQSbrHRLUZK35pU6qE+nvY2VZ/2tQCX9QMAjjERyS8NKJeVYbX/2Lh3i/4L8jQACOLc
sd/GK66ZbvVhVJXZypB8wpbIoNQHZO2k5Gm9kv+xvyNudNA4gTUKzCakF6EdOV7WEg/y+EHXSeUG
ecXFuyJ1FcUt3yYgHW+6lFg4xlQ8DxpeYtmGG6a3wi10hX5eaoY5OjLdI8+HDaEsvcA4oZxnhIEP
ZnNMquIw5vUgBgnsWy88X1d7CWxuxteEPOs9KwgvzEvisQ0Ar/7XBKX/zNAdIel1xLyYRELObqwa
0PZNiKFQmKx7uE1zp0C9CKN9T2LlmqFiYXURH3ZxV/hniv6PSyQ5iUwgbzHE6pKoqi3s677R1tcG
h40NT86U4gq6Ggz0qmX6dSBJkqtBm2xYCf9IncWZTKn2ZrI7puYNHZ/iQIDm0BiIIp2eQjlzvOvy
3HDIRcyXhJphvs0MiWkzYLPjqh9Buv7Z8LLIIRWytmuKA+dTHoqz0qWbuQ5fbi/6WOczjSpWFC4T
VYkTFhOJcsk8AV+rdAeJQ9CTkbsrjKkhSzN+XVXvZAHmUS4YssKkqSdwK3g7H9jlgZ9N587+eDjJ
KfYra9BIzijZryE36Z3FOQuWp/tXAb07gsMoNl4hF7rN44APypGWZ7XW12zFH1A6h9sCk6obtYxK
mwPXvuf5Zb2OQQamZDS0hs8eskTDS/5tb3QWlsEuLCgVqwOXXKxkBDLcjsullAJ4ehqRMof5nuK/
GTcl/0p5xSehe8WVceOrOvzKsiX9/RDqAWz9xniGBoRnjKWn9ifhlvhcILftfQkYoDXNFQVjyA2r
OwpwD2dW4xCsxUp5FvRdzKY1/wiiv1mFLi+GILi4xPuImlvWkhrDJKokHMjb7bm3dwtkHPdvWMA8
Sgop8lgfhyY3cVC+aeh2ev801AavzZW5yH7F2Oevu4V33B/7dwCfsVt7sao3pQdd1cDL7Q7tVc/c
x1tpn/ezXXMx5logqAuzTPdd2nO2CUyKWTVdJvOoxM8fb86dVdUJ9u0WxcMljmnEsr90vL5EcBKx
Oz5MEWaD27JT8ukHp9t75WNOnE5Ei7rQoiNFrJv9NDhl7pEoMAZ11WgzQvjDGW8AyN6CMV1Sj0HI
gJTtQ2y/tI5E0m+Zj5U5e2mZt1wWg2oHDR1I93zrQYIQKfnCyPau1KqyMgs1RbRYvVqFspYml9YK
nq77tWbqR4yTo2VTgIGlpBkNBLAFrNemUZuI46EK69pdwcpHZDS1qutPTRCfvLCNpZ8T00j9c8gG
cUqD1MLy+GRpwO2Apg1MVjcQfZk0eUczoWXR8cq6yfQoFBoEFJogo1oRq1xINGUZw4N7Xb4vVSEU
/ebECJNGhO+i5/V+uAoAlqAoha1aD5VqhvjPBwzMRHT6RQ/bnXkFXG13bTM06MyMpS3m0DduL6YX
k1KjDFusYANnBMicXayTBYOH3z9oa2nXFzCucZZnJSOzm0Z60W//6vLPeY0TYzn3vS/4LL/UJLJE
8UL+8sQsDfks1tUtvgib5PAywop2eNYNbmMknI4dC1Me6MhmQ/wwKTJb22Z3unEgC7qo++IkOXMF
TjBXz1U0ucPy/dYLRGrzWBkgZxC5+er89pmaFh7LHZUJCmVSZwVIr/0KkK9kc6U/LKCVSSUMzMuL
hSdo0JNNrnYGx78VwVQI/ez45oX/kA/lm/1bAEuTgCtqXvSUDcPdHBlXXrFtpLU7Jjum1w/j9sfs
OaMXYGkvupDqp2gTE7nadUQRLg0tt7BjzvYBsnG82U3ECHudBF1g4Ofy7rwryPt8IO40pziDP52S
vpmPVAMGbPKl5gVa747Ih7C8T7iwBwVMoV75m1RzTzJGmfe+t7vre4XsBKENt6FDGRPyeP1T66kM
MyziMYgvdHsXHXegRGYmRK1qPIxElz+WNeR57Xk6a6+AxaRQI5BypuTDBQq1teFJhtprrKd6DMh5
bA5/6eJlcjd323962+yl6od93bMgJME6/6dPHkEZ6yRCYp7qQHDsixms61U/CSmoTzeEcFZLWQt+
oa07Qfpbeau0uH0PxeXhkK3mMggvk+7j/Uexlcl7ONydXvknZxYiqJA0/WHpDEcxBBFg6H6R3xq3
hcmuOGkpRCon06UK2qpD8X1lwnfLjQIQkqk55M6w8cDiG/3LZtcSxEa8L6R8DmTuqadymFgbGKVs
luRBn5h8l7T7KiNxSS7SeAK3qaFNgFD6FwPpNtK94cu455d7nS4lXDvRxz68i544HjVZoS9aAlFS
jsq8tgW8MY/Q7qKDHhjfCHGdyj0ni+7RH6fPkYuND5VfupMHxbSZ8U2vD8fbAJ5A51EGi/nHsu4O
hYKCVgYlQHqgUL9FrwdLp6q7MI9N4g6t393mCBJzX90JEIDrg9zXQ0O58mhxHTBtX5WwitrwuEY/
QAnHo2M6BWiGHgD7fvyqmRSUV/aBbzu1aaB5KGpx4twgAtBO7TH0qjokWztMD+ozDV09rOCq9RPa
yV+NGko2ZAig6E/hCDOLl1bjJw1al2rj/t0pqH+ZaeWEYegltgIrxkrwx7AfHfMj36+h80GLtkzQ
L051S4Wu9IvvQaL44EMqseF3qoLSu6H6Cw/ttd3L/28vr+EG5c2lFuer2Kp6RADadjk2kFZT+biZ
3i8f7IbBo8C4exRiP1ndtGnStWhr6FZ84wFIGvimxcqNLS1kLJL02kocpdiRo/dlIrdafGwsGWNh
8AcaG0YEJW8M1YI4zUoZCXRIcVgzXM33Cu5UtkdvwsBfJbeWjHRfs3KXglGthgj/fc6Svb1Nt92T
1a8NiJMG5u/D4kwOENcmJ+ZS4YG7FjHXG1/7YG1Z/q1uGIwZqa6rCo+hE4OUjQuwgydYuzZV6Dv5
aPip8lJSnmVp28jTd8mk/xB3WgqwpOkpj1eSWRi2BspRO3k2Vk9YKDhqafmQ2iVhfU8TgtSBXvFF
ozfjtBVhPYQNzXu6zmfFPnXkkE8Xcexnmpo8PZub93ngiokcuXSHBLVcoJGiE3h2Gz7jt+y7TiKR
02eBWx2PakKiNBrwcYA1HANBQKbXrjPQoZNpMc0/Lq8eyciIOu5FTu0A34Cr0ToPL/a5p32hpaxk
aIF97yTtugWuKJJu4uCDd/UZjbgFDQDy98Br1jhcFsUHZy3DlLeQFfaJyRb5AhxBlwSVLBl7hBor
ivsE4aQ0J6JcT2ohZB6sRBZus2w332cFz93rqR3wPtVIpkLa20M5HQqcDrwnabTAqDmIySeHenz1
H0uTlsAplAG7y4kGZGxmebwlIjLU6LHFzrHy+TndbQbPbyYhwhTCiHQ0JC8p9ZWy4PBvoVEi7d9H
C37zIr6tj4UX8Ci+bqPOQTRv7kx/ZbPgreVOKeJya5qyja2qcLiO/SgdV6XT0uY/ws8Yiu3TXMfV
v0/qDyyL1+1kx6ENCEqGCsCSQrL9vKsXlAMtTeA/nMfqtBpwqnIRv9GGCu/6fIUJNNn4z7dsCBQ+
mNOIu607+XClr+vuBvKliVcIRo4GgKaZ89+78uVQlviDfZWJeumU3WFHAnccdD0k0xh5Kz9BOq4x
lPSX1T+CRF1bS1/VQ47P6yyxPe7299fS+OrZiusR//i0eBSILhZPPq6lZeB4c3kQhqW2Yt6bjuUJ
2V3o3hwk5WSvtz/WaXCAyVcHdbFk8FJ61AFQ9+aM9Ur8nucGAsxuAibYG9XVxw1ghXEs5vaHc/SB
q2zRdPNUtqRL6yZtKXSIpoY3uoDvsEgwTMrjC05cF+T0cnOKP2Rm+IPby22Na8rIAK19VEU3+YFE
GThdKQyGc0tkUK/rs8T2LyYFpiA6ASOw4XwpTSWCJx1sd9vWlUzuAaz3hWAeyN6Z3n975ahS4oJl
fPDKaWwCZpdwKdvMTKY53UTh+5EdrSxb0VgyN3j7wAw9J4vkVJfG7cKsjiLNe5ytDQzs490+lgf7
qagpzeQeINTbW6qj5PjVFJcEyba/u0DH3fHWKgWao81oILEUIs7AluR3tVBzduEpe3kU/HV8cK7+
hSvLu+Op3wISFcY9DjpgnYgWNcfUMNI/eRwol4JJJFWYHTr5Yc1/msZODQuse0AIAzSPS4NR/CiZ
rnqGzT9iOCi0rXYJdy4I+28y0KMpdlfxz9AEcUWR/w7xX/R2ArQHBBZHVhZBSgODlo6jZp5AboZM
DPpxrGbl2kGzPld5rzk9uDYLAI/mKWUZ1hYycJIQ2eREGzAN50JWjkzyQgIynI+W8BdpHzBAiWg2
jv7KIq2Ddo0q+q/+onJNGE1bpXNfIbROw847adoa2Kv6AIjbEBAGjrzlPHbCrrw/eyyiDShlJamJ
3rfBSZTxZmUtX3XVOJMcsZZ0IaItgzNH3ZBQiUnFaA0lLiETUDG1JdDQPP3chxunFwA/2Udimc0t
EtpXSsU8k6dHzZTsemxvV+GmAXL9VKXLrGT3J3R2Hitb1o5s9JceP1mQteIKtsksnfq1RzS4+O3p
rHXqn76nLXCXAKL2R16ZFaE5FppxWK++zPXrSIOou/f9BhsEaSoaIYsDB+GsX8JS2IKl0bP3vedH
1/AmTvC6I/SSBPUeyua/92orRNdzY1zr7sMwFXl2hk1+TR/pW+Bjj5uvM4JsdcpxweY+1IwTTTh4
+NXLz7vCOWngnqGBMcD/QwCADkggYY/ffwd/PAXhb/RFsit/s5APLIeFJW9JUdnJ2V1qtbIjRguj
SNLKoKmjPbfFMGuughNgoLDu7hknwSfytQ+FUdMucrdmeoj3cRPoxJvEG8KxrhjmHeBKKeT0aAky
cRRYJUomMByZL8MWzXLofGQ5iOUe5G48R1w4JOxvsx2olMXCVP+e3q26QYXVfxHRJc60K1k4jaPX
z0DrA9GxFo5obFq5WeXMBWnj/V+hJ6FpW40Lclebjbzv8ZlkGE4HDQZDupiEUSLpd7YsHSpYLsxs
fmVc6iMVRjEW/p0ZwBG8W66LfixzIAt0N78pO8QlfWumLv83FSKHWaOP5nhA3HEhxmpQFWQyGQQa
ElwWn7bxAaxHYVTCfu6rEHslSa2OZboZDY/ONGdfwBz7Owzf4fQZmcMh3un0+fD83guZWmxot/ov
aCqZVE8NovpYP4h0pmPDNhHyVNShEfK4f9JPrneFjvzcPLd6umT7CyLEwSgSYT/4FnutAtdBMBxU
rJLLSgUhhiBtF2qEaHn+ulwHeOY5ApMXYwOq4/JiKTZvkJGv4yPaw7GhAYRdEkkhMyApjUJs9xvP
ZjeNpuAjuRJhpkL4gpu74aMan+alePwxeAGLR55DkqVYGdsYTaLnGzFn2csS/9gknuA7I5wLvVfH
rtrJQKYyh7vU4Acp04/D/mZol42rGXoNS67/A5u0riwIidc++F+C6n7InD3Fvy8O8Ovr2p/km6m2
kFyWS5X/YyTzXV7hckuWzFNk/msNLMxX6z/HE60asNs56qdJ+b9PQY/JievBAmGqZ8RcRZX8OiJU
Nf7x7vITGMf7UPdbJLbyBv0J8vK9wAmpDcfJNRPkn4rqradA3LodtMCOaoZiaHDd+A9229cc7VRA
wLOloVt8VnL77cOCOT0Vb3TSYRkapTnGAzajdEktxECmFowllnniCyZeg2fg7DhteMaCl8SzRAs3
haBe0vFPU/SYDG5hs4uTYvsHzWZGLrPhlsmPfU7+xYfduymbkNe4gaTkrv9xzhiiwLIyUVmjf8LJ
ePVTVHAQ/nrtnTD7t3FeVCMw85vxgW3PUe5W6SdC5aXAQd4UvUi952uFbONCWOQP3ByUbtIoG5Xl
AIr2qt3bwa592d0V+PqnDOExC7x1ScGpTzEC6UWkHu98x7Mfzn+4N+MrimyG2Hkq0KaYEB/ymepI
TJ+876YImwzqaNJatAd7ACtyn5lpdKbc+e96eg+f8zBxGP96OchjD0+ORvPaApZZjG59xtHA3XfT
M5vRAf9AfniDDounTMIbTOtAKIi+sIJqS2a3dO5wU5t4ME48jEEEX1o3kTXF1lErv3Qc+I9QA2p7
qKn3pFwZT8vSfF/b0PWsSYI+wJnROkCGlDUpinuRMglxa5kXD9YsoQGFrxEHv0F7aOH9NP7sNkkm
1bSr/6cskFFFcUZM2BLpimdqGN6EUV+LDxKJzjNt/q9D/diEIubjt49rAtIoideLwMnFMpBCuH17
JeqiSnLEDCfNiVhQlN6yVXDSHxbR148FX8uU7NCUrXT5RUDUD8i7ckvYxcgqD40SN/SIKUX/FRAT
KeEdME99rdV58bpMg4/Kz/hQkretqF8eGqL/+EkswJQNnW7v/D+kZDHoDP/QIihD3pc2Yrtkdkf8
rOkcgjxh6PXiOg6iv4NeusYDW59lmFMZciO9GyZmPbwSUsUoCLSoM8v2fvm/YKEUisdF8CstzC7z
h1426K6JuByUIM+pIZ6REcYkU1ioLLa4HPUC3u4lXWPTIyr4LCAxErVxFUFHES+yEfG6UwnzQArZ
D+QCYuj86LaklmkYUcGnCxhpjQmiIs/MVkD6Lbg7+R7bA/Zun5TWKT0eHKsvXPCvGpSQVJTzHPxI
kc27bOdGbP7zVGuh/xeEHVFPwvdAfCO3xz2XLaViodry0sk00YGLSXDi37eC+kAN4vR2lbWjevYc
WmWmM6coOOa8E8TYgx8LKqjtCv332CgPuIOVZwVcakw2FtgjlbFybGkgI1V8Ai7X9Hkav5/lByzY
cjQxXHo53N3KvqUlY50Cs+Jh+DPNJWzoG+A0jZDyLscImGbRmGP9g/oxswqYtpCA0qaTtQKgVeHK
t2aStiR/SV4e3k5GHGyryqaTd+0Euy48SnM+k4p9qcdNeFdhSt5VR+9CNfWvxlcnLrw6E09xR0R5
vxCF8uWT3hWPrEm0WoGf9CimeRCqA2F2Ps1kfOb6gLZplM86taUE3x4HgXzRZRdha26+6SH6TkwM
Qn2YIaJRopKZe1Ucffrw92oGKR/uDYWLmg7oe2S7xOY6OIvp5SPoyFHA+dyAfCijc/mGrzeaDmkT
m1y0DF9SnwoUU/0H5JszMFUhcHwt5Ji643QBYXU0aePFImn0ifQFphH+uRFmGyVidClBDxNyyMke
bidNZmrMECuBAF7+uFdVvxosj4mA7GuPGGggS4aK5W+cUmXzBHd52RyJHQ1hWWChNj6ARBeeEmaK
3hFIt5xHWsSuBtd5BbetG5qkDQ695u8pU0g42FQwcDG6nrT1OeFb1iKz7KJqi+oF/kCY5QSDijIU
uM95q7GjiWz8twPsISWk9wfEHWWLmpzyEaeOY2lrCoxklA5G9r1+vmz4jFYWtpzZCP+jPvYAGCeV
sB0g9SHXW9zlXJ40AXBWDVfsKDKkfDf0noYLQ1utC7N7K3HpUY7hSGdfbCihmGsc0XXk0ijJWlUY
ddD/5Fhjmj+rNIMRFCyjz4T8kbfZ3pbNtXxRzbbDR11hBgARAzq8CdlCKAFKcjFcXFeR0T8ipvPl
Mmedjjptl2TQB4T0ajOaKIXo57bz+QG2TtIqKB25KyypSaZfKGzHLHe7a7oP+8rQufCh/8mUhEBb
84nObMdLPp8d9Y56hNTmysaT5D/9u4Q326SR0lRfnD3kdPOpkueOB4ZnXxKv8nRSdo8E4XHGGgPy
h2ezldwox4bknXXpNumbtSDxpGj80teHhuE6/93f7zaiFYgIzszrbFp94/9EuskvjG5yXrQMRptB
D7N1BWeNps70XUGusqRX+SME33Y68XNHVf/jU0gvkdT47YYPtHA1+rR89U7DHLMv9O3PwoMZjrE+
l/7ElbA19fEB3eRmFsZMMhlSijHBLtKXD6Qse+rTb00YEJZqfpgy0xZomkchEmy2q7gkmKuwP5wP
00poCfWYJPicevsFvLQeB98rzekhP+5YyLmkAZF3XrolUbNXcAHUqo2iMlIG8YOEEfkwX76YVC5f
DCCCOUlryQRgPzSC13WSPPIUjtYyovLKGmhU2eLNoLQlW7g1ebODUAYLWb4SHKTILVBb9Xd8K9x0
kmimUfvHAOGDjfA+LaVnlQUtHjAqqmJMVluxGn8pO/5Qaec9JDa1zZ032tI3OCLzFY6H9eFwwC61
o2mf7mTgcgpdi28wEONxleXAA/B1dEuJUkiIKPSg3MlRCQjRH5xioUabd6PJXr5O41y8PpEk2NPT
rUIoljwV9aOPMuEjRSm1rUHjQsURkX4HkvhuhMM0K6zdG9a+rZUl/qox0d4LTyOeWheoI1ps7Yvk
rX3zffsl1cVogtULJe6vie8/4IcPD5vl1u7fOtOF2VfZJGJhbk/udTLVaZj+LUb3vtBy2iHL/0oS
nZ+trPY9ORpeI3GJfypgKjvZhe1xdk9r1YCGE0gn7d7H6GGhHdJgP1qpLsCtErZ/vNNGNcTo9MdR
mnmzGCD55diO5oLOqEWysl7/pg8T30JXYRoM1FnXufks1WCdIq1NyIUw5+46MNznCZoro+0dTSKx
tLG1YKZX6rjimXV9WRsJe+0hU8eoUTFGk5X5ECp+6SU9IVF83S3u80fyAzf4B7FqoHzjhs21HUbZ
p5uxtydhcPqnbgMiJmyEJrugOVP0V2ykWjAOJpeAGS+AEzc2DnY1TXevGnNa3oCRTeeo941cWpGE
W4ZwImjNaHlRNM5dJawwaFN8cQ4xLfl8lfxgM50pXIsgGI7w/+k23YfUrP4opOdWhOtMETd2zb9s
tx86lfgWSk80qU1XktvGrimJcGEPqRaccBVKGSDwh6Lwxt7b4FeW8B49iYttb+CDvQwu4YSlMftO
iWS26WYjUBpFEt+xS1uPOO+lS79bmsHPanpQjUgbhYgJAamjKps/NHmioxepM/4Vcld7VqzkX/Sa
X+P87Ms6UVQAnGUB1P39v2Wfct43dCVgk1k4G/Mb2ZCtNjtL+NmdYpt1KKP1uCW4cEEERku7JTMT
mdzcWagbHOw0MBVLaSnZRGdvqgfnU208Yx3rDcQfULIpOk0b0sNJjbZT0NDR1oNHGQhFyK2nJEVq
ucKpFCIh0aZYVqdfCKBXhKvs5pC8W2ASb3tI5+T0dw4IjO1wOlTZqFJbItaC3DNU8jcv20UuccnT
203+yhCIjf9WAKROM5UWB6LKYJT43VTDHW6n0Etd4OCivEO2y3caJA3xWKH8FJCUWFOx7ZahSJPQ
Xk+A+sqRczaze+950rX44lB8vvZ5RjUVGhHgwwyibNbhHhDE0odKadhH6I/DTComdKLPX1WCh9O8
cCXQK/3nRFDQTakEc+QkpWwUdoo9d5CU90yyS+3XABtxIOG/Oqsy7ovTs58cUmW469EfsVTJ087B
FIqJlZt/nwMYGHhrYMZl/awbMjan0Gi4/X33lVn9Tz95GG/HSsQde/gAcV4ejxX6ftIme5fGkb8g
4IZng7hDrsgOXqzKep7owQPgy8HVXQ7EG6DKngC55phQpz45XwNEIUCEdtUu4X5v5XbmK49gm9Fe
WXHDu2guTW3mu7Y3BiVkqGD1NBEgx/XZQjELUmtcXwnIeFjJJsk/LKcARoMTNubWoKt+k2LxRvGk
clQ9snDPBxFfl0uW8K14TbZq954Z1WuXho7lZu8mVfN8U9efjO5XtL+N1L+aC7ow3tNX6SrIuDov
w8cT3opI0Jwe+ALboKdiEsi54Nmonh3YCIhX4CjJQto5HHiUB7/iNJU5H8ZQ5L+nWC7aZePVNjWc
lOJHg0l9iGuJ6Q8EvxDSusDQNYndvmPDCl6qRnKhTymsXBMArOiQlxdq0XgLMl1cmgOXz/J3sEFA
v+M5iD0HELO0kQUcOi9eBTtOs4eWwU7DcPljIth+9y2oxX0ZPhS1z2U/a21EA2J/f+Caeq7bBe5O
3lmUANqNnDr0R4WJe6PrS6QexmS7v+3g4D+H6UOUyAeivAsSgqh/VK0gwlBu9KMRtRss5hid8Jpc
nRbHAdYOpDNMy1pCuQ6JytW3SUC8/8MzvzSrOc/GGgCkPa1KpRkuusBw41FwgSOHqtw/q8PuDsd6
pbzDJbWJgeUAF1YA3mjo6G2KlyQKyX+83QmUsya/tPG3BzqPF/2mvfoTfs0ZFxKbgoF6Z3BS27mR
avIIQAHBrv/9s3arRez7VxsJ5uiOD0vLEZ2IveFPSbSKwDicPs6meQOakDt7M4DmpBuIMUvCJwqp
tk7FI56SUgR3YTUL+pfq2bY3/BvQrZSgFPvDYkHZtnIbxf6lab+aVHSCNs8pw8RyYzUFySsqTl4S
gb+zRSqb8DA4qS5KyH/a0Do6xXUZ9lVc7KtLE7KZgWyA4KKVssczv6A6Bfj27+UzkMwvn1yYaV7G
COhp7MsiUOeViLG2avDPczPxuwCBo0p06Xfr0Or5mL8KEQ3JbH4U3oZ16Fzlh6tbiRBc6RGNlrOu
OgLxsiIEsRKP7MZDY1rKlUE9YiXLzjHUvS3Wxd5tUfcRmJPYCge7gBHO8Hy6dl7B5zgAsCTK006m
FoP26Qu7itEEU0joSlSuVHJcE4htkB+XmyTwi+EF5YzMlM94SxrurcQ+5CKp5wYXIY47HS9nC0md
Y7vbwjkzcO8Cxzan72/8tn3QMXsncncU5YmB86xv7gtzk4A92eJWtNOcb8sR3e5ynDn0DPN860aE
MkV9HNatZlNs7aUn+5uE+E2D2esx0ffePrnt6+4V2uT5kXUWmyMABGiw3JOx6V3QMJH78hSFsUro
Q3JVFEqGemgDerKUZWaXIuQeFWecAKRc8A0ed64LxzI+ifoT/8KO7Owui0Xo002Zu78BAyQIQ4O4
/3OSDTk6w7k5CXZeV5ocHrXkllzhZLnelbhRxgU/YabTg+CeifbTwvtU3puovjIJKmU9ihoaJz/K
mUE9JvGcXGLKm0DspWYdgAinIS/Iz+0KuGl+5Q4p3c2ZL56ZhvBPJULPd8Ox3jqa/aBcbSqKDocq
8jk1mOv/XfE3GOaxIphUztAfmd6X9+YkjeeNJMdOZJ/ekKOUFdqbL3ShCLJijYs9ME2V8pxY4E+k
mcCJ2sA0NBEenq1QE9ShVidlFqMrTYouFc4kcISPQvEX9xHcs/f468l3qIWoWm6fejlPfrroRxEp
89XRNfllkdO94UFcrKiGGKerzlQjVDBzhzTz6sJDZ7BF3KII3gzi0Ny45quuKKlixLLE48IaLluy
othz4uixQ9714htX4DxsmFk81BkLuzV/cSrkw8goo6KiLvhYK4nHjKhwmiXGxtYhYHYdOpXfTR0u
8v4bTKt3zS6ttSqdCqhjVULwaPXNktfT+CMh/6nU0gS1nsMaKZBM+/OgbTGeuAsu7OP6G0jPtQ/e
/S5BJdCuR0WyMey0NaRTTfjybqrgOX5/2ivq+vtfLBywzJjqpLMdDjT211fis7irvUHQCzNx4Re5
zg1V/qlFa597sZy3r12AvYpzP4LEVYHew+0J4DxiuUDNH9LM/RceIcOxsRyXeISoSJUSBBrr71yR
3yUVb93/2G2vix1R6C3kLCYnLcDPRCE69n1zyh3SQ2X+NO7/MYihxYpdKeTLFRHQgZa+QLLpEo8j
T3rbb/hTha+IiY0r9uNfRYxxCvBLSV8NruhuUVGjRRlZV9wquqQe0Een6esRCHMbqDUlqYtX+rI2
jRftWj4JQs6C3Dy8EKCaub4OKtjgx2HMnyTxK67YQi/OBtAKKPP/sFRSSwKklxIKQv0fAx5irmoa
X8HGlq5BgnE7qEClNC3Zp2zZv9kilPYR+mwU/wQHp69G+TVfiJYZgBYHeGcRQtr9q8QFLf8vGQm5
H82hhxf46LeBgtKt30vTCBNxApA6csy9jxgbzOfBKXN6CXZYK+Y7tyNSTmZWBaV1FvmFnrIy6ThA
WNDy3lQ/K2IjKbNqMplBGcSvIRVzQFNZAf6vXkN/schlxkSoba3qOzt+3VTtg0yJfEDLnZPYcIXu
Oapzt1EJxw+ThKa84LuMFMeYNKlw4vNDJabhRmTFYvM9UAyPB7q4O3ZwRDeXp0ead5Khti8k6hHW
0jRbGwHI6sx955Kd0CgCZRytKxVEbyzMqv+zQGf62DNr6PL39SuSyksO3DLpWDgSmwlVL/9a7eTa
LCN8gazPQYd6x87htcvLDjHw+ZdLGlZ3WVg+Fb4TLuWzCt2wruAoErYUN2KUWKZ6ZR7d+7laZqt3
GVU3vfBTKoVnoYcXCp4xLNXhj3ao0bz8vnnKo2RfQBZ1ckzrBmmLxOJAR3lwZHUcvn5+1hU8zK0H
tASPH8QFtMMOOzytuXVtiBLh7lfwynYvO4B8QI8Yc8NautrXPuL/D/5IEHpodQz5iBG/DRQW7np3
YYkjgRqp75a0vAEjbzxntXb1B5bwIi48cHAmMAc5ZkSH7aCoSwdrUrVyQo7ek7hrFRqNjMI5AtmP
gMdiIbY47WgdjigRlPXAHoRdz2P6Bz9ehn4Q369Fpsc+vH3TMMy37LmA9Tsqe8EzjokhZT+awYaw
Qh2Jmzey1YuSjB49Zbuly9nZudDes0oXvQ/EBRve2O1k8+CDRUJQxMbSOl77ZGXC6melImUAlahx
yFKwSv0ZZ7O19zBfWp2AbXQd37yTYNw6nG34bEe8H9QwoXV0aB5C1/R2BuE0XvgkkBBijnNhNlSF
NBnOBwvrPJdJJ6YRWl6CkGwNqrSZSWf+A0vtsEQPc1nI6reu55J6yexxlQFdMETAF8fZBmh+nJYn
zpXMMYqaHI1U/utUrwCJxpPV1xZeU5p3gbBSw7ALlAduC1J7lrha/flooNe+NyGNfiKLzblkGRCW
rJyuUdUQqGTjXFo3OWPOVIuxZiuDnL9iIWZ8ndoTR65Vp4SQ3kW8x0Q+h2t6wzS2rZ4WsZccYDdY
BcSeWbUyT7IIfKDx3+Wlae7mNAuMDYQO3AKl+u0BCQ1yrw20otnxPGTRbGympvl9Cs+7/O/rbUqy
IhAvD3i0oL62tcxrUG2wgXamNipnpCekQBUN/x96Zcw7cVh4TcGrQRbjR3mOK2eokQ/En4nc+KkG
C/yFFvcJLqGDi0hlf0m2f5AXicOvc5I9k0V7qtvhY+O1BdNzsEVOOU64OoZR6rQJepLXobn0RyLN
JKLfQKCtMVsNNDtnOqs/ICwEWlJqVnMBZBQtTN2Id5D1rBePxjpPUAZ2hD2flsTfmC3+ti8ZCSFa
Q2GlXyNtHFKO3IlhaSqrg7mcwf+oHknEXI53ZcHGrzsYh6eSI8VhDnil2jvqj4FXp01UpZfnhnTW
9vEjuFXduPE8DlHgwqwhXqHtTgUQbL/VerTubEyxaJDw+ZyF3plWd98ezn84fe/JS1iKVdL+vuTh
xceLrFbkxLwMcGLhFB/XLbnrnSract06hRACG4R6VF/7gbkdS5WwpHXvhMltoDLbh/YioVydJoVl
eQNLSswDUUkhTLkKvkl/IJDEEXyZGpuW+Rv/qAFwYwl8fRAnR3e27ZvzlodNwpRsf9LLZlziIqwV
ALzxo5U5tGirhPV1xH1V1fqyPEvVf8CGO338hmgD8VDQO/Dq/7E3g5fhWg6Oq9AgjBMcS/ZYmy2P
iQ6u497fV8ZEIUsv8zd9p9w/2jxBU28qyPpcvyklEIMElQPwqujlWr4yFCDZCP+fVojTLLDILfNO
8trdIB3b7Sy2EjK4MQDYVPfvjh5+to0k0tEAHfpitX4B6RREEJDW2MbMr+5M7nHSwRAyRfBielDo
g5EiULjO5c1fikrkdj7Nq14v23dP1zSJTH/nbP4ne/VZXH0G3fbzC+g9CrqPG3uTb4DKnoGnp11M
bQK6R+R4NAdNPy/qNilA5k5oecxR87xvTXbg0HggeRVxmdf+r/sD+M5q8wy63aFCgxqIVQg6G9uX
I69Jl47sV5btOdwF6noGbbyvjx0uG52rrhVBiCrPqv1qb3wLNYrQvkbozZr/WZBaLgMMeIzP2zZ1
Y2KudCzigg2ao8dFDrpTtGsBqXgin0tLNUB81JTZHeAdJF1uHU5OEGwFodMwkyVdNxVGb+2TpAmP
ykMhw3hEKvbyqCfbpNVpQ4oeAaqw6aw+i0wIgnTBhIEjAzuZIwnVZiGFrMmrM4LdROlT2K2gc3Gu
HU3L1p4AP7pqoLNkEK6Ux+NwNdGzpH7x3ePmpo9Ape1mobAgcHzivB0vAUIMXXaqX5hVcvJGwIBY
71923qqHAwU+yHrM255oi1z7msSOEKXs6Ou9q8U0zbbXXQggRvWS4H+IkV/mw3QDpMllb7WJTTxk
1uHF2SiVQYdk7UgB2hbjZ7uYhOeNpK0WjxubSUWVOa597bemx8lw/Iu1wKujHf3iFcC7TdDEhc40
+iPqTgoY6xggQWgza38c6prtx7tqlW37Rb0OFmBxnWl8/Cf5Npq/XW1l5UgIYsDx25K6wz+XwrBP
cCAWdZeJRgeGfAYoioVB3fD76w9m5933RyT+0u/Fc++dOrXD8WhRGylyd0C/SNGLgTCl6TzbmZYL
nK355JH6OlkxW53hSyu0dfzdfNmMtFlT4a88w4UH4+7986Ypo9yshSsK3A6UGXG4sTiv9rSOM7Pz
FdXditzJ29E2H9fkOCcmHFD2kb9ciSTkYWYUuQ6fmRL9DpMqozce9rT53s1Rt3iElSQZkLminprN
JunLIgWoa7xQkrAdOnAJhA29sV+HUUOryH1L7biPbvx6rRGcXyWtJt2M22PJ2Yx4UqQyfljwpzIJ
uJNaJrdru4nFzkmxMtJzgqdqDnwhNO8ItDdE967gHEYXSIpggtFkpdfpwMrviKk7yi2WTJYoubdp
eyjM7mQRkJWM72aCVRIU9RPKk/RP68b3SSGsv4x/opyWLC1PfokCojhb2eqzuZlh8GmFqGgHsoUS
LB/a18py1cxhmxw20B1XDW7T9QRaOCb1ZRwAN0R0L9ZtgtXrg1KMzTCdkEyJV7wFIIPfScJ1EJcp
RWZW2IkskbyWlHinMnIqIPLuTkPJwQXsq9I0TjAcgPmzgM7sKkaPisj6vdYDan/4ugyoBaV0oHxV
/8KTxfSO1O+R1VWH80tBpd9j6hkKcLd8ElmIXoyu+Z87quVKYUWVY6doOS12djSvGaMvpflxSjTt
H7oqKar4s299WJMrF80kXgxHN3Jcneyv7xNqpL7bPA9/jnfCvDNUEghmHmQp8PQHrDv+k3WHgNos
3B+xeqQsXi5wiLvd6mvzmmG3MUIh8nfoE2iWug/wGv47usMxrL1eDMMy/yFo6JOdRMHnuuzCeL9m
iG+zx8HU8uhukGCanIV8NldOH0tPY44aJHCr1RhlEDABe95+WkbMxUu6ybK/u4VYHwPR1FIYjxrk
ZsAs60+pabggNEGykRplVLKk9oIpwBGZD1WdsJF2d9xjwZ+RtPq62OoSJdfTVNFUhkPqHgLDNULQ
U/J4ruLJvrTPAoPyOWXRp4Mq4gs5jaYAc0xnf5jaI322MRrVJcKCIlRIhFM+vcXuP9Mi0mjmHt30
1/3UvmRN4UzsuYzvHZAT9WjFQaS0yuXfXv/n2oIBXkQKYXloAE8aZ/00wS5i1GRBOiUwyql+YkQi
NzwE0KW0b7hC53WALafN91sRLj9mOKL8GfUmBYyorIL2zKMCcCgQTdam9/byiU21ARzS6odI4UeN
YSTZXMmwoyr1WWkZFZqy5V5qd/jp4yY4FiMjUnjQpSPLLyxtdjVx7jEePWcVrj05U58lSQQJDMeF
NYIE3/9WsF3WztKlhg8PlIAkltn9xxcA8NAqyu79swo9bR7v7pGIrJw0MBCK5vD3O2q9dSO0ytT3
iceOX/407WFFgxUsYXFX5uiij83vS1Q1iCP6DexIcW/Nw2hCBeeg1N90JNS89jBwUHVicvBeaMMg
UYH06Vm5V7fpECbAhchMI1e6l92LrZDmssDBOI4uKrsN3G8T1pS1F5MSAM2R7xCFvVDfnQxMdXhU
VEH/bg2Dmi0bOEH7Z0MiAm3kkaD1a9rJHmsDoUKwZao4KHtNAqAVaGy/G3rD8JNthCk4QGp51Knw
t4uA58xndRv/fFhJsaMqrICUK7glQxknkynSFxLBb47+RDP33MkzK/6txnFBLljkUN6QtjPJ/eSG
3aeETr9qYpjbz1h71MJVNFzxitC5I+sU/s7hQdtUzEHYfanN2veaL07NqeSCxnoZen0vS2rp7izX
s2fOPDOLvVtT8duLQ0bzfd2ngPelhAu2BIVxTnOlAnAIyHLxwBfNueaHjBL0GDaj2VGdGaCAuz4v
rNsy3ZgmD4BvY6tvhTgxnSGYbuXcdVZg3VgWbt2vsoh9wfakFw6A3gJQ/a/ULSJz45VOpVZXUtO0
4BZn4SwYjjix+XjVt6gYRzU8oKAmyklrIlJ5vLGfdAhDttZsB1Glltc8GgEUB8UWM9dIVU2rukjT
kQMGovq4j8L4m71BnOAaefkw7L9/c4j1Y3CUxewfbXBJxGFIvibTbWyBUtHq+JhXyIrXWL0iYXlS
6GMHMcQH4/yPOD2GeXH/4i8g16bvDKKOH9ErO+qrgQN2/CMCvUbza9CBz6JQBDwgqsA9rzf9N7B4
bTG9Fxj0rRXg3W3DYVlhW+Dqf+JwYF7d9tO8w6myRhIrCeRVCqL0hAoFd4KnUXj4WztoY0Xuw7YY
kQI2OL1b4Hwgygs+fp5/8rC4fSJADfWzlzBCgdY/Q9/TNkm6cLAigJ5VYJY/4CsiTEpvSg+fNNI1
HGcfJMwbNKEZ0eTToujBMDVRKt+SoApcXHN/HZnYXdEFQncTr6cvMO8H+sXEyHc41NF5WQyhoLwC
N8evU8CT/YoI/peF5G7sI1zPapqSqf4nanYP5vevLzIzQqDEBWhCureBmHOLAb+XYFELM2MdZ/wY
T5aIMxmHKHMjYYuSLAePovqjRdFDuM78OWzT62ADdl4OICIJETzOTVqulcqoH5B86uREptfggMol
EHr177ujgOz1xJ1ZGfk+IWskTLFWlRKlwZW7VsnqKQF17E9jNrwZyPlSzSsWrd/Y2eRz7B6B5eMd
hnGjYSLgEW7nc8SgSz1lm/ZHkSR08uKvnpF5KCIIlKPTZsCpmodk0OKYgIS/7g+g83xt9Vk6uL8p
b6dzVnZai9zbNsV/X1/bIDyLfupltp7Fwd+wA5KGjrWwWIt2CVxG8NVm1kfBR2F/bdArlEZ84pui
hi2fvPrMFB+I6kNawYheY49Ns3LND35dohZ6zUJhymdHUh77zleWwdN++9OfPru87nNCmaPv7FoU
OSbj4uJ1yiZ7o/fSNv8m55Y9zjPB9EKzzolNV8MS/YW3uQ5Tym2pOHjy0RE9du7myiwNTZxJDL1o
VpwpXNL+TvbOsvyHzxQOKu9hfNMAQkb/GFyI02Bc9TXsQv1q7+swEMHLLLVha9DPkEmq9fGMIrVN
Ftctyn9dJjl52sTFH/mMKpG3zaEZO517zbGJULC8K4L8VAE/e0FjzTNswZA/k8NETWQGfwvKBlKh
04q2rSX+buaWTE6cVY8LwhgmmASChlnVqXVzOvymKAjB4QGwh+sjwcq+KFR5UXo5mWb7bZoa3MPU
NU3MnhAuhCXz0eZPS1VZKEoP7Phg4SRcPDGGhNqpnwsG6wiHlTEZ9e6hmXQn9IbRqqfbKmjMbDmO
qxXlczwMhgC8oREzFkijZyaeAliE1ZQGalE0nt1fAOhCVDomG+HZUQR5FX0CCeo/hJhwHn6Q6EsG
cdrn03ltj/jlldQ3bR8kPh/dPrVlmMSHHxd2s3fxmd83GoKbyMm3EezVHZUOL+md8HbTSsDg0rxF
J8lUPBixZtdig7VBL2cRRuBL39/EXJuZSnvinSctcy5j/1dK5l1EgXF9hPs3GyPm9kW6aEdVh7hc
9Zj7DMAR90rfrh8dJr0FODzPADXvqmTPKdCLd39MKYzhvSjiQ4isam6tFb0Ja8MG2UmoMy7Hvlg9
7xidl0vbccuLkQ7/a/MMQ8KV1/fp72LbF0DHpR8FDnn94q0Kdk9vp7oW4XspJUgZaOfDFIfyGltR
5+bzK+NoIcK9GMevbA6m4yW15j3Pv07Usa53BBPrGytvib4SyCZd0Axt1EEe3bTrZHu8x0zeXVjI
Wqf2xVpItGAgQm9r5F9I4fN1wtt+PTbBlQJQubWQK+r4Tci2GZlY+ywc2k9LmfgDv4rc44lH+Hcv
m+VfnzVFXcBJI9Q2rk2dk0fYWeFqWVhM6mR7j+4k3qWlJ2Sq+otOS26tj+o5MGSJIX1ucJmaZqnB
9l536XLOtx7S53WKAM2SnwlhuOsqWnwAQ5rZPkiD1M9G/u2EINGqmnUgIrrpK9+jaMai713aNnHm
I9PRSWnPFQOEbp4eXV3Xb9ByGx/lFqhkmR8NeVKTXSXoKiOEtlEjeBU0GTDCV+/VAP2rgzibsEt8
0yLrvYf4B3PdLILta9fNemFTvRoOP6Ar3+A0Cy0e6WiqWHk64b87ix4qEmrMBK9zPn9PCk+F3bxQ
CsQf59xaGPNx/wvxqhetTmetvuZdrNIN4PmZMffvYjtosn8id7okIfbIT09vojfGmeA87DXjIUHB
8gjNfO+TvizvCcGrcvJM2l/HqRqbcs5sh2GLeeacK83Z8FwgWddMtsqZSsXGBS5hnqdXFAwtLsww
lQmioO80ZLsGjo1yRx1hi7vJRyicbVBGVObvCjoHyZ0UFowJJX9Twx/qqUXKjRaJf87uyYfgAxLL
FlHJdfVfXvc41Mpz9wMCOIwhxS7j90QurnR2aqNrNC54qMqgiKZqNxLMtzrL19DVQrhUQy3l2uyH
xjl7wRw9DBYXa6+c/JXXjD0bo33GrKC1FuESZ39FUVJVLTdlZnI9lppsQkHrKXarafM7j5HRIOlW
mcFUKi2lqPmFItR9XA/rDwDEzPr5SGJB8IeKDPBVXeNvNk+qD5Y/k0zgbOSvMi/ILLWmzntofFGx
esSPPk70oIrUudcYhXfKGtSVQRWka9Hbz2cjAhZIk2nRdwKuMvGX/MwWK28oEO4fqrmo3to5+NYB
FAb1iXQcg9S2lTPhMoS/vlt5boHqdnEMLa+xFqGpuS7lrQvgY+3mst+DG9i/XMvR/jMkqy+zqago
Cl1q4uFbjVr2EW/6Hueex29i+NAlhv8NFDWM2+QCnjEjjJOPDxyBvq4jU0wFUqDRegOYVgEECGOx
kxaimaby4Orq/yU2sy7uckjuLAILQVbFB1zKxzTF7GZPZCe9oxkZmLDcelM32xytZyy+fi/OI8Ci
KFEPOajDOTtb8ORBceYH2nGfEhA3SLpp2w/ocj/+dpoImQoc0Y53tZUZrvHI3/1zYAI8s5/ij+f9
guXHA+33Eixd7aqXI6hhUn7vyP3iWZxN/kMg9g52f0mSNx8p59nt5cL9w8+JU/v8mYdcQrj1/qUw
cqJyraj5+gMiGciJFTl5jbeIthEIQ9/m+iD3E5BEi2XID9guvzY5lorhzvMfX+aiO8A4sPiT3gXC
rTvHzUyA5QybzjqrTrS4bi0wfMw9/Im9HMuIM2dppC+iJ9YyrAwvzvng2kI6md8yVfC7bXG8evcn
CuPCWNzZtrmHQmDW0iuDxI4dTLF50A/A8WWTxR49VdOcfyLg5R1u7LFFglzZo4pF9zYm2HUX4j9H
XeUmKiWf5nnKFiljwqhQDQ2uHmMpNniZIIxyVjJKoJk4kY84gZVlpvpYjGZzjJOuxdLjV2xwjpn0
fDLtRxOamsRbxzT+fZLeywG3CL9rs6QerIvkTZgbA3qn+9lTCfCahSs7K6Ke+fSc+EL3c1uLNYMj
IzKO+StOJ8YCt7DsP+cnJtsZQArO4ziU5Oqr/3Fg32kKfgOnuNpITg1DgoYRV81GSJ292JtspEIh
RucpkEB7vBeYq8eRA3f3DXeQ2vIPUVyKBXIIgSzb6x9BtqlYvT7qqPnaaMsCiuXjU0y566nAd6n2
+87w92QVYeiqTVP03HIcETvIlQCAaEMftaJ3PIJ7QtA6m0jUgLKZZdlR4iHoKqISGPfqpvByKzWn
WLRWoQT5UrDirqEgX47z5CI9tY33QZkd2D/6PERopo4rk5P6PTuv2XgRt1OR6bIvSg8AoqrJdjWQ
L2QDWIJ6b971JTlqx4q2vtIJrHpyLaoo53aUx8gzXXVBgjY0Zgs7Kepd4Vi2oVSSn3EzY/cWtIyq
iXLK1VlgG3LxYLha4U1l7RHtqKI9lYb6ccpw18Q6fbz4g6vIMtbmzxoApTr21uFenNYOpJE1OUJ9
Wk6tcKIwdKigdQWQztu2jp2DuVXKO3Ltc0bpxK6PaRlqaj2HGr6otC3XfuVTl1TcIwzVmyvi2iJM
ooouHglnGSkBlHnrpk+9l1HzdrT6Nvg0ujDpNWcvmPIGzQzFwumWgUwCqaNE82LAaT3uqH8OnADn
eUEO3tuTqHiRetMdbQalomFgLs6+nO3pqZkiNbe8nEscWrUZAd1KDHFGnKY0eKK8d7vh4ncsh16V
U7+Ia9X9gQCgYjP9Pxx9SttmavK++4YBVsY4+QQ1eAR/Q6l17Xc3HmNkv17JRZyt2B1vH2mZoynm
w+mN44TaAc6ApEjPqPrPvA8gxzm2cgaRMjsB6byaSToixgn8iK25SuZl+9KkjYPl0jN7tIPQDat7
JlMmi+umq0+0PmLzVzxTMgikYQsqwznHVKHyXWtl++SxwddXvHXm8OsT+PUya8QcGR+z2nAg/KxS
ArP/GBznssz31ZcFOExh19LxrrGCQnBtQF6C+0S/uSo18rzCYbG921EIO5qFqV0hPxpjQbNXTIG7
mzXBMuXLPQkwKcsRKyyVWvNf5pkJYCi0Y0kRRBgfRnXHef6QA+koF+TadNKrckS1u+4KH+oGJxD7
heN6L6UtBijHSYu2RclzzohQASCd2pmJVnTj7z5HMG35r6Qu2nCcojm2bpu+mHGJOUQJyVbytqCS
wKEXDaRv3iPk3ZyahuNrzaOUTMr6iFTR4Bplo3vIIkgibiCc7af8NWjOokJP9ESTrOZSlIPTPRDG
l0tObQeGo9O/t8mYoICVr54z0JafXSojWfWFAYrsAX1N+KJkZfEvXjGFlvMAxH0zZNtDTc1Z2AW+
/sPRLs5PhhnVB4t7V5wRr9h/5BEZLAkx4dvpMf5l0OAvw1hijrP4Aap2wXg4Pz3Z/zdyOrPv8hy4
ftlZnhMWkfBf4OYUyRoDWrV6o8V68Fu3dv6rGf+tevWKMcHbQROd2Nj79T+OA+Da8DH55OjeDP3m
MpQAFIdZd1W7PEDG6FWFJynovLZTqfFZOwz4j3AUeCnrBElNQ2d/yKm9rwSSXmHPlrCTCg+3bs1X
YTZQJgTkdR4rFnODCGjn51tuS/3XXIfs0sYwEI87bYCPk/UT52Ju3I1J31M2cq80qUsrsd8rst1p
bMkdYLTc5p4Pg/nIu1uShNHHHZaI5LEZJd4239aJy9Gp5bEd7XpUWoQCwI3xMy8aVIM7fXc5zFzH
f0kS5zAPYzy/p61pzFgLdrlntgtlZQxlf7KpDpnOQsAYynK0sRnQwwiM5uCBHDqgLlIIFuUXQYUl
Zf32u5qncliPi9bb6t+bObJcj+pVwPwaxahWbFf6NNsorzPP1vCUzDNDLPH4i7+jJ9yTcYv9+aoL
zslYbRhab0MjtQXhAUtSd1DN7Bwo4hI5FFlVkmVFgq2NpoCVMJgR832RAMreqUlMTooPQKaqDHnr
zU+3TPUl5Zw71vxA1o3Mfy6zQhiDMNFtUiY6Tm5vGAea5UkNj8LzSW5LzvwtEBM1lOFcQWJ+J1mH
tUhBiggds2/a0ZOknxbLs/cMpNcuoSljW/+Agd+SlmpAo/W8pe8iT1AWn5IZAVnIewP6YLaTMtHY
dsPlZYIdr1JvNoeaEHMWG9E5MrGthtaTJsWIWvdzqTV3ffK2Rhhl/+sClZLtzpiVSAui99ibADw7
Lzcka5aDiJyp1tj+FJZWsOT/j39MDkuXrhmJt2s7V9rHhEV0wAPLz57e+PytCjYiUnIxhoitQC0j
nFQBio8Kf9JVnr3r2o5TQHr6E/TtEul9+E6Vx4wcUBpMlyYQi6OY6Zcj2dx6xJ+tn71PtB4UfzM5
sjMVNwumLhdF1G2aEyEf0tJu5QpBdOxZSCyhxGq44pld5h7gWODe4j00w1nVBtlCHqj3RXNFDDnv
oTlTXmnpi6JhsoGLQEIE86t+tKe2YfQiR04wFEDsk5LX1VRdiFVWPtsstJZiXBG1tCc5xD4ZoB7p
tg84VED0qRFiTZORmEarCml4BMUH3hASvIv1/jl6kxWMV5xmSaxKjJod6x3Tz5/0tHBBTfzKmYsh
7CaMZKeIj6008KeaL5opi9QCeW8ijZW1oRz/eZWUTl280oCKgqMu5so1/gNJ+a/pTOdHS3ueE7OQ
XhYSjAOHjJvUeP04LJeH4jiGMTpSvr3dN1fqnDYwqz9l0aaStjdZJ+LUfF+aR/a9zKUZPN+/BpLz
IOy1eWUFuRI+z2eGXOp3Ov3PDEsN0/xvR+g301zMBYycKlc8cxHX6lOQti8JkKnSXgKN1Zvu+xZs
J9tu9qd5iQhl8ktKHGqtfCkbCyetk2XtpnOue+z55gytly+KhXQRwf+GND5E2UvX5TasFfydUfLa
UOx+o0fVUHLjYCWHZzkjGB8Uds/eggJnWZWIpS7SG8RkuSiuT8xD8izouCUWWJW0x7LJIMD2U1hO
8SNK/zs00178FjqfYgxO6kYnsFIEVHWn7um/zpAtS/rw2NcEpkjbtFUEYAqpY08fqq+0pMmOA2Hq
4RPfnubgezXkMuGXIm1Je7sU3W5o64OAdA5VA4kI1GZfWx+vOFGcKM2Obq2gJHkJJDIGsfWnfo8N
t5wRbmteseP7LtWXPZmxEczO2RqwolCcluqy/T2V8HAaos7q3xUuX6CURuYCPG/tY0A2Z/GCcaXc
ch08kM58fNVzjkjv7ryX1ktN2d6PbU8KY0D0vQnlEyNLnmAEyhZrkjgwmWu76+UHV9yjk9rYQ9xI
+LnnTrKB/N4JVdRr+otQGiI87lgH+hMD7kXvOs1N+4LjUbpkBAFCdNx9/TCHl5qBpZOwwUStIRk6
y0oFxcMUwwpZFZZ6zsdZESVhHJZLLXXeJwk417cZFBj+sgpIk/79SzEjl1wcEL/7uVoLEQm17m3w
FFRye6vyT1pUap9Spto6hMyKdxoWj1ID76L9GlEElKlPY5Fyw0GIkfvIHjTzP5i/TV/wMqmZFmy6
y5TBqyIBgGGOJosmJlEprRRoTFOyWM5hnZwYXXihDC1N2nkzQZ6xad9blxOU4SxnIs4t5gURh92l
l7O1Y0AWqUcsy2HCofdFuwf2sb1P8dSVtNNqr/BsSiR6MnlBC4UJ5ycIwLt/Ifm2bN4e44nfS7cD
mPdbFH1gishn0iarv3dgj46OXi/7iLSMIGCv/rBD7D8blJculxA+2nPhsoHFjerDYISkdkQ05lCl
eVQor160ZsVlBj1/UEt/0GaIWucn/wsUagqjLuhyXrxrO2LU0ShknRiTUULgJnwRKoilZVYeOooT
VOhFNsIUkDGlRiqBMGOPLmOauZQgS0iEl5wo93FoCGTOrl87Yv/7zq/g+T8RNrqf36BkSrEMQj6N
hJmaWKZq9DV1t1wl0uaH31rtTOIIOwAdTFu1jqf62kI3VCJj32JVERknRyqXuSyjURae3WJcf3Ub
EM3JpblBqDABLk8eJ6VYlDNgBsYMNcwdixkCxKI+ussjAR7vDoCDZl4mI7YJO4h1gOO7BPwniHmA
xwUZeFwmY82PRbSUMG5ITzWErPNSGvyYKzj8Tl2Eg+QhDAdGmJ5gkQ4G/zeJ8xbNOuKJRiwQDjY5
OrbOeKEdxGn3vjpwbP/biyO+FJcIglRH8/cJsUY3zX6LVq4K131ZQw8aLU+59n6vPROO+uplW2UU
1+LuAwwiiO0f3YTtjOKw0mi9aw7U1bPI4dQNUBFHkrfyuwyN6v81kFRa7Yi2hW6z3mYWw8XY9HJs
5Ha6TLB50DqihH01I9/TWgq5pz4lXXnWhQpuTNGyGPc1utCXRCXPp0VwgpGddLpCltxkgZ52Ih6c
cqN/ClEoVqxhf70ePD0z8pc0y7wKVpSv07ZR5CCkvASZAIel20V8eEGcpBDy/OZYnu5airPotLt3
p3K8YZS/wlCy3b50N0ewBULGKIYk7GG2MGsXmPviBRvtjajTjWR/iKkA74bfW/6gIbLhl5jw/TN9
tw/6UBo+B53HM1uHmRnT+qrDIggduMKJdd+NDEuChaVjt6Y3RxKqj3RasJH1CJJEczCtQUlaHXXT
8TuHTJfSZgCwFuFH/tjVzdkJDGdlfvC+ENgnknlV/KomW0ZR1zuHt+lfaCNqf45A99BJQnDaFAVb
NLrf3AZhPS581gxh6RGkSeH4UTR1zP9F93Jq5pb/RUT8eXy7PlDtex0re/tREad0725hkj915LhS
2MvNUObACy8aHkYsDzYtcvepmi5jPivItvlSTHRV5x0lHaPiDgnbzqYwued2by4+d5jlI0lafP9k
mIo6u/Brh1m5bgUQoTbXGtNJyry/rrNlP+6/HyaSl94egJ7lvP4rcmEb0AotZWEV5O+/HKpUcixJ
v5agD6O4Ai4PuP4bKHqk9ebdA+6HhsteizoFPsNHNY4OdazqZInZZqz7KEqqC1AbNZ2mjGjPIk6J
ZgnPsplP9KqkBlyn6z1yO/G/sv4yCvp3Z2Vrbj8J0xMun0nxeMP4ZYcDHye4SsRqLG3UZBlfccmS
zhVJkps+lkCnA/7OhwdBKOD19072Tt50d9Qy9L//Xdmc9uisnwJYyoUzm1XlzvxdmFLCWiu/7IrZ
o+LiFwtsLBhSeWZ17BONGNjnXKFcJcpHQ3t53G2KUl382644t/3BGpcA7gpthLvOLKw8no9pG6+M
VS6jvtqgFqrYVmYiktHNnDNHA/c+ikcPxLVpeqd+jHspMarqswGWHzoDz5MUgvhyMPE35gTvXJ0E
3DOssPgO1/vR50jKL0Jtbnkz+JV6RE7amMS1SZsR7tOBYJSycL0yXEJKPikbpPXhdYrd6xXbBOAF
17D0XJmVs7dtK3Vv7O568rCGxUzXIgEtnOer+hWdJi4HbFp+6O1dOoM8rJpbyBAi3W5NBosKU+Qo
e9kkakyHsyHFNfzHA+dPDe/+dc3WI6wzEByXobzy3n8Re7w8IhjeER3mN63R/pAxrdll+yIa3WPt
czueZoykbB3ixzknwMok/b41twLmJE16LqozYnME6mxlz90CKA6zkWC+8Ontk9i24u5WP5vOGY5Q
sgTuHw0cGIhbOG31xCOhr4GoisnVIb969IBEvosQPfxR3gh9QtD1lz0rZhWYgGKltjqwrgjSdS1k
KvQ4d7+6dIst1pQgOp0PSbUq9sxCQFn1XutGXETIOAwpjPA2hifEfZ3tbbF92TUn49m+psb8bkl4
ExRNGhNDC5DYET/Yiyqz6ut07S1ZWV1vNSCNTcHhV0p6AvTCBXeDuT8OXiIcOb2zjNWpA7vhpcFL
e5tpxB4q+r48d6LaIKtnUtaDTWnaJZXznwJadeHI51wTPuRxHsIyhs/XM/7rS3+PFat39pncEd1h
ZgyK8A0HuvfwRE6a78Rl4OptzIj1vO9OiSSqPyGUdobxMEXLp2vOHuxsKGpdmIbKZoxdZZfpANqv
gs085tVSvsfS21cpoQOxUzjLGtd+xATi7OOBxUYt9k1QsgSVxaGG+9VsS/XQhE4s7zMsj6itQ416
mjd3quFU0IaLdkmjkMbtJ7eaR65rfj0B7kv/x6FpYOjOfgEwlGUH1hWR4CKFmR1bjopAO1j8z23q
GhSTlr3ucCVm1ZDIrHdiwheNBu9FKsZAEA7tfcOiHaza8FahfaLYmravavB9uHvZFMtH6Lq6eBTw
YKUsq5ea/hEHHaGk67v2qSbDNi+f+St2FyaZCtMJRM+q4jpCfDugWB13FhPcmY01Jc6PesRftzCN
KfI3/n9fGo7m7TbKhSS1rUIgIRNldBK0YVpDR/+ofahYeyU2ub6fPFqcAwLhhEJwsiB2EqCPNU1c
8fE4X4oUz2EywS8HA1foDgoRTHkbbYkev1Kl5ATpZbraMKW1EJm/cV66wxawyMdfkclEYg01R6gw
fXzeZ3eHdPrzvMh+KK4fokY4pC80ZsBUF//u4FE5muPFVIPJetZpWt805oJYj56ERXRKxLi2brSN
eY9o7hmJ6VOYn5edK0Dn27FVV4YuM/qRwIRmjfbwLcZDvNUZesXyYwuwnSuH3tzbeR2CwQn/BNF7
l5Z7Nv4cx/2oqp6sycWGRcYn/o5yvElmKs2jROxPiN8gPj/LAd3wFGq0ONPOSkOJ91TLcHjRYngM
OLQ+ZV6YF2XBMidn3fQcsgi4GUbN9AFGwIeSFxBsl1Qempo1Iqzug2VyqC3o0t9rBNraCPrA+Pcd
ykgxVGUAVFq57kGi3shRTa+I5z4/4Qf3bB+Y5ts+c7Im1U0U/AifUuZVoaeEyk7qc+cEb3pn1sPQ
bQVP6w4GJBQmPh5lm+7zdDzPCBvc+g8wUszJiUuBtJXux9OvfSqC/LN002Y3Em44fGL9U4KX7ffH
357QNVtC2NuTwRZQmUI9p4i2Tc2ZXRUS1Qz9QzhKaQWai783kyB+3v3r1RN+6NTY1hUKR89HB7gj
KWDHObgPH5VrVagwUteGc0p0Ku+/zKlk41akzJWahRPHsdhW0cLk/C41fwtubikwV2hHoGqFlXBc
OwLeV0M9nqZPPwzu7dOLFouSWWtVOT9XdZbXsCB5JXANY3X7ox5BnnL3efijjEcyvaoE18yhSbQc
0Mxo4ETQvIv6i19gaCpJCSJW/9bROGWT9b4ag4ofZJ5PVbpHqRPtma2zO9u0dZMVq8H/+KLqCM5H
T18Fc6Z0gZJQsepMK2G5bo3pGHmT7fI6wcfwllH0Tyt42mhFGc+4IOBPRo0uqcVpuQYtQ47N1ynF
EF8SeEFjBGhwhn5T3P7MIkoHJQ3e9uPKfLXzcL9spqENTg1LZv7ZKaZvijeJr279NJ7Fj+kqTHRo
KVWwH+bAqOpv0Elap/wxuO8k13WA/w2s8hIuRb269TWzLT5BUGOaPIsKa84sRpx1qk/UZS2807Hd
/6CEl3zky3F2x0hzrGLE5zpnBI0Q4XJBNKP6MWGEt+9fFciZ/aFS8VAyUoxs4srUatvEItj7iNAS
vbC1V/SwlNxqxYXJpaU2dP6OIEalBjsyaDkPbuiMTfxgAoGvHXF6ueCG4LY42e27Ldz9+Pd6A4yx
Hn1exltj5AZJul1v/AnxouOOkUnfepAMGorOQNs/qcm0e5Odi2531gxg86g4wFaxrmBwrDO1nGRz
KVEk7vN8Zzcu6DFvHCRrE9D52EQw36I8xLRpCmBGcL+FCHT6RrTsEhGGktSIdEYDf+EhaCxQtijG
4zowZ4kI1yKAW0dKaKzUQ8y350BOr6ISJX3k6HVGeZRr80zLl1AUl7avzCTl4aW031qKygWvGIZ9
Uz10nDUTVlvxKTnEJM1RH90jU5vty2pIilsPBNjyDwwXAuYi+eIMIQIDONGOxdjd78n0xyCf/JWM
De999ifcHVBusipP24SfCktmCSXE04V4vEmv0qqVeqPDRSMxFyEwjz4nb1QNxZ7S20fXTk5Z5/El
Hy1/mMYTyY2kdJ/R6Jg5WhYaLjKM+5hDIL31Rj7HuwMlsV2+E8iX1oHkkYiI3gRg/hdyXkyAOkMU
jZG5HK2/JyObBFBv0w5Mbbu9y65qPT0vl0X2ogI3VJgbRhX5eM/ISbNO0XqN9vF32ECC85tonfb7
VpAKCq8IX1hvomzb6qR8+EuxqQlrlcvPUQw14H55Xr8wuBZoDAhVHyUHQBaN1R3mfvvvXE+MTQ1V
ErSMx6niuICR86Th4QjQKZY0IZQoEe6hj7u4Vr/RXjfcN1Ahf8dmwe8LVdZa4W41wbBqYdk8Emt3
2CU4b/eVEc8m1BXQRoxZsVt2ETPF8Agb43iyCGyZadm1F65bkR4dxyIs8zNRABf5uveFhUcUccXB
gnquBzh8B63aeSY13bd6Ce+J/G0tKbYI5maDPDVn/2aXwR/AdtWVUU6UFKxIYIGf3TGqmDVZK0P5
ehCIlH1zE5SKqyh5p86cUlEQICWzck2W3RXVOuFipMfexKmNht/PLjk4qScfcwTcbD5mwMqWK+8S
3p/iNAvWn88ptfuTL9YQnBlhGq/Sv35UhEs452s1bAV/GbYNbzgpteHGA3mdRlvfpiOiXwlZ+aG1
14LkcyeYzoQmab8mobpC8JmXVbUqWi0qwkp/6YZo8OiXFh/ZcFIo22xJ0MWQHDJgZsxczoqLhTUP
XwRgWPuQbjX41JjHty20QJPWbyWEnGYmMKtzzN83PRfqr0nFb9z71ksjYvfBa3EsPjWtLu7ZHsaa
9XXVoQmBvA8d66pOW3Xts3BbihlYtH6fbaq36FbibnXi3ORpntJvxXRU7JkTvGqxKqu6lK55sE/5
MpydcsrUXQVLEfX+AoeMnQC+kBVchgrikmagnb4kTQFW8yKAE+VnytVhVn8OggqlsYKAXZe9mOT6
I3yG0+iNvqFnpuNsLFdxYkhGyAQTuNlxCLL7IJ8eYA96ETPP/laKXChOJ4x/tz6GIALpD03mShg0
Xj4wqVGJS9AfD8Gjk9ehKYCWRDSj9ZB/2adaQnC/rw0C2HADRj/HDAAUSizAyjtoFXOBxPyCyGoF
Ocmdq1+p8azs/WpqWiR0GEYYEFGa9BbVGzV0xvLbux6PgdXvtM1FIqMdTGnq/Gf4m/QjSRNNJ2oT
OdzBil0YasVTuM+zBbKQzaCgQTrAz9iiiJ8r27SOYRaqcVpQr8nuAuTGhgjOFoVbVWC7VCziBLSN
77Gjf45m7jZWvdD5R1HdY+Teu57RD7MuOBicYpsRi3ePnJKZ0RvpRteop3g1bz4JsRAVDAnxxf3u
7T2FwvOT1rV8vts81LG9uHLcpEbliuBKEr7uHigSoAp/l52BNKKSoZcloRxsDAHYrb3zr94DXZzZ
tgtPLBxdwd24R/qv/pyoT5iBvPDoHXIl6OZ+VSTJ1PVvc8O44RYsZOhX86kEBQci/YGzL542qCdj
SJ95MEU6Us8S4kLRJv96PhR0vAQuA9F6pXCFt5Z9tb2tpKrWBgnhyHz4KSl1UhPO+xvfwPwAtbz1
Rtqctk/8FYgUjcVC1uiD6AnbCsCJg9qkBPiC8j0NDOqjyX/z9TJ2tZXr4ez9IRif8wO8LIF/q7hW
8/RS0C+cuqmGypEYsN3CeZKH1rabNU5fFdRCiSRYO0uAnPZoT+FcVRMgIysMm+6KpvmC8ZN5M7LE
OjX5mGooQjY6fO6PY9zfQWK194o//tXG09cj9xfsIAzFlLpMipgWIBs1i0sxyy/yeyOLKYuol4IN
H6To8tVaexo0AjXsJdFQykJL75lON4J0fb4srKkTnPQelknWkryXbpXi1mAiJLxwjotfH7e+nxme
k52KDVRqlXtTOAOuXSqJ2FVeMXkkxMnUxc97gf5bL9vUGVmxjbeUG28wi8ThtqMFtJRwy+JmyV6d
9tfH9Qysdukdiqgb6wCz3Am7+1ngHCQfz3YNrERmd5j7OFUj5CycWWmIv7TNhFV5pyxuBcIGsYgG
wEwC2jLZm1+b6LTjm1CY50gWfaQqJHTfi0FFXmTmR7NXk9K5s9rNytxXXesg7h9QbcjBCOHeUwkL
n2Rtp5MQKqxiZFoTrSvR2CAmTyLiG3x2txv46z4yZUOhGctkErIsf+WRQQ8q+3SsMQtjizZt0jdF
U9ZxQp5OXYKOHKwD4AYMW7XNA/aYlvr9rVEnHlbRc/NSE8oeqR6pNUBjbDvV85je/OE48unLSTyx
KwNgSV3rS+pdAUlPMff3Mqnwwy302RvOlpsztCzGzhDbuW2+QrzIiPJmt2C2esVMY0xGcVpatqSL
fnrqwf7O69vGGejs5FrfcFUBkInFpOIZAKHKBnpu+s5MzmZaX8ZzSKEgZh9TZtSTmfbHoHXK26EN
Ev9boPHwjHL0mEmn1bcbb/lngAiYRrtpUcrNwaoc4XfSss3aU713DePU11gieW9yJTS1Q+W1qu2l
a4qXdDkgYITCvNroDyY+2cmutwZrLW0mVHAhgsEY+yzxxpSXVt5Dhu4ilFGoAjz5NAejEArKI2p9
dXS09Wh6a+Yc6Ljdzf3RywP4EHPEuXitFqMMRb1dDTxjn8REHYMfkxYzANNCs5cjvluVOjwyLYrm
OZj0RxCZNbLcTTf6GKoSii6TNTL5/iA+wBIdQX4RlYzs/rKGyrxbga/YKNCqGUu5HhKdHG7fSK4e
qrnW3wxfHfRzviCErKD9INMe4HW6ExzyWDvaZnlR05wXGa8bWtynNtDLoCAz1g2/B7TR9wdfgyKw
9yyWLjTRSnQkVlHrv+CZ0LuOaWDwd0RPsrDD7d4MrxXpw5oeCrwCbc1XlC8hCuNEGL8qUTV/QomO
Kntd0uxbZLKMnXar/bqY/H2++ABgs/i37JSv0sztWGir6dGWZYoF9Nvxh8bN2mQY++1wYbC30wH7
gia7kEI0/H6EDeTVT+ku7yrnIs50GLBSbmHRVQRhfyKRHYicXqfUQezCgTiHUoPZMmGdPd5HFTSN
JepAf40fm7jByQmOczJ0+oCM8kcqSxU27QvU9Y+NTzGIozKi5nVv2w1x1j6/XplFlWVeAYoZHeid
2/ewiVH1foApA00C1gsKQEjeAVcp4BHgxi2NatxDM8bijFtVP+eVlJjFlTlTFyLt95TuM+weRBNH
S6Ef4mhCR3yvqYF9YElf9KH1x4XxStJpCMewjsfSXBJd89qJf1NwWv/ehJzY0IOVDdaz3sqNclru
tUVMJgPib7M3mPA6apROUBtkVapif4NgUhbBVlMcAf2SXnRo79BbIDBT1Ljc8eqdked8xVwExV7M
DHMzNcMXxONQLEKM3UTh4JmI0iC8a9mrxzrVdhYtrlkBnkMjPlUgBIrT0KK9AkXvqMY0JIYTqejv
hhYE1BYnIx6jedF4sDE0UJGtuyIkenMXAAcxlfDawMUEviUmV6VMuCm5GW4A3Un5+GqpUfN/nZbO
tBsP+qWLIYgvp5c4WklXajryg3IgtTZXqVsEU1cWIIqVUcFJkvMcA/Ai1vINc5COgBG5nRaK0eSE
u8LwhKKOtMNmpzD+SzHYoziBKv58le6hn+CcHBbDysQ9nfBRQjFK9RNimttEAepkbHQr1UQxE+kX
VmSHMhXCk4Yz1eCHyqKiN2+BV8Z11PGLquInMFy0sk+ERe3iUfpajL/axnrDPNmZsZtWzSgIHu+P
oZHB78dbFui3xERyVV2ssibUr0siGF4BmFwDlvkkQkOReBjRqtt+qsxEIi8wokTr7cZZMsKV8XJ5
6sAcDkwZRWREIEUAD9iAFAX9y6SZswMU9xPIOBrW/a+uCUxl8n7/toQO7xafDYvRd7OL7ojniqsa
Yx9aaT6b6QS4Mybnwj5B+MtWwetQF6DKy1AMM0T9cm/bdK+m0M1uRJC1j2iUKwo1e4oe7JigBWk1
e/kfYTrHFm0FnEraLTdYZhlYzySU7dGRrdaaC0kIWokOaptWbbMG5k5eFgsZPDimONtgF/CQw07+
Ee62cXwSfQmTzOaVGowM57fwOU09UrWHL3n3Sb6lxsc1S0/ef+qmEJ3DDrP2To8DOhP0OeNbcoZc
ph0s85SCkC9P4OLtKpmGdkoL1+bDMZQjqBzCS3hu1Tef984zRUC0fGtZhJGXw1cCl1fb5iHCHMvb
5i5Ah+Rw7rpwcFDnSmxPUlzEyyoajWSj5IZ1BM+gI47EkIMwnPkuhJlf2JS+n/deYIwrs5+I+Hxo
xtVmlUfMU40dddz/cRUyffLJ6blPYgaRZxOMo/1cSjLq2qxZxYiKef1kcOIxyuVB1fjw7r4dvNwH
lyKVnSzfcKe69D/FBKagErsYoAOWkivnQag0qNHPBAvdVCSnTPhGNIDRm50uSOBonY1UlHD3ycDo
5GKj4locKtWdjO8r5pKLCGqIBlqoYKkYOjk3LVqVuEMfTnGPvKWcfsDMyxmCMAUYeXfUtNCxPfZ/
0LcHNRnSYCFTZWGfiQttnK0cEXUwOln91+WqQytJ/vpfd2IcuETdKh3VNMS/rCwZo3h8RKHH4pGe
2WCMZulSZTbtlfn59NKuR5RuJx3ECWlB9lH5h4CAZUrdlxDBX3fWOl6tCahcjll2jHlRD9ZZ3D+7
7ko33nl8PnmTVKjXFI3ESaLL3fh8WYrobgU+5dBJ9Dmwv9a3OqCI8L4EzJo+yYk1La3U8C8tzFVG
T2cNXise+SVOZ5ujN0f9ThToDKzOHR+BsSBlYbIesnwCYV8vVphRJ744JX1UZf5MOL63PhGkQyhT
5pcJMhLy4+OgmGRbpzPiFB0NONH5G/Q73NOD89USKwFr+hndtRuj+LAPd5yrZr7whmfKO2VCNnQN
67N+wbYbgYXXXPhGq2NLvxxmnCJMpx52hpbX/cSUjiphn2QikymV5dV17h1pVdxg0t2+eGwxGv8Q
pY0uSRbYXWN/HY7aPxrOJcSIXu1XQSjTntUnie70RAZEjH0zjxaWeiNIIUjHJ4LphaY2zrOXIUci
KgAganea+JPekuEpEJ7pdhurJzi0DKLiJ0KN0g0D/SwgxvNsHTAtXKVQBwyg1i8R8z97+koELqbj
/sqfrCdtrZfOOH+62JedHkEk+kvN9Z2BgFbd8Ee92GrqzWwBchUYrgBn69PIW40zn4KxDoIln+zK
77WxhZxY+0wZBB37fhCbxyljKJR4Fg6OUMRIBQmQBXXwMvs3ecQYkX8CM639N7+PBGVmu+efVNkx
Kc8EGux9OyR7dXUrbpIVDQVOFeNeWEHDtZnVjcb5TEJLrWgDAiOTMtvHGRqk//htYJctrrE0UJYX
GQwMaUgd1ihTFnx5heyl1zcwdN99fMKuQhp/UDFJ8fVZtycHkCBsas8YpJnWUmlWoS3yjn7wDQIO
AtIOo91vCMEl8P22YBsqUhAhZbW6ZckNL5qlzYdJeSPQQHTgtqiaf0Kw6KcL8mFyK04wRNudkFwC
w2UG+S+uwsz0Rvg+NUzjbvv3qOpeMfXQzIosXmLWRymi04iDjR0t4PF1jh7ltCUjMZ5NXH49Zqqz
rtzPmTsTwlkFv3VUKIV+LIo72y8rOCXNzfPQ675uFKVKWGmYNUdwGIjcYe87BbW2wKxQ4XdxeLc3
N8OR1fT8LtjBpI6RSf++wEzSC9gr6nTS6dz9VZ/ZMp9Z16Z7p4egVlgw1o037LQzWDsXU9ol9IRn
pHgcO/+ADe+vK4p6VUG7UhyAubIFtT9mTSHkOaii2HZzAvBbBbOc9A1msf+5ugyFaBZ18O+vHEbJ
wB3mMNS5LqOXlM2ScYz8m4gdkYV7cCJ6yekhNsORbd/Xet+gRTWF91xSLdNJHchpCiRpPIunzW5S
578XHe4Qd6ix6MjaB+zQhYb9LjnJeHMzqE9PBBctucT+eCrDNOEro5/dfFYf7XXtpMdOXeFkswyB
otRU4t9PVi7Uw/kif0RoDYYBb+hmoe5wNjg7QZ6N/EU+FZT7OTQ9I27Pt0v+ux+Gd+YiHae7KMYH
s6JmR0w/6k++Kypz3k4qXAs5ReW5O4q+kAnsCdQhwlaxIWK1bpr5iYQOWTp+MzkdL6ehmJjuVOWk
r1F2zAo9JS4YO4GRTnKytFWKJlFZZcHZGqLbk/NUGC/KouVE33Qqy6K0UG6mtWPQE1muFHA10is5
9HpF8cUzeaVpPlRW7Hq7ior1mKcQ23Bs3hgjduLAvbn6T9LhxyBdnTmYcjIAfciljB7vSZIiX4Qb
9BVelT05h+y+NQvxYwZmCK95Cp5rwYc1CeR8RzdftiZEJ6DYFCcm7qngMykprIReLn6X5f7ZMi/L
vu/VpG+Xlsrf1AcxG/xVx60d5igQ3tewWZBYY1iU71XLSn+yYKowKBS9xc3sBiQjnU3PcThDj6Cl
pWL5021Kqvm+g5rfKjMj8Ar5cIaLHd/5kNx+zm9C4S9Pe9CgH+blKv6ujdXIlVrsI4DU3Bk4U+lE
sFg2NsyXTn4ryXEdiCP/ru2kKonQdkhIfoFv543RIFWtnDYNAjPJrdA91tzm802Six/QVOZcphTD
UacXuypWfjgsVt/EIBRPOm9Kt816OJg67jVrxRsh/2iLX/ZdlASd7PeBPPyxu5yqT34BIKggd3wq
lHTPuWb37rklzT4ZERnuKqPJwVQPrChjFO+qw7URVvTVHf1JW6QFMeV8janJJnRdASanhKxBs5ew
PynqPC1gxyeIQ0eAyD2xyZrRlfcQzaSuTl2bAo0KJvP8lvfc0n6Mn2YAzr3lXF1dxojhMyDj/R2l
ipPQ+2TPqymneY+PxbfBLgFshjbVEyO0U9VmDtyI7i5bvg8YGbA0fNbW5AmWg8LQiceFF8LHGnL4
8uDVK21GEndUA7FmMkAh+6TMWDz+BOX82cCzVBcZljDYGHl5lL6W4YLpvpbX9IgNdVgQ+2Lqp2SJ
B+lwEH2+I9v7UWXhZJyWj3wrLbDky9oEGjWXyP2mgySa22yNFMlMgMh5dcoM3DciIyqbDMEZsQSk
CrtBlf0tin2XfDUK0aL+1mb9IN6TFgc4bJFtWj/PRJSQjrxHKOPhqDLjrAK73R4qAER4sANNQjAL
pgwao3siShBiShncnEn9FgSwQ4oYvUPTt4SRr7TqftiA4UkfwEJ28UBcM84hs6bifS/AeezQIdQ5
8fudDmGetx35fUM3btsIJBqOwhZlL5T3j8YehpESpD4VTvql0jZbf8owvSWV9qgpUR6ztyXLoa/u
QrICzpyk+uTRwq8HShsUOB7sa19+9NU/S73qQUt4/dQe7FKMgL+1R3FenCtfOlJW90yN8S0uZj0H
PQZIQ12zyD3FcQ4ewWg9KWMPvrXjFOiobfa8j+8OmT4fGlCAHZPFHNK9qnTuMXqBJglEetMR5jN6
6QFsDth70yuwE3h5obFyL8HcbnBOdF7W8pbzaddAhwhToCe0H2Y2saa7wRKIhu3g9p1ptyvLBmHd
oOZ/keWWVHBKjmciTjnLBNoIeMALueSTrO9ImnT01JBSkD25hWcn7pzEACxAygYaziRQO8aiu26j
jlDVcm7fnpn/m7vh6oolRzrrbfGdyEe/y3cyK7Wr2g1RLhiWtNGoyxWF3vZGmwzCd75mZOOL6Zl9
fQ4Gzshh3zl9pC6UKecRgjmXFCiyDJsJgpAYjevOHBOAhnes+qysAAMFVx+dAFdBQZ6I+Qn/cwRn
EmxhYvL4ajD/gvuOY5s8vpi7BlafSLpDVYCXOYDUeiN1zfEof8TuB0SE4hxtgB0bU25mmqXn0LBW
ICfO8CPNMoRdGZVsTvITlPYTeGR+yB3LR5Vx8DQuS/ym+4Ij3+UQ8cl1h+IYtUMom+zga1LHAGeT
gke/vgBlie9yQkERq5yh5rRSOdyYXqx6kxCBTT03y6RDfXzlJSuALelhQTI1SLSPMx18bs33BfVQ
4tFn2bWwR32kLNLipC/jvezAKVv1uItcYQCR/dND23xbljuLANyx15H2cGfEesdaVagdTfa+Dvf+
bhDfOxSjZHqlYol+3hNVQOhcabi61zAsD9b21bS0IdmWYan5zByH3FClefJpoKCL+V/x5ZOm0IaD
4aVpIf9E/izOcAVuK6Cf0OBM/t8nO+ZA41E3uPpa+x3gP6VQS5JVStWaw3oQ47zE3QN9QH5QHk5k
oQR3CJ1sbzMYrI5xPytSHXC7DfTSMp6uguJfqBfn9uwwSjA8l+ZhhF4Hwp4UjKOp4hqN/IbrH83f
cVU1bNEnsLpYfs7Q/UK3R78xL4BbA9zMsUihMSTQKTKWbqrRliCxhV3uv9ydn8vRIZXHvWVjdzsk
NBRtgoS/037b7uCR/31hMiuYRZIhYKmgGnBSzyhKSoFpr88I+WmFc+JoQTVWZLZqkOzV7/XdJVzA
mkSjvGR2qSucogjAwlZcXcGkLKTPoDQ7i39ujDPD2uJVkuIAbhlJm6UN8uNeg3mwETrZLKwCyqtp
M/eqpU6fHXnr4p/d7I3vtFxyo5RcBUH9qemS9jJLPXQkfr9+xYgA3wAI8dLt5opHaikJFyuMA7HE
jLqqu8iHO0g1+/xvHO0WNgVWqyAw/DETnxcLNkji4/3dzBrxm1rGNYnxayh2KeqoPn0RHMRpTK8Z
J5WH1TdjuXTS0wM0TT7YBZOhrtkVLK3K17Xcwqo1TOfxyWO4hHp3pvBRdofNRY5EctnQ9gdbqX3z
kepLbu1p3rITWZmPmODWFhEuNvWXWKdrhwn/XJ0KOT6qth1auMYTP5ryFfk58qMG4QqVNYoQU1o4
u7CqlbdReW99NFTFBcUvszLek6DVw6cyo3efeVqWXM4MGTddnrz0X+N/KOdB3rc4+8E+kNWvPA5g
jfSYOGwcj1qeICosqwspwQi9myDrAwl9yg2K6OqKY0eXAsajVeRuQnTlNetHRGZrhGWdsg9DBl63
TE9J2oM6WdJoMAS7/AE+4AkxVgfRi4+lalEzWs+F125GjWJ87JgEwvb7tLbEdd51Fb2UBLCnh5cy
3MuDjnbkaLBe6IM452h5iT21mtWLn9JpubCtzl5vYZLtw+vb6lXryIT++sZA/dAQcAQdrbarqalu
J3CfcinPTuKrON/e6exjBqDCP7wUkuHEwyEA8RlmpTnkH0Ye3BDUwldkQ9CbryoaHeyb2pbvCVXu
B3cpk/89+CaXavz917SMooKtQGrPWZM3oQEIJpln1z/qS4BelLbsI7S2wIZM0oaMYeDFVRuQjFB7
hMZcrAnYhj83WaBRATlc+gdYozei16RaI4oLZmCN3cP6fOcuOagTiuYllGahfJNZM7nsZgWjDya0
iXZWRNe3bQbKqIUJbs/6pmnbg3Aem5OBjod32Fn3rMrzt+NLaUBh4zutHIB41zdsSD3e6IxgToV2
fDfFMT/dtox66Oqc8x2lEIsKrCdZF5TfBknypW2X/o70BI/HKvv1hKcFIRGogewlryc++Lz71n61
bZMwo91fJv1ZkAAd+vZqhkStB73Ug9EKwFJUmJn/eflas3Y/W+e2d0Qxi1rWMoYO3cFJZAR4GSJf
NCsIT8E9Iq5KgZBPDnmvJxby6jtXmNq9fPSzcJn/WEAZWOCT2wCdNgfpCdbkOXBFwatzB3Qp7q6+
cFVFKFk9HrvVm4VNRIoKYTD4mg8HqRMvITKhdcFEVFkEmrriaRjdvQc6ZeSCmx1loyncJmoJHefE
2iMUqkUs3YpRPzfGkZLT4BwynQ23+TD9jzGmzeRmpHwxGh25FcaJO4qatzfTkeRPF+CX/7hEfpeM
2CpoSzRYk2DcclYriJc7eU2H0+v+BnV8r5v4nCVgTV7OYJp3+57t0gz7uCCQtlooc3rtPPmebeAe
nx6SeMu2oHUv8NkNYs1raWKMfg9Zwq/QUz8h8ZlIqqWd1J2BsFLTxy/pMBylY/DcRS6Jf1RyzTjb
mtQzZjTNNsi+ENe7k1V9S1sM48TsALcDie2vVMU/LrFPuEL1mP9I+ln++ij3O71Y+rkLr4JYh1sS
ETuH1/1vXRpzK+mSVikyQjSM4YlSn1TJriQl6fR9UKDcFTebu9MXDi882iMhwaf4JDWD2KzWd/h8
xXWASMDfNUUunbl8qvfqsK6QCvC+BHtsIFg7GSR7RJWUDf2neokhCdVuH4yptjqzWcOR7YkIFj/L
2zqKzNvdk00IcXcFcA4srAaD4AQDfLf85sIA1gPkXEhnJXjOpqr7fgWm9thBfUVOHq0JYHittduV
wankDPQcG5i5YhDhcwPkAWuFmvtJCgKqvRr5BX3idpNIPFTjEyPpvodLBJWqfFukgi+03KQDPgOL
lFsVgbokSlvXBqPHPGUqpHN57wOApJYZcla7rx5oYjVadzaBLgH0tSGPzTvLTVHo4nQUhzxFOfmA
+sVxm7p4xr4qNez/EiY8QYK5ew5zh8XGg+2paBQHcSLcdoHkayG2o+IrnCUjjv+jkn04ZW8AR1aK
ID9wLYe/xcj+CzZIb+gx9I7hQPrXs3pa+Cq5XLC+98KTEfBKjRC5myqAHJ569uvh1MCpFU1ZCqO5
0fkiDeiWC/CPV05630TOIUDX40QuYfzneeRlM1CohBWkl0AnlVw5fqbhPJfDzOOaM39zflpHbYZ+
ggpFIakEsX7dJhpHUqUBZ/5uR0yexYrRatXD9K0+M/5Ih8vZav4UC2KdBC7ZT0f200+3etqKlJe0
v1ZQuUIV+wmxq1JWAuF/4lUQyJIwe/zMhE0e6NtHTTW+1EO8i3dyWLcO4Y1XHhECtAoGxGx1tQ/W
ZKOe9iTSs2/cxSQXMUKUQLbM5ctwa7yMqzynTraJJTwdZgs+bDC4vGo3scsBbORAcYoYSIT0kImp
qBgwkNo2fS9+f+IKX1nupg2gozYPH70UCGCym+OXq7tPHFu1T4y5XxdOWiKl3FnetS2b2Lym8D0T
JiQIaXyL569HCPe/N+r2HxxbAwWroIzTC9pRhIgWcw31Kf9Yo5L6SeivhUxF350h23WKrdQg5Uam
sqpw4Mpr+Drw4wf6zK9RAaCVn4hfHw5fLdrqu7c8v+gWTzaIG6LjZFNYpYUL4dF9ujFDc1XNW2jG
Bl2Xuqfl0GQVPRvTXo4d0bUmoB7jxea5NoAhmj3rhNas9uJtynFjjIZ70FUbKzcgHYhSulwIlU7R
F9vJa8Rer8+lqBuJu6hrLwTA3+zbQjaKpiv/dc05ErMupWWK/XTfv+0KXcdjhrWxzl3uwUOOv6UR
pC4NTUhVIQ0Rvo7aQ+HdoQXd5sXejXOVPMnvNt/ulFu4k+Xcgim8bf2nE8zv6K8UMLc6qGJ1Z8ZS
sSagncKPALL7XXeZk0oJdsa48JSF8D5gOwmKUMNmJIXKGh8dXJ05rhPe6c/hBgxxhvc8c/SWU2Ou
vfJ8XwGAypIb9sZ8Ecoo2/ZAL+/1lrtevsUTyZ5lddNYGVUPcko4LVKUwA+1MN5BI3VewQAhtkkH
HHga82Vy49Ky71ooceTzCBXpcRPq9rL3zxTdZxNazl+0s7ccGuobIR7YApIiKAc4zOWD3lvOnMuU
+uBBpS/iSaxZ7IcV/4WoYGJPWkuyKofXIvBdDXAQPbFCczP5UW9bco/fS9Lrf1hlyO+zZZPKyCSx
4DGGJrqDZdZ6/AiSYEsxgk1eWG9/8YyU1ZudqaGA3MkODGHwUh8/AD9tsKwOPg7Ex5N0EdNCs+CY
3DNgKeHTFAXydYvkwlBJ5sKL2e3EkUZ1USvw3vi/qU2Kd4KVQq3XZawNddzLJky1loLwHyh/t2Lu
49O6d3dIn7Ls9IJ+rpSadgz89g4lGiuRbaWnpY9UHZGVoQs+Mw1xGteM8mdiOSeKd3xVcyBjFYWE
oUjem9kUMGaeIhs4dEQ5hm2mKe85wsKoAcUb4M4+RwSznYMRqiT9lA8LqOQxjyqMG1s6zsZmkXjG
rJY3Xt1XNS/txFKIKh7+cErehlqWQoPDZIZt6XtDkQRKSZa99VUIxp71bDEGqO8gFOK9kSNhCn1h
0S4M/43PDJEGA/QY72lUDB0L0aDGm6vRtaSHsqqUiEaegOsSfS+ASbm5JMMLfsagN0PRdCxM2eBT
Xu1uVZgp90IDwIQLctbMrX/BKnzD5t6WmDd+iCc3Ix8M1wpQd6hCwe1qXgC4WYmAm6ugtTqRB/8c
9YzEWrwBtrdAgaYbkikmz+a1ZjDfPGPN3egbC0235/pKi82TCYob20hyNz4eJs0TjyKRnXjAlLU1
BsKXcONDYzADdN+EDLyFYIxLCXqA985tRfUfJ2mGWPOi8HOJjxvoF+t49vTsJgS+yDogF+uNBrHy
OUaTNDQaMbts/iWJwfJbjib9NoDNSdVH6fFS3ziK1K+Kj5kRbd2IFswdHm+5wk2RIgfXatlIVDSA
joqRe4/f5GwuAEfnKfwUiUN+fYBGNIfCFCaQhOuvBHI5wafX5/3whWBseKCeNDyD5MOhNxG/sxSx
H44CUosP2R87X7+fd5fLcA8cSwsfZ1woTYuR5EVlYAU6dWLYeXis2hxopVmfLrswX9PnVQGKafRv
TgtEp7oBUh6alN82L//70vJM/dvo4m+M4bvCTWDrBWDAW6XwvVKDue8RRp28vNFBj9Mj4RJgduzp
CJGcoriaZTfFz2mXiVDeauvGL2BtuFkg5Tb7WUZjZpKXpXqVJw0Vmj7ubwoQ3KKoyOP9aAeTWORH
zeLHrYtZcpQDJzqvXQB2BMj2IqW5FI3Pb0HgI/7zhxtc4RgM8uDYOjtZY9qJeqh2D/UMK5lJMPc7
fydmue2CXxAlahcyZG7w17g/XVwQ7Q8nEwVR7NN1ICk8lTMdMIo8fXTHUz5RaZFlXioeyArdC0kZ
aOzt8AtxMRdUV9MNKwP2poNxz8K91Ch5NB9vey600PPIx7KX58RKY74MPLiX7O32XBTPs42AZsKd
vvtxinmHIQW3zbBTDFsmr8CqPiHbVFchEj95gayGc1gvtORYqBeqDFs3lX3DSgrV4kZ/w69aiU8H
qj0YZ62d65IBnrksybpWQVcAtaUmni2OsDeA0d8XitS2RPM9rF0WyjMMBQHnVc7jC1Y/6lvrHa5r
XqHiHoavUwMIhRG5eh65LNf5nhTe+VHV8XVp1+OYMt8u69lEqjlc0p4NDKKCfdRdMI47LojGCkwq
sOdJIsRXGda56c0bkhbqlngtYufdwhZlIDVhxnCj07Y2HvhctnFEpI31P2bNipojqhqxlr58zZcv
LNiRjpDyQhBMpQidwFb5qGMDw83YRJF61xxWuQ1ZtowAU1mYWR4SAyUyQbDNXvutuowZmQRLtLjZ
aPeL5EPbh2rBOETfaJv4NSF9vbhdUDi1WGLMu2L5h/CO0CpQJ9Qe2ZFXQUcGZR+slb1Bs6QdlImk
cPUmV7N0TCSP6/eRXx8RgM1hQ6dhy3NDnjAV95yVdo9PQUha49zvOgFL4JdlSGxr7zMRNl0Qh8ru
aOr0E814bmAlmdFpCD5k4axkjYILR8y5vJ/b6EHHLfs1xSf3iwcDtU6e+1qOgusqCe4X3+6ZusmU
64JFOENvCsmJqqiwdDOO8tAfebQJVEF/WYu4lXKnvCsA9OrHq69zcQ3pfOaN0BbPo5SPchEXMTft
E/vAY7PL8yXwxSHDbzAwMGXEsrsFAEnjITKaVcgttLcAAukFK0PP3fa3D3ICzs23PlbXWt5sz5+K
wkQisl57qh7Y8hn6G4k3bc2ZqISfyolQ8qSYXcsTMaDNu7bUdFWoRK/hJnX1+bmIGgtk+9Ze0Pqm
zkxLkZEZTET8Jq+FNXOlvSe4N4neCJG5i7CJ2AEepVe3JbY61EMiQLWrQNxfRXs1p2PFgfMt7Qs+
OWkzfcJv6mMHK573t6gItrqlVrLveDD6PL6FgvrkpMfckc2yiT3M37CwctQTz8wD6dEMLTo2E50W
El73qrNj5nlImKP0vUzGDYemHtcUhzqZ3nDeU4YUqU2W+LYxJ08/l6c3YxhesbhAPk8G+G3L9rXn
IMeHlbVSe5mhkJyZfjOrbZvkiLbBtTPqy2wB3LVjNGJcJPkAzCkqrKT22v+pp03Xb15lA6C0Jjfy
6vnFjdjEZBHePlXPXezebrWVd+mv2U2dD43nYHP6t/A84LYAQD75yPUlq9hZjXfPTJ+Hzxd7qhR/
MPDKCMMb9GbeQE7MsJBrzVb5paXzb5ZUNLPbwrYd2HzugRXgnIrkMBs/3jzZLP4xG7/5sPLgOWaD
kIvjEoChqUUweymzubp2cP8aNiR0z/Doy1QE5ZouwaKHXR8+P0tNlk0bQ0PJxq1SlKw60hyeAt1H
Dy6dx4qgDJzsqx9+C64OmJ7bmtaP6BIl4kB4uYEEL2yzUtC+UuBJ7lcaC4iELrTGfCxuYVboAcmN
SE7OuQsFyDTp3iw2hUsBl61AmjDH/LSb33bD/887anNMmVYjlucEYMEOdu1FYiu8QVQtQWYE3yZV
yBqqKDPKjKKGxPCyhxk036jpZmOx5xTOlSBA4LQOkAeWQSUDw6xAkzyzMf1i7+UvvNqRnJ20DrFR
bzLCHnu2FBKFbqzd+4BI4WR9qMEByY/Omo1GxJ3mzmW5SK4zSsfVe9voTVe9VdIN4QmGNKQr46SZ
U0KA4mtZWAlhmQuq2w3sOA400s93a2kH1r1IOt4v8w62tQqvc1xxGFGaJBKz6xCKmIRNFA+kAlZE
pYrzYLaXwpEty60GLOynwAtHAEzGKLKdqik+tWzRJu6+HqMexMhE9T555hZh7qxJKghBQxCcIkH6
Oqo6XEn0LdA71rsGZSeqy7LHrECWaabkrcIfUQXGK0PtWfQ3Rp5n99ZtBo0Ljy784Sy4dI1uFi4L
WY4rMpuO7zLNRVKcRW+SfZLRGS3qp7rjh+WOFlgHmbMxRC6wqcjZ6dS+iULVC9RwAZGV7n5Pv+ky
EeYPM8A7IOvuC8kahTgnuD1VuSpW9mYbPtLQlq6746DmCrMF5ENKWA7QMFmnUzqbSFYmHovHV25a
RDM5i+TAxGDMuBfeb3kTcSNmesMWtRKGThI3vpuKahoKvlzr+dPeOotDdSTGTUHZUua3p3X8KdB4
oKugCVyyeKQnJLfqqFRFtoOhGYzqSl2Q5me+8v7bOw7SSHfrgVHlVnG79GY+tEMV+sSS2LSruYE2
6R+ieAAwo+3s35JWyTEvxRalbsHBsdXYuWsGqV2OflFM1KkcFh7dVF7adCIj1p+eIIr3A6o35qUN
h0yRul7WHhNIs0iKShe/6Ht/fmzpbEFYKYa18cn2xY0IugMLPtFnC9ClL+V4m5Lf3Q0yYqNwGJxE
cV35tj4d0c0+xYVt6Gf1gi2JAYUkUywF5/FFZ8qIrVgRbsahpBrYL6UP3/6oqrhFdme3KsiIA/JC
wj3DblwUNsQlHab3utWXBBwUK4PC5bpANssYlCijwcNToaM5d4JRqP7UnbAi0NmwWayg+mUR9rhO
q/nUAQOuHRbHUzgXKshuOHOL3/Ju74RGJoK804YUtpKUCR8xUyEMcqybt+/oMPaI73IErkUdhzv6
W2Cqy0lfw+YgJRlRR0AX258z1PiI8HCCims5nn53iGK0znpp/b/jWq0Ujw3yeje8l34ksjzFRYpR
y+EifuPK2BFONKpv4VHkpppeJdLG8hpIAk4xuZ95Z5RHPNP2KSiDdeQP7onbu35TZlNEoa3mHir4
v+x0mbOWhkKABBYDVyZBsljTNIGNfuZceo7jz/g8QDaq0dw/co7gAGhQTIFVmCdDWh0p2M3ar7ig
PqP/Su6GDOM0qVHH0aKHTEl/h7u6k0mva1V8hzBzFE5SYhvJC2IOxiDDx9aZMzlCAQf1DTzMDR40
rVU+HtcfFheJnGU7InDH5CFXrPvJdXXmNkIQrrFuNmRtMtUsm/KDhlTkhfkZ3XJZiXWvJ0hZ40vR
QP6hJMWvvaEerfFrZYkSspjwFF0uzxeoip+fM5xHCGZLiO5VuOaKUn8ugRNVRlnGSCU4cED7DncK
1Vs1poEi/97VwZLlRVLroWU+uyo6qvmcq+LltjfS5gwPIfToeynptvx/35WqOdvU1j7ycYGQdAF4
MeC+EodD44gEmeWmab7r10ExuH/rQiD9ThoFb9s6nLlwwBKzAVLI0gJ4YBlTJvuiVCwsfg4C7j+J
R4rt5Ix4z4rnaVM0utLOwP2xXI2hV4FEKtBWaU3drOmVF47d++2U/CYwYFwRUtz/3Xux90vR1c5J
/Nf51DDPJwCYWVYerhH/q0/Tdu+j4eI2OR1rOo0gAUfMgvJ1gk7eZOeSrOcpkRr5FcweTAujqj70
DV/YzUvxi0nkhL98uNu+a6hPg24NURRAbiXSL1itnQo91Ie+gU9XOKuz8fqzBp+uS6n/vUWmzEEq
ivvY6fE3tfMJUtcA0VXUcYeuYL/doQ9NBjDheknRVBVNdDDy0ITSoY79oSX51sJ32gMBLRqRWQKV
2WE5s7Olof3aUAeA2fBa+7Iw714cidxiPb8o7r4QrZPxxAtkyExlHgpW2dhKySxBr/tjMoUbgqye
VXGQ3i1ByErHudNtDu6bM1z1/b6ZXjcvejUh1fQ7qAC5ehbSunx1hKv9FJQx4up2KBBGOyYc2aAd
fNERLwWCkWWWFGjWkGU58BZq+FDgceKDFXEwIOPiTmeJKTgwREqNe+tatG3Qie/cwZEZeMrJnx5U
Tkz8cNzoPIXu4pmfq/RaykuJOkecIWDWQtyr6aqDMhCS5MCCwMvcFDge7MmZcmD9Stq+q4NfC1oK
/8AD/sZdW4ABUBctTirm5jQd2i+9UtG98GCa3WsjS0w4FBOCbT0orvAA+EHKkhM+n1557weanboU
bwbo2ugXMcj41KvVcbvw9r/zbb7ycR5bxHT9VMphNjDO5EjpVI9Ihws8/fu//zoiU46BNf547FKK
TUGYE+uvKqGD1vWX/K14K9PGbnLY0bEAjX1CYn3r9SGx55j0lyVfTymOd593Lvpvjl4/1c65ITV1
e4zUpGulSt1QRHVIADN9n/mmnQXsHH3iXTFZKeYk9RJ7akkp9TWPRizDBn56Zkp4eDiHfp0b19n7
WxqMjRgJ1/M0WMB5H26tRN35nPsPmFiPV0FEf7JRX9XFFZFwedahgc9wKP6rVRHWwRbVyBg0n6pd
1BItyuscKgW9nXNSbiJpO291++SpyfqFUvnPmg1UFvM7OHMnQ/ZurI8PoUZl+yTT55Mwt6qhKRwh
Ba1S8udVYIOTX70nx34Z/ZVcmS0gKbC76d2tNqvOspeul1MWXp+1+IyQZhEpv08g7dNW5+Ze2ljt
tLlsYuAF68xvbAytg1NFX/6zVqBJtFycEoOMFPcP3GJ9TryydCK0WO+r6tdMgZFR01886eIXIppQ
VlWOr/1t11wOVA39Ht3EbtF8AiK6/dIx1cIarlp+jIfqf8u+AeoxlDgXfdU8cKeA1XUdD6aB9xY3
adIIyJcbvg3Fd/HYOb0CD5vrsk4OLn45i4ab73CtJgZnYWUXLRR26VIAXR4WL7jih00o+k4bqghP
+hky5bxZTF13powlu4h6n9FGKoJOffWa3vlsb/wxFF+1fK+mI9Sjdo2iHDT3GSZjC9Ryh+Qk85it
aOc/dGyaT6jzoM0k1z/X1dAmjdIHycC78z3JyFR8rlj/DY+HNu9j/jrDrnuLRme2oeDHz9FNmWFZ
uYvM10UYfPe2UPK2e+ifMEozC2nHzFTOoL0E6nx+1H2iO/st2u5iMqIjQw1hQ57suwN/7+ABjBxK
ejDjw0QYJCjXo3svAJfjBoZnmeflss+H+UTKQlG6AXD216qX28SOnsq+zVuH/S8cQO+OHwPzaJsT
rc7MnzcOj7pnrl22fHcPgzMP0ACduNRWdyMdAD50WvXqbKnjQRRXSc058TzNHGU9HzSQ6AGAFhhU
4nrrUV7jJmRBAlFOadqfXkL8VpojGxbodd2moqHaMwfB3hwgrU1HjSr5XVqUHyX+c68eAJ1RFK9S
4hFslkFQvog7wSxynOlmbMzNMXPTC41VDwpPWLXe3+B+kK6aFeD9cFT9k3Xh1sxWUBstmq3xbanL
Y/1t9zAWRNV/2i7N7gg9oHbIBc+fbsBTmeKauziBL5Gxlo05wKxnwaLvN2ZHtOWIOElZonqSoyME
55JIN5ZsQ7x8I/fr82HHpMRhk3aKQVlMwCensIziq7A5bWVHsiE/BGOCfXu9G0TuAwcMH994wTuP
byC9jZuS4CfvbSHv0qQTh/u7QNTMoMMiPy1pNNf1MUfMguzHkbNLr8BlxovC6dnD9QrdaPbT2OIp
FB7V5pQY8712DWUFbFQZ4M3p53bhsVHsrmOEH1M18jHHO3oHw+HFY3EmTKSvfxNmPjXiXsGEs++R
OCYW9oheTrxbeOtD0TutVJkCaU5Gd0qKL1l7a16zE8z9xy6NvkKnzXu4Ayha/OL1hPzZeJEe0JwJ
qQ8pR0PeuVBfrAIkIq+46PLAiJtLX4c19N53L1nDd4/9EXc1yTRYok8tXs601Ul6ZV51Piqo0ZCd
wR77GEjMcrQ/zaGCqRejn5sfyZM03rAc23P61kdy3VwQgnFTCgUHDh4DydvWyskU9TzvyIRqBKwi
KyX0Z7UZvmKTnYNzqoyha2I03AKQwesiCSaNWQ7t6BsIcbGMe4G3FGbhxsyUEQQv2jV1CAEL0mc5
s1l7zZMYpfyhtvm6khkUrgkNvyEmQlTLD0QwJDsD68+ymb5G0SY0A9InCo+wqsQFr9S/ygdF4Sdj
3cWBKQVgrk3t8aq2ZXrbNlnPOx0JltMVPORgMRKgCcCnjZsgCgNxh32BW+uFpoJ0E6WwN7KYlGCK
keYLyofVUjB/LS0CkcBYrIs4iaTjE/xm5uZD2SObuO+P4aGsZyFW/SqWNNwURiXTCRK/JGk2ihyj
2/V9YZ1cXyMZTWLrkxNEfIky7N4/RmkyompWEmQh84LIB8FEWR1389sYZWw17JnPQykKgy90fcLs
hVhurRzuaBw8oTy2E+nMtj8D0hzRdPAcC8keWa9r5A/ycmtYLnvwliLHuCRpl3jRNoG/rLX2neaZ
1fmvriWzpKK8+NXRF2eYw6BCfVgPC/B9zCmHDt1LEdCUuIKzmT5/CHX8+/XLu8vhpl31iqxmtvpF
zooOy0uU8IcyMFbv0Umf8chnNtqdpfpHv3cLbwB67Pajg+8e4Ts8YhFl1bclQk11oeqGqE3WgPAV
9cPxm5kImgfr/PsKZP7TU3Lqw/6U/m5keEDUe3ithmuWGSrw2oajXEtf5heRfRqiAPJiMQAFBvcz
OpY47lLnDEtv1Nk59oRhrt3vlRP5LzPV9UlXQyjYe+kaQsVn5FJ8gYhxiwFPALhLTTXfhy0wpudf
Ymptxmjsxgj3xRVhEGS2KlIz9sHI74015wJQG7+TjP+tuaZFOwj7fIZIRmKjwXN2LxXR1LIsI0qc
KeXmafavIPYINBobwpTH8Crn/1zzWv7G2B1D5h1UTLUmzN4cykugt0QIUxM05aNxjVtPc/jpTap/
UUhEdzFrNgZoM6RajjzJqW4aFTmNjQ6A9gDXAMsIAxUXjFCzsocPvBwAfJ01ykSGldBchszYopsx
TKaP0SWX4viqTyU5ActX3krWPnAnL+FAulhV8j/JTle6bud1tN0AV4AHgP4W1M0QAOqNMUVVgUH/
CUwcdwuXxEJs+XEDYAdJlPCjn5SJ/KtuIQ8FzLsYDTHI4tldHAtwT0zh9YzO8dg5KGjuWyXuuTlX
Ufqz/wF6lQ/WoQMfCGFwcxcr2TzdNWQECS3WWKpnX5Sopq1UvqV9cMtNPGlFOvmZUvqORGAO/wQu
ExxozDEurfswvgo9rNlG8TFySX8h5xtMIBfvtSqrqS+0G8oPY7tweHDBMRUqK8qZdUkifEtP0ZTB
6jPb8+qCFdTor7uixqvzU4BfUVlCkSsmdASQ50aGYVBTDHedmx4+bpLUYXsfQ4LNyiZcoTdTO34N
RfWlVYpOT2TJDwuNfFcYSwENbApux5MN7m2r9WZ+yhE6QXmImZSir3j+jO/mvkosCD8sTWzP3ufr
t+5BVS4YInUHL7QVDDDLGVyqaLirYz07Dr5+cPuhMo7SHiro2tiMgKyMwpK6QkOpLlxIdVSxKvgP
vM5TyoCRPf1WEVgHv851IHRw1XcJ+tjwn9RdtdVaiWqZTMkbvQviOZQ1P81nJQ3BRMqPCOjrVS6B
+HMkBvRafJHMzr4zQXRW4LrDy7WBbtxcdUcIAfVuXWRXTmAiCvSi9iAyFz8D0u7KkC1sYTuJ+MU4
3vurzgXo2eETwP/M/GbqvsTagn42NqsV5JTEzRXKbhbbZTJGLXs/FruIUXNGBr+/5KCnb/WYjGWp
XKW1rjztrjKkElv43Z6SO2O2ZHBoBvdrh80jwwjmOSI8FpvfDlU8YD75vU0q6s/0PyrlCfsE4HRs
uzQcHZxNtPmKsrWsX0IvAgwqgIH4yWI7nt68Ft+5izEzy/ZLZgI7KdEyO0HvUWQeQvryGc/kt4iK
fnxddK+f/jUd/eCrzrYeQLdzacoh29XQq7tUyhAangG7X5Avd8/LTQ+DjngeLQlfFa8KAQ4HlSb5
H62LtDqcZ3Mt2Cu1z2YvU1VpuVZv2EAFgZ7N34nMsuqAqV0Zg0qHMV0pHneI1kQetEbEIc7QGeaO
2I2B93sZLSbOkVl70IzUy7aHWk5cj85bydPOg5tttYmqI2oAwjvLRZCrLz2M7B2Y0gZ0i5yn6jBd
nP4aztID6i4ETgnSHnmirLtwRYHhg8pXUVkS2HurnYEIo+mEkSiwTddRLMJRv1I8f/H8FyrLWPIw
3EdaHzulFcbjsOABihYCoO1iviRjEmYK7Z0tWW/CGo/kuoeLpt4636impFMIVmH3TNofak89DELq
IwggYUi4SjW0H4PudPCFUoZBVuT69godEJCpsH+7fyf00Jc+WEyCWZanLYHJK6q60BpzaZUxi5P1
2+EhZjIJACV/aey/XXf2HjQKBzXRminkaO6ruhr0bRAwBEiIld4nnkQh6AIdlG3iM7BBYAXLTohR
O/kN3aClvn2TXF4G9cREHIpOgeh+n46yyKmCdhN5Oo6KO9ApqjuEOc4RGzlWFJzDecWYQpdRki1f
R7i+oqqkEBdIciZEyTwiPDliuI0Dp3riGa0fh9o5xa3P4JmqEN5556P+awbzmg1Ew85/4n3L7eJO
qwQztwHhWgmwCGaGSU1BWPfzXvVH3Ap8dVbWlS/WPHgVnjnbnkjjxazc8kB1p1HrvzCwuJ3BkYNQ
cNEck1B5MhxZPfX/QTcRDzxtMhHVaMfyg7VnD7WKYulbjBm8XSZvJanbuPiUq5eiq8la08IrVDmr
ttZmpJ5urwdTtL90aOWifGJu2WEACrxm16OUjDO0eWjINjWMwYxM/N4AAfSgb+/XjK5fUJH47k3B
7fo0Hwt9X46FAf50BN/rS+5jF/A0ofDNG6hflAoijgDcS1n4JmNvoXbwg8nFs8vA6w/D8c2THvzp
MH93A6/mL/SqG/eRqvrU7WWtShKDarvjK6Yg6ZJwqoP+Ge+RWxL5rLfcSPXnLwDCt2AjCWlwIZxB
y7pq4h3LdQhQaf7EcsabTVPVT10Rg8OJICQOiKGjckY4u8K9jGX0j3rWjSp6FBl7Gd5Lk2ffGT0q
gJckfgSUQJrFc1Zl3dR3p7YIDefQJMtS+3fp6ZSBiRrbQb0aVru79fKCfZs6gOxbM70YGgatoAOI
7CGQPT0JysJ/ZBb1c5L3lp0/owU1V2RlArFTSsEX+nYVUn96cSAZwnQNWdvA0WlGbB9qpg/xx+f0
6KbmSYvm4JvVD6FWN+otL0e179JJIj2KK9h5Y7X2EK/vrh7MWwNB58wI2aekYR3GWmQnVQsrJRyh
j0xnYT5/WQnXd9i5UyL+oyAZOwSFigYLLgqAs8HfCE2/UUJjac8ybUTih0MTsoJQ5vaaKBFQX+ue
wTCq45zDWmINy+V/jiwkpw91YawSPswc3SS0TCDp3HoLFAc84gGLyuQMpCe1FKLsTKWHfZ/xyhvJ
tdGiRXyMVunktXt0CG31FdGS4hijzHYjS+4tnfhil4FRZ+DkfKYPSCfZ+N+yp0a4K763AR1VTBr+
XDAW2nGfdFHbxFahmoj5wCxM3iuOxGVGWQ291WzcbRb861sZ+PXpaONmzrJsUXYbDT3e3K8zjewM
FQlM3xjSJ1/wYNbRxolpHwAPsn0PvGSkbP2xus5bsc7KTH7lCY6fQa15QoKZjltOYch498FEKeuW
X5mnqYhGOMWuqGjNk8MWHzN3/AmtQ0bBK9VspLLTlJwAAmHMLjW8b1cPLbkF7wH0S6/Bhcm1Zmp+
fHNI2gkSsDX8aXeqIi241HYVFgEmaMFWCFpNgdTwQ+NbPWjcVEaNMPqloqxrUQHwgZCfxto7VH/j
MqjtLX+prEioygHfyuiWVZIpo5goOCOQrvjLo1L/QeKq6cOlyAKdQnyXsEo+fdMLdBGmC4R3HgEt
kbqT3ZBD7iz5HpC+9SZq6ymxLiXEkrYRcmDYOB3MoWlGOE3Rz2o1VQCGIHcOjMpgqFeKHJE165pr
oa47qRriE9daoc13y0TAv8QLQATsrHqLju8x/06FIHjOGsN6DVpDc5d789ZumaSs7zDGDLI2h9hV
vvdkMQmEuVJySpyw5iYhqs/ksgq5Lffe+1AHZUDrF1dqoBkq9eRb0kfCe+92TKyuCtHBQ5c8lmYB
KD0JD90RPSlBBltor+L/FprWYN3jWQB5AdSOwzwF1RtviMnTsEpZm97vzp9sfPxeo0GKiRC255lz
YpzfM1sCj/wTO8LGODofpon5gYvgCHtt8lkSd4KtxbZpUktzddyG5T0NesF0btCJQb8O+ySiD4QA
b3pEH4wDsUwb4kB3YKn6ZSAG+LrPH6go6ROZD4Htg9XdxrT+4TUV345O/d0dODeooDkitBkSHWXF
GahYPWXdnGmXarnnj6y4qJ4qsQ7fmnc3Zv3fpXcGq6E6oeX6dUlahPMddPsz+HVbpKOYybI/zbUt
oqJHAuzKf1xfsfwqz59NmncinGpNPInRiTkLzqf6gNFmTDiYSCIcKtjf1QIvw0yCN646ajsTjVZs
S46YA2bVNGjGKYsNyqRzSSKkVmAQlV+T5lGAC2ULgpehFP5V+ubxhMTtviu/l1Cp+QDrxmYFqQxC
P3XFFjce5x+3UeiCSxvT+pR6dp6lc9P/aaWaljyhxIwJR91cWmyL/ooWvm9JaL6MnSeIMHSWkKN0
+/QOOq5evANIMRLithX6dW1f2903dAv4SfdHaTMwOcH7Y/buiBkfbGg9RoF+vfcWTgB8WODxNOQc
26uiRfsnyaw1azyqzsXIYftNLu8JyOOwehx+h2tS8QjSIMH4F98c+iQYQdvXPQ468cfnxYXwSQmp
4AB4iVdYYmv7zA+L/3DF66Bpd1x9/HrOmWqW9lrTzCI6iUlmv0IYleQ7LquD0qrhKarwAOsGMa7t
Ny0XJOTIWZAa5inFO2788tX+lA59wZ37mAjQUlPGXevsYuuSGgYamZ82uEHa7Dl7jfCTYWbmu3qJ
KNZNfLHJBDw36owOE4TXMZR/wiF7Z0BMOXLSbbMH92cRhJFwF2jaLpGE6pZf+UN5bcr9TyE2L0c2
U4hiVVtdS8l1U6pUft/2INiQf1Nv7NdW2qI/zXTh9gudQx1zjAl93gammqCm8jbaDO6TedkxU2DT
CO8NZ+HtGFQMg2gi8PtIKwdl1Fsk8tbt0FiJ3Edjphig6ogeYRDfGgjXub6LHRXOaG9tt0rUS7x0
nMNaiDaMnC2YL0N1510huXpf6ULNHnPQ8v4u2wrCDrdNsM78yLn3pl46lGANx38NFAbkIkh2I1/H
hQJro/DXZnyNFkS3LB8f4tYLQU+lHSw0aHSCD1U9K8UUXWUl7hC0gAv3WGndSM/o4Tc4kud6vV4y
ZQksjn0TSmxbMjVvOVPmE6Lvb1Nbossibak5tr1wQcFaP1EVKVN/yX6bOgt73+F5GTRzS9Oyo+CJ
3pgN33fCOv8xG0/9kc0a06z7CoiRISZw1alA70vm1uP342QzNp/um32pexyRKpvyNWT0rrzdvSV1
bv/sHuvE6gFpVRWuDHlj2UuTFLpJ/QTnuPB2OQVbd53JTcQMKG2w/b+PfmKIXFgDcHtsuwgopkuD
n4MU9Ptiua1DlLyYnCZxFXT+YxAQUESzGoNPuzjsC6nITrMTVMZBrayTZJjBTkQNn+QP8LkSoBMp
bVBo4dFySFUJa6R8veX/Iv3MMTyJQIyQ6Oxt+QGSl2yvuimYa/D5BB4Lz3Rt6M1TiNfjll8zNBAd
8NPC0u5WyMsqwvm2sAWrzC+2jgGWQLcaD0idvhjWSCblWrWkz6g+VRydbim5/ivr0nrA0oQhGrFU
OQ07SlZ6uxljWFSjd6iBpuCAhKdNzxO68LCn7tGK2UrkqBj4oKwK+n6UMW0z8hWej4a38VD6xK1Q
R8doSmnUNDBdQTh7Qidegcny6Rdvz0GeTLytsmy2jd1w3OYG2g/vGrHd3eTGDDMqwg57x2tSP5dz
cZE1yNE25x6V21T7McxBjfLQr7ZCrEHEI1/KA+SyP1j/oXBgZcvOneSOVo8G/45sU1tLjC8oveLd
Ve/1DmJzkH6dbkxATpEmTrXL7KGjkwQap9+EkY1ZYUBDwlvBg3HYYS1MHzIx2zFcc3ojsh6TMCCE
5cUs3gaq+iQxJ2qm3Iq14/0SF1zn+y+v8UQ+4zEkaG3uWiSSfhOCh8DvblpxjG5LYXdKLxXMyY44
t4leuLzqGV4O0mTwm1g8InIqL4AmNxNyx+VwYaF3rO4bnWcvadIX+qNY0t7LU4TRnREZRuwh3R8t
zAj/4uOntRXCwpM/utDv0cWYXsQpum3uvLhZ7bc9AHOhxn1KAceMh8p0eJJ93n9fa+cPKTm40Nrx
ONVMqrNRCFUGwv+8v/9SNkh9ImjUWoKBFYpgMzIZYcjI2If6K/xl7xoYNlIKC8eK6qVE6+6FnORP
mnpPrNUKFUtz+izKqeVgtCA3rnl+o+r1L5F+ZP6SzHxgBXS1Z+lGdfjDN0YD6UbQPavJDJwuOdwJ
bCaPe95Wldpl8unRx4c2ECr4VXeGRTXiDeWbs2GgbvO4iP4/cM1kG1PMg/1lcCvZdk18dgrkyosl
E0uMpUET7GdZ8wTRxvYFKtjWD2ykenMhzR7NKmlagosGxnDhiCYn5/aYvuVJPPNjxl9pgzBJN8ue
8W/B5gDxcM9HGZ7B5wZwPDc6tdyUSBwCbJwaX41N0St2Jp7EC+8kKFdvNNIXXbPdXw4nUMW7SOMk
PUsGBBF0fpt3F1e6s9EL6l/HwB4WvwZKwjDniW8rmiWr6PTPLk1xetOtWemvN8gETWTONAcSdL3r
o4bebk7IjDOvdCRcrgYiT7AK7YufUwzTLuAL9BnAGVsEhSLx4BPE3j/JzothstC5ac4H/ZKKlngA
L/0UJC5HtIGpM6IRn5lBdrurmxZq37qTplS4jSn3KM+Ulyxq7qsZwva6z+B/G5DDW53Q3Q8dogT+
oVCsEUrSTMBMwYDBEzsvBBOpO1KurDoZ8BAEF1ToVVI/mCj1z2snjlR18e/8r1OQjiytBxqPBy9n
5tSTFm5v1lEHS9g9CVF75oMC1KZ2Z6xHv7qf7dVbO1h1PWVRir9NN0Zdxgs0a1VjZpl27viVuTiV
OGAQhNr07cebs8s48lF9DdgkLaCz3fx5rPLmWfLyRp9JUFu/nShkNjSgQ3UAqwZMDSAfc4UsjGy7
VnC1BCmfRNzhwNsmRPXAAf/+Ect9ZioHVD6qysSxDRTqODP5u90sS01hAES6k8sKwjLHrPgFe1Fa
YAPsjtVd1cawj+i99smgHoA+Dix2miKY4KgEJS8IAR2vtfGRnMrLt+WoY7qtdTjI3BpuI3VUFBbI
zxwNlL3fHBFS8PPRtAWEgtHVEz2ucg+IxvPFMIfIRAQ9zdIkgkkW8YnDpvTtYKCGt0OJ29KIF5dV
o+LOtRRFGwC1OP7/8Fy29gMda5RPjQXgOZgaHLztW5vQgq7Uu420vnMf5CEZiRnw76vfkjxoIS4Y
0+msQNwy2DNk15eAl1y/ALX8FO1wnS2iW5Er7Db/ZiopP6pnaMNvj6LpoFFKcW25mRSDT1yzVKVS
C7sLBR74GDun04/w7O1J0HU1m+KfaeatIsvAXWY7/Hd6hJ8O4tkHroQR/M6U8BaYbI9vfoCGweFt
oICEmes6fFcL/+F9OyVaBGoF3H4Xpe5QYUrRWretO1VSxD4Qd8ZeuY+M40kmMH2uMcMcGT+c9iWP
J9Y0mPKJAkQH+DjuLtWHn/V4nOxjcBuib/YtykJUDyJKnYsa3badhetJsRQa8PRlMl2xDaJmPIfp
u0m2mr6Br9zjg/MdC2+zK8z+uInaZ5lVr8Ccty7uI4S5yRb2PRa5P1MaSAwY8/ddn304VmkLuzM2
DrDF6zj1dC9vju22zZMmyF0UaAvBxO/55Fs/PUVyBCA3+OlgYQuupstJ3Ym1oCh5LLrAxXIpwJqM
Q9P9QBQP0FHtqJVtcM6khW6EHL9l3eCRFa5nFjeGiEPyrwDpfQ6IOYK5hWdvUm0fnSXEdMR2FokV
AMzz7d7z2mEaFiZ3LoO72lPn6PJfJwCad2kNXfpSUWdWlfqHyJ1RK1lyDrdDgviKnhHs+3qOC2F6
0jObZZ4uUX7jK6UJCBRJgq2ETjxuv2lra2a1GRrbsWgcjJh3Pk8zmH89xodNUHDVnZ+fnR+uYqua
4S4w3lY7MqdC/YvTRtnYVN6/IsOq+ax6ryIWX/UTg4DVAhbNnBrIHLfSgfBZ3UZZ78RHBTIgc+zX
ntpRnRXveVcVo+g1gdTsY27RNF4mpB5MbvBVKdxzWOCtECTzpR9//h7F8ostBpTMufIX/DJxQAq6
RJmLIraRCIfeZKKuHa0b1qY17262+bk15Aq4gSleVwQbbx0YOAZDAtTSn4PFc/rzM5+HL3NI1mVz
V56mg0nEqDUQXehhXVFXQcvrsjG1kSW3oJ+anklPw616f6nLAHrVAbYoQqy4pGVcIM/vaBgLI8BY
0+52PUfZ0RNk4MqTz1/NTShbo4rXrxE+LQiHQ/n27FPYI9pdRH6cHgMQ4n0zdwDs5/3ylZWUvl1d
5h3kmbT9M0Nzp2r2bWYk1JG0fWawaYXEiMacy7bHxKOFOiY4jnlM29EEuAJ3k7TEipog3CH48iz4
1ov5H0jlKaXBMvOmAoJCAGbdTnsV28nXywMClreqsM44g8/O8yWzl4bKgbIvvBSABs/oalQGzjbe
3CAT4POnK6Mbm4NwtUyW9foMHH0tMCUvPaDQBaW9RZARDnuyXeFlKefDop0ELg94bpKFqT80nCov
GHdGUN4z/Y0n8wUW33QGQtjHuqoG7syWs1hXooOZb50dJnCNRH1hoFscyYgJJOTNWejRg7LM7Jw0
/f84TgrCBrFNkLY3Tx45ATHu0GZkLXAipwLn0SNoKc4+4eD7yflGdAPvtamc6upa8zMv86355957
rZjNgqbBdzHkQC9zCUsVjC6jyqtjeG0UCj5YPsWrBuHaI6r54sxzj16p5Ycw4WJ27yBq7n6Wqq6C
jqpXdK6S+a2y06ognItFlFaiyutF4zmlfrBfmSkk2UC8YJ73Jpp1/4rany66huWNrWPBnkWkdmjh
aUEQ915RdhtEI2N6ThvHoxf0tWwmPafrQbsnYBpjIbWAfUxnMIKZeCbyTQV4/nbeVlaJuE3CtPG1
n47/ZESww6TOQBxNcOETJ4Hww/fBIqcGp4RzdOLOU97SIUc5TbTu42DtGdOwxfRgnKGBB3AsfOkr
PagEs/Q+kTP6qUuBgu1HA6DFi7HBzYDrKuHCfmi8OKYr/7xZvP32dDBrWgKOz1uaRgZKmxfJzKQh
hmb+G/yRoc0t1V9zLtjY4rTcvUr/MfHXj0WQTPqrPPTC6kLGQa6N2UBHN6g+b6YnRvHmmv507QW1
vzSeou47YRg+WmldE2CprUeQ5+11AB0K9yCOoJIWLKazSjTIw/08RMcwRI5zWxdOO5tIJ3aiS063
F5TykbIbRhW3oo7ye4NBd7H2BC1swbOBnIZQuf7oPJGwA5gdEyt4qR/kT5TaHUJcrSRb9/Ceq4gu
EWtWcOlmASjrDF7X0jnwT+h3zo1DWJ6DK48fSvZ2139jjuYMSt2SBjlNLYZkX/s8wmeQTaVwLTGy
TCQSxXvdjsNyu0Wb7ZDZrwoA31nliY+U2f8K6C9OiJViViGPY+JCQhtLwBB0OdsvVlJ2P0noMomC
Tv2qb6L+aDUczvvdP5vlvSH4tsKabLDXZmc+lRNVhUgjqMQqmm5qjHhjMeqHreA9kIOqyHoDh2/0
4AgZUSrBiGcCjS77mR4TVBj0AztqwatZOxv6Da2qomk0/1eWb30oX2uFbHInQV1hbs2XCjZL3yNw
oIvtd6dcx8ZNXk++LMHBOF1+o3f2pDr/2EYKcFLedybFbBtJhwr/bZ6blrYHxgiOQlWZe4lSW5UG
L/JtNN613eDZ1cOTKMS+35Qze4KUQD2QN98dkDA++EoshQty447e2Zmu0dddogI5W/EOE4nnUPYn
puVwZybVv0eLYgU//LMkTPLwpTddtulb65Xi7Be8ZlmINaDLm+FEOy8f/oCMU2J+sFGBvhc5hNFo
zbUsriGB3Z5MpYIjkkX3SpFDVHojaI1ugDWfFQ1oC+OZg06+v4PDJ3tBJRWpDzVCnWgBceUS3bqA
O2xHQXMlgwH/n5u7NOMF0DjHRSoQcUwOZO6DqwcvZ8O2L2Fly0Q9MA09D5z9AYm9hPDJ37ab02KQ
XYNr0ZBZcG9zfpgo1dHSBG6EY0tvdVa91KQmm5J3z8f4xFF8uUTeVkJoCakVLAKk/gk5W77AC5FP
idLN+/9LK8kqnZ/qVPHGfdUdR3v74C1xJxBqYg3lnJp9ZvILc+j0jx2jY/KhumdwxUUvcxXr/roT
Wbm/0zluR7m7uiRRgCwVFgFu+CsThfZAYCn+FOq4VsKQTFTOseOs/O1fvCASYF2cbRWOihXGxFIK
SaC86sf8Yrry5HCBuqWxVnpzFbGPZB/MNLAlR5mlE0DFD0m7a5WEhz3MX9vEYdz0kGUXLvyr0+z/
YToHLK2V05WpvaL8GH9Y/mmVTOCsHYzHkh1rkqg6S1kAEMZLtFPhfCMq1yxJ2Q842D4INcf5vemc
smgtvZj2EXys636/fQPATFYnOoMRqpXncqKJeZtJmrFOUWhI+FpSa6TJJEMAdj9OfQrpOwRHfJwG
WvjY+gHLcDXfwrK9BhovYBmI7ZXBkoJerWCJVssHdAGutcWy8XXYuGEq8aj4jHI45iEX8DFSCB8C
rwTPETrqM4W4lH9IQvHYk8oJCWH26s2s4oYHuI5fuB/y96QNkrbhI9ZyX4jk7DW7uDR8sUtEp7CI
QTvHxhdlao3wLr7FEED80t0BreLAh1At5ESyQERvmz0RQsQO4VSz6pjk3LN6xhyRyrQM0IwTvcs6
mPKQSsHq8oNAOCDC6ytE29Y1sdT9MLBRRZKZva3iAU+Mq9yYKR268kDb7lINBvfSz1by70zZxA9w
PSO5es9PMW5Uhux1utBBdyf1qnjL52c/y/m3JbmztesgdtYjqZC4iKlyhiE9aSjpmd484Z+3jr6U
r2LN0E9Kz3DQF6bFIsD8vKxGR6zDnFxgntK9YBnqGGN0z8sTe9JCsrFcrNOIbcL0pl4yULtOVuPf
dZ2ZnP0fCUy0lqG3IeR8RzSHC/FCsw5un2biSEFzC8nCm9A1qXUOSBArRDrAm46LcA+H8rl9GR82
mxddsR/wQdtUyJ7GWFSi3HA89IIYAaerxY3n3lXJQXigpXEFXdbszFCLFsD4zBCWwJTTdocimoUh
kqC5hGfU18p9TDqsxzRR+xSK4lCyvy5biS7ImN9NU4mKG4p9FWJT09fhnvr3JRGcOOELzIMPNdwR
c57zzUazby2R7+8sPw6B0qmuB4omzWgW0bjb6uRQuFDAWPPCssz/i1szBHVc3qONWXqOCV5kRphB
6LB4yCLRk90LUhMZUx209nwHLatzHHazJJLQvJXOt2pqP4MnaVzYjTJodsyBoY3hnHkgb/iOP1qb
+UKAqQVNKNwVtrnfwJJJHcvEXZKFRgI0W2+3Ei3D1ITP5OqS11WoW4d3zr+VkFnNaPA4FgDIelPB
080iUk1PkojvgeU68TBARsKA2itOfZ46j7oT4bQIuicQ+6BOEoQVLMZCUUPOHQefh/zpiR3//Ec0
Ysr5XZm3dNJj6Gq+qKrFKeSnsk/j3L57rZVB8e3SRM7HF9oT5qtWWFzNaBLhn/GmpCzLrqZNhY90
GMGY2sEMd/uHTwZTZ4lLSHn5TgeMIzvSXh5fms/3fpyEZuMSi0SU87NZYCQfu/4ll7+Rcn/aMEXI
mjBCTbtfGAztKNu6afgyz1TQDjETAFaTbdFvWr6uKetjrJ9s2V/1EOpLDz7mNZ2DTSYQWx/xCcNf
dty6i3Q+jgo+mCZKChBvgNw+iMGTXFVrF0t02I+8o7Sw16/+ncKnjRxCOVt4oTjlXzg2JyVj6BuS
cpNIR4nFNShRsk7n37aOXGNYLwooztBzsv7Az1xvpZkJQT5bIe+Yued/4NGPYpTzPuuPv28nckMj
ZzscdeYnSDeFdvKXygF1x/daB7Q2p+Ze645/uF/h4jDV2fQNWxQnM4FtixPC7k9xl3qey5olwN1N
YJJY/lxCAfGEbYCS0iuHQrsP1fRk6q64ur3jfQyzwQ01LyFFSfFVVmaLarNk2dmB1Pk7c3ZgDDzA
8mq1DukvSAPD94YgPALdKF0DfaggUC72v46CMiGeXq8Q9e0vyD6srQs3GuVHyyjNRMHlgNNzCCXn
SG4HsYD+tjS2Gi8YKpGNl3HQVJViQb5ZDt1Adk/V1/sOKrPPFdzu8QhlrhJXN6vDcdX/PXBQTq+P
sxNQwxh5QR8gFEGaFqs55FIel0HM+vcs4G8rAcPU9xk2lF4UM98j9tDZfmlmVKkPT4Rj7sAj+HPD
QDGZyT9Eq3aXbB9vqSVQ9/kz64/SfcrpPHGbSmwLT2MG6IwWVQQqEBZZblXi3/61URuLCftUZfaq
uoOaPS5OA7ehK+O2FMdshOk5rnlKPdEDQvVu8FscOmJOLrEruVw7U0m0AT8waeTMDwuT7aNEaHdy
gS2PAT7MYSs9Xer5YMMtwUoY+rbQq+bLkF6E8XKUocH1lUC9zvn83FKXOv9q7DxThP64uyZz2U9J
eZ4kK6vMSlC+Uw0t5MsACCkZCQle5J0L8cTwJ7N9q6V26k/F7KrA0g913T/OehPG286euuvRqU4m
Br4skOM3njzuBoGEQ1RX+qWclTZGwwXhC7XHYOhiIq/6tbmJEZsriJSsyY3Nq1Qru0L1ko4MaiyH
JfoAucr3FTILdUnKpIrkGPm7HknzMvCrT+KC0d7V3jYecD6EuXCrgLnPBVNUT0A7Il2gdfRGvwAc
+gp+2fiBnxBBOmezas6owzXZxoYKr9JOcsmFwJ+w43MM6gGMsDkPyZP2W4FSFbV+cicRrB2cF1R3
gdJKEMFdpbOV4n+234RXFeE6ePFcruKE3cQP0RhVCkM+68NtlEtT0EedEr5u3Zzr6UwpiJyTJctz
kbqY88egg1SNkqOn9AKOrKLUnzvmXhbE14slyxYm/2dKQY/Qgwvxg8WMVR+IhIGWksjC35EeE1eM
m92KcXDanamWLmITmoDUef4ovCUjC2wrIlwMJ9BJKuhTyZdGAh85mwtFTM8Ab75yHrHokJYkmw1/
rd/hZWnXdQuNuf+B8qYrXGdeSgzZgIxaKX+jHm1c4QfUhdICa5+CQzAmoOUkOjqqBVUylNg1q+SA
c4nywfR3+M/xmI012MMsxEVPl2yL2/1RYkNMyl4Kwk9210hNdBUiNbOuFn2e1kjvjERlzNcHzTZR
l9xFgiMIeaeUzWU5HPEAL7cE9JZEVA9s6XmJc9nd5jOJrL57mGJuPG6FP3Ss+K4yU4R51gZyGA7T
cDw0ZKEMCC95gMKqXKppXRSsavpthMmSYsC8iIw3SFyJXdZSb64cN0k+n7Vi4KZqTUlhDa8n6jnK
jWi0SW4zrZ54S3+gnyloK83KvwDV8HopevOJJlMcH6L5JhMZcNMthGwUqA72XBkUrh7c00ZxWuif
4IxKFx/3Er5yf/ec9ovIC4MEKBZmb4KjCSM+1PkjRRTISGm7MNPpTWiPmeBauuXCo0PsD16rZ5mH
Fwii9jMAMLcZBFftxXWWurOljZSuE9ynEaRFCXe0veD2h2ZvJL233IVt3HsDm1xt+xmhVmmOiKW5
sghbOljMdC//yPjlTiehKwuKaKdr51yfELmnFDpRegi8G5+Z/Z0EHTRHO1VofOMEMkdPFyJ/Uwe7
qqaiz8M1h8h7Y+8U6dwROG+T85F/Etn/sAGtUzlzY+2Q6E6NJccXxZ9HpxnGwGapNrZ2jBhzl1+c
td9FWX9j1BHJfFYPxGFhbRvpcKAJJ5vf/JWjs/SqBQVfC0WxqD+IuT41hCg3DrmaCPozmAsO4Sku
l/rA54i7tmwgrngJQeaQ4syPbfgBXiTiIhOTKw8VtcGBuawTJE+g6ZyvkKRUD92tzmV2HexqaMmk
91v/lAu7ZxJH9DJgBWJv5mrEn1AG8jhZZLh58w+7Zlttj5JM3YBJm23noArkbVIjMFRfzUlyYODX
lZH7dLr/rDe3iX7EJAKlQnP4/H218PHV82p6hNGmCkH4KuFsdImUJm/Q5Y+1L8co9TePXlaIrUTR
S97OYcxp9kgc90C1zw5cuhDPJklFFh3kq13dI2i+FQvCDMre8CiY8+Ub6QoFsJpQHv2nvJdcLNE7
6p5MT6hDx8OOQCraanMhm4UrFIA7Fm+8UzKQieO8YavsYNDWiA9EwCTRiQ9olATkxjbTpDdj2MEb
8IATa6iKG1H4oCTzPB8uh6vDLTibmKKwSHftrVRcJij+m9EyLEOuLgOOSblBhoRw35a5ya9T+7Ra
HIDoTMvmvruSkHCNZ6/mN7GSccMAWR4HiyHWv1koYQQZFIX5AcnJ1xJ/k2ad/L6xJqEZ5i79fYu1
OVpfxMGm3Oxm4N6Zx1oaoht7dj6MrJx8WDgq3S48xLs+B/T1zG7cJ3yc4/12QeU9w5q9eBe0tjIF
0en/14+D8p8eety9lfF15VfeX/wt47miHzGVpREtLjz1UaWHjWhOdvQbdRI1YHeGWdb+27mRZcGs
2jOJFb5tcZ8tW6HgOG0uLIp/+PVJ9oJIPK9lhh0fG+V+jcoh1dPSjxEyjai4aI4aat0bo0kB5WDf
npJVwZPDc9+yUMjRUPIO0/hxwdddQabSI2wrFmKI3Vxg42wTC0EItEu0re7z/nWf4xWtyMQcFRyr
gUz1MNLraUV2jCLWYJJLW01qzaZr5s1YkOBBlD6CrrBBkKlgB4d+HsdnXUKJWE1rQO6yQCN7CbZ5
H/3vuAPkO41jXMjAMOOkVgVtgASbRrEUqzJb1Gg7LLYAIL4yNcUp9lv8EJpm1Bteu9Q1ShBo6g3H
pohqKIbEbQzizBiF7W3WVhS51yIJlQG8uFqtgBgvNiOH0HymqsVstypnp2tbGu96l4HYy8AMzFtR
y8lPs+uzMhS3iS2CMKPPxhLWzDIcqNtc7bcPLy8SV0hIaC4CeyPM2HklwpSuEhunQcWimPbhXjOd
PVpxlN9lW0HEYgO7mPLltF0ldoy8nyQwcu3L5yCG7qHWMt/CaPZSjKKm3SqegzlHFKb0po4aKWCR
bC5BvpP+FnWBPF6SnHK1+DwoQteYX1y4fcaa6v+Ia9mRFZGr0Kj7qwRuXaSGyZflBrbNlxYswoFv
PFmbKMmGRn+Cs5xGaQzO+mUnnIG54FZpGxO4F+lqOowQI6ZlNLhMYywpjuMB0IZ4sYAjHxt26L6/
VCIJu3K5ezUKiUHdGEPdJgX4FYv+w4yXNX/prceukOiqhTTJ/R0WP7dv5DZmOwD1mQlkT6gMfXZY
KqkDLMRtSc4GU/+JsnafNVVTCox4SK35XgtMZs99ChaOzXALrFu0r65AU4szGmj0+KN0S1X2L2i0
QkGaJ4EkGbe+zldkIqhUAP8aeWeWmXxDcK5uNsG5wpDAhYh6RZ+dKb+WMVwJHlbY2wcDAQeXKkTV
8yBGjxO8ZEKEwp5j/QjDM52b0WqE+xCIGbqISAQ0H/xYkIpPl4w9a5TmNdOdiuhs/wm09A1cr9Tq
M80+TZ/fhn7gDjaWWeH5egBPDnVYAh2oMcQMniRO5++abvU5Ji25DHPeBj0R0nsFR9YC1l4RZ14q
omHuD9cGAGzNyMYtX3UnP+auLbF1OXkugrKn60iEl1wgFg3YMKtB3nePNmoU77G/tQIIN4RfLbng
MsUfZoqKLpv+6L0kcWYZ+8/iWskD+OUQR3y5V62GEVBhD57i5e3N2zPsA5/EoCLHmBczhQw+2/PJ
FRmt0ppfPBNKRW5RV2u9LoyV1e+3dY5aGj//FPLCJyUmYtq81gLHDCUaIIyqLGx4Ao9SYVHB7LAb
x0QpC3uiGe5ZeUvLDmgzg+ZjN4+pC18akxxmFTjjvyuTnsHijPegeuxDp+GqnAXlsSVa8UXXRJcq
nDe7Pf+fnKI4MstpZcNlCbKHllbolR+QTTMP546bxmgzn7uA/1tZ3vlR6OW1kV9IwvA1FVqBH1le
W16QGr+Z6F3sCnEPsg/dVNxP1HwGp7i+cnbpD0TnrH5wAznKSSG2j3ugGxiJE95L3QzllYwFENFa
iLYtgwlWF+LF9YAezbCfkEqOaVayxVEjUy3NTIBHGPRSNu54i/Fmji++ToTz4nX+gOhnbBtNu3Wi
yetG0jjNHm8d8K63n31nTm9Dx7tbyoklh6aSSU3vRBG7jieGE0Djk1bVBM38EiTmWGcIpwYlaJ7+
1EN6BJnd2APWnI5B/QW4iXyiw82wO8Fd93o2HEAB7iPWpRTED1ulaEg0zPXMl3fYyUJgpY7MBqkq
jF7ztZ4/9HTmfinyrf3C5auss3yLrAz9EISSql6mvzGYozKNCa5YytKfj/V9duZxGsHul1PoQhyn
8aKkEos2brujWND28JnfQvUhqouMIcl3MC4p8v8gmv5cdHfHjimlomN0D8k5K90sbwqM40ZLNjdq
NM77bGh8c0w9ZL0dfi0uCgknY/lWD+PWyPhMrAi6eTfMlq01aKZmHm6BAAC29DUqeTsXOTxP7wr+
SyO1Qzbjp+iXXoV7Sw9A+Xy7i5WBTumzrcHtgKwQ4cxgBWX2xqSvMRvz5Ax8PeizmNImY9EWHFUA
cT6eOC2kUN14ojpJnDF/OMmwJzB/fjK5DHl0tq/ZhXxI6nGwcaOc6usqBNaf6ikDs01n/BgX7FrJ
517Y4GywSDv+uNA2dMPa90SkSv/fWpTkIJSfTn5eDunxfSziGpiON2CjnEj8F4GbApLv9N6iTSLN
kq8nhYveGnVmBfu5Bw22GbFlBSuORRjSPHekbNEWJv+LM8o1Ry/pab9FHsIV7iuoUZ5MhG1n3Q6f
U6YbDIC0J3X2GKj/wCyZfu3DYJIBbFSsQok6v1t5868oXxHXwFbqcz39xZ3RgUXe0wm4qqmeyscA
zNUtQpNRW5Ull99X+7eXBHctxGbwffI75bVIGo4K9EU2kSvylSA8crQCCa6hxMdXW0vQRWQLIfYL
dZWLkABoSfc4p6WUh5LN2fNOH7jxsVASBTAnjuPE9Kzs8k3lZVL14PtBHj+PdanSW+YMC/AmOMCb
t8uEST9E5y8lMjPhFl1M6OrmUGyQ9jFazt/uTnFZiGlu2XkQ1gjQ2pys09EygYpsqK4oderheV5J
9lD7KgCSQ2Gy/QYEYAJvxdNI85v3C4p85E73RjvxMQZcfnYIopyWPe/OtmG0mU4J9MkbU2Lc39dq
lEwmYTiu7O8x00UYvHpIBhDwO7r1+o4p1AfHOA4pDgRmxTq8fcPI95rJ8jc0Thr9UIH9sJ3mv3UW
7NW0x6xYf1vLRVsjoqwjdAU7hY0f17E4QR6WYhg9k2otM9xEhXFMWZ8OXOXYU3souWXFIMie0ETP
1jMO1Hmvz/GBPTP0o6p7rm1VoylXFIUEUI3e4CyHmGh7bsXtSmACDhG4tQwqfjR0I6Rp6xTzbOiz
bfnZYG+gzBevlaTMh3YrVksovwOG4mNorBpNt73tpnRyAsFxzV7T5o0H6EAXH1s1a2TrzCJu2xfo
XL6JA73I94YbhHX7gwfqb77e3r65Nlpe05ew68lXET0IMIgURXqbAHeihabaQjCNl5DVtrmfrwJG
UZgP2mK3BKP9fN66Hde3q/jjHAH57wvja7QAUHfPWfylFEsFRzrqx75UsQO/l/b/exbGw27B7AeX
I15J1BJu4ZDpH0z1tFBlK0j+C9yP1mmMzv4ij7fYlSB3NqbuhcneDO0AWe9AuCQBYGG4oIkr/Q7x
q7ZoSsH9sXNGXEA/jBCjslNfbsSlUwiOmC2E+7AUAWeJr4BpR0G4WkWDXNdx4oiAOcQnS0iixUyA
qdoDTFv1IHq6J25C/j917/t7Co+87AaUwYoFt8ELCcn+LLxNy29hEUESSHZVVsJlucussUC6Im15
bCmXV52ArqHmjYaXUxvPbyoqZeq4V54fUpjlkOt9QbNfXgrfQgzRVHIAPn/gkZhK5AbuNbppLfL5
2nx67W5eSxjJ9FKo9RpqpnNcBp4gUwhvpf2E7YtKHY1BPk2BBT3TIR97yIG0C0dv1kxsX06GtEKh
tW7WLnJz+TUCQtFR1JHyrkrecS1/11irdgbnrrqQsifqsQ1vWiX2EPbFHajClogrSXRx1/xs6dzY
JalLA693fXPoNdFgsgb5KkW1ETdtRHzL+6eRkRZbT4rL3wMcYzLyZpv2s7fhbre3/hpvle77I6aC
khfDt/4kYtfVB7gif3VVZEwOQyMBmoEu4fVc90v5Zi0m8a8mN2ZyA6zYFXEm6v8vuuYHWT1A8tmP
uufB2VRBG4rF1kXLgEVc0L1OqoBrDqbaLfD/uw2e8564nCueIvAYBjNsizXNrj5n+u29rGh1upms
QeSriMpJ3pl3FqK9VJ3iXWxz5oHtfw+McOjiFmqv0f+GrVbd9r6xCic/YkGb5SFRV/yNb2dT74W/
0qqMiedMufiVQr5J9UgeUIoCai5NT/T75GIjFim0/FvrCTsqJcJ681I9BUHPw3OtHualubyXdzq1
qhmHhMEgrmgdihBvhiIY0atJMO9O994H+7KXZT6IQp9A0rgWTBaoCk6Co8T+E+5XOWau9P/j28lq
+cUnd0sNjg6/IojvZAh85lkpQMz1xZnF4lTApPCMGlGm7icyFRBvDsqqWAiGOLMjagbivtl5JDc/
jaM1NZYeEC2BtxMBGbmlSfic7hisL78mIOyp1I6Yzk4mZUuwkelI5EwfbW1nxLlgFw7Z3/5S7OSh
EItLr3tM1uE7urXDCMGmJoNpC9/+imPBBM0+oNK24j8gyP6L31iI4fzbhot0KM7lR6CER3yxGmMA
a33aW8zGaFO4hwoUWaC1CvIpn5ar/ubnTGKWO9kHZXPmX+3TfAJUTXz29JyP1gJLfZBNlXQd0zMS
eA0dEkduJm0e5fn0REvq32w/nePeYgwff+CbO2Rybn1QMpTw+hpgWZsWEuAcbXtPuyFj7NE04kCg
yb+ZZd0gPeaTCEh6zQoal+8TWlaWfDH3y70apvth41hRyebdFUM16nQgny7KpZmE4uSaqpaSvgkX
2W4bpd2HQ8qe5FHsDnmZk3xBbxmDbOg0o0VEHxPjmfsUJ7/U67AYoJ4lzC0fJFYtVgtJ4THr4hdO
X0WhyQGnSCTYxXgsOa+s8dVnb6jOvH0Sq7ginlVD15eSeECc2iszvOyp7Nt8MAqXrqVFBuf21fb4
DCtnuEUWhQPstpW8edDLVufC4Od0jx+EhSfnPE2TQhqfiqlU9q7/V0pHy8gF6hgPhNdwJY8/PE24
ujC4z/d9mHrulZGRf/IGmMVM8bdzmBK9sBqZOZaBxO7rF6z9fBpuh8unfONpMWKVk7eZe+XKsmii
zCv8jZH1gX7+UnqpwSw5rZ6Mm7A4XU7z1p9RedfybQxW2KuZGO4ETUwgTpwGxLNrf4Xk1OkCUq+G
dYtAxCgkl6EidZeZUHlzLN6Eo1S16tWTz2CDFBjUgbglZGKl+3G0dwReK7mWEokTEyLIv8B3JFXP
pJibHAgs4O+P5JzSEMqkbsGy2DbWIt3Yh+vfZHUTu4V6EOkTm28bXYrqURE8Hm2vUnHUZBqYLK/3
SXwthUgDadbjzlgR7AU28uUif0iK12dy0DAz1rpI6u/qeFwmWM5tH/K3VwLphPvs0wXbeaFFF2up
Tpe3bAyjQFsVPVqn6HNktiJt/ZUUr17uVT8x940p+EqmpNOOYx3uHDZlNqbO2HC0XPzpk3Mamz9X
w/xQuVw3WSW6Q7OiW+6mITy4UVFM5aRQIDeSx4KEZQgRaTGt6LpAiHtTsXfprwM95m+QN+kMhhKM
eYT4vQCKjQRBIw6gkJQFrP77ddDg+ShcSrwdRkkNztWzwk4fudXNZi5xUS+ozTHraw9i5xvIkap8
FPVE2uTJluNBLK5CUhdj2T+DH/hJa45YXQV9Y3JQfUHWFn4AnccQ+q3yEb+Z4JKP44K4wzY1KNGC
ShDUDC2ftSTIHnngQ3xiAJoQMgib4g+4/bCIVKa8XSyiVBSWR+zV8HL5iihIydgeoPB2NMD4P03E
qEnhvcI0gsFseewefjmqa4/8LuP+4umb7tEVLZAGKn/j6MH/GVRMQcYhkN6V68Pexeys3/Bixawq
vlX3PMbWDVYlYyL1FnD75iM0yhRmZyOvPVnsCLgoTI7O1tsZ3YHgRg4bq6YFDOBkmgW1nQH2yJan
GhkPRuvtEFOdgobD+/13YgOas+nxiwn04fkscVSHJdrWYxYujzAinWPy4COfeM8JhpXBpYZr7y/K
EQarwyJlaFLPoWykQJQgHvJMUmwmx3PWSa14+4y10SIIRBAXNjmQaZ/8HNjt1jHLNGj5qNOfP0LI
T+YDB1aWV5Fu/JaBEmBviAPVI9MGT27nmxSJ7Qf/GSlm7tcnNHSXQxKHEWmRM4Y4Zp3BbsXzCxxy
LeUKGOck7vkJzW+sCTMuLtgg+qkRdvyCscVXdz9+PZLtzgy1BV1CRL+wk2F7Fs0zYBkYn8KV4EM9
ZstgNNVK7ezHbmLkEs4TDOZSpGV1vLbkEWsukIKWXvwY8Y7RltCufaFee1lzWpyE1w/eRWvF2byV
+ZhOiKv5CttfcskGb+2+gsx8qtiSomZDfRfHqXui7ZxwFWm48hHm8OMKwdBF2Ggwq08WmEHlr0Sx
eEquyxGheUVoC13Gebfu2Ot53cINy80yJWV+q14e2KinDuFzO4OTdzWafiETwaKlq9+Ir2SbUjju
xjSHs9NYug3aP+nEQAUW/0fjEZJ/Wh/+3n5cVXshZMXn/w1h778K9fmKSe23DPDYTnYLA7sYkMR2
PatrXG9sU0n89y6uK06fQf0xH0wOLS48aPYqWwBVHo2zUa204XDAiWVkGq0WwGQOrbVR05Q5I+9E
BRKbnsK5+aNzWl3hnpqLkgJRtFmrFS3YXrc08V5h8gbe8JlV1HLqO07EK8r9/8X4btpdQZWq6Mk7
vQYWHbd1OTWPKbUEmIdys+KLSoX2pFcIY2gUOV0FSclsw9m9P/7FYuaCNVjNVsmxN6bouylmD1r/
Y2LTgjJktGIhASx7OQZQXd5LI/Db+kCORnseYeofooNy1RSzE2VedjZLgaYXcSe0elyGlQMUqBZj
PGSMHS7i+oTsDx6YZgGYblD93pzTPAfQQz+xtXraRR2uZEMHzSOUye0ePSigkLSLT9dV/0VCZsxM
hBonMgb/lIdkG5jC/OGvJYWZHG5uGeyOnBphWV6Rzno5MkcJFCDvVpFibx7PTYkUJP6FjRuzTRvE
tY2ppeA4uP36guJft/JkkkT8GAcceov8aOUZkg3ezetNp+SWZA898l82oSJhw0Va+WkKfKDyT3Z+
9n90Sqp2JH/pTFUXRp0xKpy1OQSZZDEWEPvQ7JJJCFwFS9KupFExiMN5lc2NzvKy8VfnZsDWuzwy
cakHCPMv+3/MkNiy7KYz4sMIADxzATosUpQi/oLpeWZ9mFOps+HbiDQO6QIU5x5kSYWYqnYFk7kz
r0JjUW0NU+RpUOjPa2BX2yKCvulMaa0GwhKpWFZnvHXHzV3H1/kYDkZv7ofdRxgE/h+uJRiWiNw0
j0YG4o3fyWRkeu5TKdCztF7sNCwYaJ36PCQxX7ewGvPgnY68eJeqFX3R6vZiIm5jxAMl65ouk5Mr
ZM1O0FbbgYC4mDZcG6np9iMeG96qVd/Auam/wlF13eUya5KXoVQtEeUxUDfFGwrAACbAxSx4Jy06
HZWy5DSwHraObzejtA8/yMXpir7xJouOpkbEFUhO0qNrbuvU7r7IUwVcxu6dHJN3I9KfUZUpgTCv
mAru/y7KxBR9g16/vZF/UbWBn9GhyeNvzu824KpgWGei3KAR9zwHzEjVGjHS9l7t4LPypO6w74/K
hKiMctV88Hodpr63UI/cRD16pCFyLFexLWuHMcogqjhF6yjtsbK8v0+Lq6U4IVFKY4tR9NxRan6M
EQlaqCLaqGelCBdRRhOIACyChEGaG+kOksG5RLTDkYhiOPFnkoxkz0/xOqyL7Qe29kLxI3cBxe7M
9WVp1bn1xpX9LbX7TA/XxJzQ0t5VL+RD58/+36bXicVS1T97p+HKtZQDz2JRB7EvQTG7Q5km1mis
FyrbqAVnAJRLqn0SaKaeI1SN6ANggJ5y+aPvEKmC9jcCNx532n0GsJcua+oqncFic9acunIKez6S
8Htz6EW9t//SUjvoBhc2+XI8eKkZX4sfWm96TaJ/GT7cusxkUyRpizm6LzE3X6rzUaoQclB9bDo+
np53DgF0uaQQEaqFiyqq/0eYWJeW73cgKXg4opber2Mhx5MW0DJ1Y4sr5iklPmgQ9+cx9mAsaYHZ
0nE/y9YKubbn9o1bARJI2/q28acv7Mug2wnTNMczplUYVii9L79u86gAXBkmooel+20y3wH5RAVJ
YWyymeAdbAssy9puzfnB2qU+i9le+Brqyu0VwE6jGi2DOLnqT4Y26szG5JvmB4msZcExbDL6KClY
w6F3fXL6j9/WYpdMHlHvGH134D0d1jw/hkyjHZEV4M04uVb1TgEYUMVLcK84t3p9I4tv+EBdsdMV
p0zDW/hKwecLY0MpqEKgpU+n8X7eULl1ZrJ9M7f3iJ5PsmLSboHCvFdFYPB7qhWOisbzDoSeRuSL
rdOVcRw2E3dgKFb06UMcl0J5b1TBoazj72hGjw0C4GShO/6jmIr55L1lnMGyFEjz+L5O4E1+18vB
l+KEH/DtdiGVCwWmKrd/9ypyBLOXjdPLcXJPXDY01G3eJKaSDpHeySlqGWERm70Bp8+erANCLSLT
y0/gtZLvGvLtOFL7bTaXqHtK8vml9IjEgXMnRTNj/na7jbS2aDZrg+AysrG7vlsgA0a9Jc5CJ+GU
zHTRy/NJIrt4Ff3236XQGSr9duC/4+V6jpQtTH1QcSjqFO/dZcfey8Kqzz/itRFp41ccK2MW4FdC
lXD+JIEUjrVn+qTW0anUoh1MTVZgdWbvkUrvbF44RsBJqyUXy2YHAkr7yeCcFB6jwT9uVQffqBhL
5Zt+jt0Z7obE2XiACkA47eNDtx923OEK18o9sTPOPLRTKa+D28An0HLfAzWAA088QVeJoYuRWe3o
qUFDBfK3BEtj4/72VdBdPbweY/oaq+ksxCyhlU2Ldzr3W6pvtTUB3KQ8SzuVBrN7trsFzRAglGwX
awEWucziPH5XBOBu4nVd8VBOBKWDvAQPna2QwmricbyGJ6I6R5jRttUzJpimm81D9nru6k8DDdiS
xaM69MWZhHBkkPJadZH3M9cuRgeW+vCTQC3589rWrZEXh9tm+O4ehec9Uaf8VUKxzIW8yz1RmeId
+j7mUBmKcvPVAjWQ2jyl1T/YBcWLGd7C+LR+Q56A54A1ALLGdF2eMUA8lFXCCm0O1HlQhVZz7LKM
iaUtd8z0LPaypz7N3rmBm0wVVALHp3e0Hmikk49TsrlWsn5i3yTepT3x3obOKaotXpwtl3mVDlz5
0fyy+1OTlrGjOeXKOr+FT/fgtFEgEwZR3WngVqnmtO0s2jJ3aREFoGHwRo2QQ4APhFuJDz/6CDsH
wa/q/Olg9GiwXae+quz6YJ6tKrIETQYOYNjPX+9zXkd02C3noAqkmUmR8wBtSXxXOpZygYEIURgm
dXmRmsCZIC0T+WX61a1tR3udd5LwsLtu+wKBH+rcr4JkntS559nnVusdJCgmWjpnFF0wzn+xhkNV
gv5LQafIltZ3zLUNZ5ncQtZip1rs2S5aoJ8XpdvJzgERwKylPlmjPv4GYkma4eiq2krHLpYEimnz
bR0RCd9S7Mlspp++30C0ri7xtVDZM/i7DuovLqJHdY22lhoZQbV8yu5p+V1Wuxsg9Ku9p2Cd9k59
OlUTP/Mms4BaXpWB4RLYliCcSNfIA0/olzPM1J+WCha9ZVZ0jp9n2yJXq1RL3UAqnqU6ruvw570K
NhRiO+ZM/fhmOq3/vtPNXBwv/mpmixueZSIBYIoONfR3Bfbzw3bjZaPexMLjoIs5Sj9LL61IZ3nd
/r6jRxTXk9UHqDlr5Cnnde8R+XQxAmLOC/jzFD0vB3GoQpunswKy7sfhvMFCNpmGkd5gKFG6oWhr
81Ft0dRTjqfNzZK/T0QRqcdjJuM10pMU1vS5BxHaQ+GwSD7Ih4Ua/8irtGo9paBRTgUacWvRh2+B
8ka17QEBCPirXp/O61MKH0rPxISbeZBOkluh0cDEqMMa9TrhfQO5iRRDXX2M8sEqz6pDQWbVbM92
Cf0Fh1E8mij26jS4ZrNc1fCcc5j2sodB4xxXB+7nXlgV8c4+ik8y4zSeGde09P20QTpddzClhP9/
PWRXRHdk4uq8LUabFIhccUtOnLrR7NVEcYzUjZsiQF3vjThOLqG6q5PWRliqTt8Fo1mkjnQzEhoP
TyyKBorfFAK/xTge59UB3SdQu8pCoeeMOOG5+UTIE5sEiRjFGzXIwEdAoZAdzlI/VqGUJJfC3Zo+
fPSdcmJneIxzizNKSUTboQ4Y9r7iV4MNVqK2BfoZxD91o4UG1NJrYRt06Pa5skEhONWFwnrZRZH8
gSnmMCzsHXUpcBH3afJLjyWmue6fOxIT9tul6G2qro5u4YCjcIdqgef/FT8heshDPEsYkse5231z
IWUv64Xapf5r2LN5J0r6bT1zlTDsFx2iQTVOmqUmaL1qTQCEZyXg3IOumRKfGfpwGDSZGPhdQkGf
ikPMTN2W0cukW4PvSFBnnn8HRl1B5cg1xnnZpfoW6G/JSlTWLRisYq250uPOCgoGL02/BF3hhMQ4
MLnf9fn25BNbU5ASvh4KHjKV8WX2Kykk7a1ArhZaLvdxjfLzrOfk8D3gJDAqBBqnydAqGvdaoktE
U0pvkU2XBmgkD6GsFUipqznlsgsrw8MXFAUmJ2L9Y+aihaFOXEfsnkN7z4zge5Ei1JAHDmuewqNd
9mTt98JZCXHIDt0djsfxOSqofb2Nk3OW2UrXW/jrQqN0WeBBJbSk5fi4yKXTDEV/B2XtptOPzws2
8yNU8w4xcvTvsNuwlx5wvL7N8oaq5DNtom7uHCW9/KLeXWDJj7LhzTKMQI/HIFCQ892loz3RJMtj
YOeQPD+MoqJmYER4j7N1Uni3dSvdDzWvRFd08ouH2j8KC14TRFg8aoJjfo/ORKYufjTN2l8O6atI
BKmyDikuXvvNt2gD6KXKiQsnT//IBqa1D7AYp5De2carNL/38slPVbqyWHQhZez1d+zfTrPQoXfC
MeUFiRe4RouRlqsvpttd/yWdR2p+Qs1fP3IX6G2YVB3PuOCoQ9Kjd44UR2dkjW168U3LVS67Sf6o
mW06J8QZSsYX+ywr3lGCR7Rzjd5rkHUvf1fMb+w6p1K7Oqg6DrG9kDt4JXFQF9QCNo/JAhghhob0
iepXbl263QhRYduCAWVQE0+2DBZvvmErsrAyiL26yiDooOx/rKiajVDWCcGmgeZnty6NWPjIl4Bf
E4jkaUnk52oiA2V8znx7H0x0y1M70Ghdq0CTH2MZ3F5TXtgP6s1MylTucRfPem5WDYN/d+yLUymt
ehktN3nN3a561qBXvE0bzWe+ud5xSHzeChf/5NBqYDkMOOJEizk9QMoS12Uv12VJGRBfmHUdVLpy
hvn5j0jVSAwpRlTq5rTiXoaypfO3hIhfz9OqC48IkPh/1L1VEJ+smiH9EHVtjL6OJOGkQW6f+khY
yaz0OuSfxtI25aB6auXoWNTQSpgKhPlQAk2Shr3jENE5ikIMYM81f/0dcm6vcd1rIhuEhQrAhMRA
QRzML5foEMFgQKYvZokqlu8OlTZhKZPMj/tYTye0ey1ZIIDjZq9QO+KOUnQ0M3pp+wTaldiWMcqP
XxvywyTbRvnH2g92BQwbySZL91/bto6Cp1wOGfoX1BESmTXLJBakqdd1a3CDwQGFGqN2IY3xX6wd
tyQF1MJvx9mAaKFmgk8HTe9L5yRsZNQ9g+q2uABVE62n6jBZX//KbJFdaWh5og685ARxzZYsTqY5
eFvcd9Hrehj9K2Qm+ETqOO5uZg3jXQ4a6IEcsdR86DKZx5Vil/VsXXxlvPU/S+T4dv5m7L76jeK6
ZIitMzVxVasG29RBXbvhbs2yksrb24jx3sxym/eBEcmDPFJlgg+VeCe6RjPsIM3Wk28GkmBW9Xg4
gsqKbwAYmHAsILyF43Up+gGDK2diMj2NAW9gDiMZUjVBa0vzO8zHKigEnMak4PQljppZkOhbEQHV
DhRzCYcpLYBhebI4f08DOL0jzoby4Hg0c3gfwr+AGj4t4USfE0CYBjzn+4Be2n74vRn+IRLmNqfu
AEjoBCAjGkLGNOJbiXOOuqBqM7gcemSIsVV3F/ZX5K7sTlZRFiBc+dCwO2yUE9KboBYJp/qH9TH1
r4BCqtCyfXr23gNJF7iK3m+xDHs1kE8ovrDtFXmlDhsiocDAiLx6YkXCUDweZmZny0JJXsqDSy13
HYUsMBf2PrHySZ6g3LzK5FHkUtEzK/Kg0yfWSWdOPIvOBpudKZolxg4YdYfr513SKeFMyZdorZFL
HB4FcV/+azp4/qNplXwTFpZ6T7815dDeOy3uzVMuOvvOp0+9C2r/wCBterPT69zuydnbqI3JCjVe
teAkNM4phxea40f94lgTWJttWC6K/xuOVbF20opeX/0VGvNHba7g/p/wgISFBMaX0+pRQG+oQ8H7
toD4jOH8kjfQMF8wiIpTfYyyxGu0lmqpm0iM7qxo6pcP3LK1USDu5TqH72ENyyhmlRMSnMk0dj91
VATnxiC/OPzDxdim3q6HZRcAEQsfSoAP4NLR3l3XLWJHe19d4kSWMSv5mVnLlZfYAx5kzLZcjatq
fqvN8/2E5jnwG22YehdAq4CbGwp9Zv+Wwzt6I0oSF3ckFTVpWa2oufls/NMUu4wSNHUrth5VcFOv
5oFGEyTv+Yas1mPaEqDueHj6C+Sln+HylvAG0TNc2jAFCn4sLyWILcc9KaKO+UJxoYPdMzJp6hcM
p+S/7LSiXZ5rZhidsB6KjANQfXKQYq+b3FpOaweXx9/DXuYcFePBbk2tpiJr2VGvd9VnnQlQBBlW
30+w4lNGid/vD8wWF/FSpF91mGO00SlOJA8jwzt4kNOpTsKUD5aVxusU2Lb4LewP56xcvCKlczG0
ZDHGeL9j7HQL31YDnPOJ6FDQ5P4Iny/KEEdat/wLjpU/Jx4G60+7xcNUZN8BQrgrauvHAnZO1TUQ
nLpXT0jY/5u/45Ze3wxxyCAUUviECfkMM/SGv1pPKs9IL0enDekUkhu/3l4YJ/o1O08QmwGvlI5F
WMVNcFz7dhxryBo84cAuB/DyPLwtGVO8T842+rSp0zOWJY5PUbOUc2HWf8pEfiDQ/LU/ZLNO1TV8
5XaNTS9uJKkdf4Z2NS0T07ypDLKKNvW5Mt9ka0fLXD8jm/aLFU1bnGLOfIXapLBC7wQWpfB/ulDY
oYOv0hiVGkR9ToQ+97qBoVhkwFQmYLeAKOhL84PvJfRAjAoe6yhF1mLakbBN5PWYGhBBlAqBZlsl
7VBl5HWZtuXFbwGtodVC/kGZyu5ufpum30yLb1vHpIxXcn0kvbNaekSjm54w3eaNKOKxLk/k8GKd
LGy5UXn5IaEMeH0Yki/AMtftSg3RAfVOqjEPw1TLOZJ4y88DHLJBM2ompU8CGkQs3fGj4o/g0gvY
f/vL1qKQMRk83fX/kMf/vaZQKb4XzI+dstrkbx33+VWLdZty7Rh72xvix1rDYHqAxfmc9gKRO5v0
sYS4txcwXw7xTxnVx1FvgJ9QfsOMiA/mVQBHJW5FYsSA6ZucqZd5jgq+cJ4ROIa0ZRQZP4s2/1BP
quidAe5X5ybhKmyWQa9I8mUt8PBXjtSMxljYPfFI08av/919XFD0v9I+Ivw99iR86xi7ZzbauDsT
3PYED9hXxFmUWLnUNdr5oLS9wDlcJXLiaa9TEVuOt+lj49TxEJoZiBaPHSSwIbppn+5eJhmPjHhP
qmLVK2GmUAesLSlYheP9x9PKGMPqkcJxw2SNK6rD/+t6ixFrADiVCC1yp0u0Bil+Ux8BaPaBmBl0
jzhDvd9F+jsEh4B/aDdZ8XTaQZgjcZ2fNTpEu7y4DgkzhVYGMct3dfgq3muRXQnRcUvIL114wcuy
d+DsNOlF3VCjNazXi8Kk8SeZN7bq+qRI4GodU5gWbyCp0E21M43/RrBpJFOyV7Uv6hmeOyiPiiuS
uqXb+eBfpQUr9ijhvGjyDHbw/GbGdF3zbCwBUt3oxxkOnaRaII6Rh5j2vHAdDFXR/u5/mbBG9jS5
OQwOJnxP8Z8rZFchbNL2w0+x4oSg/kfxQy5V0F0jS21oRRF/vm1A8n3sGVV5fTE+++UBKOBOBu0Z
arkGcAoSLqFJIsyK1UT3ujdAREIz0QuqPyQGRfB3hEBfTpfCyo4f7GiZfh6fPMj+qmTHLtPyIcSy
sHeTRtDHmhMeL32goFeSSP+pDGML2LSD0+CsQKesRy/D9AkyEcDlKnsF6kfCxSvJxZpvoVDR1uaC
uHGW0CI8PekFyc3rzW7ThxmlTKoJnB1EzFSTITvYHPbii4Fq75V0rJkJdH1WOYYtS8ZgCQffZK/m
wXV7Sdr+L/C8+Mgi7K8mqD58sqwY1l1sij75SuA59Wei0gxgpz2bcoTx5fvEcWDymMPWR8Wus+gd
iJNioO71DEiTsHqQ299piDnDctsjfuP/SvoEchxuxa0x1jaU1EmJKpsglocOHtOzFQqOP/Yytlxd
6/5+PwWcIoFF+99Uj6zKNJywgkrTWUxeelh7tNb2GzDI4y3QtXYYLnq0wwGF4dbqxtezlrbcCuUt
Z5USbseYs5xBIVCoLT7GWlYPxbZBb3IEQm0EzKxhAzJwlNh2Z0ovorbjWHO8lNSWnUfW1/Tv6AP7
GcAHccP82pNc4s9KmFYR6ScC1MyMwZepoPxhxwUhflcUjxRRiuyG5pkt0ywWvP+ydtNrKd3DhDxU
fBgzLqcXlk6dVlm9VhFh68EOaxd7ailoY8khBuINgF+sj+ObkSdSlOSto5VDOFwteS2922NDLKJp
B7UXAJ8UXKWFiY3H8ytbZIAmYW1GJ5ldIPkEWnBmA7bCXzT9I9yo3dtDnFuLnY/B8VvBhEBK9MfY
S06+13Z5ffKbfK0ZM+9acmXMku8mQJo9nXBjneYnEagPsWbqqgvLmZlMJyQGU281Qu/GY2JcS25v
KF42+zNkiPE/EjK3qI9QvvG/GtNA1X8UjfCC37ZoRKIzjo1IfVeyoKXlrfc+uqXn57g1v2padmNE
2XHx9GR77bwT5rSqyHV9l+vbxICN8auq7H2/sH0lzx/i3H/AS+GQO9yH1aKtpVhT12BHzBIc/ZEQ
ZG8rWKFGqzlkp1k1IYVQvV5aFt9VdNSRKbsqvaA1AwIQkf6jgWl5znZ2L8ZSbiapC9+1lHMXleaV
JxWSkg3S6ekgqV/TlqleMwvAnaOPwJ5dezA/oK3KuME/zHAzgOIUv/qdNs7zaZeMU9yJb1kVcYa4
haQ8Vu52VPZ0MJtrbrqe5vxkneW/CVy6Ux5TiHAs/FPuMvaY7ho3PpfpOx36ZAbNSsg57qDu5zxV
XriYXJnJJFtvPWO/x+g35SsCxbWg/V6q/db6o7VbyOehHEM/tG2d1pX64mGvhsuddKlJK1UPlApa
6HmRdtj696FHBY6RCvaV3unCd7H+FNFVsZ/zyRz6ek3T7lQBcVuivueKoauo/xKmanGw4YJrO+6I
uJAa5gj/3qxheAnyouZKr2ZzCFAEnetVvrHVIuXZMZ/Vqj21ojoGEqDTR66ofD9bIRjdyvDhPCDm
or67Coo5wXYcrZjnDY3+tMkiWOb+504RHCax/to/Ww9+etcN182Cx4Nrn8jeFh+UjT5q1WhZs9rf
bPXkRDAE6EcSSJ9+gDvq/unRSxComl6KxkXzU5Yg4qCh1mtvsN+wOvfNL2CS5bWnBYlnvsQ9Y5IR
Y6yPBhDbcDccZi4cJsrC21yyVGb7qZG1tyHCW11hZ30vV2lpgxb7NBS/n6yLCW0MRkavX9epw0Nm
6T5FaJ/+DRehsXNb9y1d7ID0jz/Kd4hd5+vT0vibSUz8S2sd7L1jm0b57vohg/qp/s6MsKYq2ytL
M/wsXcmKioXQ7EELU87cpDY/MEHnRvGExY+uhRpMZmUk9rUjSz3uE+6YcyZ6Yothsi+7nVt9T1GC
FAfBULZzl3P81VH2USif533K7nV8IM04QxMyrXQydlb/yMhxvv3yTWW3uZ+hUrWdVBbJkIkHhDTI
zdUQXIbAwEEAMP/dHyrhvXnP7JZPdm4XO8HanrD83FqOHw6IGItQ046VaKkRibRCo027i7KteZGS
0oDU8eqMMRQ/xPV07f5/Dp8ZF4SgIeKM02+lJNOpzg/p2KaIXlKrKyRAoU59P2vj02cPaFJWyl9Y
OmuEaRugcNCd2Dv+ENHmP+lV+dz8WKbKbAQVMUZNWMr4hCAlYlcXE+AIY1JOa+hAMcv1luMZU/jr
mSrj2IIb3XLE91qcx4zdaQMo7HjuzdJDuOTVFFmuaa1e9T6n0ovl0XR1XIWMXKKW6vB4+mQemQMg
L7BFUn96tzh61lzcG2/KwO6w5KtDOZoK/FIU3K9m5MfVFUxRTZj/PmnvrVQDJjJI6rLhwAaGzOB8
hJWX63dZZ2CjBuIYQgef7jf3KNOqVjDH5EYtPxARIsJijGorxjSkmSXGnrgxG/sy3Z8V03/D+V1O
vmOOu5eE1M1Dzl2x2vhJcaW2gZUdMIjFdsQojxDbGMqOopKhBUeuxMuVc6ZuOEK7ApHuJ90OoXhd
MgCEQcIzCb0QlGqsQvW5z3ROxk0kX1qtrP84juA6DDmZNIYo3yLZWWA6bbUh+crV7nER3WTXuI9k
B8uCfRfnNSALZK7nvS6H23WXpaTCwG57ymJvvVksHbNVOqL4vDvvaFKWXAFrxt6Up1q3k2p8Nh3t
n1b+uqhQ+rE05fldEIAYXOzdgHLnAwxMksh08cOiLNIlJbZJ8b+ROoHlw55+vun8NLMmc6b+bL7x
FGB5M3xvWif+3SZPuPbqht5FLmCJ+7m/OgcGFnIaB0La9Au3XFdPVP07CGyUK7bhM/b4PNBaEJzc
90zb4mQNraTNNrvwSZ5kutkfV92Bg6nolovrg6lrIBXPgYf/xzGGl892I9nydnxrSms27OLima6Q
cRZwj59j/CvcTYU5qNvMj28f5opBy/79k3zdIkSBAeoAnsIQtz6J363Oyv/Fa90LjqkIG/IO3WSG
sSD+wz5GIzjzOGYsqlvON2dRPrpSpuEjD9TwC/4bf85vqp6Z4nP1Vw5tNm0pZRDkhO9rWc9yRPhA
5dxueVqtSXUIwEObaJJvkQzX5BFUqsyn9CKkFCu8OUuQqCPJtu6Od4/laGInocgj9Nd5RDQbQ8zF
1OGYzsO/isyjmQJrghjlOrWe00kkPpQxCDDqQY1TpNfzuuOyjYDiCn7dZPxyEHGFYOu1UfVsZD1y
hHah38Fc0lEU53Ki7NQONVLVkXHlKl/WTh1c4PwBdmv+m0kWCqTOkIQdogNwE4vFsA+sRekMMla1
yPB5k+W52XWI2fQWTzVvZcY9HOIkR/10P0RKsnBql45GqdGTy+KiuF61mVNmjPUL9PqPoG67ux1m
0spzbmAyno8i53+v1jI1K3OXG7hmjxiwpMIlKFrGY/MxdO2peiAQJpf1fNRGxXEt6RrJcUQZ+8Dg
IPQrnaAI1E0vWJv/IphzdRiggZ6i6jcjgjEgoyuzcLC5F02ePo5u9wwLhjSNE1Ei6RB/65qhrWI6
hiWuRYzThKmgzdvDLFjO+POdzSO84UH+SEode4eWeHHUvpRwsA6gTWXCDUIxPUf2ceyrf4SXac5s
BoPlJDiyN6LQq0aDiJEGpaIEmuHRYSRTVXDFUwQ5dq2HmWnWKPQO0pkAf1xv9NM8wAe9oNQNmJCn
xWlKWRHRj6L6zqYxRghP8WNgkuIVznCPYz5Y9yynj9LWRbQLPm8f8CYuxIm31m/dbKQHTG91w65d
dMLvrgoy/Zs3Y7GkpdR5wOhg9ZHcUPcFOQ/KE3hYaQvP2QLQxkjlWhmts02gY3GgyEqXx5ru9NJ9
bwg0hLHd2j3Ry6gACLyCkTUz/ntExsHEMhb0fW2Ui5mOn3fmRUcWHFKZ9NC5+PrwchWr2V/8Myka
x8CgtilqaFfZnzBCIzAb6uKZZBtgsAHjW/+EknIFr6wOT7fbtvWFGcLSex7q8ooyW0KkFXZJZYcl
FCrjmikYOI6ojEJAyBWfDVrPXpqjGpwcRC1wE/afKVbqiZ3QAjpBq155Qt8iASjpngY0bkX/57fg
k5bL9efOEI3+INNjj7ze59UnX7dQ8KTWmiX/nkI099ELx+wo2Kn+9TUsck/moQmd056VtGg28y2o
Z/RcJoB7OsBKoAjvCMqPALxRzCGo752rspx+jyh3o3UdCLR8WLRfwHnZHHTIzzgswkk6iQIPqNXb
kdbTb9F81ecFh6YDlGFqGvPLet/Eg/kXICOWlziIZdRFrM8J9gL8LJUsEPRr9UrJOjEFk+yVGff/
7aWjbpEw+tQOE+HeSGPe7UMoSQm7ZpDyjrzGKqznFPp0lC7qNAmWIzHN9EdSTkQKLw/2upqSoHab
j0IDEwWX2WBIRVT44qgwv1ejJ+SIWykd8I0mJgO9pI0tcLblrgLEyd9ogaq+NXwkhYleB8c53swz
LLRkEaylIziO0CxRwqn9HwS1ZHh7LjxOBpIh80AWK/pNCZ3NUPlT8ZdVQ5vcLEvyxSHVx5iCmWxw
zJi/HL2+tbyPaxkrK08OcBgONKXnH8b9bTXunMQMGXw6gl+ZQjfqer0PkDVxY9S1yxoYLjqhD/YJ
YHqFdNJPRJzuCb7oyDp8+3BH8QpkRz5G2jsx9Ksjnv3yAm97ieWw2oOqMM+YWfohGtKVI8Ll196B
ioOc9Bc41EFzW0zTWRHwKpANFkmEjy8esKnSuWOj2XYF9C+uLMdk6M3Cq0m89FjriNyUaBbdVXTV
UAY3xXZCZvHKhVOsRjjIBYBqGRbjkTeO/7IC48HTrj8iP1Nb+E9lgI5CzBOAGbi/tVZiQxWBrYou
MygvBzGm3boDWbDFtplPi3yz1wO45ZjObE4yoXaNI7BUnH9bqfD2l3tHhOgXxWnqb5jITabB9uT0
4rBR+0bP1F56xEYbhIGZvDj6vlVfOc4CgQ5yt5EpJfuW6rteb41I2Fbb4B20rg1sZgoQUasRB2NX
O0D2Z6oPLCZy0bQpq0bTRcWjmVkAVkD2Va2DSgG+ae4f0yOG9bAfYvJWulEtsDpxWk06UjuTQ6N3
KG9Q5VQtvjNYAG3lb0iPsvxuw6vIf5a0+uA6Sp9EkNsCHTT64sUQQlgiCHIdq0L3M6Tqo62UyMcD
RD7LAiGIngcctVrJ+rP1ivgjcm56cQc7ld+MzNSHMkENRm+LllmW0pUvxPcJ7VIfiVGy80rJj2SF
mVQ7Uzcy/+Haov2vkXGejDfd9tZBBEdI09Q+GQmJGbOOY10WbLnaPe5Ubm8TaPSX1S73W5MdiABz
0rzpheIueLwYZtgWh0WJ31MxQ8rooVZILgA0OEhYfmfmx5Wqn3GOBj8muucADIkPKVJvodpreTp5
oqEB0pLNnOHMP8sRte7vMofufolr04aPE8dt6Oj4k1oa261Kei/0wsNycg4J6XJnHTemw6UCpQvR
mtFA3f6S6+UFxNCFrE3TYizXvHjgz+zPWkPQSjjmYj92Q0yiOv2e+SDOgczXsD03gZopfUSmeYk7
I16vmVN2duGajdpHhGRe171BBbadB5KbvkcgRzsYcZO8YUQT6bLIMNXYBOB619L8yOx3jzzwh/cn
GYmnn1D/KzePixmgg1VTodld9Y5NE+NBPgPskA1n+i5WgL8JxoxvYAdBI0+cmqECCV1NumVV/GU0
fjfUxdpsr/DZL7JLrpjbJ42GZvs9JglJbffZk0BEwMrK4rcrmixgejo1bkJyA2hhlNNnredxZb7v
e4LWIn2IN+FbdYRL3WoP78GybvxDi87InboD1HTBLXIwiBBNuQVUy8ZCQ9TG1e55kGD8rcCELizn
sN7GNjyoTRjAbusEDiTxgQOrgQVm9UnfOoltQHmU2vkeBh4Dc0G5w1JVGpyI/BlZA/cJcp8Oodt+
JM165FdsT2Ij1IRuUtYYE1ULTrzcGqvbmTQ2YB3q+NB/S1/fY9/nY1oN48Xeq/5fLosGg/BAXVAx
KVXbaSyrRG+0SSQ5b4utz7cpctM6yFmt0W0N8zzF13PO6oIDiyQraHdyO0t+nLsizz/Wn3jwo6sB
R/w5xq1fdym5JAHisIMcRpRdzKT/NPzMDQMgCJ7AorrNEQw9kR1gE/yEc3WZ+S6Pt8uLvxBir8YQ
sLjfw3QKD1TTw5SC89UIJ4HHNGFDX2prjoO7Cmq7h7WI31Hqi4iolgMw+CrsHAdT1acA2+lPwxgo
O0M98nHUQpBGhNQiMEFtDg+KecsI3QlSYjGdC/8X7XpSHeZapfudvho6gBlnsyxAIhS7CPsq7HdO
1ADcM5deVU8WW35PsHviTcgASFi3oBa6NiQ/ru5AWk2xaSl6OSpVPe+WQRUmoVglG+tot2i1UyRE
dPwZn3BpheeFgbejA87baxhDcp2NQl+3pAnRGeCDtMgHWEhnnnY/BbvzDDqACQZn3fYq9Jq3cS9x
WJBEXWWELDj0lJXd3PJsh7gNg91UdMXfK+dNrLpVxR++G2g0dreDTP6IdzVYBUGGX9SYyOWLGJX4
jyux/ym69VIYhOqo2S4vH04KhQhgevCmF3ooqLZ/ggSw0TR5yWPW+k2MMwZ69ocL07G/5ABu6MSe
ZjoxgiINrKtFw6OaxhMpehCS3LyzHN/wHl7M0HIIwh6XY12hE1TyHF+jRAovB57pG64mThdMd43n
RNXWCMwJktELBTdVi52PvFUJsQn2KuQ4SF6Y85LEsM6KQ2RKt3Z1HBD7/L/GcO1wfTqSQxBm1iy0
LaxE3yg67YZVE0yR2lK5m5BIK1CiAl4hJ1UMMwS37RZQ3GhuRGXcfGW1c3kwtN82Wa5kk4iIn+mn
1gCgeAIVAs7iMOR5QFoFVYQu7cgTQg/jHzx9ZOgZrN3Sc5b4Y2sjnxEPdVAT3y3DQEX1fvyNxdGz
w6GjNxqE3jQQCsC9TR5ydg/uNHNqTPL4Gt5MiNgwBgAGTxiIWCJ9JWsBfCgMCKqTifbxzEviEPH8
Vaa8d5NoO24qi10ctGDT3g4adYvX5c/cpYCEUKFFXGJ6WkbTBKBYzeIZPbkZkGUYsAvt+gKTPNrV
OmU9NqD5Fzh8UnstrNbpOa8Lxw2Ifklj7+ekoIaCoY4dHOvPc1QQWyj/ENQ9BUvQBkXnY3/m8F9/
aR2x/MvzhUBufxe1FTB0ltd+wONg6ybfXFSYrKgrs7ILsZJuFlC/aF1bzoY1kfwcqmqUog5uEB9N
XUHNcoSMBx9L7z6oTMt7vnj9CPM8crOe2EakyCHgXtVm9zuGAsH2zJrrJDs/HdKehNdQFe3PHYHD
EQw014k4QAgVs4R7Kw42fs1vnvbSS9w8U8hegAF6S3g3n3GQ8pG3CunijpTp11HU8QXm/u4IVsm/
1z5YJmnE7LyNYBacVIeaCNrE/0ard686uB83lhHl3RXp/7yTWP8QuyJ4AkpkhHDJ/2cJdNf+2cEW
ziM/2xpPfe9L3zjXVUGnX/tfbfTNsfjI1fCesqAbMr4/3snipLcKkZuR6/oy2S16ZuXZfTbCn4Oz
YNBOFrLtwmdiPzbzYnusyzpGDrMYCP+r/G5NGF3uL0cfVqwxjhsMH4HnHdGvCX0OxVi7ttofUZo/
05xdtDZMM1/VuvXQctAW0Ns6c3lnjQW1CGVEPwebhLb+ZO9/sx6pJIJUpqV02cCSltpQzl66yPrn
l17llV7NHvStEbVcYAoI6dx6xh/YAqbak1ZlXo8hogasVa5cpBXL0stKWkAMaa+G0DHaNU2nDrBv
B7ZDUNCcRKFPhyMQJJS7dOI7F/YrjrGokCxFq9weJSEphZppLnEa2qzFNcoHXfjoTiUvTLU3srLS
+IYfRpuFB2MxVue44OkrN0zWCvg12rP1v+8+syMHWD6kXId8hb7zgl+itRD14V4qmxCgetkIFhrH
LuduaQwruBeXhtSoRGqn1CZMw9UK05ou1RjyjZHHjVINuKNw44S7MjYh7qflUdmmpQ8xnRnp+ddv
GyYSilPdsr2BlVhZY0I8fSHnPEc7gOV3yZIorrnoP/iviwuPfeSrdYceGd6yvsax0Rd6/v8teWCN
VhxGM29a6rev1SUIDAMxqhrXqKDqKUbw5ukO5MJHJFIUf5iv8w+noFO1aCxIoKv0/wL73fHQB8KQ
a/o1TboyghBAqhF3MZ6hriyYiHVhhv3JoAU1Rt5rTUTvOPaIuLio9UTXEC/T2VP9O9U1GFq+sld7
RnNnZD0UUoCR5asITvCBsPUcBSHxWuaEfTCO4jMu8lJZBCuaFo2GYPGx9FYWbaDENnnO0Zrg71gJ
tVtFn07yrSgbbgW1YK7h0vD0htqpDovgFrL5iSWEKqIL0S3iNHm3GUd8/93jcma9kJBnw8vw4iQa
kbxBudrN9xoc+Fg6Bl0pV9rshI9IHzHyQQROEJYiEeCnTbjZkI+bui589fdkflX40CXdk2X92PzJ
FF6xEM8OIcq4VXxNEOz9llnw7RECN3QDHWeP/JdLVICtFujNayR1udQ94W5g9hGQgyNvUQ2kXyO7
GMDMenY0RvMHhBspH8K3kgjkgFr851IGMA4o+K3pjyUk9rskXFyFFBax56UY+Qh2AHlwawadaG5W
xHBSucuhrVDPWLm/oUEbYNdt1CIUSzhIwMdu2rSDTENmsyjNQsWARGJBPPL0h6LOFZihOrZHu5ux
6W0ZjC0vxIfIF6xPbmmPhLqw01tZNAjJ2lx9pzn4YQrVDAOugsKEf1seoisQ8Syh18d6hl2F5zCZ
MJ3JCOwuD7SXNpo1dqwb/wC8H6az7Bssdcq9hXvILDaBJgzNUuXfapIimGmOiNI/w8ukVUpKuPLu
KrgvmAiMGn5xVz9qezn9hnUJoWHlA2Jh9N+djl/lO1UYfXXHalFn9iDvZpyhPAGQmo6VZhVcZu9e
m5VVWDgkyqjZBO35nkR8MQBvgx5o5xXkASwvvi2/2Rhd3hYgw3qGhmfCMXQfgRr3pKuPTWhnN4W9
zXpA1HZD875QJyyyORD5uPFtgEsd1GLXoNOrk6r0ZBCj+vRcAXXBLhBLWq/+N2g5pgDiRZu1DWaM
04Ln4X/ydMOHGL0ufGtYOSUiZ86mg/CcnBXW3DDhBtTqkBUBrklA/hwJbLRXHNNMDXPxRC8+m5Zp
2FxVdQbKztBtcDc2vKdaV3pAK9iN2yKyg3BJzSe2duma+mwsGejDRifp5PJWqv9Tu2P4o+VDvRHv
h8o0k64Zh4KOslCFlvvcTGq1+jxijjg/A/67DIkPdUEasFxXcjvMJ6sfYTSMhhfXhtrEkIv0SHhl
nOVFreM6q9b22x730gBIoDSVqWbhqIo8LKFEhHzvNaATdy92rk5AgWHWtIseGqtvRORPAOKU6XCi
SCPrN78guJCFjHXa8ddLiz9ElHPcxfrC9ejL2KTPRcdaIMN99usF8OYOkXa3ht188ZVHELfyMyle
nnkk0KkT5xFmXEL64XgSgYjcu9/Lj5J3PtixYH2v0rfFHX1FfYgqdr3WYYU8cXxkON6uUizeMOD0
7LQf23DSYO3i/sR3M3ttQADeME8OO4CcEQr1kscvSBOW5lIpMxOrdEeJqwDa4xmvn0NXUn8+z78p
H06Z+bJCozvpTVLIYJD4MRKoSS/PxoNrwgyT0oTDuOBuQWMIyKChxOyzEohciiGvIt2HrR62V25E
bceM4cZBZSE4trB9XvlH9lK34TIq3PoHq6A2CpglSs+xQvcNsXfnhjTOffU12tSri4B6THzivFAh
GtoKMgaD/x+BSzdYvGV4tdro+JXAjK9oWHk0hQI82D2JjEiaLa4chpIw4s96XWQtUEc9BotZKUIm
YyNMOAMN8Us41CS4y2sKfte0p1p3fJyJchvyYQ48IxS82Dzu1+G0kdajktFLbYrH+knypj09xZk8
u83X6Eb0BhHViLCAqfUIoILdGKGrThEANSJEaTZM/nL3CIaGFM+FVXxM4PIzuUL31cMXB/MFiTXB
MSk0YODWcpwTT8pK+yA7c3XKPUDq9ByfzvXDwd+G17NUsZLjEwBqaaFIGqmFcwHA+qtj25su/cXi
zXPs/jdHsCX8t8igWh3Ah5kGvrizmM3P8OSDQp5gqGh3F9X/joEVXPpuJh7uO1xBRApDHdUvh9m3
mf5byCXqAQ7+YXGOmGtna1MPkI0pTHJfzuybNWMtj6TjU3hWsIBgqhsJrnJ7kylbbYCtVU3KIcMt
/dbxMOv6ildoXQOMMIqA1cK9bYizDIjdHAGe47xQR4gJ9+8366d0hsE0SfsJmW1le0+h1h/AQw5r
TLPTlzWUJNnvmELAsWpd3qeftgXSSO2tSslr8pKv9/sygSk/o8vnPrPJfopWNMPWqSt3NO13eSF8
2O4Tuf24w5VcY/aR7V9WzJhXu8j9tK1bAcdCkutXomsMgFrjaca9qLuPzuP3zhHfThdSNCqkr/rh
HdXCbx+0R6UYiB0lmTeRJgLMwMBh6JSYjdzivlf3DA+hKtj3U0N0BGe19s5vj7MDIWqnDMbzx+8i
0BS2/kSC0PpIqmEahv3B44M9ey3UEsCo78TWvpw9Nabzbyx1TWrRpWHc/cTgvb4tdh3Qb5e9d8hE
E1WORe4ct3nh3cGaOSSKmtfTFfzPHCKwOu8eGEZdouCbRXN/PdZ0t+01IZT2zPQIdI2aON09FaLD
y0MW+fgUkl9lYLUs7ju+uZXVaMhXsbP9eyaF5Bq/k2ZHLShGZ6z0R5cZ4Qyx3QmEIAv5nPE2x/Aj
JaWr17/lirBFvPZBRt2gPRKCHl9Mco8BRCMcbPySyEZP3gtvOYbeKp8X0gDCV8nBfTTsP2iI0a/y
zV2mfaf+yU92PRVAhH/8M8sCQfzH6SBO/rHfQBBhdeSGmqrt1GXVDAremmTAqYbCjdRb0d47HiYO
pW07L7MuUD5evElab5kW/vP8bsa1TCZyUy1CMX04HMYYvvKSdRD8UDHdwdE1tDzjgI3czv0FQySW
14yrGDIlEYqx508v3mqdAOJFweFNFAGVL2XXjvBEUg626OC09MSGersMmFjbCHxBJTWGnrgroyYy
t/rqeH11VJCK788qJb+Bb/i8s5UGu2SPVFB241143d8gb59ifFSj3zxqBepa2mrshEPpXdjLZJXE
WWVxmEVUv90iRqwOQCCc+8zEZgLFHzGHZSb6kDe4qbujR97kGt2cSFqurH3yeZQ9qup24+cS8JBP
VbsmCGGYh57W/iubrWkto0Vnwzh48yG1ZOa15Guujiq+B7F6oWIRsJHdxTGC1ycbLPwr/L4KgCLz
zNu/NmlQ3avsPjYjJjnHNSmpgfsW+BHHT+NWRCFzQQioAcnFAM/lUQuy22L3/0kNyV1xuQb2Go7o
2fixfdcEyAZCD6mPcZBXoUjOMMX9myHx1ds3xknEfDC6YS4m42VDF79vJGbY/EBMxRPVrk8SSXi2
s0+KmKo29PQrxW6HhLTpSfVpdJC4VSH3vTiv4T0OX4Re8UmOFrx7dYJ74HsraW4vW0ey35+2nF45
TMTsJhiEEIyfHVu5ZBde5so/QP3PcLsMNPk4Qg0ynKDBRRLpwmLuFHGECtZzYXXTznCmft9NoNWi
wdwzjqjf+aSpyx2NRSvFIZ94JhsIiJTA1UVJCVBRL7IsPYCmuYBVxGFOzzhKQkjZDClmpzX8/kcR
ocEHB/1+BXxAgiBeZ4bCPj5ANfjWVc+LSHCf6W1XrkbAnKTJKrwO9E0V3BzGpMYc0sAOfZe31oJ+
UQ36g5bggar5QbERurTVJMtwSe50vMVSH+3h8yfN7M3knAB5dUzfpks6qKIEjlR09hLysnGlH+PB
WjH8P9iePRznjPiHQvYEob2039rf7j+uUlmeL94iH3NdIUyOg831VnTQQBKo8z4rDDRnAsRbggsv
byIORy4Y/+4WE34m6drLXJhj+Lv3IjVUXNY4ErZcEitxEGfK5FxRGP2hArFMkNZ0WXA/fCynbfRx
JtHmDiaQZYfT7fyZTyTdLXgd3X6OowGOLAkgiFuGwe+TYVa/FMryEnbzsfjfLWgEl9us23s04Djc
kEBNGpVQs7gKyt8kAxRJ3V/f1AApBkRHlJ6Jo8Y18gYYC2ir3aaf1Q9ELzhw1Cf3gBISwmfS27Bx
RqbprP2BGpMOmbK6IPG9S6/OH9jyL//Cyba4zVGhHYDj4CbF2Hl/v6SS6JPZm3KR6kq+DBW2oitD
tH2oesIvx/0/pZ4i5n7ubY5jBFt9ynIoDT6DG+fNX5p5PoNVkagqiBp4FoRqCWblpuvu7WW0PHp7
zKESUJIpxKvdGt+kDIJmy8EFBu6Ph8h6Ea8xRSSVOqgi5ZYzh/lM+hiQ6VHJLL82PYczizxhbiBy
JgAUczXe+uHszhIGyVCxuKVQK48GzlD3nsGXbt4kbtEyLlOLsNSkJa7CtIFa82tFgIg6YV6KQFFo
fcmgKxG6Za5FbtxRu/+RK/4tYh0kaggd4w2HuMItrk4pYhVFfzjEzS7bbmKJaCeX9SE6ntfwJqMW
22OUzteFEScNU8qmcAUva3iAAxtVcoPfL6HE27UlK4NBcrFlZVA72iXWKVq5WmE057kF8Rk5oLZz
B8oFmaAp69J/KBrUk6kjJ6NumcCAeAJHU91TCWA84v8i3gBPbBHRf7uWrIe1GUM8M2OKZSx+gIy8
CuonN2kQPw7P7uh1tpGbAggvjcjcdgu15dZfPn2Uj4UeTDYDAIYSwUZpDJViNKWWZSLY0rHKzqd+
/FLjywzH6kqXTVVY6Cu33Nt1Ls/mcsqx+UfxNsS7wLg2wTaFjRj3m9k6viwS6g+3ET6fyi0SL5MI
pE50u9xmSV5s0GfPY6J5lgAUVM2SqxU0ivD9UrUmLTg3UOsXO+Gq8JqmNOFCY4gwSjoP4XYMiHiv
OjQbRrOfiX2paaBnZn3NbgYVEPv0abOiO/WfUs6z8g1GULdBcBt05QdT1twEznbGQYw3flNJCC3E
rlwK5TEasiWv6P6WAnMgcWMBLz2pOrY4UVlDqLKXLUGI7ywMd2qDtlSCUcXRKdVgTagzd+mG+TNL
gCOQgP0GnMLv7lfYLU88K045MLJaXp1QbesFLJGjPXoii1Vo/3BaFgMczvAFF7OkMrDAUUiyOMBi
NyW8+RSfJ6J8IvN+p45M2CDx0cvjShLzBUoXeTsrecoOMBV7raq4grpVfmmlFe/Vs8VepfZS+sl5
HidF7XNCml8H4SfHELoLJCggzEiHMB+yy82+Et/i2CinBlXxDEQ65PK7NrA13PEnyv1ZCwr9ItHH
NLuUifhwy2UCLUXkyAMNhZBKi89gew46DXuDRWkdmKHKnjKas7/cPSJBhB1E3Z6zeM3i40FqOL6A
M0VkccjB3wxBLqgI+0c/X9WaHgU4PLuS18j0ZGwWLoaMLsIs7LKGM2Q01opgfCwhZD59fYmivaot
ltQW7ByrVTyekJS64F/LNNyWIYGbJPNIW6V6MS5Es+5+FjEYVfQiJgEtNlsw/E3IWVyijvLMfsLw
+VuFepPcohE9IG9xgF6ikoOBUiCkSOIYb8X0dVCbTbh4mNnskLdN7W3Ek72Yx/AeX3gcYXwK0pJ1
T+iO0SSO5juimrQH9r9QyViVbXBuq99SGUO2ccPKQXgjnoti842l2sbVPWY85654aJun3OkgBQWG
4uSfPKJpeqXjntSv9dyOoKblbTb38JbGcc604jScG4Os5vdYA564/Fm04TlK4I4Qd9U9BDiuQPbz
85RnHQ4YlW/8rgBM++ceJLm3VXapzP7FMY+vWeoU1ltOjSCw43Ij5bEW8Sged0sYFKGsrMZ3i3lN
8ouAYmIsxuPHLiUsd3Ga7ihju+AYEICyn44oqfXgTGepMJm1HkT5hLWULD2psL4/ndfQ/hG3mdkI
tG3Mjwet7nl74m18DtsCvFj+aejw2HylVWLnJtANo9ocBGzfifHl8F8XG5+iXS+Y/c48O78wWvoY
fH/uKZyVibJhWh5KxP4IHLlvnL80Yq+hFrI2Cj9bdo1YkhiaV0znjb1fKKXMjOcX0pdZF3xGP+eU
5PhIA1q+bpfJzluwIFPPbsOZD3xPEQzTYw3P1rEN38jE6Wx/gCMpa0jo9YDBU6LdjCkJhDiONAEd
92eZf+mdqK5VytD17EmDvGNOD0FzhwgwJm73rpVA1Nrz2PBXeKW2PrXW9KD+RgwQgg+tCfWy5Vo6
wjnNZQyovftOP2+N+qrresE6TQ0l/I/VH3JqXS5wo+l3rCOFrEr0Hl9QxgF53fSYK48SNr/JrmWe
WnMeU73JalwDzpmTeU7jecrTIvErFJZT92w3La0UEHxYg97p0fsH7EI9hxoMCAjqitRCI0Iy4yke
o1ZRpkbdyWWQGz1lCvCevAfCt89pFEoraHKs9L7O34EnAdxr0Z8LUTiF18vjLut9gBF7qk6wWAmZ
SnTO5fsashsNRIagVroEqv+RoENGop49D1zrhPBKp0M3i2/L9nHVNAwBdudINw9jIREz9BrhWVeN
F+YjiJELuZWE5ELr8EenMxDRXg4NhUVC7A6EE0eQ3o3G6bGf8dCXMDcBqnYz0PIWIlZy8nz28d06
ttXeS9OlAAWtekl15lcAufOimZ6F/2OsSL4WP2Awacsxee+6Ahxys8kx6rL3Yklcyk/Dv9auwm2t
/MNAeq+8eXpObBl51XXTbC0rZR6o/6konpcmR6+qxSA7PfD4ivr/6oXwcd5jF+0GHwc13MFzul6C
4rdrHKEdlJzlnxQBivOzAepxhn7c5g125OFogxwbWdyui8bxuA8FaGgID/OvtiNSnyOgonCLtCbu
/JGojlKF+w6oMDlUrd3WcenBUPttMHn+c7TQ42RvnaE7CkaZFzIcs31sgx4LTq3CNHk/18mm04R2
YRkxJ1NdtSLtqqjHc75oRBgmkdIo9bvH/LSC1TljZktbLvaVqBzKsTyGXluFp0+GWk8Oq3C/WEUK
rJLniLtwsygJR75Nt7QZoPx6va/QjwSUVw2zqEsJPv5u50dl7+3kiWhfSZrRd91mYUeP3HscdQUK
ALK3fQUlGJF2MSUWbUvyjtxCnZXl0M74+rY2L3jjl3D+WvP5CgeSmksK0+w3y06ULBpVGFk7X4o0
aWIJZzqjW5PIsfCfdYww6u8aKGmAiVtTo4DB7Jo/ioyzG+D8N1avDK9j6Y8tGRiWPayAvPedxFu/
tpmOOcB2o8nlaB+73C7DRSzds2bVPVjhV0c9sb+PmfA0dfMhNJ9O9Gpg64ZY0f1rEOtMX0DdRziX
I6NDtFkvloNOkRWircZH6s/Pq0L07j6BV6L4C57dz1zz1g5zhSxcUKkBVEbTxIYOGLwbaJ0opmXB
TpfdJ+wa1S+x3M2aXBJOxnIAIBiv2hc2CccT7onN8M1VnMRjWkmmx62Iqe3dhNapj2/HBPrFQmbC
/iD+h2abZnYiMIElWwe3lATzUr+s+1VcBCp9op3AArc4OGOAyxgpM2KEujSoh4MS1RHs9tlF89Bs
FznvsQvSyv4OZb90F9IItxv+7QsqYi8snoHKY9uEujhZTKIKxw6OFD5BY2D7K5pZxYyddbvuiHe9
SaIH+zs1lb8Sor1MmPZCoAWVO50t3P2wbbFqEI/vaIOfys2sNSoILN3p/VuFJ180wmFJZZz63rKE
p909DVhp/gkje8KbNEUIZzzmmdWH9YwJMQFkAWg4JDrr/HyLJXrFfQI3Lb3X6lx67hpyddkbpiYc
bCAnJ4X6zd0uV1wVWwb03ll0eqcSI++cXU2XVMHc8DFm7azf2//sEN3Hj1TD7tdNQ9rR1H+AJqs+
L9poCrvH4X5o5zygPynwpko+JwAfPSAJCg4hxTnJXsGZZVbXoqzMfhcwNFgW69+RcBJz1AfM6iSH
DsCrSc3z1FK2E9tN19MD0naEDHCoOzqa86Y+AxsAiCEzfUvDsGE+TpvPAdguvtDfxrgcDMj7pBE0
fGWDvtGS4lxBo56PQPUHJ/7rQRY4crb/OtOubH1gSbPcVlT4SaMpyp7PLyB9ubws8xrGNrCij41d
mJvexwlmkVQ5ZUD4iajTXEtWrE7+12WUwakMEKutuKPvLRhKh0iKE7EQH6oF2/vr8APxm6N1si0B
9fJP6lPkTJDLutEskT32O8O9Hxzl2HjHWjqD5JIkpR/7nXbgK1GYoxpoEnoA20/2G6ru8aqEXYBN
UWauhi9wbKXK/wDHsXSkqWUczL51vORaFiWwG1LvPAs7EByO56PMeZBiZ7e9z9qo3veDNlDG3NXU
9SvkVKQX0Jvr1wREDVuuSihl6c/8+MelL1KGCYoasdYhfZqzRx9dTHwpRyoZygaGZqC3+7H73Iep
mdsQYeg+M6V/EehGJUL8c/JK3qCawb9y9XTRQYfVPGzkv5FjmbQcrGbMe4imM/Iyh5vHEoU025pZ
3gp9NGgCExHJ6n1ZkDHBJL0BMBAiQqKTary+Tv9wVwKLcWNnH7TyudMOqMlDDkDq8I/IkmxlU2vc
iiPbzzOtHg36tMdwlPjNOsPIWX5t2BtsKKAVNTRgY53k+0RUagAT7vkfAU8KIq3zxK8EF6zJ4IF8
p4hZ3Il152qwCtM1OKlNZN4u/dfIEDtItUANsF3SQwGqSQL4S4JbEkdSsWFEmjzCycHbDJCSWmFf
dqQ+LkN9iC62DjGZmOUac2YAvxrnxw9eMpYQBBbD/0wbyrgFjuEkaUp/Tr96WljMbFEkWprp5Mf2
H2UJlTcBHlN987osI3yy1YtRZdeXmfxoDEja0EohVU7DWyA9kM2FQ0vXRFsR9B/F8H967hUH5MbG
7v921eFrV99IXK05Cyw0fniKCBcgXJNliJuGfaWD4Q7WAs9ISRI0hHZfziq8TDcqAH2FnxGDfZuC
TTbwWhEF1w2b5KjVN6kV6FcjLmNWKVPJ/TqW4DwL46farc56cRaBk5cPq/v3ZaE+wu99WeBgNpwx
9DPJ/iE9EQ6vog8C2jEJwV5w+93Br8JaFcMuYNnCnBCr+tQuAcZv+L4qG/8UQyWveAPEXVVb/OB5
TAyBjJdPjQ3TMCT3cdRI9dRraWRzZdkpbLek8zIwsCGXgi4bVybDDb/NOOklshk+hvalkLVAqk64
546gAlnY/DWFd0X57v7SmoCcZBTGfytfK+hTjNvjhRNwtq+v7t6VEMFJfIU056KEoPa3yL4oPy6u
ucQtLWqQZQEL24l2U2fjDeojdERNZVF2IirRSWm06sn2cE2Rivf6rIY3XEwK3p7XNgUEL2Ywqx0O
qkjfm4n0LKaKP1PJ8XbF0QirHVgIGxe8keO0Rs8IhgmbT2uOVz521d6VFvOKVyJ6Rf9m5cQoABRd
1ztebJXVlQzxMEmt+r3PM/djcU5FsFiyA10fXwCj8NZYYNTT4flcuNVoCPdxbl2ZL+n556EFjlcn
mpV0TTnyN4/hZdt8fN0ntuYuqjLFkn1gghc13phGPb6fUuKNM+AV6q7QScEvZlcly/329JuRRTOo
/t3xIzciG5UulGa46erFmjwg17ZocW0ptBUitOnS4JyLyPduvOK5kxozE3Gnbpzd+VOMlbvozC5v
JKHTtLb1C7l5TBos3xb99rQBD6WtYbiXb+guDgpYcPnC/EBa0S4q7sk/tJCzF75qWLsmJeRf151R
hA5MTLjjixlWQhODwUGBrq9CDIXtdIyElYCHMesiSHDd5KCweM7fLGbTOUvrwQrhCydv86iz8Wis
1FbmtfXxVP0g7ucf4Q0VLfkhTYc6Vc5jGJkW46K0MpeY6MYRKq7P7t7qZP61qfXNUrZeI6tsjqaD
RjuKHoUhRLWAoyG9NS4xPEFirUv8kr6LNe32rOpNgwTJcX4KeDjQ+KMRCYts3OqkTPitfqQ9nrnD
CkNp09A3PdiuftEjTpVHU/9xVGK996vEBcvKCCkWcS7vn2ryWDl5S9UxS5LlyKwcqxIP+8n1SfSK
Re3Ac/dbsvvqxuBBWOoZls+nfsaGvDTi+7Lt8CfBGjmbiCyKtVJmpbXAw4zg44rzcmMzbGTzRy32
IuNeZABCdWR8kTyDqFMBlHI+twHcra130Od0oRe7zVMSWMB2pL2NV7t6vYUqy0CijW0KVRDm80K3
SHSqWqjZorfj0Gwax22FC/ydk0Sh9WDUGDhJIhDCZS9v/a0Tp7lxMKJhkYdvrap7DJt2cW9phNOx
c5QYfuUIvwbWfKIgi7ehG5fiWuusT9FNLQWgqw7MOGmKbG0ci0pXQw/KgC/t3aHmNmNGUNqHJcjq
YY39TpHzHrNNxlp8/bpKmjx0/Cbf8n5yZfBNY4OTXBr7sJrQoed/5vNfVKo6HDFzu9RV+fwBsyW3
iqLIshd9TVOF7M8U3djGhHBOf6EArqZNl4Xzxv6uu7v3Vb7AZr79UQE1SPT770lR2qe7iHSO2h25
HF9BD3VJpxGKByHidv00I6ojqNKWrmsS3zkbUTxpGEPKIuM5N9FN9KDlH4/Kf0E3mi3m0shnmn9Z
0sshhRBAAX24nI9ayTAbOv09rDBjNQfpZjZxYPnarbAV+qbCmnHms0jw+Cy3wTvjka3z3HXXFirz
Ah0bADTeUK4WmFPFAmNzlS50eSYKliQumnF8mznMjoVZNNEdlp2ky8pVdVkr6zGv1BLjM1S4uJqY
gJ241dxtSeFB12SoyUjCkStrau8M5WRgL+erVYk9YFfK83HgLXls5Zkfsu73lmKp8hTkFeNajHVG
P/Nn5r1D/DeEdFtuCB5TM9W3h2EaftcSjFlUHn2XUbuHYfNex8oGODI8dFtc242MGsyNyU8CD5ih
RTYdFYZq7ArIl5P/mdLj4UBgf8aWr6zOiyq+XZVms7gi1fEi00XW5gZLEc3+f0wKQARWINcuEJOY
75kFqbcAkFJo3eDs/i3al4SYAR/cZwMpzAI4TcwqOVkS1HxF+54WpyIFwbbBDjqEclyQyAhBMejG
5epQnLmcvgEZjfp9pq4R1p3CZoER0TXe2Z6XjIGyNgEygGyEPZxLDF0qoG7op+E8kt0Dcq5qprgT
q43JAxexCyNhg2qITJ3B3j+joj1FxtKoNktucLxhgkQdH6eiK4pwoh/tr8xxGvmNGP/nDAhhsbNG
mn8Z1Jv4iX3gblf1xwY93xCgHxp7UVqUgnt9E5aHCfvctXa/lYPutlmsNcPQKi7mj4bXe6I3ICs3
OEKVFt6o7wwhjUymlvnTNdI3O2nhy9wl7+lDNWE3dGq3e6dvOedQci5pWqGc+yRWoY9ne+vaorV/
KgbXrCp6aBlcqJunOdF017VP6wmF1IxZMoL/rD2aWopxMpioarNIFRiyyfcbWYnRSgPGm7PepqEg
jaUUVRSVHAmKN2yTUsrGAYYoQnwUiPeis8DsEOHeCiA/nR1FU6glOXvYoRicC4nUBdCayLgCoBHm
RcgMQpm/o9Dx2FsBv07yfdsPv93iyGPMINtzCRrJbobRJwAqVLUHa1Y5+gvvqWFC9hTzIsVpsLQg
/LtMs10JS1ro3cVYwW6xNVAvi1CoNejVHBxKfogWlwIk+9yPHpXCgZx2KBEJ1JxrNHRRCoe0sdjl
GH0uvaZ6b7rQ1ipD4coyI85zxUHmcAtmK7tRu5LB65yozqJAWZ1lJbHiO3/6k0Lhx0A7t2XCUNPH
YdS/s++M3u8wyUzG7L/JcQxe1SA7CwqTQU7InssMkCEZLlgey8kqFM1zekdqMqe2Fv76sSpXN3Er
QylyO0WqHWES2ZFEeOvxaPAqJlXcffqagOnK20kFBtsxhhaAG7CHVlDU3VE+/o46lG7YdIgjd+dE
eVuSSK1i+28GvWr5z1BeSrnAZKdJru7nfTDlCLzjyKbGNJlNRjB4JJ5yquxfS8ad587S+JZTP+Rq
bKM8DW8zs8OkQx2wUJIWfM0eMxCbltAkMW3u+jO/83nEjjgO26I/fwDDXVkM6ex8ABbtlMzRvAA4
IB13Vcs6ETyGa/RzpwpZiLTTOFR2Rcw7rwiC11J7r3Ay4uANFM2r0ZlpZIHPamSEQ2knesOt4GO5
1pwRDjJ76cePUqDq4weNwyiYNAgGUSRd6/R9COynHTn/9sOSrmViFq7ScsfR13MN9i1z8d0X1kfd
k/fVJ3X9QNCQ81EzPUEJqqkh/Lsa96CWvvkOQexxpw+SSaVVLR37hRbEtl/8zj9DjyKyfQ6e+47I
wf5Z5XO4UAsKBH6nNhnsPra/kKMfG9OPLtIFvK+Y7z4CiE6CEdMs9NosRPUIcZswQfkmnqEkmQGk
pmO6pdv42LeyaGln/t0xCsoWPsTo1q6PSrpGfnJ0irhN389oYCzdCzx7R8n/BkQ7LVW3xmwFP2uM
vVjU41b+C2K/q0A4aanK5a4d6ecsu6Nyx+Pl/8LTPwtuf1jZwEhwkPrEolcbCNAcDIOFT2VYs61x
VLMdEhSCZNoctV6t2hdktzApehe1xw/kHaPs8Q9auC973O5wLGdsk0/TgSo1ZGcbbGvodMVnhHzQ
N5yL6fqQ5ck6EVc+CS/RKKQmCkuuZ20X5wLpkYOVxVpG0++Bkl14+rjhUVzci074tNCNcQE42Kjy
4ZDLXy+8eapcu/Vtcb8fYDeWgqRo7dJwrip31IjtsD32x5157OWQ2Q32jdG17mDl0IPgbKT0xVeL
gCG4p3s9v3WV7a+ViXgzsk8S9IZJdD6WFyJ66hzaqYWQZZliqYDs6RXKLhokZdmGeKLOMZLw1ZiC
+KKzooW7iADK5Yg30r0muxTikYKJIbbPINj/EMxmGxcbOKp22Mse54BpN+0/fDpr2nR2/c+BjY0b
LUYg/MqZAdBjrWSm2GnSaXbViXSuDkHAkGffKywQshu/SFtSARTLHlLWAzM9yhzFpBZSRMVKTMKz
i1eiU+QfglhLBhKmtiMdUd8E7w/2xCz/h4ZD+fzftrvb/l9vB2Pi6c6iICXUOkJjqRIiLdz6K/NG
BMZohPa1bkjLwQE3AImxOy+58/wuqtmFTd90dY06smgDEf1zZwMu5AzRAsa1i3zfAzRfM/VH8RcK
4V6C03wKfdhbXBKqVv9VEn2Ocd7E5lmddX33fdoFndSdhKCiZChDWOeWIbQoIA10ylKCodeNKxkm
cFP2BVoqzmlnC/RmmsME9Cnv8pBwPeopDHu+3U9AGN05CkhpCu74Sw2UhbwY89Mg6zpCDYbpp87B
SLpGsA2HMhVJ49HldAHlotggorRQkoVpo60pIg7UYahs1uCSoRQidbhhwVSjmzI/29y2xlRcbN6I
BlLu7Zf7ak7SUngHxe0jIYZ8ymXcWdykvDgfdMS/pYim+dfila5vd/hlw0QiIOtUMvhnF4Dd66q4
XH2v50c5TAwVMj/8oHWDnvfMzmiczxl2oHBS2rlzg4dSe5rkX6IVkWPH4X9KMUHdw21QxvtjXFt3
OGPtRBUr5bVUa9HfAvLOnZRJ47qqU9rtMvPoCjfF/wMndYPsXL6TeFz+ITQua0vHReJrPrBEvzNL
0BkQcMIYZIX1qnySvWFVG6JR5XcN3P0q3q+eNVGUSTz7kyiX3hG61O7RC8/C4yJxxAtNCcwFi9Kb
DT2GG+bbrU0tYKK95o4/mFeY8Hz2wxNa1g+UwbbJSQFwiv3v9bx8ZgUJf/PlgWkQDnSZ0Eq3NYYV
6+zzZwZG7jZfrzgjbmXoAldacJas19S39R+gyEvF+AU00LErqPVdOonpcr5ubRDlKbfYqt8zQtbl
9vnIcdMugy/hSS65+HYbBG5OEU0Lk4kzQ1tbpffwPcJvVncxRjAcNZ+KBO/ofHaU9b04oVdoPGY7
L45NtqwcJbHRgOZQgKphmNe1Mt8J29azbKdvuWxP6DMKDb+kEHxYVcLzXWJSZYIOj7f0EwnZNYbi
lsOeiYs/f8Bxig6bPcOIs/5hINsL9euYbgUOub5MsFvkT7pQH7cpv5Afj4E1Rf9zRSGwYtm71CrW
uBvYZ8zBtrs1OVzvuiGmIymWm99KJyeduJzHrV46sCzdsyDgRJ0J7DjkTINUUPaX4PBsmJhMxs1v
yVP2drWsZAXRygJZVzRhhYeg3HvgDC7uIhqAhtVbN2zP6GS/M78zoGF2A3qHBfCa3jbOPklb/az4
Vkj444Fx5eLboMmZj+gEyYtlM3PROpTqZpM1xWZ3icyvpzIA7c2Q7iODWE3Ymr9Ieno4hJEj98Rt
pTVlY9yOs26m1I/HqugIwv4RjYaXHAP20lj5U7ZQW/0e+B7Q/6BBPFNTOgXPkcObOF+1WIZ8HzS9
64OZdwcgp2TkWuDkjTTFyExxEdM7nzE0QiOOKt/HAmVoRsii7r5sTwdoxnAeO4B1BHttz1axrmbW
sfun64iRxbM2EKIWzM5ePEUTuaut4mcYgpqprQo8ETLx1dlRCRK0n9LDD358lmc/rkol25FcGIYw
Aenfwl9xLdUL7E7+I8Bu4+EzkuOx4lGyy5vFkRXPUdyVyE3Q0JrWRu42zg63uBaqdWVgonXJl40R
jWBvC9ZcmxiC/74Y8Hv/M4I5LXxL2UcV1RWEUJtog9bPgwxlwPoIk79udNazH2xirbpze1WWnIii
8Bvx9p3xOuJcXOMXsqKumJzPOFJJyCTIYh5yn+SW5oJMgOVlG2qJGIfjhhONZsr0aMi5gUHzIJz6
q3Zk8sq1eV+5f2ZSVYJ8boZqh7u82rqFVZCRZvCIzOqlL2XtYQP+DOf2R/5u5eFHOESHiAS8xBto
uEPGRRlPrYVW5Y20I++k1cTgANKX4weXp4aS+fPiFGqnmGJ2kMYEP7xcklQU59ktC4qHFzI7IjdJ
RcCTR3Somcn31nBaxBO/QK6u/03VYYWVtv1bByo2ELFq0dedjg4qBmuvyzBPqiDxxq8tDkjdnoD6
OW9osxtEYN53Cz7lmyDL00t5+x1gdF52PsNDetELkgCRGljS80I2iefQZGf1Tv1G0ivl8BzSICim
p60SNWE5PARG5lAEm8QjXPDnDmuCbYbvYDRSROK2Ah7OOvd7F78QwiA1b2SVngjO8DAE+cnkThXP
nq1FosP+LwQPPoMQ3k1FK/pBXVG2ghG2Iq+66q2QfLrEykeTwIAcj0ESfgwppgMD9Pb20Hjg+XE1
Tz7GhIoYbOuXtZ4shA66DsL/0ib0Zw749aigmhZPN6UZat2oXLpaCn4jjLaiFC8h5ncxblfE8yMK
E5YW+ufBAPAD4Hy3AMQckAp6Fl0iOampUHu/lcp61lme3ejQz+XJFnxU6rgSJXbeFfgtemrAwOaJ
ZNAJwVEhm7mG04JtRwcBmvTWeAFURP/swyPZ5CuU/VTc5Yx2Vh3RK9a1mEHOCruvU1udUqBtES1B
UNTW+d2skM8NpzfxNP8HVtdD+Tuki9gfufdwom2x2VveZzxxWhubw+yVijzsDbB/wwhx271gejLE
e3drPZ82RuY9VU8crmjXfToxzqMTVonzenW0p04praxjnx9Z29pWBeJeFhzw6beoLB0xwDiXxZHu
sFmoYIUb/FCLMkEOiYVkwfuVJTt5WlqVrkoW2bWCqg0tVy113rDnaWclEhXU1HqqTxDcYZkvuhow
AtC4+VThYt9muOdRM+hh6bpr9utuEFFOjS9jFoaPiBelnp4GDgwgyA4IvLbHv08lc1vYr3uLVxAP
XxXjFmT6nQ+14oJl8NaaMpH1E9I72MFUE46p8DkhoZrzITgt7EYjk0ITG6dIb6/JR0BOGjlLopup
v6+wZRHFzUXJP5aefe9JFrznt6Uk/QYJwZbme9bihRwn8xyIiV4lPF5dT115MlBCr3usuYa7dXHU
HpzU5AKG5DWWjQLzQMCi0Chl60OinIkkqBaJvgAPdtXjC2pXug5PsvwqpivJ0mC4oM//BuGL2cQm
VWrd7kkG0nfkIBLhTS1XKSbkvny853n+HxAg4Q7K5EyXd5IjEDUHJdeOvOfB2YiX9U6S4IE2HhNj
d67tYzEwpcySoyqZSxFuTn387STx6GuMLeA3IrwGoayMRqz9ngZM2wkcqDe6PvTgyqiJq3ahUEPG
nkDBWJNc3JNB32xEhBr0QV6FgTkk9/0np7snLFSLPZbpwn7t9X4mEvo0Ag1IHoRXoVHe2B0xZuhi
HTUiRbCvC8f/ooLM/RZi3gt2t8eS1ViLAdqojrcV3G4x8sDSOmTIsrWW7l+Qs/fomieIa4R8iW2X
qpB64jO1rS/DGcNdIxklFoHtRFyxTeQ1sSrPpCSqS2oa0f+fC6RCdeTZ2MDDx+yP1vMuwFjLvTec
jyZXfgqNpeHKExYO+Fe2PjbG4MT+5/lLy5z04S47bFNBkfd4OxZ/vza0ed96K9/34uNutvs7CIHI
sRtDhvfX1j7QE/yMv04pcoGsJYOEYTShkgDRvlKM3FHZnl7eBRJ2sE8a64aKXyR2ZMgUKNImiRJM
NKhKO+Y+H9gkkispaj7fRBEl2Yvj8hV4F5xqyYj6BJJ8Jx7gIRf1S5sYf26JUfYY406/l629mQdP
r5FR3CYqhzGJSyXFke4PH9jGHc2IEMfsPpG4lccEC2ZtiwybWbPPaT9dZq9YUXiXL6IjGQjtLjl1
yM9GQwy8s5alaRy7SovUrLeeaRILAdwRSutcSFS/hFkWA478EBncNsnHg/98oKso0c3xnsgiyYm9
n/6k4aKqIEFJHaml4j2lOqTSBQVGH9FDVH68bPLI4F7W/vsF/A2Vapy3pyb8kbdOhhwc4Mu5fuhY
MxrwWofz2vwJk6LxvMOSDe0hfqPhuz9v5O4IC8ErsYrraTJcKucNa+q2rUwYZOERvdGVqUN0G5XA
oSEw9i93dgHePPClLEO68FDXXkdar8xM3/kGFsI4xtjwAAA8zkghwO2HIFW+sO1I/3tSW+60RMSg
RNhOw/A3kSJqJWVjnyOHNEc2968dvIBskxt5jWryIHguOQNtkUkHy949OHtGttm9zFI/O3Mf1fiB
Pe6caIXO9gG8Mg8IDxPQ8UAZUvLpl2gWsYWoOZt0bg+YIlzwj5INe3bt80UyQlpK6Du1tqAKjbZx
RYwxd3TPSvjyZRYYSYlhm30hilc1oVlobBXOvsiIEMGXKJulIyag8OGStcH0+Z1X+EGDo0OM0a8U
wTDbGAbnfo8lOL79KiMn8Trtp4uN9NIfc1jtSdnTZyNLXi3b4jdNmfWDmN3V9mt7s/9KK60uQ5Ov
Nj9egWI4g7lh6jVVNX2kIYQVbUjuJAXuZobEhq/Ee8seLSOwe2jPLHvmyMcYWV9bVxlnTnQ9fAAq
X+NTIzj8x+Nt8qCb5eNqZtkqVSteHWruLP7UCqHMXzU5lQny1u6X+z0V91cw00Nkun3ClQTeyDBc
DUzhospz49Mb0yb1Qtp0dW9+q1s1k15ty4zOAi0flNcAMgvYd7zZw+4xPuupsb6E1zzqSW6myDCv
5XsEh/XpEk7Ch3GdpwO6cWC+cxitt1FFxM1qggv8RvYNLhA8K/j2r1igo9UHK+eao/LvAvcw4CjI
0z2kk/imsoWaYtI/FPd5oGBSIjzWecqXgfOqKUGD0YAfk9WHZJLEKpY4c/l3wZwn3Qr+OGB+MXcO
+W9ILmLTUWQkTmr6wYRHHJ7sfifVriqY1w1cfD5aySvTIHWv50YLmq3wTEFNjPq0IublbokN6aTK
/5PkAG/Is8yMIuksyMHzp9lQty4aUCsXs2w1gnXcHNcLKjC6y1MjjtO0P84pz8pUo4SAQNKOjkgc
KQduPz/zMUZ6Unm+EuLYp9DHdR4hEiVyky7oBtool0PU5fmkUOoxeKTdHVN18pFxKiAQCcjSuAmk
m663n+vkv9CrVt6F2mXkmObdsUUj/oLbQ9A8504S8WIJddSHnDP63yBseJ3GjFl0yGpU81o046aK
Tvw1OjGOrohtkmqWtSbbhLx3JxJsv0Ev+Nrwb/kn8a0KuZOPKoxsLH7qaITnHP4neKYiWEJacsmN
X8r9vygCHd1oELVcz1t2tO6FomSvFQJ4cH+xv0wwRrK0MDySr0evSjKKdbA13e9zwIe/WKOjeVAM
1nMOoq8RqHxCDxxeAb62M2jUpPM6y+sEZY0Zeeciof0vWqB0J14BUvl51ALBNl5/3VTpiyS8HNkj
xL9J8nxfg/stXmpfoDuAG5vMDdb/8XpdlQUuk+oHW46V2B0N4ymya2CtmZ0M2zMADqZG8IQ+OLLe
20lPoKL9xQMRZAyML2PYxQye2HmVHvKT8GEGKBllx7ynam5/wrSTqvw2sjasoR/TrgTqrXIMsun+
ec35sLXQZJii1jcTaKKphcsljys0MvL2MkYzNpJwXWFOgjZEcQpQczGqXkU6EFjiFKvgXpew7D+U
0EdA1WZOFCEpZwxkVPGmE8oPeLIr2UmEqEPfGMu5ipitzshfwiR4kDw4ejGPN2QLlZZi2ieI/BP1
Fl27UIWHy60/sKPPKuMOiKQIVuvkHGca/pZy0zOkwmLdnVvV/RnsDR2+bnuxY2PVbQu5W5yjB0/9
KrWtp+Le7amIAvZlrUomCSR0DNL/uty47ts53FQQAucCKjnufzpoL4FD60cbEQrAedtCUuBElRxQ
ixZ4femga6r1koBffK5knZJfW0OhjV87mPj7lJ5bSCsy5RJwidW+Bj8mpYhBFxX/BF+prASkFTAP
85YNyW3xgSjTCL9UckFxgLtO0rBvcxD/3ptGcYgVRKPZ7IXMU+SM9bwElk2e7WtYwWxapgHSG0xm
0+5Y14pUYgyakQaZxBz2ZGCKsjEmsDEK4pAcnVLMagiZXjr6YD9cbS00dRiSPAi+0ZQ4d3WNPJzN
UwwDJz1+3bWWoWgTmHzkQ3zZK8KuXSMmzpdQPAV6JG081Ux6HbQCfbcR9nTP8TAvbInNly9hHmfU
XcfJ+z0qQduYhQ5RxxjHPj74Mk89+6p6bw610pDvaDgGRRFNwMkkW+0sqiOjqQduFrUeQ3wjp1/I
U/pIJTltO5aY1G+csg0TnpSTIO4pZKxZKh6YGoxAwZP6OJnqIOi32SmMrQMOy8aNOa5TZ2ux2fvl
Dt78RaZKnB5Q0099ixx3WhBp9FimLs2e50yngurgwGEnVzRXObWr2TLCupQw55T968zJtp3h2Wn0
wR3cCxm43cWBwtkIqjX9q/AtOZFqX5JA5qmOfV4YogKHUgs8VDMXLWV7e+wXVrtdZPx5W5esDLrS
aEUZ9Xw6EmNuUWvvGVVnw0fPlDG/8zaMHS22tjPWfKqPDNbGi1X44iO+VoIAqKp42+q2yfn8U6pZ
+VSHemqXsrhEBReTbFW8Sbnpm68FMQSF3zbvQ+QX/66J5GBn9E71p89f3r1RB5g1kXA9xE0oKH+l
TiNuBDbQnIobOctqTiL0IgTEgAfEx9XVvTONWpLtEbKPwZmpG934+G0DiQsDLpgzdqHGtbcxOFUz
DdXrKEU1pYlAPqyP5iLkucn5B4pJvWluR6MwctLMU6fzLsk9WDmWnxkjoWpN1wNjonmum+afGZb/
Wr1Oe6Uz9dfwimhKdbr9tbw2AVZQmFF7evhPl0ExOBSW4aZx4Ts14El7wwYTtabCvKku5gt98yek
k+HAvHGDRvQ+UkOJ6sSKs8ZXa37VGrf8EthwXbhz1tGF6T+ve41sP0H6pGlcO1ftDLdiU+t3aYZj
B35BITxFO6mNuPAZFJ9fUU9z+u7VhxxnebbxviebBn85WocbUMhHqssyJjFbCVSr+8uSKHlN1Hfe
J7cd+h49qKPjksg1B9FzP9Xo5BSr59A+fZnA8WgwGsfP85KwA3+tGAZaMGbhrbm7Tx8FHdZBHUsI
AI6aqqoVOB5ZEMb9rIilol5lp6Mc0a0Tg9gVY10RBxeuvGun5/qr6basT4nbtzbAFYGvehVe0DnR
dVxYbwvd9Hcj4TSbmDa+VKpLRUcu7aPMlWFL2q5BmAiOD2DI1r6fgIO22ygAIwSXqoShEKqco1yV
9Bc2fHgKFZH4Vp4yy6zAvRL+jFLDHZ0YRwdUCWgd0a2Ob5px+omYmL3iuKgf4x4dPVo0sMGFs69g
QhGTm6D3/BsHNzMBdQBpaDGtBrNuhcl0g3S+pM6y4wjnf6utxtar0Fa2i4ecs7qRoiz66TtfgbrC
UtIuwoF71epXpXtAvPK+dOKT7CQn3nLZf6/pVzuf2hBMK+j19OJwGmGqnkomhMIswljn66VNS9zL
F3vYFyhz1/HWrV7LkjKYUcHnzoeOgu8OGiePc4XyfCZxIL7QL5q3M7Ah0kN3S8UfhbPYW0kmPmyC
bI8gGx4v9P+BwpOsReE2E3H92OM/BeTawlVs7MS7vEaPdgWlP9eCb4HnL5e0fwvspaGZVGghEjh3
QpxWGfcQK3JxZe5eRMGD080sAWY49/PH/+6Scgss3DHDB8V8JrzLkP0w3GxNnaiN6eOhuDPPLFX6
NA9dfVkoxA55Ai1Nt9jBL6y8MsAsUWIlPfCZzwkLBmlcrsgPRe3pxjDr0LAuq2vD31lnEY4Fux9k
YR6KRbJQQc1VN+XH75j7lwz4XxgsVn9UIRymFGTcIwYJWbr43hlT81/0e147yDJ5rpgRj16mM4KT
diWUnUzxzd8NKgDPQ4i+DPhRVZHWvqnlB6pCvRwjy/OXfgKgM/V2380U8bUN3cKxJNJubEn3CgUv
eEX0IPYwVQOQdYAuokPWbALfLf+X1RKxqnQZzGAQxLI361dMQ1+KATfG6M/6ucyYPU2NK/Cjm1Lb
ELiHMxxbavetu3sPz99AqWSoUw5R3Rcx+/sNvE839MJ60wfXkKYyljq0NXKo/1/Kay18/FnJPcqT
ho+QEloj+16HGDQuKrYvjePRIBI6CNIwBlAuBLD0f5loJVLDsMnkngk89DqD0FczdU0IInO+7/7R
M6T11iIIDP35Z04TttOi5Pw6XJFcAoOpjLUAOkyFAX7bCdMx1lI+oF7PL1hJ6v+jLyP4DUbI9+sC
JSdK1LYr/j4jAcBRRw9ODygHQDVqPuLUVD+EvWdOJOlDIm8hjQYEAAWAqaoMOP+eQxNoZ7RXMweF
VQ1B6tRGW5FppYXU5n5QRiQDRqr05KV12rVmb4gHEX8NnuPCD7GkA7OO1Pwg22fdBlnCQ3e8fa7t
2K7a18q/5U8dIexPR09w+fDrTyRGTbovif8IrtHRggXbngNFXgQWdQ8k2RPvFvSO0kfMRaft1+p1
F0BsjcMhd6z5MjDc84bVp9WsBnPw6Q/3FJUrG3EtzoWHAGSIFUtwzeJrJJ5xODKsDdFt8t3VkibW
1DYKLvpIMTXtOQdrDmY9XcK8PXJDWvds/j1bdFxnBCXjFjcx8meYtMDkQEqqa8E9kLtwyC3PhziL
y/IN5SePl4msu5voQcN4BfXt8qLIyo4kuFjz4XeFU8N37aaAjn2nQ7mPx0FUhKKyEKC3gcUCZMx5
zxyqBMaOBkYWDGcqDIOW5PC8bQGtp+WOn/EElTUJU1AwwrhWx4QTPjf0GIYO9Co99csD4bl7E57e
Lba8xoHyLbWFTPvS8F7m/z+DXDxIX4fSk8B6AGQGquRGVVIkz5g1vp9ArCl6v7YdknehTCa3LOKB
GC0pey7sW5hOjKJnYABKDvveVM75v+Vt8aEWWCrAkFj6bovjdIqtSL+b3EAfSRMxptefraQFHKQN
BYlrBYN9kXiAlrBOFx9lTjxxUgpjYj2+O2EAMG2o4y4g17876oYz9YMM+aS8BVdrJoPObuCndKal
LLG3HXs6vAqzRkbNU3IA9SJLC+NRizGrq3yuYzFAlkgId7/xCKLRAVJjtwYYqNAZK2J46pLg54ka
OHtr9XW7eMxOcDje1Yvv95pyanqAshBfx2SgZWyNI+lxSj4+WbZAkLtvQlxMB5z6Q33pgeXQSnTS
8sHP7NZg3Y/SnaLStODVDfE6Ac2qcPMDCgQt/4dJJ5JEK+1w9GVYE7RmckcyckHAI/1VlzBXRWUo
Ci6tSIvLpG+fU+BuEYKEqPkoJbmUbs+OIknR2CL4fYM5tLSzBwfE3DDL9Sg/FEmDgMlm7ZpzVT1w
jzz4sIB7zAHjgk4W5bGxa+Po0b6Cxld9DiHNAWOEuB9ovvK5RdpiCXtb2PevByl3uMxLmwcsvyIq
icqDQrLzkX499MCKkSxtpt4oTdoQ1JLtJO+6NsFYX7aAe+xkQmJIReoi56Z0os/atfNllcqhSuh8
oaZm0gk2qnbFhNJoC56OHAiZLyI9JpLFZwg7AGqVSoKGubPE5tTwios7DGlDWU9OKb2yU2emfSMm
lqhToehXnbKibN2lSimkjb+VJY7GnE47PH+s5lftbBUF6Cc1tM6pANeXqiXRphgdp+m/p/eyGk8d
921PDUcm3tsnH4cVEwK5Q/CDZlWUpzlvtN3x2tOAsHUJ6KejEtgRAWd/4SSPr4qdw6Yvo7KWFM6c
ncj46Z9N3PfPLkqR9p9eGbDkmqF8ZAwS8OwXvqBHfnrB1gGe4cb8grPynh4FiVXjLs51q2bHBQdR
U9xH+64Z6OPhKV6fWlmPADkNoDeEot1YmYgryh4bIQYGR/JD4eSC9NDJJhYvafI6QaJYsAfvWAVI
pmRX78Gz8ul0VrWP9I9fYEAyxXvQSy0LlZyFuoDM9J5GEkJDhqaHiKyL9uSZjK6OCLEoMFEwmUQZ
ICyu3z4VhUKvBu89+n4AZwhkLOlVHenDAdMT4YA7hVbJNPjVBewZqCJovlLA4PdzJU73RWwG4NEX
pOlnA5kXPaogZG78Ot7Qz90pH5ZNokkQxucZicNZNQ8+FrnVY3Wh0+HO/Y5eN6UcFXaqsx/iyqdD
bsn/6plxQ2zO0etk/xKXiw/rUVXmNxT4MpXkK+a40t3rBFAWcl+vYdWWgF66yBhERLajNUMMk1gD
TSxnOaO6xLy1tGWXVom+NUiLmLlJY59HwwLGfFGiEGWflkKRf6HOiAs/7B5rcmMNiawsdKdZXg1S
OfxG39lDLLLn75wIfyhu0SWdtrKRPIk/2AFrgFzYyLRYUxz640/vk7R7yi9eTKfHsUo3PSlTX3HE
J+rZwLosDWMraxougn5SQLBB9eQWvbp9rt0FtK8On6PplcxOy2GtNXhJN8wywGsGWP1s43/ZRee3
Gp0w4llb2E7NjFwlWRmFcfOZc/jMKYECcLv/q5hgyPfXWK0w01tYzz60hb/EYKlrDnmP1adkaQgJ
ztnKa5tiihXn8aZfHdL9kSGR5ghT2fSG/x9iLPkOHbxr+jTKBgZQMlwTgrFMryY4TR/IoRy7Xofh
QaNZZIZBbBiMrBQ842wH5Ex285ql20mDiTj1aVgM9rdrpyIeCP4vhE8P1gxxNAp9eWMGHkBG+epy
0rybiFS7zXO6P2iMt8dIltCddJ2TJ/mI4N1fr5P17yEAu4mm5oBf+X/eDv4mOouCCvNMRh3Hv999
/kWVIQ5TP8O1VtikhUsiOk+XevsbdRuVUHRMDlhg4QI2gaV8CjEJiMMnuSlzdnLGoAPLx+jNkjZl
5pg5GvbaL+h14KVUTClNQ+SD8YVC13uLG50JUM7mbn/25AFT5wxTRjerUudYBRR6ttxyxav2lkaw
/k3XUghIc+SNjSCoazy684RDufGPIabQBWSgVTeqr8ppPVI4EPoMHsGTlMQznouj7kIYhL+mONNR
qXaTrJv83JRbor0DX113uZpn2p3Mg/Z+G+b93yKLLF3tJKb70zwqjIQnMRXhkMH+SyJtRQ5kE4+S
AN9uviaB9QgpasgtZH2tvRNSvVaB39ES7lEVxsMr8++teOmBIDHTDCjFR6xI+KXYld3viRs2o8nR
M49VKBeB7SOl22wdQgKnX9BCO0dgPSsPpXlrv9Kq9auF4MlRYuwmtcv8djXTExnh+rx7JTmDMrI7
tmqrzlpI+gbLaUAntb+rcnomGOXE4KcBx3psjrz5HkWmhcgKEWVbXr86DZoSY3YYtxmE00538O4m
dhUC4sEhkl6qphiEsWBrVL+ydFuKAdSxZHsCDCb+FiD42t+0jdqIngSOH7McYOAKPqHBAxfhsmgp
sUXJ9lgHEQlgVP6nctodQjpLqMYKQVJ5rnr/bmG9Ltf33ESX2zu/bvBT/DHb4lqgxzgODXjw49jE
DjwjtaE8hk8WuRrYr9/SjvKhDXQsCZ2Lrl2o5FBUv2Zkj6B6tIVCyrkFavJTDyql8kxpEHfZq7si
vXIQexunw64oVAjwyyvc6Hk3A76heJXPwDqeq1SABPjaEVK5jlGnNgi4ByuqV0yqV0wjkXox7nDw
fmRfGlQ7yFIRdBbydqj0dGR4Vvf+9iTe60Tl82Owi5lCVYu7lmCsqbX27bM/Izmr5gT1+/bMUU9D
eRdsTHyLV8M9BxIW7dbXuQgWWQIYSWf1cDlqba6czmfJ+9xm/FGYMyMDMq0Y6z1Uc4vQHxsAY6q6
hA7rq3SsWZRxZZDac7VhdoXPyStUBsWFH+d3oJGHRWEd5lWHDLyGJJURXAjF52wIoQGMOr/YJLtP
cV6fzP09axX46qoUHIgMzLTuZ3ZGDq97BtEtdQhSNxb6u0VsUpwyjUQd0xs8uM7HSsfh84yZfggc
mjh1VnPp2QJm+N9Q9w93yzhBwwFKOp2BVhOZ2b02NhQfjcWzM7IS28Jg/A6UKMLJoNZ24qScXZiA
rJ9ByljR6m0llksXnmEt1UQrH3hqHPW3nTV3XKIaMqOyUg1LhYoqw+ExchMvInYDJk+JEsLLku3L
KysNbG+dbgxfvFkdv3zm8HcjEOzHHFos33peqHqnvaaUnwM/3bkAyaVB+diJyFoVH1fJbXlHuhxu
nQ+Isb6qHmzyzMwenDhc49FAYYe7Wkx0utMeeVRBDwP4dJWL5MLPYLYK5akWZiL3QeGfXBOvkhSJ
ZqG6Aed6/JTJJmgJ2hkWPJOuaRqUDM3moAm5V8Bf+8Nx+Ul6CYCg8tT7L76ev1kpfW2YHEnHRZY4
luCbKxIAzxY4OKhCtBF7wS0tWkIfS9EQkB4iIM2djfpg8f4sNZXZTJrK801Dnv6BUciAI34ZoTr6
471kEL+SuSGopiyst/IxPd5WQh+iY872Ke3gST8lH5wND+izAleEraUmctSivY/YQp4gxrQHUWiO
NLCfitJw8ghUoaHIKIq7ZRLWZjMtLQX8EEq3h7gXOcFmB4m9JUA5jMVMHWaFVIRe8OeKUE02H1f3
UNVaoj8Iu5JYRCrLpEUFCYo7GMq3pnwcaZT7fXofwcFDSuTFKiuo910VHgiEcLpn4dHunrk1bwFx
UusFn1+wlpZvBSECSiLkfpY/jKPUwBKks2ZdEiLkhbqiJApxG1BNB0rMYdnE387RyMSi/058Eo7O
T9IHdG8oBP0GwfLA8AtJWRaZopA5M0ijWTlKRmU8y0XBC71oIc2akTAWXjLPc2EAy73HMIGETdFa
/fP5v9uPYNEcKmJSu5Fk9hG7Krx3p78N2h+DA3c1f/OLrrCcqbzdtdEtLOekeBNFozMFzNKyPwAZ
aKsQcGmB7cD6K2dAjVem8lJeG8q4Cgad8k23RApKunf8GZaCVhKFXPxduPwmpRI4DzyU1YUpJxmN
Cqmsxl1n+MCiY2bhXCCKOAqydIjO4tMrI8hoQgExV74JF38MZPXeuBcbfQcI6vfIC3dwsKj0wI0S
lhGXHZV9bNg0HLpcO0Szt6Pu3wTxwThodw9M1k2e2y4mtsqzxds82gDnGW67UqDXv5X8WRG656AY
qgfEKE0j1f8PAZPRnUWiu9ydDYbgsxV0dk7AttqE6fM0fzaZIGaeK0du+IWvJK0tySmZ2GHkV7Su
mtr283/TNCSAb88C3WWI9FBwXqxFUUexbgF8dpJ2EyPiKxRLEsZOrmg1+XAEtL78GaSuX/1v+qqY
sxaPvFPl1NNAiTpX3iC6tsClTC/kcuGSAXFEEoENxhl9bSZIOJze4WVJWKcqQK/rJAehuzfedhrs
DDrNCWdDdiPXMzAMbakqUWRoC21Lw7na5L4UTrx5MLoXuvfScVw044CsoJidxGPyscf73PGeWS8m
BAjGitKpwOmazcWYv8JPuRxNAj7MUh5G+aoEdz9d4lKdHtacZP5XYvWVDcbV1150arR50rafBoAd
vzRPNMnWGlTfElPQjd+j6vvcnIY4uaj1T2ROXh/IUI/BczR6+vcF5V0Rz98DY+ERTdCmIY5aJMNk
GrPtrqK4xeYWVQdgALrEMWdQaY/FptKA61lJhZgZa2KmsFiK+tLCWaqBzfx8WYsDA4EGVSAzx8Zx
khu24eeMnuEYyORLLzPoyAhYB2y9Pa2pLcRqJd/tFIXha39mWD6RylCd23SXbTRG/6OdPw4qqprf
tikvspQ0IlmnQ9il3HCoLAbvylEPuWbkPn+tf3MUG5/yY1hw85paWspiQ3XMcl9X0qtqghi7JUQ4
KqVMsSoFvqjQthzFBHG1OBRfi9EyqJxSLwQppgPFvGCzi43DDfyd4OVNYuPt1aVun+pY5b9pm2Mj
2YJPGt2ms5Kq2UOnjHG8zjZkYlk4hDhvECs+V3M+iHiUbIRAQytXET+DKnlJ6ukJ3XKsCc7b70kd
TANB18rACbIg1pQzZ2N1T+W463Ic76qwsRsuo3lhu7obW6cDepvJ5ksBb36rB50Ju5ePXh5Hphba
W5zijayVdeymmaNt1QAp2WjMhZCdjdNkWj36ZZHMaOATvZhvv6604OftF1Q3wCEqw/03HY32febS
QQpKj3lJCATCBm0a/7Dq2zKshtN/1oZnmpyginBBZYn2woSFOabobYgQ6ToXQYMQ1eQSVOEshE9H
nLIGVtlcpfiFkb/SNqwce0s4ljv4WDzyj1jCcPj7VL5GiWJd1zSZP6/yjPFA4xLIOM0tnpmQEPxH
ayECgIOBZZzE/gdO9wc611o/pr/d/VwAyBqChxlL8PXmK2UAOAtxoiMfLTjVOLHtgiw9Pc6M1bTr
7A1LmX63Mv4kbQMMMKs0JRD9OXhomv0xAHScKHpRcNxYwVPcYapcC1I04aPtk6ukc2EkLXHCxnzS
mALGgdJxD/OZr44M5ozmL3L279yiq3eaKAvT9r1U39Ss394y2kMmvh/8NKggNqjAXm9pJ4aAH60T
GHELY0emsihNRLL27V+PzxXSNRctCIqAzbYyMxkF2xNoUSPQqTxCV9S31eCqShnJxm0cfBgtr23s
2hITMrTaJYTjMqG2qm8EQKYqP06Np7N6itnwRSbrVIBcvz2Okkg/R1j57NU1zptwgvQ3nyWdtncv
EZDmzK39UzVzcHd19GNvOR/MyxAXU74/yuEbJNQZ2N0EvziX4RFZKRaD5D2NWlafsTn7M5NJBcKE
drtWqtFiGZqCD2l36fKxzlbFf10sJsMauiDSBG9suOjLn2NHAeGl1UXNAYbc0L8xFnujmSm4y93t
aYKSQust8x2rYuWzx+bY/spQPp/YNe/LtqUmt/LDiwN6MBXCiFRBIhzuVetZy0apyOZwqzqspJIq
RlexXEdsSkhNOLS2/EozVMjV7FbhOIq7Rv/9FDm0wI3S/W0ypzkM0EUjDMREs3r1TWEm18g8GDzO
hndEZfLprY4bMYpXNRtv1+uO8+8wsHxIVLzdoTA6AjAsFzM7yvGa/F5DYHA7K5ye0nZBXDm4XJht
/TKZD+OEQvRwtZxTSkZMgby3gsy/m6vjPkLksbKcWg6ma8jY8wxFXQr28taMm3ue/Sv80b1hr8j7
vyHpuNQyW4CiCU7jc6k/Z+xQTW/MnrOR2LJIMrUt0xGechb5hhaimgBZX7UEa3A1idrQqkPoB/Ee
teIszW7f5M5FuR7bJC0TUkSleoKojsdZnI9Nns/FCezm/6VhJa9NhKc1+eRA4jGFbOCK6jp17QD/
zvuWIJ0isaq8uVgmxrxPOkoUzrwsBMJYuy+/JJmwGhiJxgG6MVoTxPCnVntbhKaFLEwos3Cpb8pY
ofuT+EAz3OcR5pGsh5mE/7mhnoSzPc+Ngc9wffpLXKzL2mpnMJxwH5S0MPcYHLU0eJLmpZUzYTEM
867jc3iPRJ9fNlGbcLZbQyO9kO0UZlsLgfOkSReXdMryUBrADIuj8bGdDKwaaNhacZ0vld5UjTra
B/Qttr053LDGNJU4CwEGUZEEwXHg9k7n4bqILhGC7p7jYeRm6E5pwZjRPASBpYdPvMAJL5/Hommp
skbQbVwP2O+3InOQkmohq3BBAHXqVtwuWQGbEunlNSX7B1nz8++NzzPIL2vpaq1ZemCCW3jpmYR+
YvSkuRSE8M+BqbVyaIfcMqLRZOHdCVGI+qY+UV9vQQRU9YHZ4flVdoSpPII54cjfkUXR9zIZlkFO
n9vt2fTkO1trvguV48RKuOi1vRB0E3SmTw+WWsQgtXM2dknzqklMJEY0JIWf41UW0kthX9q+/EEn
fjUVJpUBA6c7SYIMGAdbwoOGXV9AnoGQvjTKljfPdTYha/2B7YUT6VxxZt8JZYbjSnVCAve4LLrm
mfrgHPqfCPvhU/lXAFaExFmzbXIKLgse2l5j44GGSrvt1r7FhL5UdleocW3ou3UelvBq1S2ICw9P
Rhmz+bPXBRGfKvmxjb/UhLxw5f3ziFiMGLHQ/7aR4WqNKneg/HIxMvZCQuWgJcpJ6L+CodhfJ1OS
rVwQBdrUZ+N3dYcZv6IT+h6zyfEBhpr863FyaR3WiNI4sAfTqAhIAQM2n/rmdFbQpMnri+WUKV9I
C1hiOoahwuQI6+AbnezR3WJSXDQFdpTxudCu2QTvU/77YQiu7/cyO9B8mQKnjKY8S5auyn8fJPTs
FL2QeBrNP/sq92/CSzSerHFvkKDLmOZzMC+Km2lno9pWGkzFlCh+FsG0su6kU1FxxpSEHxnnrC1G
dWyL9NXl/R4wLxghBz9zISzrDjX3gvFipZ65Uut996OY3YWt576bqolimuZTiqgD+OExTLJmVsV2
f8qsP9w97npGkAU8wwss//dvL93RBldjfiVSIuL6ljoownf9aCIlmeH9uZgeAYFRmjKnp29bA1Jz
3KOtbEvNuo5ew7I0JoE4340/04wvBtm+PoXCRxzen0knyI7Za8WlDfhXtO4uzW1E3KjNTb7mRYMb
yLn/f9h5RMgMizeRSDHkNCVGYPErPsdoKK0vOWWU36OOLZVwOin24L3hR/BfK3l5RxbU0PgtMocm
L0Dm6VQPVQIgTU0lTQm+WzSX6FRiQVqR3tIqrMHvQey2I0LTLswWRIrR6T+OYviqiBoPb1i/KyMO
qM/AeICCEmvMqsMLzt9AYldVxoUiPOmw3aXJprWzac8eJDUGbX4y431hD1dqQgfLpx++TrQiD6Lj
/tt8KtrZOM9PsE3poPc6+LPxHhbeUYc/baN0EW7FC0m0buiTl36/ZHaxwzcRVNjFLMvd1QhZ7lce
Aal17qVjzPFHCFxfNXJN418QjO4GsV05CxpX0zfagqPogdHcE1CpEh/VtyOqpK+XjX2QPpGpY0kc
DXOT+TsWPDXHSHTisl1aRoQeWqohWgA2viuN27Ve2bOZAAbxlO0/QblVoFJuHsYBdoDyc6fHKqL9
mvFGqqwFix4pEarpNyS3+qJRu9OL+wVsKy5Fr/pSvZdES6Jxf7okp7nPyg+fsXQ7iHL7yZ6PBu66
0sDH59Q6K6r8csQhT6LfdEbxUDnfakAie5FX1MkUfH4lU3C3K72pA87rp9Vr6rx2laDD67HGN+O2
f9OAnAmSx2C7Igyhw2SToG4UiI9k8sU3B1Hcp+WepToIeUBlqX+ehK12Jtoh8BIqLjfPgm7UFLii
ndyEeTsQ0PMla4GDSLHA1PSZzuPFrh9dxNu3h3sMnJsSsXUpdJ3MaHVfYll4Ijre7tvNNQ9Nkd/A
H+GCkpJguSL1jQJJEHBHPf8TLOy8zweZOcWyw58AVxrd4Xf2NwhzM88FVTq5CLmJg5EfRk9/zLyZ
TKPwSsj9lNckfE50CKwHEmntKHqS7txgthV0AXLQDR25DcUjJMV8fYtnDwKuJiOnVYB5pBPnkTDD
e0DKBmG8Xygb/gCDBD4n0y3+DygTfBRERj6IH1ihbJsVJ6l4nCktnJc2uBFaG0WOYvwDAFAyqQr7
ifov/G96NQwkl+BRPSW82uNDPIlwPvsl4KfmF221/KEWOsbb+vmhggjR93GPz5s2q1EgMF9pbxGS
dtfi2fD/ZvzXC+VvErWpK6ishm9O2OHhsq5uus6CVFyawtReSZzoKLXRLaRzyXZdfCCBQbV8jqwq
GUUkzrvaFEF4rNOdytmeiNtm4hUCzcUTVT/g7O0dFIh8RJ5W+9MhACkHPkhLiOh8ri6S/vlHfcbI
44gUvQdFbtzALhh/0sSMACTNxhMUkf4JN3XvOdT8onfrQYKs3R/yBh1Hm8YIIrnv8P9g3UQ51yIU
2P9zB4OS1IJEveH5tseybmz+9Kir/K7QCwNPTcAisWjKF9Cacs9ovTjY5MnoIrd1gYfhUz1qzLyp
pSRgg9RXx0gB9gFZIvnyk3MMzcv8L3W1MMb2/ArBzzyUE+EgGu7C5SaTJ8lHTEwc9NdobgdNCRNb
aXPkfSGcRDTOI7pLL4R2cMMeeyn4SIGau4hEg9BUIahdHPWRKYz0E46mAAMqaH26a7ukkDEAGM4/
JRRVQo52hOcXQiC7iVKG0V7/a+SSYV+Qoa7MYSbRrtsNya6MHRBEhPA0VTe7mY5Tugkw2WBVwHop
er1e5VHnMVcjV6yovrS/anvMDqNTZbKH+DTimZP8WApi1+R4Yy4CUBjFcivbZ1jycE5MqWdhJr57
G1MsqlcO7nyYHM6rfQ7N7re04oq7RBwZmaAfK3WEtUxbJt7Nn0VvRCAL45+AibME9EeehczSKDCG
qUtb7Y156OaYWB+zTk0v6/QHvN5HyR1b2Y8EMhpmKrIsx99hGd80yWod9JvUkYZgEjirWwMduu1K
dIY9OcC62xe5Kpm1WLDbWOUBFu2aMSfzvjHrSu0adocj7trukR7Fw0fyGpeseOr1wd5fgySfBPuy
To5leiBHVZEwAJT7c76dar6nLG4sDQKuiuzU5bF0iO/TY0NKXA7TX+gaB30szcpV3KvFIlxeux30
cF+Sxcy7tRpdo3/s/epFg3ctN7Zyo9Sj+pqU1JIUqfOqJ9eyqDgTc0Li46ThLoXY/5nvysny+X+k
D0MzjXb1RRray8Zv92KtZ2QaBUJi8PvjRQ1+W0os2FwyJ2b/UFPV50GOji9JACE7vwT8YRyclnNy
fGLOeYA7KBUiWAj8owcqWwU85oaCwZGH61cBH6DnHQ1cR3VI5DjrBrtHhADTlPqRpOE82Jb0hiyF
GAb05A6sq66SIvFX4R3vG/vjv7kEmwKwazrO8ngP0bRFiiat+MCzRRgGId8E0B07brwDwayUBASM
gsJb+nBdKfDBcnFhftLH7w+OyQf2/zXr1fdkl2BWQwuThAfWl/IWBQcLU/lyOKw3o5JuGdi8LfMI
YXJtoZbcEAaXcSKklVay2BpER8pUo0ic4qQC9ry0gnhjXRArkDChw/YECB1+63w7at3lnGEnbKQA
wHTch0tEy/ByVDSli0EO+PnDbs23y/VqltYVF1ut1OHhIHWHPPW3ZGxktqHSFDDA6CUx28ESLUpu
FU7caAE89Qshp/zNlQxKNZslbwCK4n+B/HU3vXzrCjGlFF5jD9C+SE7Hge8Kz6FyunEUUC6YzLqc
lyQqJ4yyoKxi7onFj3zMU7+ZCAYJEEaoOz3QsT9Vf4TYDSm7Xv6K2AaxQJ2hxSuYLIXRWI3hinqW
xJOYKdwpncVD5bUk+etNzSjUqCZxqgUI0lVSB7B927swg3NW2DDO9JRh4CaKXQQXapJDOSV+mFSB
9SvYU6pby8woO2BidzQO+GYOKRVa+bljLz66q5/djbgBscXtnGLHc6SMMJDA0iKf2Mbsz5aLPHuM
8hbFSz1gp/d2XrLiKIbeGWcrQeyCmzc0FumKnsZMHgoM0GN58MK39VDnKgKeTdHvAMZJlMvT0JO6
GqoT3O9wMZKvHRpumS3yKrav/fhqbFjOtdeQlEM6Pw+ZvcVWeWtSSrnmo4WMKaqzK9Zeug+gCB4W
eflClxUY518z8MdR0bP4s9CyRWe4fHijquz+uavQR2Y2LVcbI1inrnuSKurK9BiFsTT8cTf+uALX
169lYwm6NasqRmTMcOAXeFDd6DjHWUPRkif4cyoACFmHgki2CHiNhd5ktURpdaA6mNwJwsZYS718
2TqWqmj6s0Jtoqq6heBwWJppNsM/k46ZewLRKH6hEr97SIsZhkhXkvbZdDRTieqLR59a47jQNYLf
Ofr9qIkbffc7XiT2eS5CI+BMvatYxiBNDUvJs1Xe8vPVVsbcsDx9uPk4IFA1Lj7okrPNY/lcQKam
ZK6PqZkpSvxUnBcDH+qIG3VRyFXWs/7lbmF1Iv7A1T6QZPTniaVjx9DpuOIG4q03SHXII6fJGYwL
ARVHQcWP4CSHlwmHK8OgB+wR3dGsvQZTe6Og24bjvFoHxTG2bLI0vCZ9QqvVL0P3CQdFLzKXbAsU
t5LZypwJh0UQ+5BA00+CrlKUUOaKqwpk8M5nY5pRWGX5xoO46fmtMDHOtHJjJszYzyZb6WXrx4bl
WdSuK7pUgj9yk1wddNK/oR2av5kGsYglohRTbA0lAoX1+bF29JeM5dw14FPXjyLipAuCNV4tXfrs
Fh4FLL2kJWOMkXJf39GhjGEZVmU+vqmXRmMxB9dfXUnyjSgkbg/NgKy6SXBbZ1zn+b44r2ayz5XZ
+AzKZTB/sp7Rn2rvoYoNJF36f+xOQ50/7JHmc7Xy0bd61wDV0x0h3Or9Uff+9QWu/caeBC0fMpNH
fex7mgr/EyT04ygthFh7hJkxe3EVAJZFh0kOMj2UZqODWQ3BDjr2T1kQmD4j7wD+TANJEcT7O6dN
ArTdxtf+5coXBvcFyTKLTZuDKePBEWnLwbKeCbEpDyFEENI++hSWG+RWy7y+Am5FzpaZul0JpTjV
3ohCb2IQkLPIlBk7knijkt7rVbF0Cd1MC0KgtNQHp6EcZbvF5ggqdJ3TtRlZEIj6Mir5gfoHONw+
0nb+tvZI9Ux27xgNakr4KT1SHeZRhwIzd0XDqEcCG/l1hdEQHH7a3joFX/OlxuyPsd+mb9DOLOIw
hS116GPA0kb2MtGjwaqljyTXm7vGj4eHDdZxZWhJgwc3n17JNHa3ve2qE8sjkboxg5HOBfEkVX9L
XF/k6n/gRnuFoUzTviThLJeZAJovAvpUKQdWp9lLFfJvzzQ0FoRRctCiaaAiviKRrtpgLxTHxLnk
ku2XkrQhU2ooFF2xFcOyiNYYXwGNdPYgEqSDDdPbPAi053Pvp7t7wJSNliweeKyW7Y8ePeAeatug
IzhWTfqTs/+AZ3CLlSMlu+F5xcB8thPGWkowMggCBeDXxg/KZ4PukH5cRT/Y69ewk9H7X/mej7Hf
IUYudJa/B1mt/eOLIkbth6AyPLlDUYwhx1sH0YwY4fqk50jt479/KBawZwYKgbTbpuW1QS1GN6c6
x0BrgxFiLsRu9DCtTMUoW+IzGtf52AaXPUk0YkHSn6rReBvYIlMlanhkysFmIR0dRbY9X7/aI3Wi
P4UEzxt4WKdVl0Aa5gWZmxhaBh4WReje4VrN526AwrgpFJ/53z8PLHOe0g6dq5HgVfNFrb8ScKy+
l930mcaF4BHfXOfCCCK0dG/x1aKh98cz3qyDJZvLn0z2+ovHkUveteErTNPk1G9AwBvoTdjsTUXh
fQ3WlagaK9HIIO92ki2u4AoyE7oO9GqUiGeyC2T97+1YIR6EU39E4cHHvKyIat2Ti/Hw2Swzahjn
305z/grfn1nchenssxuvzcRmvd7OuW4ZPR3CznQbaO2QAU+pqAB6fV/LEpg/LMCBqTu56qqBIEfM
1cH2t8Mx5en0FijqBDlBFXBnelYFfFiVRH7muceoSXDpm6MOjC3vdz9M53/RiyKKITfZcJkQT1dd
Nt2xJcRZBdt33d1sxegsIRpFAGXM2+kT8+IEu4E1fBt066Oubp4gFETjcnqVeEtgjR8yewtE7uZG
v1dJwEMCwjU39loIavap5OhmKRRJ0g4MjtusciHq59in1CWa15+PBzjAK84Xk0060xj6LTmpWBUW
TjusISPRaZr8xP8DsOB8LJmPDkuzOgAo04yUnCY6TIkZB8ic2KUQffMfDSkXm8Dasn+Ir9qYIo4x
5JSSOtCxtajxA5hz0KY7UFOjwgSBv88pOGcoHYNntSgbx/pj1qGvCtf1VSA8GHEcbIGlkBUjju1v
lYpjpTW9Aqr5jcSqUknUrNfHQ0KWIcT+l8SqVPbBs1lxfLDxnA1uhAg+haomCYoAQIv+fttK04JV
iA7eFUfoH28tS9eMC3fgCiNudIlJLpjW6rjKK/Ix6wZ1iOceiRqNqn0+0H4ZpQb4Kdcdv4EJuwHR
gar0/bLwpu3Iv79sssi4YElU0H/vRYvpvb6kyjAMRbT9V8lhyfKhs2i5+MBeWozx82dqo1vpbLhG
8TxJVAvtUH5O2hZkj3jpF+hR8MOirh1nTF/djtJ3+XG4QqIga1cLCi9yMKPk5uwRnB2OHriq2BDX
e7xGkJ6U8XFOwRq3HpWwCBDkT85YPEnhW5wPPmTyNNuEqAgbC6GnJFoLlJAMC6VEjOn07QKYeX2U
oVH3Kr/q9ovfzvZavCd632d6L+AWb5Gee0Qj6oh/bwvsdFo90pBnXMgAsUL4v/GDUwSYooEa9wzn
/dT1R27ENwQCPgpfV9EiOeZeiWOscJXH6AXWZNsBBBFSp+m57XrD2D+MnJZ6tNP/CTTmQbyDZfrC
Kf1elWvYHcbhQB8p+tVkpS2fE2oKhVGoClugDHE2p/Hdva2jKBR/K8AAtoJC6D1pSCYImvkKqkhy
Set0cS/ukuexQ+TXTKgwlczt8t0EKchujUrhUcv8kRooopTAlqYbKn/pySRgwQPxmvDv3WYu7qXY
Xpbe8KQatuPgTBGmUzv/FF8i+JkIkkIME1l0Z9CnPpRVauPRBVvsWJuhqAaOqCNNEGeYpNAEA5dT
SkAEEJfUT2bMtH6sZ7tiLiU9V/2GTQuwFSbqnd9d9mUVRTI91O2myn2R+nY/fV6cDV1eNig6MiQa
totmHXEEiByxSfuMzQzwBIkjk0B6f0n9YJN8As/fvU+j+nYGp8qWC22ejGgOHN3CNle8k1gUBhcx
yJ81uSrBVbEV9ffPBz+0RJ3DlRRdo9grQ48LZAgCcT601hs0NerNzcEGjODXenMNj8Rg7klFTY4r
FgzKDEfnbE6OKqG7F+NiKqulQbBWdHAiSRoWyLoW7UHaaiI/nWGll3c3Q6Gt0qIBjof0ggz5dG6m
HDD9pd8tJR4UqKX5Rx5UK00DwJpYqEAqxjvR3CdtutysZqPCt591+K40JLA1ltLXl82Vg0EMRvzn
MQCFefTqeke2b70b65TYYZfnfhy87ynfYr4tVU/Bfg9s1BypflfWmM7gbYwaFFF/k+0PmcVpxByN
SBHG7zqo+4dJcjVuqw8xejnZ4IeD/VeN3Cgh5myJrtN+5nV9PNiGW4TE/2cG/xAiFJ1o/jc7bekg
SLJekIwJ0WFuYVB4HvdIGEPCJpefadvcMERO5ng5mX38nmKRLFWQ4geJo9QS2BVxuAh42JPavk0y
9IkrBOztIw3P2sBY51WAf1x0GSKM6Mg4ZgWbSp1SEhZYiFiLOQmmtf3MAAQyTMulsFA9+Mm1dCUP
Ew1LcPjvccA5hc4Zqm/0+QA9IbpMi4geRd8wVweTkxL7ax7l2zxTL4pDtUA3LIqa5XtUw2ocSrbv
GCagpImVbJ6ySHwHjAlG005JZjJO7Ni5F1O2i0HnsGqbDzDafNUM+1EU6coALR6nxdGlegaSIwRS
tnf3LjJklt9jnbLSjAZkThiItlxUhvOUvF2HmPkdc0DdCKjnI6Y8Sr5Tayu2H2ZFVmly0vPrnKmG
DCvoAHvmLFrhlBg1Pmj+HmH6SKeD1dRwP0iq7jZ1RA+btPSjvZrelEThOIcfR4PMwpzhnbfKgTcy
0SG/b/BRI0I4ttASdtd+zVqLWpIToXdBak9FKDQzCTDEFuGMlgtTm5dm7jqMSwZRI5jukE9xtT/3
HQ9RS9J7R9jqrlLnCzgdnkdjGLbHqRzEqp9E+9WaUSJlql3ZtzK1IcTU8oQBR6PCuiRVZw1sqOGR
nR924r8ShzycJeeFXoUP3tZXvqLB6oELkSUikQ6dtFm1lykxz5OnGEnetDInJGVFkSruMjT+UV9o
kJCjDO0JEbxO11wOjOO2JNaaSEqAxru3uhnyADmRZCXvHa86wRv8lvJEtQExtVogALSS7NZV4WoW
nd5O1dXxQ6CrIyjVXl7AdFpqE2h/+hv2H4RZp2ttRLMTpEEG1EM6o3a5mLReMxQFWng+PeNUlGJe
0JVmt9on9D6XaNO337pT1i+FNposdX9hdO2UkE8tZ3VqcvCRso1lU2W1ZfnRoDibNdSAXyIMJ/4E
NoHcSQUw8lDeoXOHft77Q1tMQmCE2TwuyFjSX1HkJZCwg4r32xGjwyHmcAI/ifRslU+8siMpfqfY
pxJ4ssleBRnvcQenhxOPqJc/+a+eSp4axOmib9ZRkWBGnu9D1odhV4NsrLeNTcjXoIhTmsb/ZxYE
Uv9U0yF6UQETG8A/4ERP2SOlGTR+FDEBpJocIhHvLSvgNGxnrZfzbHdOJVItfxmB5INwt2838jYc
Kj4J8/7KsSR0Sh3BUpxA1SISrCHiEGvrRxNvvtFZXOaqJoxGQqiCtb0Z0BvBc9ARJK4eVT8BOVJb
m59OliD/Bns9CGeu2KemmvOkJ80Lphq561+UpxKPQAPlomO2OGghMjw9aVC4RHnblfps2SeyZP+G
LSBWbAgM8f6STIk1PmiCI/C3qRwK39xcps/GSF1AxuVpHGbIIJtUcQKPR9QxdPLBwSW7DQ+9Nhga
muzsEtw4KgU3jYPjAdEvmESwmszy99OswjX6OovTgCIg1B9XAh1XNtYcrQWSDsxWvfPWL/wNWKu3
TmdlcODU0AF4pMmbheyHkx8H+tjAveAM1KV9bepH2OCQxwyIXU+bqsqGCVvP0MWavE+YzHuMGXuC
BRZX9PIWWVDu8tPpbbDCdDKJqGg5/l6TjriiBUXxKLdIV033vom5XrvMXqZRcAcvtUbhdO1m//Kl
89ts704Lw1xHG+P7PyXuoCmt6/ojmb98nKarAvl5F78hlyoSUogeV5XcwN1z7ufx6Nzp+7vATd6V
sdLlLCFiyOWYgsjlaCtEuntaXJWATFACscX/GHcvv6DpzikLB+651dmS7/iXvSnQ6IW2pj7dI9Io
oOoLO8cjfv3BUKGn46q9LtnuaNdN8pBR+BmqO5WGjJnGkuqYBxKFLTxyryIvyfUmXOw5SS+8E0Bk
Ox8TpqIdEYIdXbS2YOjstUTD0MFxLRceT68914756TbT7R6mKvQBt5gq39xMRNL2bZRkyFQPvqu7
o0fvXzitDZX0/soVqBXhnnBksyMVJPnwNpWdw3E6wjFiMDiCMPIxiIQgYO1/qo6PwQeSQqZ7tr0B
if3mKMDCkXks14qCNFIK7vAWu/zSYmCo+Xjm8Ad0EOYY8tpcS/lUOEqgPznBlY4eZsTUFJs45MjR
VIV9rgLsT1gBpLrOaP9fe3f2gFfIZsuNJY3wD2NThkF+5lQ2hAFnYI1XI1htgOf1gnKTFSJga3mh
uc38vS0RSNXjKr6rxDg7VIF5kPEeGBatzlHEZ6uBW9yo0hIBuk9x/YLiJdCXOiUmlquSc+eqYqC7
62/ozRRJj9WDK9tEgz9K2e2PKMnZL6j4GgnVYMv0MfJORQuBTKYh4rZ+kKPedj9LK9PPN+Aj5ji8
rCAcVm6fu18WC9jaB0V7emSwe3EEHqu6g88uXkTLEv6jX0XoppkMPrR6Io6hBTOG51q7LMc7bu49
4dCdoYYp6shJ5xcGcX9/Gtcz29fT2epvaCVQQyGbU4l2dXKaapoiRZ8lF8p7w4FQCAa05kqD+C0J
SG8/74gpq5/WAwU4CZ8xcbECrkR13mWWyEIq8IEYTbp9LF7sF0Kzl4pJYX7dFcf8TBVpW49d/oX+
qv+ZtO1wU2D15fSLzXf9jLUY698PgUFgXvL4dG8q+eUXPuka2ZLyLxMKoHA9T88Is0gMOkSo7V48
US8+74rp2DCXnTAVlf0Zk3CgMUiQnPvawpp+orXd/eskSICK/7Y/TdNiujb22upY1uZNMMycVwgX
1A5jq2w4/XtU/R97o9gKQDn03lT0k8vEpggOKDUQIFOuSNqQYgYdtKUyGJnTMHA56LOnetI3Suv6
qiT2bwtU7LstqKllgGYJqodkB0aFRWQkfM/vQOkwnqPKmAOTIN3gl3UmmqRJQk3sw5CqIv1XS4BK
XP2CVLBgwKUdMZB31CUvazFYHEgKg7eU4wPmE0LhHHnb5zODjRV4ddvoLBf9p/XOd8q4Tor3ppUM
ThV9beT/EcoOq51wuTTwibPN2u1Y4FV4TOiNjN666rzZOxOlkmvKhQP87BPpc8y9iZnDbFmb3U41
OzzoBZl2WokaQFWJvQNThXxR5Bhi0aOQq0rEcAngBw9XesGUPO/V7QwYyZl1gMfV/kwZWqvc+bKw
ByMY0JJzqGWkgjonnqpSxHepAdwA2Squc3z4VeHcxYhjP3savtY/8lcrDHXFF6ylNo9qAk4lAd8f
lUKJXZi6W+Locj41JhTNS9CNsA2cO8jUzERgaTF81q8dQofKEi7Y/Vr5uvDgjdAosGpu7xdXOg/T
oB5XGV7qz/pFR7cbImqLOBO2mVaDB/NlM22wHGQkdv4Hq/VxSlXsbec4odwAFUmjrg3dSWpaEgvG
R0d0aC/l7t+cFt4kNfdapETw998+wrAg8gv+4ZSBoizESCY7qQYhmgCknxkaFH0DfR99mptVxzw3
rT8pW7Nhu3E3PdLTJXpkoddG+YkUP1SO7oqCM5kwTsvzRq6gbqb35M0YtSz1gDOZfN1NdwI43wPz
MltR70C/L9v0VSWF4wC7bYr7aSAS9k5bSrVIpU2T1JF62HCWuOgqWcn2OENMr3VLygMxlsmgFLXX
RStyaQdgN6plZtFs//ERjaoE/oHJpi3uwvUFEgEKlCJIuC4sSGiyYNzHPF3fUCswApbNjjbNe0sN
9pt/c1q9oP/jDIulVPn1MdgWPir2ntVKTC/IIXSMoInFmZFVzmJtl5LW+sRZ4NQ1/3PPNoykXBQN
GksEBwzRVk6dfnoc4gC+AgKK1B6qJGQgOCpYgpHPzB8hzUvvYsTOB8d5cYeb4pAqINIQDpFjoKtK
2a/WG4qFtsEAUZ8dHvS2KRFg2DV56NCIKYmzc9bCHHq0uqR2qWWJdsbejO23MM+KT0goS02H/X2E
QoIBIv9dCoqFM4yczJve5qlTaURG+HtfSe/hkBD+6EwV4+neCtjUAFDVhuNr0Culg2cux5u2Gm0v
3ZImRn2ySzxo4rEwgaFNhMxOJclusJDNlx/b6Q0zM1OQEEVSzWEDAexbh8fHYvUKzlpGBku7pycP
eNse3FW4UONskHkb+rkxyVoaHoQqZy4tWCNYAvKtvSgZq3935myTF/jMi07CesltY/VDVxMj+CE8
eOUudHSzk3uhuVO4OFzkhZXdGCcgUhOodR1E5GgPeHEBKVQTs8czb0cMdCZCr1wNC0l+LDt17V5h
6VRyN2r9SGJxIguJS48BWxdtpjyEXORpN9VZADTOqwPdn8X/B7k6DnOQZVa/aAOG41uQyd30fG40
PBL0moKwmXJL0qiG0KOREDhmA4dZsua9Iy3OtBk0DFChmTvm16AQNygBr0zigHGmTJH6h53wUYMj
F81lVoRTXPf34rEkYFvZvgY2gYinp17z+ZsYoqsDBKcTlgafqotq2zKz/V0gplq2/kYAIJAzsEiq
1Ll7bS4PoEVWt7zEfIEjrMOcIooviq4BJ5G4DzC8INbq+qQNxAj0BGgpbLbADyPY2w60etCJo5oq
tQCf0T/MCCE8y2e8fKdFMMtMc8UmWnGNPQKD3Oz80TYXe+0/cjor/NlaEySaIsTUIzb9fys3pAvk
HgMuSYAzxtnosqPcxrGDL15EtR8pFhz/RLkDEMe8eElxeH88URNHlq3RbOuaMwAA9zdY8eMdPpwI
vePNwLjDWi5vp8Mz9yBFV6KirEzDtLOSdIw1E/KCed7CTjoZVjZ0LgalNfDlZVJbs7sEoy3nEHFy
Tbw5ZoCvsWQXQC8sS0O83UhQQRzJfADIMYJuwSA7D6ArEH5dmyAo8OIzVe4wYJeFx7f1XbzZgiNE
D+wJB1pL9p+bk6hOLm80UK0xtgnVncwHR3kE/eXR/725tnj6FBwgDqs8SVurJKfmgRAg51lWpY56
mdnrsNJ0sojLmd1rmDGOgP44O+Ls3wB18WrxgeS3ziEy6D8ovyYqkBAfrbRHBisy8pQtcWPVOUC1
8Rs3AEGEYNTAHXq9zE8egJIZT1ACaawevBzGctsfieDsbrxiynPDu2NgCqB5IADXd22hV+vdMlN1
5mkjwOyvAZMH8x6EElHr36UiEwIPdJbNynikEHEr/MesXschHp/Fp6d791drDFh7mZoahu1zcYyq
b9id23Y6SRNQOf5me+2/oFKF+RTMSgbEDehD4Z3z6L9eR9IbR1N9tqwN9esWv8umxlggwmQM+5hH
2KESO2iYzNuQxPmg5ioedCg7BZDuIZu649fFJvFwx+twoyn/m5b+hw+7nMMCaCjSnQS3iR9fgmcR
VyVKLKEeo6o3vCeC5dlm57PCLSoPc90U/k+Z1vo/Z0r29KKMUd4LLdC9Vxhns2DJjUcHNlSpeknK
WOi3V9/sXXbIrT27W/SZMaXfcZfwozGCklRNoHgmSSWAampki4JaRQIJqytWW5KK3R34C4MEzwGL
LfDWRsPeI4RQA9BpWoa6RA7iDe04g64QDZlUIqWWwOy1yvjWaPxN26WAb1FHm1UMzzPjT+MkHk8L
Zrj7CcZCT076KplZXFxZwd/02UY2Kka8uXLfmIOJhmQrw+XWGQOOM0KhTzGbRTg4kmiVQEioXAzN
zl5h5M1MIkA5ur5mDe/kJp0JywDuQ5Eqo83gVMm/gxC5rg4Q0moQIqYyLVHtvAdeuyay9CQvqQ/D
ZlpcBlJFXYrL0V+7mnoz0Wl4OVz4PgpLumNZ24nzoSzV6hZmWZZOYQD1NkLyS9eyT3B6UGaQAlNX
a/FkmIsSCrA1/VOLZ5ZjA0v+Zhg7owJKePdjz1TB3kQAfSr8a+IoNRZFSWvj+PKjP7tyKiDj4m0o
sYWqoeFXC6vChpsEwhIGseKXqSkFmiwx6p+SEYpb6cXEvz2yg721Kd7fIfWmPK4gBqTeQNSOUtXO
hH9P4vy+8cbel9/kehotpACWtxduvy4IfZ94X05oKNZylfTkLna+R2Pgp+zsU5J+ltTIP8fk851E
RuZyBLB51AMRSfUZWukeh6m/rkIKlcHs5kzf9vEiNCImhvM4J67MEP7BgP4AfCYmHk3wM00VEiwZ
SyfjecKbO5bs4X4I6HDdbdO8MSmoX6mGcj4AmHtF+Ja/3DfVSCHGm/089pxJ/l13+40eUfQkVs14
yPhhwd3DAY9QpcciTzX0gcVMpeh/8b1WMIbUqp/XrZusrMi2Cy5QQ0MpwKxX/eRmXDWKD0ow9Lww
xjZn3woitWJN/+GucH5FsZ8wVoqvAAbA3OP5VvG9NWLq1rpDyOgoPZdnayCcBnaLTMvy9O2UUqJT
5ZGUEW+XxqcehKcpus+bEWNQzI1upR0Z9tSbrsQx+n1KBclwwY1y9QufsltwmoJ+bYCD+a8yTGHv
2zutgqVpqeLZ+c8FGkWLQUugmvm4R1u+04RojZ72BvECaVhop2kazhkFwvw5CH9Tne/WzVwG30mK
oqPe6Z2ra7If9j2HeZXrPIL26s6p616aGUU79dy9ojxTStIFp1rJPvXF5dfzKnBVNgUb6bcxQCOr
GzZzMXRlSqVp9lv2WDcBdwFwnJrn9mdN37jqBFcwrQt8REt+WWbM3AKRt+Qw3kO9ejIlo0CuWVWf
IFb2LgegcjkuAHMOgY0U4HjNfsmQF5l9irNhCINUoqyueqfpYZHzy6XY6OZSB7WWksTuNYA1J2PQ
bWFMSkS/aZtK/T4RBdGmrNh3J8Rrd74Tr9XyQiYkft9cTtmQml0GKfbrfvdulIKnZ2sLzHfir4JQ
vhrUr2O+r17/CVbcslwSVbvaarLrA4g7mA3k6OMsbobjDLhOZR3eLL0vEE/vYS6Qho9+htVuhd6Y
dB3PQcK4Rz9xmlBGKenGi9IcWSu1LdIs/TVcR9JdqsBrd9SAN6ymgdN2212WkHC4YxWGJKdbSOAD
6rw8aSXWUMISFMr3co41mZ63e24M64VYyGOiBnfKxAv0w5R/F4U4v5aGGSLjZK1ZKm69zb8Wmdwd
8O+GLTZmOhyAMwjWUPYL9oKvCw/BW3PBwIiZTErbw+LhKbOLL4ZuLJ9YroThtOKFNBf+6UqgBCAm
/bmUS6lznJyHBoWRLdrM+6ydKHynLp/zlS7b0ntPm1disoeAO5W4ihKAwx7Ir1myNut8XW5Ti9L3
P9PJBxTKDlvoyzvEZoJF8yIZELLyIrro7wD5Vb84TW/3SDyRQU9X+3zrecOiUfB30ib5n43Oqy89
aIBbk3a5YduwvctPZTHitdIWibpoyrBcJrA3zbWpf/00tfKP0uyeczFehnJfgvS6wPV+qnvZQJQI
Xa8W7/CuzEowzrp6rhCkMiBaqNRI/OYtxicPhHzStDpTMkWXUVx5KWbjjiuJRa/iXZvSuhcwJl4r
Huxq/WrgdxURLOHVy8zDbpCVZOu5Z3QmYzeTbokb0gyynV1ZAGw33m2qFK1cYCRnUbvp2VLmRhH4
k7wxylD+Cg9T6pVYPXYO8znFpYx8wnNoViYRGoaPn8dUAEv5ofRgiB4higJWWKFw31fovq3cVytb
pwQ2Hzs+92EaLsqsLw87+txutF9yfe6rYYvAahBx5J6NNCGJQpLA/RyGLeHTvldZf8FGpiD0HquZ
APh3Pg199ReMBBiJM28uRpQI+pOl5DpTuG9Yg9WJ18soKuInEbaOoLlY/Z3LruOc6IsFCJiseP6b
lh7hNJFI9t4D+fSOideJtyP91WnGkgADNHqgkTauU8unkHlgS9hfsY8MDpQD5VUqjmgTfxvZ72YY
aTfbukMc39iNTkJaSBDqoEfwK0OpFLD4YV/y1Oinmtch27FKyM4k1E//UbaOQQxbSJUj4B377j2W
bAS2yGPW6FqzKPtni7DZ49zEBBjwgzUJbD1Y1pw0nqSEVdLFe+Nc8DuJfW2QIR1Iy3xL1wzOnh/t
BgAVJDWJ44QSlOvnefhNH13xkzvh4R4R6iWoOdTrEIkSa/+HJgb0wFmEOPxyVhzglg1qh+mQRxNc
cBgSJ4zaXU3wvscGsFh9j+Y4rQt+0m9/JnBdCR/t0DDG/sWphplxku2kvdOe7eR2GG/5OBKSTGYr
RvFpwAp+gt+0vYglVeMxdTeMMSR9XuknFg9j1GwYDMtxmXXQAKOk3sYSvb8zX+SVwG0CiouVScY+
SXKTBjmd8FMAeWHqyxhO9Dg/8laqx0QEOIcZV1Is/lQZniG41uH8w4iEENPZjt1uvZizdOYREWjY
GUxiJuSFW7BqvuhOdBXLk9trKDKAKSGcAhPvyWhv3/va6qQl5OnqS/gHZSIxvhZP4kjTPnC2aI96
MxVTvfY4OCEnD6Dtchc1ebiyUXPfIId32a60xHBXi1Jz/y1hfDH4dMSq02hxcXbYsaA9jOkWNuki
orS2czFQ1pxpMLUp+ecsOTEj1miv/J81i9xpQgsxTYioCv7pH1WoHYd4QcT4JthFi/VrqUT9gh7u
lE/70KpnbfUGhsCySxfYmKIJyfQ7eP/X2Ev0vrlJVhXPUPgXSC2huj7tgJmiFz2AT5Phnxfi6OFW
plxYwaGmlFg2/YDLr+vANmWgeSoAe6o0Q7utEyRAdQE/ViwAh/XDiLQ6LQDsMb2iXX3qQKrsh7mW
hsZbZoYpxMdUh0CDnUQgo/q0f1DqS+3+/RWrUv6IfTYonbpTfQKs+F4uuqKejGjAc954AA2EmZT1
K/EOrL8/ouGF7EqadNqp0+8jonhyajd5U6OLRotlioYDdIBlqtvXDVL5bYowMO5e4A22+N+yop3U
L6jd9XSEPNXm6A9BV+eH9OUMaC5eSWd1kRLunlcm0S3RJAgT52/ZiIozbGdrab4H7xyQ8PQkaiOD
Pvcz3h7suEe7NnfptDnpueqTNyseGgS/eREeeE206rsgBpeimpiEylokV9RZY3C/W7FokBGlY4uQ
xzgtqyuHVy5Lr5PbBBE6MXc/LxFxA0xioUR8iUtF5n2etnwiYvzxc7LQmInZ76682FXXd8N/kEyF
tlqJneCr3LnNy+/ODnqm0iybZ4KDlftPdR9OAllFXTQkfJRZln7hPd3HmGGb2slBU7FzvH6tRNs/
HT9Tvpr7tWgeugKf8Wo1Gs+ebxSktMVBxlU6u7lFrftZ0yZYWYBJ7skj+Jz/sPy2h8ZTkRuK9FLL
NsojY/XQ9fwRHyzDHnA4Hq5Z13w7l/ndL2OTuuP2U66oQ6yJtBaVWx10eogfFHH1OGok2qt5ezJJ
2n+u/FCeXQ738K0DpUjKBdsM7N1L4NZ9C32CqUAZXwVQg2brBgTQFcdgJA+DDcaPwbX0r4nzpx9Y
F4ztuAx2XlLbm57kRwwZqlzKX4DOLNlO6ib0FeQIdB95k1/m7EuZg1j7A1N1+NZTIyNcLl7ZNwaM
e27+l4dzlRUO+OwfchboyCyvGEV7vOXWJ8fetgHzQP7b+Dw3b65FWKqipXMNW35MBM/bcpoB3yaa
F2PeDZEk5G7qPgGMUobdRe5gUy5Y5Q1g1t+jP36a+EEHr0paJEtmv40ELd9PT4vN3WQuZZ6N2dGl
4sOxnzHNimyW12oF0Tg1ci6wJyGcL/KrTKPaG0+Buvh50hJfV5zuPNg9jaFKLQtFeIXipscIbDdB
Ajp/Ctry3pxqoNOPUEKKpM7TXwTMLO14EsOJA3YQhEMCESLBk3cYNrqa2Yie2wHhEoYSpaeIwnBh
c7ldH9SArWFujRjqPh01FkYwA58vIiVpBatgbcQYcLyrgkn3drTWBe6x9F+/LKj+x1m64RlCEtQH
MWAq1xKXon05BzFaPlyKvP6/go+jGLmfwMUmFpoPCQWYlGZUBV66pixDGGzoAMEOMDBIRP1HYK1f
xOs5rup/jR5AuYQjYN6ejc+bFA09ETfhB8/E3KDsM7kRlVqG0jKWb00rJFf6+QNCn2YTxG49naZ8
k7u//87VZxQRBlb1OqprES92W0cXZX/bxAw2OhYHgHA7Rrivj5NcdzNE00gbggZ/qoe6vmMH5G9o
i7Tz5ctjdMUKaTCQ1x1QCCjJaGQeGD+nuOeL6Ehzju9dNwpY8f7q+WXKLYcJTUzFrKaOfhL6CyOa
jvCTPXXlcjoR7VZCl8U/Te68jVNyfzgeuHFKdgjCiSvkNozA5gxmClsnyMG++zqfVmfrBHjUIBEO
6pcuFsAXpHJqvcZOXp8+zZ9J6RHQO884kZCORlmysp57iHWHS771DV9gI8O3wgNrrjjZO5a0Qs3M
Gywyk2J66I+wna7xVqFr2HmRIcZVDghhwd05oC4MCdhi/kf/QI7ObkX5VQUtTB/plsHbgZoAwlHx
kJ1F61Nv3vAvmAsGyA95jc/gH0l/dq8C1UgZHrcQEkZ1Zw/WI2jkiYTV0iYnXd0kW+4hEVvknw3z
pP080TXJJJQWUzcp2csgrvhD36CK8axfDnAULr6NVPLjftMFL7B+4TUckVLUvbIBrz1yFmZOhYQY
g9DxTzACzXlI/5Q8qq8EdGzuNULdqQXvSMCdrfOb/UsRv+ozhaGdFxbQPT9p30qnF3gVHfLMjjzJ
UiynwaRa+XzxUSqq6rgs2HxF1OW0WDmHBQ9+sBv92kiATlFE06UMk9I0ZPBHxgwxuZEKiVK49N4t
fqlLvnaZ3yUHY3aNbmLEIdY0ysyB54l4pu8ypDF4yHs0UB8/Menw1vW3J032j0ws8pWDYrUkaH9V
70qYFow8eQ5lC8na/D1tJO+2p2526HbrzQmFZbUGfaNW9KikTEHW+2fmUo4q3ZO7nxDXAB34qevi
OaM4tG84cf9BtAjfBWiMNY7n0kkRCwLDW3cCDkvNwIoLREju5jOnHzbVMW94k7qcnglV6OtGvXq9
tZfwXLWgu/LLtCb1owtBckW1ADZ+OPH+VrViVvDnpvTfr1R7u1ob3sq+I8n8+VsVcw36kxjY1U1N
DV6c/thX3lBikHsz/x/EBRStu6sE7Zjy3Uaw0t2s/5p3jLa/ttIDrUpH4ICAFCwwawemMdXBRu4e
EKq7xcUwI1xhB9CskZNNuVNGwD3H2w/QyWOK19IO1ze6BZB+geo1u7Ev0YQK9FhEQGMCgWVqteOj
/aI3wYb05VdV4mVBqhOSuFNO14o7541Rk/CNM6gevGr0tbrOYtkVGWdUGbGSXagojuRoWLlCYL+G
9TL3HuWZI0QhyWSitycuQWSSb3JPaknAK/iysWWOFIprbg2qjdHZfby9tJ34/YNWSfQcjz1Njbdx
ZdanIXciUAfzjJ+O3VPzf9GEx9n1BlzrzvanY/5GUKpcqaIBeM9g9om6tEuqd8TaBE7Rq+SngB39
YInhBRuPrVNgY830oAnpdmnDS3/zWtPixVUW3lA2+MayiwVMMZOAcbkK+axn0gy7SAW9M6cM1Jcf
5xzMyxznD/lDK3V9yb2iSIPSjH2iqMA1xIP8Mi/tVDjERTSf2oB17iQ6GZ+sBtmspBs/cSzetbk9
gz5RYaUA6CnYdv62JOwbwbPFYwpwRetsGGjwRHv/hJ+QO9g1ADr338proUCUU+8mBsu380/oYqmK
E1B+u52wepNrRtV4a/Lc3zqlEz9CfoMU8Ew3uLT+VYLhPEtDLZl6DB0mfXsKG5oRd9sgL/Qh9+z3
PepZQ5ZBaGFGYhluPmI7nHTpg4rfaQOmfvP1Jzm0hJkia2uNwnoEFMZpORsQmhtAAvkd/vLSMMWf
WNunE2SEQvLmqx8dvuYxs3UBbZVBBEvHGLwZnvUIQvWhjhk+bSZw3j1ZhYbzflwoc1oMiHDsB9t1
NP0jSqo0Q7rfiV1jgKn9giHOMB0ZGrdij/8fVND2lofiktdjLGsc3X0DuA/+n1cKf2fKRF0a5OEV
diDy5fitgBD3SwPe4z+KFgOXn8gtZNtUxy/G8pA4kZivqJuon+YqAVqifmefPKpwzjMUA3VT5uzR
yyGwLiLGuGU5/pSKkzFJNvyVL6DBrWdbtntTMvKjoXQysJqKhOhmDK3xZj1ZXfwTdJZsF5DmUg7M
yE2b2dQQlJ/QUpCLwRY+bwXWQ//zWlwA2f3rIhrjK4heNUt1REB7eovh8w9Md5k+NKIz1vy3eQ7H
C4bOMAlAr1ORgrW7YgxuOSRcBkKDM+3lam72fR1dqrIWErhT28v7qJ8fZumqkUSyWUpDZAO0gji7
2FNQ7nzFoHB+zsaoSp0r7FGVBZXA/V8enc2Q9TZaLDKRS1PLPS78kVFb7a+9njqw4gzuljK8JHNA
MIR7m1OkRY8cT9ZAwAf/zsU8ICR0lhYd79z0I+bygo+nqD55XR9ez6JzBmGbFEJzYkOKxwQWKOem
vEi5fu1a+c8sxF5ceRTOcNCLcaDSDDkOLUfRSiJezsjqtMWpYSzfPm7gAQN4gXji3g2v0B49GCfy
WDLEtz6zRWNW5uNhXx0JzL4fX5m69i+Ogv4ziLAAZ+mr2aL7B1FE0wFRONMnvf3agmrIFAYFUYWU
vOIl8PaXNesCYN5LjZr7/epuOjVCPYm5x4nsWFiCWb2ODD7rAIcYMFjmF0GqfBAAuyZXkmhyJdG9
JOFpxasDqe7JFw1tDHuLSk0uMF9RnIp09ojnzRlJzyttwGUiqyseWMN9vTVzovt9RT8SJIFlDyVf
ndPteFdgH7uKh1H4vmWotgjx/U9fAOwmIl1Ua5DCyy2cM4d4TTsTwYtZBULv+ax4msBSkx8h3zyk
AycCo1kS6EJOQKUMm7HhUFesVCMkOyUJF4SNiehSKCGF7Duhasfe/L9xisZFQLR+wLshR0FaFyOT
qyfAN82z5N3k1MhJucuZyBxemw2NT9XuVu3Enuuw1mEjA6qKDTP4t/CfrAQRpl40G1nEOO9liOFw
BVPUeMOy8OK6NPVd32eE/psbkhGZ7fgBGRUm2MySvJbV8wxLJjt8bE+EsfBdALtp1jc5re2YqU5v
EM2a4pR1OCmZgH41aESRavpaXhs1pRWDIizyKycb3QkgnIiPAmcF9HW/NY/HFh7fI7lkQFnbKnYD
wQSJzG/2FYjNfHLNebEGqQlcAFYbcoZXgAYjaJL38ftLLxVxL0Rnaz5wecd1WzaDjj9ElCNsf1LW
ykZs7jpSbx5fOxXXxKPvaLeFS1dx60os87fLYhAeKR0uVKu1JbPuQtNK7tfHyZPDSsaAwPEAy9Ct
iiZSX3COrC5giXEuzr6EZl3hxM810FL0OW9LOF179Uf3yXziHr3rz7qrZXZXYD8HQjXD+V+auo1z
Wd/83uE0J02FDGeZWQK+hu6jkFycA/S1TKhs5y2ILJfGCBAZKxdnQltCvl113Yf9avx5q68pn8l7
pVT/N07XeAdStZ/9tNfzdyIgts4CgfHBlZrKmhYW2bVkmZoxR9EcjscCq8ZKIjhrfyKG72c8FkLi
mpkWuC28L7Lm4yeIMslb3oQSmY2YVliT1c1pCCZzYR0z3axtTq7SGl2Mq9PWD/bQcLbLA5neHz4E
IV2Whterebe+KaDR3ZBg/CpjIM3pMfVsOWRv28jwzGgq2ZNWfjos8re7jXrMcxGl4iatqEVabGJp
xbBgjl5fhdjwaAFfL+PjKl2UpMFqq19n/+vmTxPm8z7V4MF2OdXA8hDnrSybvVemcnVBTRVYabso
1DHFLfH5cs0eBu/9HK3rl7QkOZlrl18kE5hUOrdMaCm5DECVXZDcad8cBzi5P7eathOEyj5q4H+N
zxzkb15hfoC2wlGXAjj4ppxTNZImX3Hc82iptML0RPiQU5YwBINTQ5BJceT3fklgxDTKiGJU98TO
kpNVljZMwXhsDsDGBKu0ZIyPmU7jwtI4kAaQ2Uw3manCLJgEuCkoIgk6XtNAkzCikBcdIBAoCvw+
BvomfDU1Di+iK5ZKHWbVzX7CnOll90URuiTPVLuXvgRQjDG+SBlmQt7aBgminDkqVT68XloNPV6v
yxFjFI9jvuZN3CpFmx18udHB/hVW6spDwx9TS1YxidQ8dQ2Q9F4RtywH0/FysM1h0+EevN43oo2k
FgJRnIkZzCQl0stYOOTXORycphLmAumaWOdLywXrdizdwgxrnjmEldxTgdTHmUrQIS5cYzY9U6Ey
MdN8qKkpLwe040UjdmacxkuMjDICOkb4VUjhtpVjRkF1Ejojy/As8gX2kNwMnhPSfyNq9eXdb779
TqbMCegoehoKCApXAlfe7zgtecV00cMP76ymAjnFwfK+I6yFaUdEqvF2iuhu9ssix8ppzea7fweN
ynrSr00zAOv2Sj54nXWubOD9S2o+MsRiLos5OOyaBA3AeLWehCpv4InAl7eGKmnAVKTtgPjQTkeK
ifjronzBaATPjHNrjIRl+RBBrQwDGE5jwH8tPvz0G4gAoFnOLERN3GwHdvRAsNp/iJ1Lpm/d5hU0
XRz0zyDK403ErTf3mG2Rsp6tzrFyJfly4JMMp+fZf/OHDjLZ/PB5c7+9ZlyRR/RW2yY2rGJTwrC9
sz+N41y1tX60uzX0uX+9KQBATKhPtRVs5utnabhtUDUMP2omH5wPYJ2IUFVamI3vwpBUn73OMns9
lW4IIKESWpUHLZ7vJNzc2RBL16LasIiydrSX/ZZ/BOXxCB3WGQ2dnOHPdZYbOCk1qe9oFuGlRdeX
twyTe9d2pWctvkTsVqgx/uSlO2ZcvCqZHVmDKyFwHsxdNUC1tAQJIfUMW+aDWwvLuUN09MPepkxt
l1YTYdXuI+I4HiS2p06gjJSEzdAJKBGZ+7jG3JDFcQyZA6AOOjDB0MYLuBVZl4FkA+sfXUZfDbEC
w9rDjIvRAG5swUb0jGGJU/B8FKs4l91Lx8q6iPXuw/rWkFfRW/GxgvrEJy5vVaiE8eg1GjeNvN9c
dQzS4IkmM8Pek1A5psaI07ePeVzAI3Ga5t7Zfj2KxS74ygMeuqFkvRF6XXI0NpyLgS+SdgQxWW1s
Lf79clWeM+3SfI5QoWlXTbntGaH3eJFqCGZZvWuDS/KDKcOqKlHro7cFhSLI1+GJG0dybqhExEHz
AGDY/aHVWYeNyJNcJ22PUGPl9P9NYJCIxmfiKm05PQBMBzzESY/EntjflTOYL2czm1o3e9BgeBng
j2Wy+z791uf8WOJVYn5Ok/ih6Wcjza4AmCTP1ekMHtDScAVLIzjhES9fZRZW3eXiuADkM9B17Jrl
31q2JTVUFvX9I2/83HXV9a4L5CjMFjD8oxDlDRQku04GfVvIq7yRSKiCvxPXZth6VS85bHGT8r7s
Kr/o1gu4vl/fIANI2lu3yTE9vkfYkrJ9mX3XxB4bjF/QR8drm0EqEbFLCQR9Zhwk08QaiU3x36gs
S8FjaQqi1z7avyf0lDrzOktBK0nIcMqmd3qpEjvdGvB0TEr/QI9EFfBvGKpkx3dS1em1kd6ZMuDH
OJR9obcIaqW/2W0P8wEPnpRhR+QoHlkTZMIdQ660Fw0P/sS2NnEzF2WhyMV+DGGJITli+DJ9Rx4F
/kkVtsxceHwlZoUXuNrOc5Ta+4BzBNJzhquWfsPTQMN7hJRzIriuRFTDDFYJc5oEJTQOQP9WB+jN
ElftLv7B7EpJo1Yc26K7dwBWRpo5a4wjw8Wxz3u+wI0cAnT36GXEydZ20TZXX1UsDFQ9O/4fqCPy
rhTfjOv5uaHRPTsWfPkY82yICveuFiG7s1OuHXiKT/wGZg3t08ZBNc66BZijvnutRqLNdRkIYOx7
GTl5kLKAM9Rgi3CXLPkRrZqvfG4p16MROhGhrywCFINnOlSuGwQ2rxeoW1Q4qK3iI8sP+CRC494W
bIxo8AFUv/nTINTaIQL/r9Quss4jAMDPkLDUewCAkQ3G/xoY2RmjmgwG4lesUjP6tS/UhK/5YcSe
P3g9x6VxNsKyUqFOlxW3gcXoNYsBaIOCqGadNLC2SvjZMLNGMrKULi2oxfnZqJVSP4ierc9cr86u
pM7G6YSZne14rv0sQHGUTFkt/X1wSiKH90jN/CckJ54Th5dL1maMTMie7W5X4VhyYh3EYbI5W3O/
P/Slw12WxdI7AhUnuvVQVwv9BFvpEsNrkBZCj9KI1PgQrUbjn/57hwKc6H74o0PihmlqnD46anAz
JWA81CMCRVLF0NnhwT6gMYVe/YsM+if3rbQPVJqkfl0eO31mG+/YEtR7x95cCkbdaCCu7Q3jYZ2r
xRsvOiTrB84w12Y/ErZdVIkf7bSNioRVKylRwmAJLRyDC9RB72pB9ncQiMZOn3Y1ZU5uo2o5Nphw
u3cBmVrivlo/EtwM+u5R1+bFpEUDG4bMiLCzCCJ0cqm1hIGKJu6WDnbl0SQq7mZt5ENR7lpT8doV
cYwoVZaYAOD/DQla8T1E3YPDSnHBuoSfX2N4R2ai45WnROQrfRIwl6qZXGpbuGcAZmIGF2D6dCig
wmarDEky+KMQb6FG1fZOp5bklgYxltChG2Fo3F0qeIUnRDdPabfdSlk0J/EenC8wqQa5l4wN3XFs
ukk2VDjIQtPiK8JY6/QE9aTYCkWmFB9MMbBIPqx9xzlbn4N9erh57dC7zXN3SZtn4o7fgGYtA/w3
WMD8nDueLcN+WKi/XES4u7mckOhNSTGVm9XpKjDMDdYJA8p7KVU6MZLSzV7zpi//z0VjahyzXjSc
Fgp39HEeffOi2lq8ABcMyAC7F3njhQH4j+vcx+ICtE6iV0qrP9C8rGMZtBfjdOcj7bdWX0DSu+Ia
qhzD8uFFsG6sYF8ua894trIZuobLzAbRfva7FsSu6tP43brJPhWfObojgK34iNvWv9qWXIBlt2dw
B+0OkmiXCjaJhNZnkryYW86XbcPKgh7XEeH/S6rwtZVD2+uImkjHiHCz1d1bGBPze0E5aSy41sT0
7t3ylYgeWzoGaDX8LANwCWxpi037nBVNg0MA4zRWzPZQ2qZ0Z5cFCcXPWucb6iYq6KY6r8EZGt20
EeNdY/i2lDNokbta8IthpHhdQ4m62j4Wf31oPGod4h1U6Qwxym6RKEsNo6HH7DdGGM2+aZGTOdEs
vKKy80yssinIkXESTNj8iLILc2j156m9evT0OpmCT77y/6wQ878tuCj4Vwkcrf5DJ4P5ys7b5Hyw
l06OJ8OwIVpaRc2DPsAtf9vH8oMYz1oiFa3IGiEvF78iis9yGCTGP/+Hj3RbWJb//8J4lt/SI/ir
tkVvDCcg3xBBMZ7pq5WcbCwhH0NluqoKlBUZRYJ6OtXNclSGZzyu6z2NdUMoPjnDPtJNZ17Q7Md2
OIFh1MlJmfU5kGl1DCWFaAPeiIZqSSEm9pDHgrWmzi/Az8ql+O4+oRq24TN2TabzrFE1GLq6PXAt
SkaWckB6PJYyaNCqPWnNO8tctThVCpQxIhGNk2OnKNjdGuc2V2Y8qaLcSC6uYJJA4InhigOMf0KO
05ZLTtvHTfx6jDgRvfaO9K3AzCjGhTf5junHEctMQWXDUHDv+9wSSefrQh8t7ypxqwg/QeE+1YtH
stlIb97wXvEc3zK1bjbwZ64JVbzc07dhP4F/4WqYbv0i/jau3eqtSVbvfYh6CNL4UIPxZcUsV1Sw
xD3b/CbmTRmeNvMCjlxQrJKV7q4BsihSByPnsnWGN2BkPCAT4PP9VczSIpUGjs2Yy7ip+fdCuFvB
pUkEJKL4a5gOxAtYP2EUzJewYq8WgLYdOE1YU4SFdyLd9R6+YDrquhsAMeOs7IsvAA7+zTXxt5z1
KQqBy4cFe4d3A/kG8XWAOTHLP1D8BD34PrA/BD+1QCXICqR0TSSGVBtjlIs7Zp69n4Q+aP5RtznX
313/Tg13VRkQY/K2zQgde9Et9xz1yDHjtwqBptpG827BopS4J/8vWxahgvsVy6KDwhn9tgFIqRXP
cPRso/IgsHN50eCMJwWIJcm0aRUA+X3V7JUgTZ6UdN8bUtdEN92SshplNmBebvvj7sbGIstA0K7k
IXUA0f5BkrZXuXG87bq5312q/5K9Ap6duOYvnLixRc2GKRth3zClKSG7jcXTSh/DlfIau4K43XXT
LZCsGzHMldIl6fa3B+UniiDwPa5Hs0JcMaHdHvSUcpg44y7RQv33kz64d9tmPYx5dpQMpJ0MkdEX
1yGkV1Vt6rb615/whNwxnAYqTPixBZc9xnssqCeKsaThJBwlu0P8ufQofzYNIqrHiXw2YE/Gnfjr
+nXWU5DbszzCY+iOrZ6eBae2pNrSfFv8aE27Ek2MRsrenQdSUlQjyJDRqc3QtdNbG5JJ5M3CUfIS
391RrAeXsvcCzv2CxOUiNOmIo8BQOYgr8f525S/iEeT229MdQxrky/d36r/HS5d9OdAHrv0HFpFq
9Yl5JDUUws9XergKOoDAn4a70e5BZ9cfDXwAfPKJuwvf3wbfkKDgAugHZTdOkXYbyCcoDCgNzz8M
Jkuz4Uh7vcO6k8nacEfZM2n5zCITu3C7WWtpEbeRulPFW5/zl1L+Uvnh2houPfQX7N7fercUTJcY
Bgj3OSTUoZcUUlcG+BIZ90KUgGOUiTBy5jP6Exx122QJWoBrPafqpdYRCUxfpr0NF6GA4I6ysFff
vU2nm6L/XESO4alA2tEk4YVnNKjFWfAqxb03rck34Sv3PM9ws1wwloDpjrdNvK6s31a//lAC1Dkr
oH2TW0PPkchCNEyxPeKNOdimSTZ5fb1fXiazOqrsgtIi4vepyZRv5KeU3Wgden3zzCdHGXQInQVe
rBSvvWcI5N6RFMuxfQNbDYMk9ux9P7fg3O7E2MKjS7fEJ7KYdZb9dDAkoz5rhOA6ftfFYlLGHpOD
i4/tFw1vQQ9f2qKr8i4QPluq/WkIWMG6r570njI0EvZg81hmoABU6aE+ojxucU/lzgi22V0EvoEY
bUJukFzEqOa4NS+24GjOKm+82aG578n2kXBKMxtHTywhxHeHWG0xVRU+xAKy/TPBmJBRk9WuSRfx
h0GT9mB4zOzUT2EFpxo4+wKIG5lhaH5Bx8hcbimMRFYJUqEmnGS+j0IljlsjZizX2h9iiFMjFGSC
qU/hw/mxu985PyqtdGzqtAzRSWKk5vmVg3V/RkZTBI7toHUCSph1teJm0JTJC8259qnzpemGz/eO
cNcZpkLdhRLLiJfm4dzOdMBlv6hdQsVb3QlUx8Faj5fYwfW6UD7oH0bYElwYwFb01g1m6jg0zBz3
1d8kRKl6Zzh0G6lecB0ROWc/eUpbPXaY0cyoaPnYbO3Myx6cf0idDvazGk6c9HCs6Q6A/LmNYIp8
fugDNcQ7bXwKPJqyvyuO75E/phqz8rK8PhahM7AxmoQCeoawjHSiCL20b7ZvY/zRGhWh7gKHq4+2
WSO9fqU+qrzb2/OO9ig9qaJF/NDU/8c26pTfizMPE/t6vihHQpRO9MiVptA0El/PVBRkCHrsmOem
+gKjT7MIOQBuGjimWllYQEiEmMzJLq7JutToQeKR8/p+h61dHSQTjEp8IQcnE6rt9xIgjTX8C7Lb
veKe+0TcOqBANyHGmD/ojOA/EbdkGnemH2FzuyaXIvkJRZHrgdY50Vvhq7x/Z7WhUOPvvXFiwBv8
rdp33OyzWi/NePuvU0lUnJqd79BK27N7K9NQZnZwmOsm/r/07RnPll7KlyRdLlt8eF6XirDv2DTm
DxU0pJwGWvNAPfjUzwcIrHVLl+Bi+wXStudOihXLr9DlL84XXSe8K0drKFZ84J/yf/iIst+JztRK
AgC0w97IciAUSjhsswUobbyKVB3+tQAdfb4YYr8uRTfBDcdilDXY6MiCt/ZCDeKhjLnx0FoD6vdt
JvTeizOBSS06qytrzVeP49FY2xJJeQ3c0NF8Si1Biud5UZj1Fskld2cQGGKayc3DGEE8lBCZthBb
WL3xEK6qFWHB9l8arhtJKmAF8d1jitkbiZ5vH+u9bZPSkuxJjFYku0Z4y9uSlZMTsIZHUKfj0HVD
We0C8E9Yl4Zw5EiJ89C0oeX7JfjaNcg1e0IdqUJ+tUHbvJF6XWvHa8XBud1s995qLW4ZCySS9+d1
c84FjFGV84Sztu7lByqBmtp8YmA/edwmShhhH4Mm+0mBEC99cQC9WIP1xs8aihUSeAUrB6Qf97nA
kJ1IC84bL1QXvRCij7g5y8zByTQGZHogynwVUoNrdRyrxWpRd4YKz5TrIATLdgvvCD90H9cC1aXA
cR6AyorDjse6t9cpkUtozXFsGF6C+ZPbGKcOT3MH4DPbKTR5MKHEw4DTTUfEV6yYMrOyuBanqz2W
TVvBLBQjqZTrTvzOa2vY5NSaIWvxpGJYZXr3Ayu4yxBFE5YppQwKlOYDwCKwgGnAVeVKBjgM6G4K
RNdgM9HL0gHzKDZgTivFt0IYAvx+brmCr8gg3dmPEX4ydT4A/b78V5tqlfu6TR73DIcCV+jDelQi
/Zo6df/shCQCvvWvc/t2RXZzvMIzSm8w/NxD7flRED8qupsnRpd2ekQ46PxoebfwG0f0yNsSOJ6k
oULuRj80/C6WweBXhTKVwKogmCghatwpo63lrsXRX15Bd4ZKRs5sffAC23f+d+D9aB+2PnGjQhFK
ZzWNG6jXj1cph5ERw71UGF6tAN2Eq1fJRXMOTRHndxT6usp+yuWrweUQ/qhpSmPLs/Frmq1Wr0Kg
ZHF6pkoYhhr7cXnZRQUpaBlw/G2YB4OokSR8s8SddbSVOI84aQHxD9M7VB35nSE2VQWMc4Gvr6O4
kOEVQvGUruwmKJ7EQQZcvwevH3VxYGEiww1GO/Cls0whAU+h0QrcX04apcIi7OSATLvjFVD+QYat
2ZOFQaCUA/eLSuri4czdl5MLlq9HW1Qy4vCFUIP4lNXiJfZxvbnFddXRfK5uw9o0cEx7r467VRs5
OXMJxmMswdNUqfPWdRNnrvAmfjfi6vjtmX2F9FmUdf7EkW3QFpmeGLWJ02YE5CHHm+bM5HLMEaJg
olD3/VrDgfVw0Kmyk2iJndryBl9eLc/z/S2hIZsFUm0vH8woGN7kB17XMcIvOOawSI0VVkVvhSs/
0l/XH4dXV76vkHNkxtu6oKMY5qf0hN1cG4lvBc1nutzBnWXVd6oM8d4MHFPhEUHl9xEYdyFZ1NEp
yr5ChE3fXb8tV3czm5RPZoXs9iYuc/+rTmLbISbDBooTZ5o8HGGvFiwQ01+eYh7MYtxpZY8UFodG
nsAkUxjleI91SfiCDbIih92xM701kuqDPaJXiA/++5Xlh13wD/DG7VVN7uFk43yhB3rcLDbxwg61
UYO+XVdc0FWfDaxUa88zKvZLzhbU6WpwMocKJr9Qwueh3GjkV3t6RpXfBq8vzT42dHMna7uARdMu
SSktH87EyCN6VxTGkr89cPFsANQXepCH1hdxe7aIVpuGpT3vo5z2oOJgrF1a4/kvi8kD1pFh0fXO
5YjFDYC2OlzaKfMRtymnkr5JQbvF/gXeHyq+BNZSexqGMVop5CsMK0eH/qmh2Cpv1wxY1YMSXOkL
94StiCTI/eAp/SlJvRWzPgD12I/8qqUvEFmJkwLHHDoCE3lcq2eyiQTUBR820CcvHEm1a9RNFppK
/gHU5SzFyPIPPKA5koOhFvY4dvBQVTP37OtiOy9iy0bETB8m3EnwDod2VIsJ4Ehkz3Wf9otiCAGj
BPcO6L3GK2MHGbfO9HItg6RfH6+oYW8QlLuE7dOMyCtRnihFgt7SUaGxVyRFEVXgiuSErKoXrU/C
uxP2Gs1lsE+78xkpuLcLXMwXDtwLiuCd9g5XeHBMuz+pPzxOdvsBaWDVZQ6GpsFsO0Ft5PGsBZ86
DyoDoTtzj7Lya2PJm7z2n+4dUE33+M4iWI72zX0wS5/tvweXOOautgiLee2GO/qobbSOqNoQAtEp
jFBBwefEUxNiIZ3/X5bAziq4pxq+XzONYuqAEqT6tMRorvXI0rMMuvsUPJf45cROT6WEKkfOhFuz
aUxP0xJpMhaAU1aUyUxuRNUxvzErP8ED/vcyxiWDHujWygf6k2E9igMKjx4uwLYQ9Ui796Uq3UuP
cI3XUfc7JjOkZMtwUoD689oNAV5MWTIPT9aV8oJlRYZjthyP6Ur0H93B0XoEtuLLNFtxXYEOSMrw
4MFHJCl1Hkxb81VvMnJYSOpaxcf/XmKy0OQ9BHVi6uaVPelIoN5WYY2uxnPycyMQShqEVNmvdFSD
ZrP6DBN4NmnCfF+M7w9W1AxmcLSklg41jQ108xFUYHuTLBemf/ABW92L0c6ZzSISf8g025FTgGnE
fsL12JOLpz+xf52Kcv0VjMnCxzkoAm18FxoMvv2yV+itsHJ4Hqa6d7M57CsBsdqxAzWCKziPIeNz
5gjeA/JRtVevdIflFssa0+hIwDafKPmV6WwkvxAjI1hoIPgHn+aHoNTVTqzqA/vx/8CT+dxOKTQS
iCaHVqZ93HtYFQS64jqFBDU+QRBt0ktzgJyVdIZFlTQywIQUOu3dXjVxAMJvG9P0OGKZ9sKOY5Sd
u+Jp2CkVX1IkdR/iaxmkpJM+cbbIsD8reJ63MP6zBxJEfk9I79FAr18FmCf0dWMB96gFBVnHrl46
QY3onJKDboziv1VvoRO3oIDfw/wysRCoCpg1YAtoney+CMfPttAinn7q6Elt6pi/B6nwbtW51J7s
VThG2dCxd2oM3IzO8KJiiKC831fLVlpXRdoXP2nhlKSsDDDFxeMqHpVyLU8CQ16g/pdMSe7EpM4S
lqYz/74INKzFRednirc7m7cJsRu72RRTcGyG2tiPA3D9ove2ZgPIeAKle9XyHf7o0HRYPkPuNE/S
OunNFM4wJKsLO61U5MMJDVJcRa3eDkx76qSV9wbh7StSpvVE9ym/zkiIQG4u/glrLcWodmJJYTW/
ts3qv7K33lqobuRDf+jEbcNqLTNHIIOIt7BZpRpIHrc7N6jj0nlfvQ1PIoDC7t/jiTReQTNcxu9T
QhP05ET/+z2ZvtLuPz4/TJZT+PeqiJE5K4D62+vnc0ubBiIt5jNS5brA2XqL/mMPnJ+c/9IsbehN
Pt1x5ChuxIyIQfonFfx9b8/16riAlV4yCs09fJC/T0LvufYlYAYmp6l4p5iYuvHyGaSSukMwKTf3
SVqFctZrZ/9xm6gokU560JeTtP7fvak4GXcR1gwDpwAyyCXCXJQuhoPYrjnQ/o6Txv0h2+B2oEvI
GQASJo/P5yEjSXf/MSM9vEIBAjblEf+gwK7xmBZw0JhlUVYM07YDl8rf21fuv00N2i+eOphhHax5
TTj4j6i4JjnRDfxg3MQYKK16B2MTYMQNWoVvQCbPGQyK33o6/rIAXRu0y14TTFTcF/HXq1bWWxfg
g907a05Ip69nGGOtWHHB8rYfxK9PxmTvQrieI7B5DwLczeBywmzOqIcemIQofPdi8UdBPFQm+kvX
q3rk4hTOx0aWO2+iYTY3dSt/Y+uBxA+eLCA050NFZhxzC5+E+nAU+RjrRKIAW1p4pb4ytOCeYqFp
g+bKw6E4ZOH+b0iLRLxq47CHmb0v9zPRMU7ZF7hfnGqXjt1fCnAT1TTF11KmH5gMACOEBoAKzgL6
KsumR0JflDiLLb2kiWMUgRWb20IQfdKOt8RACfA3BYZoOkYXmvPlEKI7wSa/by6vsh+Md9FkFrZN
6L4WhSIFpcl0hlhJyUf21TcpILuD4sy3jtRMF0rMxgY/Ff7da6rbDrzNCfItDQbyA+h4s1NAN6ul
03N2fRr8tC02DidQfZnH3ptxNATXTp4mUhxvFtNKXq3ejiyF5GvF666Fg/muUuCsuM6C0XCH3EPh
4Xln/D1QYENN3ulMLof4CGPhqVGKhwGjjzJ4z8eOS5V78CORs87hY9jZPghDRULJelhWroVkGzo6
ju9jjsDW6P5jdiBqRDnYBAfpImBD8K6GmY8fWUbSvRocSAmpag6nbfE1Z/MuMH29bqpSknOlS2E8
l91lzAdpOgp3sNmWrcwj0lP5EcfZnL799mx2QgKrBAAs/sCccihhQHQB3yyCxCg0QmTidHUvMiwH
UxeQ/HJJj6uPZloHiV+78EN8qQNVHgwBsCv2DGUYevEh489h/IDpz8yOyOi8dcdC5UfJ6icwL9ln
5NXx+P48th231J6Lig8Y1Zek0Atv3lPOdtdGfL9kotrYEQSBTNXYqgZs9l5KIIwEphCjU4pQkfSs
mH/doKtmTI5WHGkAWBHxytCUgynrGPUOLidbncprp7hCO4gOhG50wJvG3tMIGxyRftG0HC+lkifl
Yx9Vhl1OOkZAeRZ4eyYwJqEHrhK7KGCMGStn4BHogH7oQHsoOZhz+JO+K0XzM+gXwrZXjg9deGKc
Kh1spA0V2CNNs/pZZXMCLhmaE2pide8OEBFIsHzsjTk9NIyJNvB8c79h6VrP+oEExarM6s1Ldxnr
Jdvpw+buXpSQddt3a6X3+bntYIaVJsmjj6TIcYhT3bxuLXxb4qf4EeaPgLFCsP0VQOBJapGaTE5E
gt7qhzOJkNUy2pNJA5hq3ZIKr0vKN59o5maxEgWMCmYjUy1cv8wttQu5P98wEtLGWrYAdc09YGJs
Ym3jqNZnzGUgcfSP7F+yOnFYYARmMzTaXmUlNFDev5jKyowSJIAhpbdIwyNQkbTr8DvyU6d5rDb1
vuL3d4sTLFLQfE24gzYXtofjdf/m8TKgi12Rrw92Cujqa3ARcB03IzOLnql/hS30wHqgPiwJfBPP
5829KZ0JF++cdV/nmAs4QBiDkkF6laHi6AFIKO/VEnCyRYxpzxyt9SDpxIu0cDo6GJEsSBPOGTJ6
/OG/d2Quhwt4WnDcT+GQt2cbRHfpdBaMnRWIrSTJlv+EJ1mElR3AzwWte9Toaz3/0DGX8rVsku5h
HYkU7wVnfRHpl8F52h/4rwghqiyRmrciEag2Usac1xjovAHhkGF0n41deXgFtXFhH8pOdzRko5IV
q7475yUfK3f0brD6/E5fzPK91HnX1GW2n4VuVJUUrOlDUf1vtAmrfB1Ga1UIoKLMme1iVN/M8fa3
Nb3dPElno8CIw6kBTNgUCWTCdyyOkxiXhedB0U7P3aCJgnJN2QEOvWFujREIdBM8Mur5jzwhaidw
P5srWQHcpAflY6iTaO3d/VPTrhWBpCeVAozJqGYkoR40sZVETTDJeRyvomUZWMcB/2GIOoQK0KTB
WyPg4tvn1S1XzNj6VyiNOyE+DCJCjw+gsi7CTDE3PEOFJex/uTUhBTAIqdhAFE/CpRs8N7ppmENT
O7h4pq99xT2FLfrztkjAinZDZln4+M0kC9rv4DfusU1SWoTWxozx4bsinCntMnwc88EiTmnyI5uC
8XMAtYcVwSbeV7kmgXw5E0RVbI31tQIn7jy/77g0Zp7trQ0rXe9bYveUdk9Pjrq3AN6mRCCzHZDd
q9QhxER6Gh8HMVY4VF0I1+B7h3hOok73bWy2oqZCZRX+TndgSHuEbW6QMOJejdmYm4NOrGzTiiPl
IjluZLqHWxJQ8WXlybrYF+JGemJweHooSYUBGmrLLTeEpYwOQijvhlVBbtwtvgoOGP2Nc0Dip7DM
FKUDt3y5e6npW7aSRXzib2MLPuKbfYlz5AMon506KZWulnr8oNt++wlPxz+N2NvAginGsywZUDgO
Q0LAN9CU00KOjwdN1xoasWdA/6aAxuijW6NMKixE0RkeLXN+WMm9aUS7Ct9nPkuZCzR06SijkbZE
YNWumk/eowtnDDkfwO4fayHTdlh7WyTbFeFMcMzXj0lUNEa7VvWbcLzDG2TZEoYWz12P2ikWq0qF
laIlyJmphWM14Ym14AhJAgTVbFjkv/s0UFB9NSOQLv2lc/x87OH9ZPVTHwIO5Y+0PWNVcknaOsZ4
/8DItb3dDZhlx/VYgv8WfJIj43mYk3MNQVR5rKjwhC53siUptRy76zPDRZGuVr96rYfDP/0dXO55
fzUWt9Kq3sUU0WGEWTS+1iX5Z0mRuwutTIm0Y9ay//7TmqBSqnvFi3rFPrBKNd0+0ABiNDUMOLr8
DOFFAUoVJUpeLhSEhGEEATzGT8hvehayvNRWSsgr/g2Nnd2QYvF06vbZpDIsjA1d+vk6Ryl95sgy
kdMafrOVnOnKQuk8c4o91swEkgk08PWgXf4PYmLf9cceaCBb6FlKmfSqq2ncfS0pCd7mk2WsVbFC
NjiGbphqBA2IKTqrqat02E+2g7+DFcg8HeOVixh7hOli28un3qZqkTZS/tZb2YpNfcGXOad18jyQ
ZTWDaFeTCUgsCCIByh3k6hhPlRUG5ltG+dS1SLjHfkeMdgd3DChQWTk4pVLpsdV2pVZgAyaHQQle
TyYA1DasWE4YThCCm8ltTKn+VuwiLb/Mfi8Pn9Y+v1EDqBlzl8XelZX2KGoj74W51MEe3m73gvm3
TpOtHUDIHPdh+T5gs3FlckHy8AJq2v99nAWJ/Ko8DifmovG218i2VmRR7ZEx+MxMaT4zK+XbubEW
f5Npti5a40DCByYjEXSFM9S5Jr0O/fuJqjVMZlJo2SBg0/3FkWHs39VNVZoe2FBYSGXaK8jkRd6I
56qKcHxVeLv8c8uW6D8Iqw10baAwntdRZXzNPn8ItwPHbmikLJYvyKbLY/8329AwzvyZf32Xh9Qc
LC/atH0Ltle+ZP3yrK7kezIukfLFxrScilVIaA5AFGnTyQW+bKyXU8vHD2Jm4CpkXf8zVdIxH5zM
u3evu5wc4SR4cP1uC6YZ+0U5UGfmWTK3jRj5oRF3I86W9QdxrIOpPtCCQVgUHPF0BpdEwHsTbgz2
zabdVM7txP8XZ8j7SpmwjBDP/WA+dvHT/suNk2ueFFN2Q5/BmjTfzvuyX3X/8HLd3vKPFp20StBZ
F4PZ2dennnCVqaN/avuOtNk9fwK5/a22yuUxed278XJxMnWrhnU5EYJ1Cx7ZakIgOfM/2RsEM3zW
5i97ai+WBJ89V9pA6vgoX7IwwNj3TyioJ56T8/DACD6ojtbwilvPHsj5fy9QT3DuMRWrnS79K9dn
lFfNT8EhN1xA7U902xH5YjAVf7vHnqLWIjfFqbJol0TPpBTGCH4xB+ayFn4l/pscNbjmXzm10Bhv
iekZrxsvl0mCoV62KaR0ZudyiD6bulKJiIfP37491hVOuQfcuFs0ZZYm+5VjC/zb0oc6aECTWlbZ
dr+v8Wb9Sh2LqoOtwe5ivq0iv1pQ2xQrktqpf4W0weQ2Bc7SvNeTaqA/5PlMF7BKX0hbmcl8nS2u
gx1pond0NMd1pPxmozO4VGT+FeujgXAC0fv8nwQROR0bjWvaxTD8k7MMlIpBdXrjDExIiKadzwoS
Mm+FfMyZTCDFeugIp9X14kxzWIS4bGWV8UsP29AWjy/B3rFHyDaPQbsskrULuaccWfkVBCN6KXXH
5xMxNyQWdDhRzbaX+WMb9urQBGjS39oqbhe4Q9MrHunV802i/ueNvn/Eyon1YtvUMOADdxdscK+T
0EDt2fYPlEyPhbxf8fxRM0Cj0FEWc1vb0s+TmxdBWIe72guTfyCwmJFvoNJbuDxP0xa6fbJw61m1
1Bf1OqFCZ+1uXSmn6WlmjOz88cVB95HhBZq/jN0Z55wO6vuoARqfQWr3ma9Jc5+YxreHEVnkcdSi
kXYF2CqGUHVGFatUUmSf9L4xEhlUxeUJrULeFEApN6rpz37Z/eC025GJ5Qtfq0EUuR9IRVAYCiJn
rm4sVnioABXrGdYvFJXmSjNmYqF3JglZ6XWK2xzzZbwKW9isFvutUC0sQSK1uojwYnM2G6EFhJ1H
iYCvqrSBQ3/ZfQUOYmUZkOIc8Fty1h5rO84hCR0xjkZ4lQuU//OfUnXydSbz97FPXf5Viz9zRO6m
sJlHbgvB2Sw7rCLCn80x6TtZfL7K8/34IyYb9JFM04p3hxFIM9206zjvoKnueOrcR3VRlunk9SXN
zEDQ0EMlya39V0DRzP9tV2t8kU9pYrPWdnxD8R3FCX67qWHCwTbvdZiQjK8NLHPQ6sqFjrEzzkl/
2XOIzR6xWRYecirkolkGzBxnYCZL6l+qIC04Vor65AUfATjGCChdZHa4L40sAWej11qzwXOvXH2L
rGR8syRZGimgnOGFM62ikp2zLKMz4ed9FvAK9nqrPmb53Y3U397NGSBvlcG4gqbnYDO9Asmenx3Z
iuDrex6Haom/IevmnOR91alXHRCXPXjaeSGK/aI3LavEofFzUGYULwWYiHxMdH3JYYOENXQYPxKI
S/fCc568TTrOGByhPv7vgk8ZmEublL2JW1x/oOT8loMxbq4bVUNo/yJP9MMShTDIJG71cV+asEZ5
RO+7IhDnqzU3Q9dGKqifDHKLpQ4KSAOZYNEGnBv5sod/8/b1jO7kOenFYkHw0UjcbIQCz+30EAu+
aKe//GKyKmbJ3loUz6+yJ18/gItcydYrX74ADh/RLhfpjY7UqmUfOdblW9xe09QaLCojrslzKxcZ
x6whaMp82poi59U3Sb6ZJ+8wjCIjVVeas40RdQ8htby2LDYp08Q55yX8KmXu8dhIwFADtqMzmskQ
nn+CBMIwDpyVGJcOqKF6d9bUj8M/4Ak998DiAaBRPLLV1mU4cBQQzw47ZC7dW9JFgTQV9vj6M6Rw
YEQ85nUO0PEqKroXeQoOKODIZrvU7QryukM/v46kwpXt0RUpXFj2PKTexWcBMDHu+nI/n1E4caCf
6g22r1uaTsktpp1M0mFRUsVVF5s68JPJLqKVzjVxZZJjCT5WRThrMsLdo2IYPWT1PGXw+xupu1qi
c7iCgQTAXFbBTklsVFg+X5qc1cnNF8qMxSgskzQ9V09cuTr8GOZrVZ2BA6ZvpaprzCSHhskTcjXs
l6FMtGsCSvP4+bosbJvMabF7ss7mu1fWw57dlF+mITei3uGWyYV9MPjX+M+2AgxSZx90LNfoA6Ij
gIzPRgy0/3UwXHeFyGZmS8IN9d2JfdUTf5xh3iwMM1aERRZrzBhPipeaHeJ3Y4G5gKTe1trt9oJv
ng/2HoFWLVvGv+O/ojBNxVlrnXEmI85GRe6CN7n3vj2DLeXn1wYtLhxPpPw07d7VB0bHBWbwnizV
nSwpHBxnNFhN7M3kSLfoClwMTmcsrTESYU4mMWBICw8dnDBonk+OuDhogLeh73DQwljq1rLiwp/c
ZfAu1XXHeFs+zMEfUUnUp7g4ztTynqPMF7ZvyDBmz4Pn6YlDFiY7v/0Lrowr9a340nUvSgvjiLAE
CA7TYYxl4zYhuTOWZLPj+dhFCc4m/KY91eIQLaeONXfor0KWtvtUyHv6Km0X/Rgg79Mwr5mLo7wM
rsAQn4rDt4Zy7WA0kcNxpTBAJKGyygdLLglvmFqh01+Ajg7gF5NWMr1Q87oFsgMW68JST3+ZwyRc
YMBfevse8CENLePDh3KRYbYpYMOEDA1jb4wr8c8MCuZTDo1cImGe4s+qaEsp1FaBDOumFSGN/+/+
M62Dgsx9h1Lo6VVFTrVbWIAc5eDXwhxxcd/nqSiJJolLvTlRC0TSA359R9DSr99Q11jGLpnq8aYD
v0zPZzS7TfG8O4nztk+YDuD218iFG1awfCMEbkLis8E42zA4PjXqJUc/+BSVzzcmJFDJX0hpBMCZ
YeZvp0K1Jj5s9rbjwrHRx4FjFkyFlRLnu3+UqHmwpP6Xlaaiifo6x1aucpFLJsmnwrmnFVf97MCE
S6DOs59BqrzJd9+M/fIPpDVJPYp4yN41oSYLIyaz4k/LybAjNerouVxgWcfC9oqIW7s6dQNmEjSl
BxAreMNLMJOr5mf4WDH0oumj1R9uT8YfwtnqTAN5+dvOB1xHGZD1YCwGyHRF1Hf2M8/j+swspHIz
DV1J8V6+ZbAiOJuyJkT7wRECf+pkl0rwpDho+Y0grvYKymVtmzl9sJEZclOTel9GuZOTb9mAZ03c
toTGNDpwdjJqFlGxt30iZWBclsaXoa0Hv4s1SnwTWNbd4yS8cgT2WOiy2WV28e7b4f1VRZevZZoL
aL9myMpe8dGhtuc3Qam5n7XuhyXJVAsTOHDUjSZSQAOiiG2tGtZxUDQUFxEAiPbdjHoBXpeDNODE
I1+e7q8Cf/8UoevUyG0K8nIFl4AOf6pHloJrWC0fC7aTUwlzFE9ajWqJ8WVm5AesVl+RiEPuVtaK
YngWy4AwVipHZrZxG4gLiUlTu88X6jOp8ybdd/2LzhSWMxRg8O+OcxFUODOs0Z4HStjc5YPJx3Hd
3DivUwj4ZNomnxwz/+mFXkR6IxLjLlFgaMzaxxcmz1IHfxS7DlDZPJYT7PaK90FG79r1cGwH529u
/Nci3mTr2/uqv9C1ZfjwovTGmfxi8x+wv6HA0qMXdmr6y62aKUjEvdoJLZBm2JDgRjaDh2GpSKBE
zHw2RueFlGTVf8Nq6rusCtsguZz6MgQMZzZ5m1RAyzt7VfykJQ3gywAE4epRgx06M7L59niEUt2t
x760c20TcbEE3eNaBBD9URXrehuz07q5w5Oyh/6kAxPSiX5zYUEWhubdNesrEBKprQWrbPM6oTtE
tkYd7SW+s/NxWCWGQR1LDbpPMqX7AF0SwSp8Ho/Nk7Xrz+RydN8WQmvybYtsUKwJTYBZwRv7QrGI
/JsGxPtyc2GAZvbYHzc8iwJNWraDpc2FIaW2EZX6auhEfFgFVPKnb3RVpTqZzDrV3As3D/877rl2
x3plWJLkjtmzuXhOsWlgahlG24Z5gYlMUPoz6SzYaFui1uLiNlaeS67xsEJYPurJrntK6piODElL
0rRoYAxdWYmvQDtW3M2nW5BJkgce2CoGiVOqTb/FJbhd6ZId6HRHep+Ibr02b/lNaBDcT8dqm3+J
aVA0VvfxPGful1W3yu/qMe98SmMfxkvg5nI3vMgyAtMpx9qI+rlFW9Ko2lvsT2ZnsOWArG8HVYpi
l/dGc49EQ5twjS4x6MQV84Qs8zK45/Womn83WaWb+6Z6d/rDAxQM2fOdYg73+8rI1lup4uUS+rYC
9SP0vluX0NLfSdFno5MHTZ4Y3J8g6k/muc6AndBowe/F8uTYpiFfIKYlXd9kIKaKL7qcHQmjDYct
PBwvZ9O5rvCkVemiEDnNlqkCbPtyqsZ5m+Vj5I1PSM5WZKW5khgcjRjwbvKf1PurpVPo11fGd9z1
ROAOHYbzHzF35qHVcAE4vRTy0wT54mtT34j1Gqp31gTwjjrtBk8AWyoAoZZqcTcqITbnrSQbjNlM
XqPfST6mOeiZfWBX/tDmtWfiZRg7uwgYniOnAWagsKaFY0uSfeY58CMr9ziyWym9anIDGQR3j20J
Al8Jza6Ti4ez7PgrkQEKAmEyi8XCOQAE4Wb7pKUM5nbAx2p2Zks5Z71Drqb8oEv7OYa5Z66hnUlK
tTdYh3UX4QxiEs9m6M+x56N4yW6Nfir/LYRUy9QTgH83WcpByb5QOyYVSv5UJzhfT/tJXzcmTfm0
4x65NH8H60nmCUt2hin0f5iHC3BlOjurzTt9acviki0Xj0Thzt8t8XtXxNzCVamwvtRwO2XLWhej
RhP3jVUMcGLZKpSv1TsuaOtEAiHn+51qJ8xET+0rSs2Q2e1F8V1dbQjPO9dm0/90OMWA4UgmJR/2
y+8F6KUCirolYzWnG8bzH67bMQXFiXScSbAPOAXBeq5WjQRlckj29obl1jKBce5LR+ktPoNQ42kO
VacTCzpp6wZN5sqOb0/4SguBx/bLR4zOXRJ9IGv26dEWEFPluQZhyN0TJ1LgvHi6bkkS2liI7cNi
gem0xo6dMq8Gw7++2+WU+KirtSC/KyMcVvp4bqfzjn6IV+Sy6rymlQ5Zri7AUroodgnmVZQYMvy/
ClAXqXRUT9OhG4/Ve5goqXwi8d9cYZUF3LuLAP7ODelbaXPBZICRa4dEwWamS3J0OiA6uwTVrHmb
xiF+gDbaJwacUi7fP9zCtyjxClkWROy6C9EGFGogZ9U877vzJGhOQEABDJhRjf/H1e5iuNig8cWh
B20z7pn15Ofhgggu0LEVuPM5DrHO3/Nv1DjZKEvICBdLyPuy4Vang0ZJUdOKKGZAmiDqER7M3wFJ
r0qDyR9o2K1OfETLM/kTWZs3lp6i6CMNPr4h6Qln1LtAolj0MuVG9BcDTlPomliCsOD8oWGx6Vsi
IS9AWYm46o6+6tmWmlpLmdXhPS1nOOw1+s803++iWr94kE44mAC7gTHl9Rseuo17KHd6cy3Fexp5
sqtoXpOcPurXDEx6ng2umWuBP5+U9rAjx+1n1/5V7Q7jfboA4Ffxo5pZxrJPUeBPlqm15UT5LD6y
iAiAlqnMSEXPpns39BhtSU9XMWIej672vbh+0poaAEBJzHuU5mduWoW2g93LijI5OYcumiJSTBzl
PQRHItFFCNR8Yyi9TBFs0WIHSGyRdFTMUBx3E4WwI0Mhm9//arXNHnDHdkzBpaXtgqmuBLT+vOHY
43rY2EsaXl21tDUaECet6YgxJW+5AZ8auQ4wauhGVyI0XivKP+aoVsHWpEFn13f6b7flY/NfzMF4
7MAIZzIg3L/KlRUOpftAj/jOennlHfWSEkyVBnR8P2I73wL2nKgRpXmaOElZzG0//RPmAmGc3HqU
GN09DOK8UDz+iEga3SSowHKcHV3tZC4vyr0soFMQCYPCoI1Es/LHe1PnCxGVRLztuSpQoqQ5uhQV
nf/RPSiZKWSLsw9DzPUG42Oii5qWV95iWjg0kYLN/llsQcisTQ3BWab0qHhYrskYZjaEO982koY/
kXmsGi6i9ICDKMkTw46TKC/cx1rknWdgqDbf0OdeNMi2SjmTG7SxyilJbBfQZWehhBlrpUYv502b
q6lesvg/rr4J+HTFwnU=
`protect end_protected

